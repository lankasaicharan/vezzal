magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 1490 1975
<< nwell >>
rect -38 332 230 704
<< pwell >>
rect 1 49 191 248
rect 0 0 192 49
<< ndiff >>
rect 27 116 165 222
rect 27 82 43 116
rect 77 82 115 116
rect 149 82 165 116
rect 27 74 165 82
<< pdiff >>
rect 27 584 165 592
rect 27 550 43 584
rect 77 550 115 584
rect 149 550 165 584
rect 27 368 165 550
<< ndiffc >>
rect 43 82 77 116
rect 115 82 149 116
<< pdiffc >>
rect 43 550 77 584
rect 115 550 149 584
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 27 584 165 649
rect 27 550 43 584
rect 77 550 115 584
rect 149 550 165 584
rect 27 82 43 116
rect 77 82 115 116
rect 149 82 165 116
rect 27 17 165 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 31 -17 65 17
rect 127 -17 161 17
<< metal1 >>
rect 0 683 192 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 0 617 192 649
rect 0 17 192 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
rect 0 -49 192 -17
<< labels >>
flabel pwell s 0 0 192 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew ground bidirectional
flabel nwell s 0 617 192 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sky130_fd_sc_hs__fill_2
flabel metal1 s 0 617 192 666 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
flabel metal1 s 0 0 192 49 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
<< properties >>
string LEFsite unit
string LEFclass CORE SPACER
string FIXED_BBOX 0 0 192 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 1264858
string GDS_START 1262908
<< end >>
