magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2494 1852
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 880 157 1186 203
rect 1 21 1186 157
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 131
rect 183 47 213 131
rect 381 47 411 131
rect 469 47 499 131
rect 577 47 607 119
rect 665 47 695 119
rect 760 47 790 131
rect 968 47 998 177
rect 1064 47 1094 177
<< scpmoshvt >>
rect 81 363 117 491
rect 175 363 211 491
rect 373 369 409 497
rect 467 369 503 497
rect 572 413 608 497
rect 680 413 716 497
rect 762 413 798 497
rect 960 297 996 497
rect 1056 297 1092 497
<< ndiff >>
rect 27 119 89 131
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 93 183 131
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 119 265 131
rect 213 85 223 119
rect 257 85 265 119
rect 213 47 265 85
rect 319 119 381 131
rect 319 85 327 119
rect 361 85 381 119
rect 319 47 381 85
rect 411 89 469 131
rect 411 55 421 89
rect 455 55 469 89
rect 411 47 469 55
rect 499 119 549 131
rect 906 133 968 177
rect 710 119 760 131
rect 499 47 577 119
rect 607 107 665 119
rect 607 73 617 107
rect 651 73 665 107
rect 607 47 665 73
rect 695 47 760 119
rect 790 106 852 131
rect 790 72 810 106
rect 844 72 852 106
rect 790 47 852 72
rect 906 99 914 133
rect 948 99 968 133
rect 906 47 968 99
rect 998 127 1064 177
rect 998 93 1008 127
rect 1042 93 1064 127
rect 998 47 1064 93
rect 1094 133 1160 177
rect 1094 99 1118 133
rect 1152 99 1160 133
rect 1094 47 1160 99
<< pdiff >>
rect 27 477 81 491
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 363 81 375
rect 117 461 175 491
rect 117 427 129 461
rect 163 427 175 461
rect 117 363 175 427
rect 211 477 265 491
rect 211 443 223 477
rect 257 443 265 477
rect 211 409 265 443
rect 211 375 223 409
rect 257 375 265 409
rect 211 363 265 375
rect 319 483 373 497
rect 319 449 327 483
rect 361 449 373 483
rect 319 415 373 449
rect 319 381 327 415
rect 361 381 373 415
rect 319 369 373 381
rect 409 485 467 497
rect 409 451 421 485
rect 455 451 467 485
rect 409 417 467 451
rect 409 383 421 417
rect 455 383 467 417
rect 409 369 467 383
rect 503 413 572 497
rect 608 485 680 497
rect 608 451 620 485
rect 654 451 680 485
rect 608 413 680 451
rect 716 413 762 497
rect 798 477 852 497
rect 798 443 810 477
rect 844 443 852 477
rect 798 413 852 443
rect 906 471 960 497
rect 906 437 914 471
rect 948 437 960 471
rect 503 369 555 413
rect 906 368 960 437
rect 906 334 914 368
rect 948 334 960 368
rect 906 297 960 334
rect 996 484 1056 497
rect 996 450 1008 484
rect 1042 450 1056 484
rect 996 364 1056 450
rect 996 330 1008 364
rect 1042 330 1056 364
rect 996 297 1056 330
rect 1092 475 1160 497
rect 1092 441 1118 475
rect 1152 441 1160 475
rect 1092 384 1160 441
rect 1092 350 1118 384
rect 1152 350 1160 384
rect 1092 297 1160 350
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 327 85 361 119
rect 421 55 455 89
rect 617 73 651 107
rect 810 72 844 106
rect 914 99 948 133
rect 1008 93 1042 127
rect 1118 99 1152 133
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 427 163 461
rect 223 443 257 477
rect 223 375 257 409
rect 327 449 361 483
rect 327 381 361 415
rect 421 451 455 485
rect 421 383 455 417
rect 620 451 654 485
rect 810 443 844 477
rect 914 437 948 471
rect 914 334 948 368
rect 1008 450 1042 484
rect 1008 330 1042 364
rect 1118 441 1152 475
rect 1118 350 1152 384
<< poly >>
rect 81 491 117 517
rect 175 491 211 517
rect 373 497 409 523
rect 467 497 503 523
rect 572 497 608 523
rect 680 497 716 523
rect 762 497 798 523
rect 960 497 996 523
rect 1056 497 1092 523
rect 572 398 608 413
rect 680 398 716 413
rect 762 398 798 413
rect 81 348 117 363
rect 175 348 211 363
rect 373 354 409 369
rect 467 354 503 369
rect 46 318 119 348
rect 46 280 76 318
rect 21 264 76 280
rect 173 274 213 348
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 128 264 213 274
rect 128 230 144 264
rect 178 230 213 264
rect 371 241 411 354
rect 128 220 213 230
rect 46 176 76 214
rect 46 146 119 176
rect 89 131 119 146
rect 183 131 213 220
rect 318 225 411 241
rect 318 191 328 225
rect 362 191 411 225
rect 465 219 505 354
rect 570 337 610 398
rect 678 375 718 398
rect 547 321 610 337
rect 652 365 718 375
rect 652 331 668 365
rect 702 331 718 365
rect 652 321 718 331
rect 760 373 800 398
rect 760 357 858 373
rect 760 323 814 357
rect 848 323 858 357
rect 547 287 557 321
rect 591 287 610 321
rect 547 279 610 287
rect 760 307 858 323
rect 547 271 695 279
rect 571 249 695 271
rect 318 175 411 191
rect 381 131 411 175
rect 454 203 508 219
rect 454 169 464 203
rect 498 169 508 203
rect 454 153 508 169
rect 567 191 621 207
rect 567 157 577 191
rect 611 157 621 191
rect 469 131 499 153
rect 567 141 621 157
rect 577 119 607 141
rect 665 119 695 249
rect 760 131 790 307
rect 960 282 996 297
rect 1056 282 1092 297
rect 958 265 998 282
rect 1054 265 1094 282
rect 842 249 998 265
rect 842 215 852 249
rect 886 215 998 249
rect 842 199 998 215
rect 1040 249 1094 265
rect 1040 215 1050 249
rect 1084 215 1094 249
rect 1040 199 1094 215
rect 968 177 998 199
rect 1064 177 1094 199
rect 89 21 119 47
rect 183 21 213 47
rect 381 21 411 47
rect 469 21 499 47
rect 577 21 607 47
rect 665 21 695 47
rect 760 21 790 47
rect 968 21 998 47
rect 1064 21 1094 47
<< polycont >>
rect 32 230 66 264
rect 144 230 178 264
rect 328 191 362 225
rect 668 331 702 365
rect 814 323 848 357
rect 557 287 591 321
rect 464 169 498 203
rect 577 157 611 191
rect 852 215 886 249
rect 1050 215 1084 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 179 527
rect 103 427 129 461
rect 163 427 179 461
rect 223 477 268 493
rect 421 485 484 527
rect 257 443 268 477
rect 223 409 268 443
rect 69 375 166 393
rect 35 359 166 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 132 323 166 359
rect 132 280 166 289
rect 257 391 268 409
rect 223 357 234 375
rect 223 337 268 357
rect 311 449 327 483
rect 361 449 377 483
rect 311 415 377 449
rect 311 381 327 415
rect 361 381 377 415
rect 132 264 178 280
rect 132 230 144 264
rect 132 214 178 230
rect 132 161 166 214
rect 35 127 166 161
rect 35 119 69 127
rect 223 119 257 337
rect 311 333 377 381
rect 455 451 484 485
rect 604 451 620 485
rect 654 451 770 485
rect 421 417 484 451
rect 455 383 484 417
rect 421 367 484 383
rect 534 391 591 401
rect 568 357 591 391
rect 311 299 458 333
rect 293 225 378 265
rect 293 191 328 225
rect 362 191 378 225
rect 424 219 458 299
rect 534 321 591 357
rect 534 287 557 321
rect 534 271 591 287
rect 634 365 702 399
rect 634 331 668 365
rect 634 323 702 331
rect 634 289 635 323
rect 669 289 702 323
rect 634 283 702 289
rect 424 203 508 219
rect 634 207 668 283
rect 424 169 464 203
rect 498 169 508 203
rect 424 157 508 169
rect 35 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 223 69 257 85
rect 327 153 508 157
rect 577 191 668 207
rect 611 157 668 191
rect 327 123 458 153
rect 577 141 668 157
rect 736 265 770 451
rect 810 477 870 527
rect 844 443 870 477
rect 810 427 870 443
rect 914 471 958 487
rect 948 437 958 471
rect 914 373 958 437
rect 814 368 958 373
rect 814 357 914 368
rect 848 334 914 357
rect 948 334 958 368
rect 848 323 958 334
rect 814 307 958 323
rect 924 265 958 307
rect 1004 484 1058 527
rect 1004 450 1008 484
rect 1042 450 1058 484
rect 1004 364 1058 450
rect 1004 330 1008 364
rect 1042 330 1058 364
rect 1004 299 1058 330
rect 1118 475 1175 491
rect 1152 441 1175 475
rect 1118 384 1175 441
rect 1152 350 1175 384
rect 736 249 886 265
rect 736 215 852 249
rect 736 199 886 215
rect 924 249 1084 265
rect 924 215 1050 249
rect 924 199 1084 215
rect 327 119 361 123
rect 736 107 770 199
rect 924 165 958 199
rect 327 69 361 85
rect 103 17 179 59
rect 395 55 421 89
rect 455 55 471 89
rect 601 73 617 107
rect 651 73 770 107
rect 804 106 860 165
rect 395 17 471 55
rect 804 72 810 106
rect 844 72 860 106
rect 914 133 958 165
rect 948 99 958 133
rect 914 83 958 99
rect 1004 127 1058 165
rect 1004 93 1008 127
rect 1042 93 1058 127
rect 804 17 860 72
rect 1004 17 1058 93
rect 1118 133 1175 350
rect 1152 99 1175 133
rect 1118 83 1175 99
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 132 289 166 323
rect 234 375 257 391
rect 257 375 268 391
rect 234 357 268 375
rect 534 357 568 391
rect 635 289 669 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 222 391 280 397
rect 222 357 234 391
rect 268 388 280 391
rect 522 391 580 397
rect 522 388 534 391
rect 268 360 534 388
rect 268 357 280 360
rect 222 351 280 357
rect 522 357 534 360
rect 568 357 580 391
rect 522 351 580 357
rect 120 323 178 329
rect 120 289 132 323
rect 166 320 178 323
rect 623 323 681 329
rect 623 320 635 323
rect 166 292 635 320
rect 166 289 178 292
rect 120 283 178 289
rect 623 289 635 292
rect 669 289 681 323
rect 623 283 681 289
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlxtn_1
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel locali s 1129 85 1163 119 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1129 425 1163 459 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew signal input
flabel locali s 1129 357 1163 391 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew signal input
flabel locali s 309 221 343 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1203608
string GDS_START 1193790
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
