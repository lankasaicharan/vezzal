magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 230 157 856 241
rect 125 49 856 157
rect 0 0 864 49
<< scnmos >>
rect 204 47 234 131
rect 309 47 339 215
rect 395 47 425 215
rect 489 47 519 215
rect 575 47 605 215
rect 661 47 691 215
rect 747 47 777 215
<< scpmoshvt >>
rect 80 496 110 580
rect 309 367 339 619
rect 381 367 411 619
rect 489 367 519 619
rect 575 367 605 619
rect 661 367 691 619
rect 747 367 777 619
<< ndiff >>
rect 256 179 309 215
rect 256 145 264 179
rect 298 145 309 179
rect 256 131 309 145
rect 151 105 204 131
rect 151 71 159 105
rect 193 71 204 105
rect 151 47 204 71
rect 234 93 309 131
rect 234 59 264 93
rect 298 59 309 93
rect 234 47 309 59
rect 339 203 395 215
rect 339 169 350 203
rect 384 169 395 203
rect 339 101 395 169
rect 339 67 350 101
rect 384 67 395 101
rect 339 47 395 67
rect 425 165 489 215
rect 425 131 436 165
rect 470 131 489 165
rect 425 93 489 131
rect 425 59 436 93
rect 470 59 489 93
rect 425 47 489 59
rect 519 181 575 215
rect 519 147 530 181
rect 564 147 575 181
rect 519 101 575 147
rect 519 67 530 101
rect 564 67 575 101
rect 519 47 575 67
rect 605 106 661 215
rect 605 72 616 106
rect 650 72 661 106
rect 605 47 661 72
rect 691 203 747 215
rect 691 169 702 203
rect 736 169 747 203
rect 691 101 747 169
rect 691 67 702 101
rect 736 67 747 101
rect 691 47 747 67
rect 777 179 830 215
rect 777 145 788 179
rect 822 145 830 179
rect 777 93 830 145
rect 777 59 788 93
rect 822 59 830 93
rect 777 47 830 59
<< pdiff >>
rect 256 607 309 619
rect 27 555 80 580
rect 27 521 35 555
rect 69 521 80 555
rect 27 496 80 521
rect 110 566 163 580
rect 110 532 121 566
rect 155 532 163 566
rect 110 496 163 532
rect 256 573 264 607
rect 298 573 309 607
rect 256 517 309 573
rect 256 483 264 517
rect 298 483 309 517
rect 256 427 309 483
rect 256 393 264 427
rect 298 393 309 427
rect 256 367 309 393
rect 339 367 381 619
rect 411 607 489 619
rect 411 573 432 607
rect 466 573 489 607
rect 411 513 489 573
rect 411 479 432 513
rect 466 479 489 513
rect 411 420 489 479
rect 411 386 432 420
rect 466 386 489 420
rect 411 367 489 386
rect 519 599 575 619
rect 519 565 530 599
rect 564 565 575 599
rect 519 508 575 565
rect 519 474 530 508
rect 564 474 575 508
rect 519 413 575 474
rect 519 379 530 413
rect 564 379 575 413
rect 519 367 575 379
rect 605 611 661 619
rect 605 577 616 611
rect 650 577 661 611
rect 605 534 661 577
rect 605 500 616 534
rect 650 500 661 534
rect 605 457 661 500
rect 605 423 616 457
rect 650 423 661 457
rect 605 367 661 423
rect 691 599 747 619
rect 691 565 702 599
rect 736 565 747 599
rect 691 508 747 565
rect 691 474 702 508
rect 736 474 747 508
rect 691 413 747 474
rect 691 379 702 413
rect 736 379 747 413
rect 691 367 747 379
rect 777 611 834 619
rect 777 577 788 611
rect 822 577 834 611
rect 777 534 834 577
rect 777 500 788 534
rect 822 500 834 534
rect 777 457 834 500
rect 777 423 788 457
rect 822 423 834 457
rect 777 367 834 423
<< ndiffc >>
rect 264 145 298 179
rect 159 71 193 105
rect 264 59 298 93
rect 350 169 384 203
rect 350 67 384 101
rect 436 131 470 165
rect 436 59 470 93
rect 530 147 564 181
rect 530 67 564 101
rect 616 72 650 106
rect 702 169 736 203
rect 702 67 736 101
rect 788 145 822 179
rect 788 59 822 93
<< pdiffc >>
rect 35 521 69 555
rect 121 532 155 566
rect 264 573 298 607
rect 264 483 298 517
rect 264 393 298 427
rect 432 573 466 607
rect 432 479 466 513
rect 432 386 466 420
rect 530 565 564 599
rect 530 474 564 508
rect 530 379 564 413
rect 616 577 650 611
rect 616 500 650 534
rect 616 423 650 457
rect 702 565 736 599
rect 702 474 736 508
rect 702 379 736 413
rect 788 577 822 611
rect 788 500 822 534
rect 788 423 822 457
<< poly >>
rect 309 619 339 645
rect 381 619 411 645
rect 489 619 519 645
rect 575 619 605 645
rect 661 619 691 645
rect 747 619 777 645
rect 80 580 110 606
rect 80 287 110 496
rect 44 271 110 287
rect 44 237 60 271
rect 94 237 110 271
rect 158 355 224 371
rect 158 321 174 355
rect 208 321 224 355
rect 158 287 224 321
rect 158 253 174 287
rect 208 267 224 287
rect 309 267 339 367
rect 381 335 411 367
rect 381 319 447 335
rect 381 285 397 319
rect 431 285 447 319
rect 381 269 447 285
rect 489 333 519 367
rect 575 333 605 367
rect 661 333 691 367
rect 747 333 777 367
rect 489 317 777 333
rect 489 283 505 317
rect 539 283 573 317
rect 607 283 641 317
rect 675 283 709 317
rect 743 283 777 317
rect 208 253 339 267
rect 158 237 339 253
rect 44 203 110 237
rect 309 215 339 237
rect 395 215 425 269
rect 489 267 777 283
rect 489 215 519 267
rect 575 215 605 267
rect 661 215 691 267
rect 747 215 777 267
rect 44 169 60 203
rect 94 183 110 203
rect 94 169 234 183
rect 44 153 234 169
rect 204 131 234 153
rect 204 21 234 47
rect 309 21 339 47
rect 395 21 425 47
rect 489 21 519 47
rect 575 21 605 47
rect 661 21 691 47
rect 747 21 777 47
<< polycont >>
rect 60 237 94 271
rect 174 321 208 355
rect 174 253 208 287
rect 397 285 431 319
rect 505 283 539 317
rect 573 283 607 317
rect 641 283 675 317
rect 709 283 743 317
rect 60 169 94 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 19 555 71 583
rect 19 521 35 555
rect 69 521 71 555
rect 105 566 171 649
rect 105 532 121 566
rect 155 532 171 566
rect 105 528 171 532
rect 248 607 314 615
rect 248 573 264 607
rect 298 573 314 607
rect 19 494 71 521
rect 248 517 314 573
rect 19 460 209 494
rect 17 271 109 426
rect 17 237 60 271
rect 94 237 109 271
rect 17 203 109 237
rect 17 169 60 203
rect 94 169 109 203
rect 17 59 109 169
rect 143 355 209 460
rect 143 321 174 355
rect 208 321 209 355
rect 143 287 209 321
rect 143 253 174 287
rect 208 253 209 287
rect 143 105 209 253
rect 248 483 264 517
rect 298 483 314 517
rect 248 427 314 483
rect 248 393 264 427
rect 298 393 314 427
rect 248 386 314 393
rect 416 607 482 649
rect 416 573 432 607
rect 466 573 482 607
rect 416 513 482 573
rect 416 479 432 513
rect 466 479 482 513
rect 416 420 482 479
rect 416 386 432 420
rect 466 386 482 420
rect 516 599 566 615
rect 516 565 530 599
rect 564 565 566 599
rect 516 508 566 565
rect 516 474 530 508
rect 564 474 566 508
rect 516 413 566 474
rect 600 611 666 649
rect 600 577 616 611
rect 650 577 666 611
rect 600 534 666 577
rect 600 500 616 534
rect 650 500 666 534
rect 600 457 666 500
rect 600 423 616 457
rect 650 423 666 457
rect 700 599 738 615
rect 700 565 702 599
rect 736 565 738 599
rect 700 508 738 565
rect 700 474 702 508
rect 736 474 738 508
rect 248 251 283 386
rect 516 379 530 413
rect 564 389 566 413
rect 700 413 738 474
rect 772 611 838 649
rect 772 577 788 611
rect 822 577 838 611
rect 772 534 838 577
rect 772 500 788 534
rect 822 500 838 534
rect 772 457 838 500
rect 772 423 788 457
rect 822 423 838 457
rect 700 389 702 413
rect 564 379 702 389
rect 736 389 738 413
rect 736 379 847 389
rect 317 319 455 352
rect 516 351 847 379
rect 317 285 397 319
rect 431 285 455 319
rect 489 283 505 317
rect 539 283 573 317
rect 607 283 641 317
rect 675 283 709 317
rect 743 283 759 317
rect 489 251 558 283
rect 248 215 558 251
rect 793 249 847 351
rect 348 203 393 215
rect 143 71 159 105
rect 193 71 209 105
rect 143 51 209 71
rect 248 179 314 181
rect 248 145 264 179
rect 298 145 314 179
rect 248 93 314 145
rect 248 59 264 93
rect 298 59 314 93
rect 248 17 314 59
rect 348 169 350 203
rect 384 169 393 203
rect 592 213 847 249
rect 592 203 738 213
rect 592 181 702 203
rect 348 101 393 169
rect 348 67 350 101
rect 384 67 393 101
rect 348 51 393 67
rect 427 165 480 181
rect 427 131 436 165
rect 470 131 480 165
rect 427 93 480 131
rect 427 59 436 93
rect 470 59 480 93
rect 427 17 480 59
rect 514 147 530 181
rect 564 169 702 181
rect 736 169 738 203
rect 564 147 738 169
rect 514 101 566 147
rect 514 67 530 101
rect 564 67 566 101
rect 514 51 566 67
rect 600 106 666 113
rect 600 72 616 106
rect 650 72 666 106
rect 600 17 666 72
rect 700 101 738 147
rect 700 67 702 101
rect 736 67 738 101
rect 700 51 738 67
rect 772 145 788 179
rect 822 145 838 179
rect 772 93 838 145
rect 772 59 788 93
rect 822 59 838 93
rect 772 17 838 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or2b_4
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2259634
string GDS_START 2251486
<< end >>
