magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 293 157 570 241
rect 15 49 570 157
rect 0 0 576 49
<< scnmos >>
rect 94 47 124 131
rect 166 47 196 131
rect 238 47 268 131
rect 372 47 402 215
rect 458 47 488 215
<< scpmoshvt >>
rect 80 385 110 469
rect 166 385 196 469
rect 267 385 297 469
rect 372 367 402 619
rect 458 367 488 619
<< ndiff >>
rect 319 131 372 215
rect 41 101 94 131
rect 41 67 49 101
rect 83 67 94 101
rect 41 47 94 67
rect 124 47 166 131
rect 196 47 238 131
rect 268 93 372 131
rect 268 59 305 93
rect 339 59 372 93
rect 268 47 372 59
rect 402 203 458 215
rect 402 169 413 203
rect 447 169 458 203
rect 402 101 458 169
rect 402 67 413 101
rect 447 67 458 101
rect 402 47 458 67
rect 488 201 544 215
rect 488 167 502 201
rect 536 167 544 201
rect 488 93 544 167
rect 488 59 502 93
rect 536 59 544 93
rect 488 47 544 59
<< pdiff >>
rect 319 607 372 619
rect 319 573 327 607
rect 361 573 372 607
rect 319 527 372 573
rect 319 493 327 527
rect 361 493 372 527
rect 319 469 372 493
rect 27 444 80 469
rect 27 410 35 444
rect 69 410 80 444
rect 27 385 80 410
rect 110 459 166 469
rect 110 425 121 459
rect 155 425 166 459
rect 110 385 166 425
rect 196 444 267 469
rect 196 410 214 444
rect 248 410 267 444
rect 196 385 267 410
rect 297 443 372 469
rect 297 409 308 443
rect 342 409 372 443
rect 297 385 372 409
rect 319 367 372 385
rect 402 599 458 619
rect 402 565 413 599
rect 447 565 458 599
rect 402 505 458 565
rect 402 471 413 505
rect 447 471 458 505
rect 402 413 458 471
rect 402 379 413 413
rect 447 379 458 413
rect 402 367 458 379
rect 488 607 544 619
rect 488 573 502 607
rect 536 573 544 607
rect 488 509 544 573
rect 488 475 502 509
rect 536 475 544 509
rect 488 413 544 475
rect 488 379 502 413
rect 536 379 544 413
rect 488 367 544 379
<< ndiffc >>
rect 49 67 83 101
rect 305 59 339 93
rect 413 169 447 203
rect 413 67 447 101
rect 502 167 536 201
rect 502 59 536 93
<< pdiffc >>
rect 327 573 361 607
rect 327 493 361 527
rect 35 410 69 444
rect 121 425 155 459
rect 214 410 248 444
rect 308 409 342 443
rect 413 565 447 599
rect 413 471 447 505
rect 413 379 447 413
rect 502 573 536 607
rect 502 475 536 509
rect 502 379 536 413
<< poly >>
rect 372 619 402 645
rect 458 619 488 645
rect 80 469 110 495
rect 166 469 196 495
rect 267 469 297 495
rect 80 363 110 385
rect 58 333 110 363
rect 58 321 88 333
rect 22 305 88 321
rect 22 271 38 305
rect 72 271 88 305
rect 166 291 196 385
rect 267 303 297 385
rect 372 321 402 367
rect 346 305 412 321
rect 22 237 88 271
rect 22 203 38 237
rect 72 203 88 237
rect 130 275 196 291
rect 130 241 146 275
rect 180 241 196 275
rect 130 225 196 241
rect 22 183 88 203
rect 22 153 124 183
rect 94 131 124 153
rect 166 131 196 225
rect 238 287 304 303
rect 238 253 254 287
rect 288 253 304 287
rect 346 271 362 305
rect 396 285 412 305
rect 458 285 488 367
rect 396 271 488 285
rect 346 255 488 271
rect 238 237 304 253
rect 238 131 268 237
rect 372 215 402 255
rect 458 215 488 255
rect 94 21 124 47
rect 166 21 196 47
rect 238 21 268 47
rect 372 21 402 47
rect 458 21 488 47
<< polycont >>
rect 38 271 72 305
rect 38 203 72 237
rect 146 241 180 275
rect 254 253 288 287
rect 362 271 396 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 19 444 78 460
rect 19 410 35 444
rect 69 410 78 444
rect 19 375 78 410
rect 112 459 164 649
rect 292 607 371 649
rect 292 573 327 607
rect 361 573 371 607
rect 292 527 371 573
rect 292 493 327 527
rect 361 493 371 527
rect 112 425 121 459
rect 155 425 164 459
rect 112 409 164 425
rect 198 444 258 460
rect 198 410 214 444
rect 248 410 258 444
rect 198 375 258 410
rect 292 443 371 493
rect 292 409 308 443
rect 342 409 371 443
rect 407 599 466 615
rect 407 565 413 599
rect 447 565 466 599
rect 407 505 466 565
rect 407 471 413 505
rect 447 471 466 505
rect 407 413 466 471
rect 407 379 413 413
rect 447 379 466 413
rect 19 341 373 375
rect 407 363 466 379
rect 500 607 552 649
rect 500 573 502 607
rect 536 573 552 607
rect 500 509 552 573
rect 500 475 502 509
rect 536 475 552 509
rect 500 413 552 475
rect 500 379 502 413
rect 536 379 552 413
rect 500 363 552 379
rect 339 321 373 341
rect 339 305 396 321
rect 22 271 38 305
rect 72 271 88 305
rect 22 237 88 271
rect 22 203 38 237
rect 72 203 88 237
rect 127 275 180 291
rect 127 241 146 275
rect 127 225 180 241
rect 223 287 288 303
rect 223 253 254 287
rect 223 237 288 253
rect 339 271 362 305
rect 339 255 396 271
rect 339 169 373 255
rect 430 219 466 363
rect 33 135 373 169
rect 413 203 466 219
rect 447 169 466 203
rect 33 101 99 135
rect 413 101 466 169
rect 33 67 49 101
rect 83 67 99 101
rect 33 51 99 67
rect 289 93 355 101
rect 289 59 305 93
rect 339 59 355 93
rect 289 17 355 59
rect 447 67 466 101
rect 413 51 466 67
rect 500 201 552 217
rect 500 167 502 201
rect 536 167 552 201
rect 500 93 552 167
rect 500 59 502 93
rect 536 59 552 93
rect 500 17 552 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and3_2
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5107638
string GDS_START 5101942
<< end >>
