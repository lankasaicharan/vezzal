magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 183 261 201
rect 1 49 681 183
rect 0 0 768 49
<< scnmos >>
rect 80 47 110 175
rect 152 47 182 175
rect 342 47 372 157
rect 414 47 444 157
rect 500 47 530 157
rect 572 47 602 157
<< scpmoshvt >>
rect 80 417 130 617
rect 186 417 236 617
rect 292 417 342 617
rect 398 417 448 617
rect 504 417 554 617
rect 610 417 660 617
<< ndiff >>
rect 27 163 80 175
rect 27 129 35 163
rect 69 129 80 163
rect 27 95 80 129
rect 27 61 35 95
rect 69 61 80 95
rect 27 47 80 61
rect 110 47 152 175
rect 182 163 235 175
rect 182 129 193 163
rect 227 129 235 163
rect 182 95 235 129
rect 182 61 193 95
rect 227 61 235 95
rect 182 47 235 61
rect 289 115 342 157
rect 289 81 297 115
rect 331 81 342 115
rect 289 47 342 81
rect 372 47 414 157
rect 444 115 500 157
rect 444 81 455 115
rect 489 81 500 115
rect 444 47 500 81
rect 530 47 572 157
rect 602 115 655 157
rect 602 81 613 115
rect 647 81 655 115
rect 602 47 655 81
<< pdiff >>
rect 27 599 80 617
rect 27 565 35 599
rect 69 565 80 599
rect 27 531 80 565
rect 27 497 35 531
rect 69 497 80 531
rect 27 463 80 497
rect 27 429 35 463
rect 69 429 80 463
rect 27 417 80 429
rect 130 599 186 617
rect 130 565 141 599
rect 175 565 186 599
rect 130 531 186 565
rect 130 497 141 531
rect 175 497 186 531
rect 130 463 186 497
rect 130 429 141 463
rect 175 429 186 463
rect 130 417 186 429
rect 236 599 292 617
rect 236 565 247 599
rect 281 565 292 599
rect 236 531 292 565
rect 236 497 247 531
rect 281 497 292 531
rect 236 463 292 497
rect 236 429 247 463
rect 281 429 292 463
rect 236 417 292 429
rect 342 599 398 617
rect 342 565 353 599
rect 387 565 398 599
rect 342 531 398 565
rect 342 497 353 531
rect 387 497 398 531
rect 342 463 398 497
rect 342 429 353 463
rect 387 429 398 463
rect 342 417 398 429
rect 448 599 504 617
rect 448 565 459 599
rect 493 565 504 599
rect 448 531 504 565
rect 448 497 459 531
rect 493 497 504 531
rect 448 463 504 497
rect 448 429 459 463
rect 493 429 504 463
rect 448 417 504 429
rect 554 599 610 617
rect 554 565 565 599
rect 599 565 610 599
rect 554 531 610 565
rect 554 497 565 531
rect 599 497 610 531
rect 554 463 610 497
rect 554 429 565 463
rect 599 429 610 463
rect 554 417 610 429
rect 660 599 713 617
rect 660 565 671 599
rect 705 565 713 599
rect 660 531 713 565
rect 660 497 671 531
rect 705 497 713 531
rect 660 463 713 497
rect 660 429 671 463
rect 705 429 713 463
rect 660 417 713 429
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 193 129 227 163
rect 193 61 227 95
rect 297 81 331 115
rect 455 81 489 115
rect 613 81 647 115
<< pdiffc >>
rect 35 565 69 599
rect 35 497 69 531
rect 35 429 69 463
rect 141 565 175 599
rect 141 497 175 531
rect 141 429 175 463
rect 247 565 281 599
rect 247 497 281 531
rect 247 429 281 463
rect 353 565 387 599
rect 353 497 387 531
rect 353 429 387 463
rect 459 565 493 599
rect 459 497 493 531
rect 459 429 493 463
rect 565 565 599 599
rect 565 497 599 531
rect 565 429 599 463
rect 671 565 705 599
rect 671 497 705 531
rect 671 429 705 463
<< poly >>
rect 80 617 130 645
rect 186 617 236 645
rect 292 617 342 645
rect 398 617 448 645
rect 504 617 554 645
rect 610 617 660 645
rect 80 313 130 417
rect 186 313 236 417
rect 80 297 236 313
rect 80 263 96 297
rect 130 263 236 297
rect 80 247 236 263
rect 292 309 342 417
rect 398 309 448 417
rect 504 309 554 417
rect 610 309 660 417
rect 292 291 660 309
rect 292 257 308 291
rect 342 257 376 291
rect 410 257 660 291
rect 80 175 110 247
rect 152 175 182 247
rect 292 241 660 257
rect 342 157 372 241
rect 414 157 444 241
rect 500 157 530 241
rect 572 157 602 241
rect 80 21 110 47
rect 152 21 182 47
rect 342 21 372 47
rect 414 21 444 47
rect 500 21 530 47
rect 572 21 602 47
<< polycont >>
rect 96 263 130 297
rect 308 257 342 291
rect 376 257 410 291
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 25 599 85 649
rect 25 565 35 599
rect 69 565 85 599
rect 25 531 85 565
rect 25 497 35 531
rect 69 497 85 531
rect 25 463 85 497
rect 25 429 35 463
rect 69 429 85 463
rect 25 413 85 429
rect 125 599 211 615
rect 125 565 141 599
rect 175 565 211 599
rect 125 531 211 565
rect 125 497 141 531
rect 175 497 211 531
rect 125 463 211 497
rect 125 429 141 463
rect 175 429 211 463
rect 125 413 211 429
rect 245 599 297 649
rect 245 565 247 599
rect 281 565 297 599
rect 245 531 297 565
rect 245 497 247 531
rect 281 497 297 531
rect 245 463 297 497
rect 245 429 247 463
rect 281 429 297 463
rect 245 413 297 429
rect 337 599 403 615
rect 337 565 353 599
rect 387 565 403 599
rect 337 531 403 565
rect 337 497 353 531
rect 387 497 403 531
rect 337 463 403 497
rect 337 429 353 463
rect 387 429 403 463
rect 25 313 82 356
rect 25 297 143 313
rect 25 263 96 297
rect 130 263 143 297
rect 25 227 143 263
rect 177 307 211 413
rect 337 375 403 429
rect 443 599 509 649
rect 443 565 459 599
rect 493 565 509 599
rect 443 531 509 565
rect 443 497 459 531
rect 493 497 509 531
rect 443 463 509 497
rect 443 429 459 463
rect 493 429 509 463
rect 443 417 509 429
rect 549 599 615 615
rect 549 565 565 599
rect 599 565 615 599
rect 549 531 615 565
rect 549 497 565 531
rect 599 497 615 531
rect 549 463 615 497
rect 549 429 565 463
rect 599 429 615 463
rect 549 375 615 429
rect 655 599 721 649
rect 655 565 671 599
rect 705 565 721 599
rect 655 531 721 565
rect 655 497 671 531
rect 705 497 721 531
rect 655 463 721 497
rect 655 429 671 463
rect 705 429 721 463
rect 655 417 721 429
rect 337 358 615 375
rect 337 341 748 358
rect 177 291 426 307
rect 177 257 308 291
rect 342 257 376 291
rect 410 257 426 291
rect 177 241 426 257
rect 25 163 85 179
rect 25 129 35 163
rect 69 129 85 163
rect 25 95 85 129
rect 25 61 35 95
rect 69 61 85 95
rect 25 17 85 61
rect 177 163 246 241
rect 177 129 193 163
rect 227 129 246 163
rect 471 234 748 341
rect 471 131 555 234
rect 177 95 246 129
rect 177 61 193 95
rect 227 61 246 95
rect 177 51 246 61
rect 281 115 347 131
rect 281 81 297 115
rect 331 81 347 115
rect 281 17 347 81
rect 439 115 555 131
rect 439 81 455 115
rect 489 81 555 115
rect 439 65 555 81
rect 597 115 663 131
rect 597 81 613 115
rect 647 81 663 115
rect 597 17 663 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkbuflp_4
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5400720
string GDS_START 5393956
<< end >>
