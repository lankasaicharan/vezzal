magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 556 159 863 243
rect 41 49 863 159
rect 0 0 864 49
<< scnmos >>
rect 124 49 154 133
rect 202 49 232 133
rect 288 49 318 133
rect 366 49 396 133
rect 452 49 482 133
rect 530 49 560 133
rect 632 49 662 217
rect 718 49 748 217
<< scpmoshvt >>
rect 116 491 146 619
rect 194 491 224 619
rect 280 491 310 619
rect 358 491 388 619
rect 444 491 474 619
rect 522 491 552 619
rect 664 367 694 619
rect 750 367 780 619
<< ndiff >>
rect 582 133 632 217
rect 67 112 124 133
rect 67 78 79 112
rect 113 78 124 112
rect 67 49 124 78
rect 154 49 202 133
rect 232 108 288 133
rect 232 74 243 108
rect 277 74 288 108
rect 232 49 288 74
rect 318 49 366 133
rect 396 112 452 133
rect 396 78 407 112
rect 441 78 452 112
rect 396 49 452 78
rect 482 49 530 133
rect 560 108 632 133
rect 560 74 571 108
rect 605 74 632 108
rect 560 49 632 74
rect 662 205 718 217
rect 662 171 673 205
rect 707 171 718 205
rect 662 103 718 171
rect 662 69 673 103
rect 707 69 718 103
rect 662 49 718 69
rect 748 205 837 217
rect 748 171 791 205
rect 825 171 837 205
rect 748 95 837 171
rect 748 61 791 95
rect 825 61 837 95
rect 748 49 837 61
<< pdiff >>
rect 59 565 116 619
rect 59 531 71 565
rect 105 531 116 565
rect 59 491 116 531
rect 146 491 194 619
rect 224 603 280 619
rect 224 569 235 603
rect 269 569 280 603
rect 224 491 280 569
rect 310 491 358 619
rect 388 565 444 619
rect 388 531 399 565
rect 433 531 444 565
rect 388 491 444 531
rect 474 491 522 619
rect 552 603 664 619
rect 552 569 563 603
rect 597 569 664 603
rect 552 533 664 569
rect 552 499 563 533
rect 597 499 664 533
rect 552 491 664 499
rect 614 367 664 491
rect 694 597 750 619
rect 694 563 705 597
rect 739 563 750 597
rect 694 503 750 563
rect 694 469 705 503
rect 739 469 750 503
rect 694 409 750 469
rect 694 375 705 409
rect 739 375 750 409
rect 694 367 750 375
rect 780 603 837 619
rect 780 569 791 603
rect 825 569 837 603
rect 780 506 837 569
rect 780 472 791 506
rect 825 472 837 506
rect 780 409 837 472
rect 780 375 791 409
rect 825 375 837 409
rect 780 367 837 375
<< ndiffc >>
rect 79 78 113 112
rect 243 74 277 108
rect 407 78 441 112
rect 571 74 605 108
rect 673 171 707 205
rect 673 69 707 103
rect 791 171 825 205
rect 791 61 825 95
<< pdiffc >>
rect 71 531 105 565
rect 235 569 269 603
rect 399 531 433 565
rect 563 569 597 603
rect 563 499 597 533
rect 705 563 739 597
rect 705 469 739 503
rect 705 375 739 409
rect 791 569 825 603
rect 791 472 825 506
rect 791 375 825 409
<< poly >>
rect 116 619 146 645
rect 194 619 224 645
rect 280 619 310 645
rect 358 619 388 645
rect 444 619 474 645
rect 522 619 552 645
rect 664 619 694 645
rect 750 619 780 645
rect 116 387 146 491
rect 194 465 224 491
rect 194 435 232 465
rect 88 371 154 387
rect 88 337 104 371
rect 138 337 154 371
rect 88 303 154 337
rect 88 269 104 303
rect 138 269 154 303
rect 88 253 154 269
rect 124 133 154 253
rect 202 377 232 435
rect 280 377 310 491
rect 202 361 310 377
rect 202 327 233 361
rect 267 327 310 361
rect 358 377 388 491
rect 444 377 474 491
rect 522 447 552 491
rect 516 431 582 447
rect 516 397 532 431
rect 566 397 582 431
rect 516 381 582 397
rect 358 361 474 377
rect 358 347 412 361
rect 202 293 310 327
rect 202 259 233 293
rect 267 273 310 293
rect 366 327 412 347
rect 446 327 474 361
rect 366 293 474 327
rect 267 259 318 273
rect 202 243 318 259
rect 202 133 232 243
rect 288 133 318 243
rect 366 259 412 293
rect 446 273 474 293
rect 446 259 482 273
rect 366 243 482 259
rect 366 133 396 243
rect 452 133 482 243
rect 530 133 560 381
rect 664 323 694 367
rect 619 307 694 323
rect 619 273 635 307
rect 669 287 694 307
rect 750 287 780 367
rect 669 273 780 287
rect 619 257 780 273
rect 632 217 662 257
rect 718 217 748 257
rect 124 23 154 49
rect 202 23 232 49
rect 288 23 318 49
rect 366 23 396 49
rect 452 23 482 49
rect 530 23 560 49
rect 632 23 662 49
rect 718 23 748 49
<< polycont >>
rect 104 337 138 371
rect 104 269 138 303
rect 233 327 267 361
rect 532 397 566 431
rect 233 259 267 293
rect 412 327 446 361
rect 412 259 446 293
rect 635 273 669 307
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 18 565 121 613
rect 18 531 71 565
rect 105 531 121 565
rect 219 603 285 649
rect 219 569 235 603
rect 269 569 285 603
rect 219 553 285 569
rect 383 565 449 613
rect 18 517 121 531
rect 383 531 399 565
rect 433 531 449 565
rect 383 517 449 531
rect 18 483 449 517
rect 547 603 613 649
rect 547 569 563 603
rect 597 569 613 603
rect 547 533 613 569
rect 547 499 563 533
rect 597 499 613 533
rect 547 483 613 499
rect 689 597 755 613
rect 689 563 705 597
rect 739 563 755 597
rect 689 503 755 563
rect 18 207 52 483
rect 689 469 705 503
rect 739 469 755 503
rect 88 431 647 447
rect 88 413 532 431
rect 88 371 154 413
rect 505 397 532 413
rect 566 397 647 431
rect 505 381 647 397
rect 689 409 755 469
rect 88 337 104 371
rect 138 337 154 371
rect 88 303 154 337
rect 88 269 104 303
rect 138 269 154 303
rect 88 253 154 269
rect 217 361 359 377
rect 217 327 233 361
rect 267 327 359 361
rect 217 293 359 327
rect 217 259 233 293
rect 267 259 359 293
rect 217 243 359 259
rect 396 361 462 377
rect 396 327 412 361
rect 446 327 462 361
rect 689 375 705 409
rect 739 375 755 409
rect 689 359 755 375
rect 791 603 841 649
rect 825 569 841 603
rect 791 506 841 569
rect 825 472 841 506
rect 791 409 841 472
rect 825 375 841 409
rect 791 359 841 375
rect 396 293 462 327
rect 396 259 412 293
rect 446 259 462 293
rect 396 243 462 259
rect 587 307 685 323
rect 587 273 635 307
rect 669 273 685 307
rect 587 257 685 273
rect 587 207 621 257
rect 721 221 755 359
rect 18 173 621 207
rect 657 205 755 221
rect 63 112 129 173
rect 63 78 79 112
rect 113 78 129 112
rect 63 53 129 78
rect 227 108 293 137
rect 227 74 243 108
rect 277 74 293 108
rect 227 17 293 74
rect 391 112 457 173
rect 657 171 673 205
rect 707 171 755 205
rect 391 78 407 112
rect 441 78 457 112
rect 391 53 457 78
rect 555 108 621 137
rect 555 74 571 108
rect 605 74 621 108
rect 555 17 621 74
rect 657 103 755 171
rect 657 69 673 103
rect 707 69 755 103
rect 657 53 755 69
rect 791 205 841 221
rect 825 171 841 205
rect 791 95 841 171
rect 825 61 841 95
rect 791 17 841 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 maj3_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6766388
string GDS_START 6759446
<< end >>
