magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 5138 1975
<< nwell >>
rect -38 455 3878 704
rect -38 331 187 455
rect 1145 331 3878 455
rect 2952 321 3398 331
<< pwell >>
rect 229 329 669 371
rect 993 329 1103 401
rect 229 235 1103 329
rect 2102 251 2314 273
rect 2102 241 2866 251
rect 3390 241 3839 247
rect 229 157 277 235
rect 3 49 277 157
rect 662 229 1103 235
rect 1548 229 3839 241
rect 662 49 3839 229
rect 0 0 3840 49
<< scnmos >>
rect 312 261 342 345
rect 398 261 428 345
rect 470 261 500 345
rect 556 261 586 345
rect 86 47 116 131
rect 164 47 194 131
rect 881 219 911 303
rect 967 219 997 303
rect 753 66 783 150
rect 1273 119 1303 203
rect 1351 119 1381 203
rect 1631 87 1661 215
rect 1709 87 1739 215
rect 1850 47 1880 215
rect 1928 47 1958 215
rect 2201 119 2231 247
rect 2310 141 2340 225
rect 2388 141 2418 225
rect 2652 141 2682 225
rect 2730 141 2760 225
rect 3045 47 3075 215
rect 3117 47 3147 215
rect 3203 47 3233 215
rect 3275 47 3305 215
rect 3473 137 3503 221
rect 3545 137 3575 221
rect 3654 53 3684 221
rect 3726 53 3756 221
<< scpmoshvt >>
rect 95 491 125 619
rect 167 491 197 619
rect 312 491 342 619
rect 390 491 420 619
rect 476 491 506 619
rect 554 491 584 619
rect 705 491 735 619
rect 783 491 813 619
rect 881 491 911 575
rect 990 491 1020 575
rect 1147 535 1177 619
rect 1345 535 1375 619
rect 1417 535 1447 619
rect 1643 375 1673 543
rect 1715 375 1745 543
rect 1840 367 1870 619
rect 1912 367 1942 619
rect 2138 439 2168 523
rect 2247 387 2277 555
rect 2458 535 2488 619
rect 2689 518 2719 602
rect 2761 518 2791 602
rect 2847 518 2877 602
rect 2580 397 2610 481
rect 3045 357 3075 609
rect 3117 357 3147 609
rect 3203 357 3233 609
rect 3275 357 3305 609
rect 3473 367 3503 495
rect 3545 367 3575 495
rect 3654 367 3684 619
rect 3726 367 3756 619
<< ndiff >>
rect 255 333 312 345
rect 255 299 267 333
rect 301 299 312 333
rect 255 261 312 299
rect 342 307 398 345
rect 342 273 353 307
rect 387 273 398 307
rect 342 261 398 273
rect 428 261 470 345
rect 500 307 556 345
rect 500 273 511 307
rect 545 273 556 307
rect 500 261 556 273
rect 586 333 643 345
rect 586 299 597 333
rect 631 299 643 333
rect 586 261 643 299
rect 29 111 86 131
rect 29 77 41 111
rect 75 77 86 111
rect 29 47 86 77
rect 116 47 164 131
rect 194 100 251 131
rect 1019 367 1077 375
rect 1019 333 1031 367
rect 1065 333 1077 367
rect 1019 303 1077 333
rect 824 273 881 303
rect 824 239 836 273
rect 870 239 881 273
rect 824 219 881 239
rect 911 289 967 303
rect 911 255 922 289
rect 956 255 967 289
rect 911 219 967 255
rect 997 219 1077 303
rect 1216 177 1273 203
rect 194 66 205 100
rect 239 66 251 100
rect 194 47 251 66
rect 688 93 753 150
rect 688 59 696 93
rect 730 66 753 93
rect 783 118 840 150
rect 783 84 794 118
rect 828 84 840 118
rect 1216 143 1228 177
rect 1262 143 1273 177
rect 1216 119 1273 143
rect 1303 119 1351 203
rect 1381 119 1461 203
rect 783 66 840 84
rect 730 59 738 66
rect 688 43 738 59
rect 1403 91 1461 119
rect 1403 57 1415 91
rect 1449 57 1461 91
rect 1574 188 1631 215
rect 1574 154 1586 188
rect 1620 154 1631 188
rect 1574 87 1631 154
rect 1661 87 1709 215
rect 1739 87 1850 215
rect 1777 77 1850 87
rect 1403 45 1461 57
rect 1777 43 1789 77
rect 1823 47 1850 77
rect 1880 47 1928 215
rect 1958 203 2015 215
rect 1958 169 1969 203
rect 2003 169 2015 203
rect 1958 103 2015 169
rect 1958 69 1969 103
rect 2003 69 2015 103
rect 1958 47 2015 69
rect 2128 235 2201 247
rect 2128 201 2140 235
rect 2174 201 2201 235
rect 2128 165 2201 201
rect 2128 131 2140 165
rect 2174 131 2201 165
rect 2128 119 2201 131
rect 2231 225 2288 247
rect 2231 165 2310 225
rect 2231 131 2242 165
rect 2276 141 2310 165
rect 2340 141 2388 225
rect 2418 158 2652 225
rect 2418 141 2452 158
rect 2276 131 2288 141
rect 2231 119 2288 131
rect 2440 124 2452 141
rect 2486 141 2652 158
rect 2682 141 2730 225
rect 2760 191 2840 225
rect 2760 157 2794 191
rect 2828 157 2840 191
rect 2760 141 2840 157
rect 2486 124 2498 141
rect 2440 112 2498 124
rect 1823 43 1835 47
rect 1777 31 1835 43
rect 2988 114 3045 215
rect 2988 80 3000 114
rect 3034 80 3045 114
rect 2988 47 3045 80
rect 3075 47 3117 215
rect 3147 109 3203 215
rect 3147 75 3158 109
rect 3192 75 3203 109
rect 3147 47 3203 75
rect 3233 47 3275 215
rect 3305 199 3362 215
rect 3305 165 3316 199
rect 3350 165 3362 199
rect 3305 103 3362 165
rect 3416 196 3473 221
rect 3416 162 3428 196
rect 3462 162 3473 196
rect 3416 137 3473 162
rect 3503 137 3545 221
rect 3575 209 3654 221
rect 3575 175 3609 209
rect 3643 175 3654 209
rect 3575 137 3654 175
rect 3305 69 3316 103
rect 3350 69 3362 103
rect 3305 47 3362 69
rect 3597 99 3654 137
rect 3597 65 3609 99
rect 3643 65 3654 99
rect 3597 53 3654 65
rect 3684 53 3726 221
rect 3756 209 3813 221
rect 3756 175 3767 209
rect 3801 175 3813 209
rect 3756 103 3813 175
rect 3756 69 3767 103
rect 3801 69 3813 103
rect 3756 53 3813 69
<< pdiff >>
rect 38 567 95 619
rect 38 533 50 567
rect 84 533 95 567
rect 38 491 95 533
rect 125 491 167 619
rect 197 578 312 619
rect 197 544 208 578
rect 242 544 312 578
rect 197 491 312 544
rect 342 491 390 619
rect 420 567 476 619
rect 420 533 431 567
rect 465 533 476 567
rect 420 491 476 533
rect 506 491 554 619
rect 584 578 705 619
rect 584 544 595 578
rect 629 544 705 578
rect 584 491 705 544
rect 735 491 783 619
rect 813 575 866 619
rect 1035 575 1147 619
rect 813 541 824 575
rect 858 541 881 575
rect 813 491 881 541
rect 911 550 990 575
rect 911 516 945 550
rect 979 516 990 550
rect 911 491 990 516
rect 1020 535 1147 575
rect 1177 601 1345 619
rect 1177 567 1188 601
rect 1222 567 1345 601
rect 1177 535 1345 567
rect 1375 535 1417 619
rect 1447 593 1504 619
rect 1447 559 1458 593
rect 1492 559 1504 593
rect 1783 607 1840 619
rect 1783 573 1795 607
rect 1829 573 1840 607
rect 1447 535 1504 559
rect 1783 543 1840 573
rect 1020 491 1125 535
rect 1586 527 1643 543
rect 1586 493 1598 527
rect 1632 493 1643 527
rect 1586 421 1643 493
rect 1586 387 1598 421
rect 1632 387 1643 421
rect 1586 375 1643 387
rect 1673 375 1715 543
rect 1745 514 1840 543
rect 1745 480 1795 514
rect 1829 480 1840 514
rect 1745 421 1840 480
rect 1745 387 1795 421
rect 1829 387 1840 421
rect 1745 375 1840 387
rect 1783 367 1840 375
rect 1870 367 1912 619
rect 1942 527 1999 619
rect 1942 493 1953 527
rect 1987 493 1999 527
rect 1942 413 1999 493
rect 1942 379 1953 413
rect 1987 379 1999 413
rect 1942 367 1999 379
rect 2401 600 2458 619
rect 2401 566 2413 600
rect 2447 566 2458 600
rect 2190 531 2247 555
rect 2190 523 2202 531
rect 2081 510 2138 523
rect 2081 476 2093 510
rect 2127 476 2138 510
rect 2081 439 2138 476
rect 2168 497 2202 523
rect 2236 497 2247 531
rect 2168 439 2247 497
rect 2190 387 2247 439
rect 2277 433 2334 555
rect 2401 535 2458 566
rect 2488 600 2561 619
rect 2488 566 2515 600
rect 2549 566 2561 600
rect 2488 535 2561 566
rect 2625 577 2689 602
rect 2625 543 2644 577
rect 2678 543 2689 577
rect 2625 518 2689 543
rect 2719 518 2761 602
rect 2791 590 2847 602
rect 2791 556 2802 590
rect 2836 556 2847 590
rect 2791 518 2847 556
rect 2877 590 2934 602
rect 2877 556 2888 590
rect 2922 556 2934 590
rect 2877 518 2934 556
rect 2988 597 3045 609
rect 2988 563 3000 597
rect 3034 563 3045 597
rect 2277 399 2288 433
rect 2322 399 2334 433
rect 2277 387 2334 399
rect 2625 481 2662 518
rect 2523 453 2580 481
rect 2523 419 2535 453
rect 2569 419 2580 453
rect 2523 397 2580 419
rect 2610 397 2662 481
rect 2988 500 3045 563
rect 2988 466 3000 500
rect 3034 466 3045 500
rect 2988 403 3045 466
rect 2988 369 3000 403
rect 3034 369 3045 403
rect 2988 357 3045 369
rect 3075 357 3117 609
rect 3147 597 3203 609
rect 3147 563 3158 597
rect 3192 563 3203 597
rect 3147 519 3203 563
rect 3147 485 3158 519
rect 3192 485 3203 519
rect 3147 442 3203 485
rect 3147 408 3158 442
rect 3192 408 3203 442
rect 3147 357 3203 408
rect 3233 357 3275 609
rect 3305 597 3362 609
rect 3305 563 3316 597
rect 3350 563 3362 597
rect 3305 500 3362 563
rect 3597 607 3654 619
rect 3597 573 3609 607
rect 3643 573 3654 607
rect 3305 466 3316 500
rect 3350 466 3362 500
rect 3597 510 3654 573
rect 3597 495 3609 510
rect 3305 403 3362 466
rect 3305 369 3316 403
rect 3350 369 3362 403
rect 3305 357 3362 369
rect 3416 483 3473 495
rect 3416 449 3428 483
rect 3462 449 3473 483
rect 3416 413 3473 449
rect 3416 379 3428 413
rect 3462 379 3473 413
rect 3416 367 3473 379
rect 3503 367 3545 495
rect 3575 476 3609 495
rect 3643 476 3654 510
rect 3575 413 3654 476
rect 3575 379 3609 413
rect 3643 379 3654 413
rect 3575 367 3654 379
rect 3684 367 3726 619
rect 3756 597 3813 619
rect 3756 563 3767 597
rect 3801 563 3813 597
rect 3756 505 3813 563
rect 3756 471 3767 505
rect 3801 471 3813 505
rect 3756 413 3813 471
rect 3756 379 3767 413
rect 3801 379 3813 413
rect 3756 367 3813 379
<< ndiffc >>
rect 267 299 301 333
rect 353 273 387 307
rect 511 273 545 307
rect 597 299 631 333
rect 41 77 75 111
rect 1031 333 1065 367
rect 836 239 870 273
rect 922 255 956 289
rect 205 66 239 100
rect 696 59 730 93
rect 794 84 828 118
rect 1228 143 1262 177
rect 1415 57 1449 91
rect 1586 154 1620 188
rect 1789 43 1823 77
rect 1969 169 2003 203
rect 1969 69 2003 103
rect 2140 201 2174 235
rect 2140 131 2174 165
rect 2242 131 2276 165
rect 2452 124 2486 158
rect 2794 157 2828 191
rect 3000 80 3034 114
rect 3158 75 3192 109
rect 3316 165 3350 199
rect 3428 162 3462 196
rect 3609 175 3643 209
rect 3316 69 3350 103
rect 3609 65 3643 99
rect 3767 175 3801 209
rect 3767 69 3801 103
<< pdiffc >>
rect 50 533 84 567
rect 208 544 242 578
rect 431 533 465 567
rect 595 544 629 578
rect 824 541 858 575
rect 945 516 979 550
rect 1188 567 1222 601
rect 1458 559 1492 593
rect 1795 573 1829 607
rect 1598 493 1632 527
rect 1598 387 1632 421
rect 1795 480 1829 514
rect 1795 387 1829 421
rect 1953 493 1987 527
rect 1953 379 1987 413
rect 2413 566 2447 600
rect 2093 476 2127 510
rect 2202 497 2236 531
rect 2515 566 2549 600
rect 2644 543 2678 577
rect 2802 556 2836 590
rect 2888 556 2922 590
rect 3000 563 3034 597
rect 2288 399 2322 433
rect 2535 419 2569 453
rect 3000 466 3034 500
rect 3000 369 3034 403
rect 3158 563 3192 597
rect 3158 485 3192 519
rect 3158 408 3192 442
rect 3316 563 3350 597
rect 3609 573 3643 607
rect 3316 466 3350 500
rect 3316 369 3350 403
rect 3428 449 3462 483
rect 3428 379 3462 413
rect 3609 476 3643 510
rect 3609 379 3643 413
rect 3767 563 3801 597
rect 3767 471 3801 505
rect 3767 379 3801 413
<< poly >>
rect 95 619 125 645
rect 167 619 197 645
rect 312 619 342 645
rect 390 619 420 645
rect 476 619 506 645
rect 554 619 584 645
rect 705 619 735 645
rect 783 619 813 645
rect 1147 619 1177 645
rect 1345 619 1375 645
rect 1417 619 1447 645
rect 1840 619 1870 645
rect 1912 619 1942 645
rect 881 575 911 601
rect 990 575 1020 601
rect 1643 543 1673 569
rect 1715 543 1745 569
rect 1147 520 1177 535
rect 95 397 125 491
rect 167 397 197 491
rect 312 397 342 491
rect 95 381 342 397
rect 95 347 111 381
rect 145 367 342 381
rect 390 397 420 491
rect 476 397 506 491
rect 390 367 428 397
rect 145 347 194 367
rect 95 313 194 347
rect 312 345 342 367
rect 398 345 428 367
rect 470 367 506 397
rect 554 397 584 491
rect 705 469 735 491
rect 783 469 813 491
rect 705 443 839 469
rect 705 439 789 443
rect 773 409 789 439
rect 823 409 839 443
rect 554 377 731 397
rect 554 367 681 377
rect 470 345 500 367
rect 556 345 586 367
rect 95 293 111 313
rect 86 279 111 293
rect 145 279 194 313
rect 86 263 194 279
rect 86 131 116 263
rect 164 131 194 263
rect 665 343 681 367
rect 715 343 731 377
rect 665 327 731 343
rect 773 375 839 409
rect 773 341 789 375
rect 823 341 839 375
rect 773 325 839 341
rect 312 235 342 261
rect 398 113 428 261
rect 470 183 500 261
rect 556 235 586 261
rect 773 195 803 325
rect 881 303 911 491
rect 990 448 1020 491
rect 1147 490 1303 520
rect 990 439 1231 448
rect 967 427 1231 439
rect 967 409 1181 427
rect 967 303 997 409
rect 1165 393 1181 409
rect 1215 393 1231 427
rect 1165 377 1231 393
rect 1273 291 1303 490
rect 1345 503 1375 535
rect 1417 503 1447 535
rect 1345 487 1447 503
rect 1345 473 1367 487
rect 1237 275 1303 291
rect 1237 241 1253 275
rect 1287 241 1303 275
rect 1237 225 1303 241
rect 470 167 536 183
rect 470 133 486 167
rect 520 133 536 167
rect 753 165 803 195
rect 753 150 783 165
rect 881 159 911 219
rect 967 193 997 219
rect 1273 203 1303 225
rect 1351 453 1367 473
rect 1401 453 1447 487
rect 1351 437 1447 453
rect 1351 203 1381 437
rect 1496 327 1562 343
rect 1496 293 1512 327
rect 1546 307 1562 327
rect 1643 307 1673 375
rect 1715 307 1745 375
rect 2036 597 2277 627
rect 2458 619 2488 645
rect 1840 335 1870 367
rect 1912 335 1942 367
rect 1546 293 1745 307
rect 1496 277 1745 293
rect 1787 319 1942 335
rect 1787 285 1803 319
rect 1837 299 1942 319
rect 2036 299 2066 597
rect 2247 555 2277 597
rect 2138 523 2168 549
rect 2138 353 2168 439
rect 2689 602 2719 628
rect 2761 602 2791 628
rect 2847 602 2877 628
rect 3045 609 3075 635
rect 3117 609 3147 635
rect 3203 609 3233 635
rect 3275 609 3305 635
rect 3654 619 3684 645
rect 3726 619 3756 645
rect 2458 503 2488 535
rect 2422 487 2488 503
rect 2422 453 2438 487
rect 2472 453 2488 487
rect 2580 481 2610 507
rect 2422 437 2488 453
rect 2247 361 2277 387
rect 1837 285 2066 299
rect 1631 215 1661 277
rect 1709 215 1739 277
rect 1787 269 2066 285
rect 2114 337 2180 353
rect 2114 303 2130 337
rect 2164 313 2180 337
rect 2422 313 2452 437
rect 2689 486 2719 518
rect 2761 486 2791 518
rect 2689 470 2799 486
rect 2689 436 2749 470
rect 2783 436 2799 470
rect 2689 420 2799 436
rect 2580 365 2610 397
rect 2544 349 2610 365
rect 2689 355 2719 420
rect 2544 315 2560 349
rect 2594 315 2610 349
rect 2164 303 2231 313
rect 2114 283 2231 303
rect 1850 215 1880 269
rect 1928 215 1958 269
rect 470 117 536 133
rect 356 97 428 113
rect 356 63 372 97
rect 406 83 428 97
rect 406 63 422 83
rect 356 47 422 63
rect 876 143 942 159
rect 876 109 892 143
rect 926 109 942 143
rect 876 93 942 109
rect 1273 93 1303 119
rect 86 21 116 47
rect 164 21 194 47
rect 753 51 783 66
rect 1351 51 1381 119
rect 753 21 1381 51
rect 1631 61 1661 87
rect 1709 61 1739 87
rect 2036 51 2066 269
rect 2201 247 2231 283
rect 2422 297 2494 313
rect 2544 299 2610 315
rect 2652 325 2719 355
rect 2422 277 2444 297
rect 2388 263 2444 277
rect 2478 263 2494 297
rect 2310 225 2340 251
rect 2388 247 2494 263
rect 2388 225 2418 247
rect 2652 225 2682 325
rect 2847 314 2877 518
rect 3473 495 3503 521
rect 3545 495 3575 521
rect 3045 325 3075 357
rect 3117 325 3147 357
rect 2811 298 2877 314
rect 2811 277 2827 298
rect 2730 264 2827 277
rect 2861 264 2877 298
rect 2730 247 2877 264
rect 2937 298 3003 314
rect 2937 264 2953 298
rect 2987 264 3003 298
rect 2937 248 3003 264
rect 3045 309 3152 325
rect 3045 275 3102 309
rect 3136 275 3152 309
rect 3045 259 3152 275
rect 3203 317 3233 357
rect 3275 317 3305 357
rect 3203 301 3305 317
rect 3203 267 3219 301
rect 3253 281 3305 301
rect 3473 281 3503 367
rect 3545 281 3575 367
rect 3654 327 3684 367
rect 3726 327 3756 367
rect 3253 267 3575 281
rect 2730 225 2760 247
rect 2201 93 2231 119
rect 2310 51 2340 141
rect 2388 115 2418 141
rect 2538 103 2604 119
rect 2652 115 2682 141
rect 2730 115 2760 141
rect 2937 119 2967 248
rect 3045 215 3075 259
rect 3117 215 3147 259
rect 3203 251 3575 267
rect 3649 311 3756 327
rect 3649 277 3665 311
rect 3699 277 3756 311
rect 3649 261 3756 277
rect 3203 215 3233 251
rect 3275 215 3305 251
rect 3473 221 3503 251
rect 3545 221 3575 251
rect 3654 221 3684 261
rect 3726 221 3756 261
rect 2538 69 2554 103
rect 2588 69 2604 103
rect 2538 51 2604 69
rect 2900 103 2967 119
rect 2900 69 2916 103
rect 2950 69 2967 103
rect 2900 51 2967 69
rect 1850 21 1880 47
rect 1928 21 1958 47
rect 2036 21 2967 51
rect 3473 111 3503 137
rect 3545 111 3575 137
rect 3045 21 3075 47
rect 3117 21 3147 47
rect 3203 21 3233 47
rect 3275 21 3305 47
rect 3654 27 3684 53
rect 3726 27 3756 53
<< polycont >>
rect 111 347 145 381
rect 789 409 823 443
rect 111 279 145 313
rect 681 343 715 377
rect 789 341 823 375
rect 1181 393 1215 427
rect 1253 241 1287 275
rect 486 133 520 167
rect 1367 453 1401 487
rect 1512 293 1546 327
rect 1803 285 1837 319
rect 2438 453 2472 487
rect 2130 303 2164 337
rect 2749 436 2783 470
rect 2560 315 2594 349
rect 372 63 406 97
rect 892 109 926 143
rect 2444 263 2478 297
rect 2827 264 2861 298
rect 2953 264 2987 298
rect 3102 275 3136 309
rect 3219 267 3253 301
rect 3665 277 3699 311
rect 2554 69 2588 103
rect 2916 69 2950 103
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3775 683
rect 3809 649 3840 683
rect 25 567 100 613
rect 25 533 50 567
rect 84 533 100 567
rect 25 487 100 533
rect 192 578 258 649
rect 192 544 208 578
rect 242 544 258 578
rect 192 499 258 544
rect 415 567 481 613
rect 415 533 431 567
rect 465 533 481 567
rect 25 177 59 487
rect 415 463 481 533
rect 579 578 645 649
rect 1172 601 1238 649
rect 579 544 595 578
rect 629 544 645 578
rect 579 499 645 544
rect 681 575 909 595
rect 681 541 824 575
rect 858 541 909 575
rect 681 540 909 541
rect 681 463 715 540
rect 95 381 161 430
rect 95 347 111 381
rect 145 347 161 381
rect 95 313 161 347
rect 95 279 111 313
rect 145 279 161 313
rect 95 236 161 279
rect 197 429 715 463
rect 773 498 839 504
rect 773 464 799 498
rect 833 464 839 498
rect 773 443 839 464
rect 197 247 231 429
rect 773 409 789 443
rect 823 409 839 443
rect 267 359 631 393
rect 267 333 301 359
rect 581 333 631 359
rect 267 283 301 299
rect 337 307 403 323
rect 337 273 353 307
rect 387 273 403 307
rect 337 247 403 273
rect 197 213 403 247
rect 495 307 545 323
rect 495 273 511 307
rect 581 299 597 333
rect 667 377 737 393
rect 667 343 681 377
rect 715 343 737 377
rect 667 310 737 343
rect 773 375 839 409
rect 875 439 909 540
rect 943 550 981 579
rect 943 516 945 550
rect 979 516 981 550
rect 1172 567 1188 601
rect 1222 567 1238 601
rect 1442 593 1492 613
rect 1442 574 1458 593
rect 1172 547 1238 567
rect 1274 559 1458 574
rect 943 511 981 516
rect 1274 540 1492 559
rect 1528 579 1718 613
rect 1274 511 1308 540
rect 943 477 1308 511
rect 1351 498 1417 504
rect 1351 487 1375 498
rect 875 405 1065 439
rect 773 341 789 375
rect 823 341 839 375
rect 773 325 839 341
rect 1015 367 1065 405
rect 1015 333 1031 367
rect 1015 317 1065 333
rect 1101 343 1135 477
rect 1351 453 1367 487
rect 1409 464 1417 498
rect 1401 453 1417 464
rect 1351 445 1417 453
rect 1171 427 1231 443
rect 1171 393 1181 427
rect 1215 411 1231 427
rect 1528 411 1562 579
rect 1215 393 1562 411
rect 1171 377 1562 393
rect 1598 527 1648 543
rect 1632 493 1648 527
rect 1598 421 1648 493
rect 1632 387 1648 421
rect 1101 327 1562 343
rect 1101 309 1512 327
rect 581 283 631 299
rect 906 289 972 307
rect 495 247 545 273
rect 820 273 870 289
rect 495 213 717 247
rect 820 239 836 273
rect 906 255 922 289
rect 956 281 972 289
rect 1101 281 1135 309
rect 1496 293 1512 309
rect 1546 293 1562 327
rect 1496 283 1562 293
rect 956 255 1135 281
rect 906 247 1135 255
rect 820 215 870 239
rect 683 179 717 213
rect 836 211 870 215
rect 1237 241 1253 275
rect 1287 247 1303 275
rect 1598 247 1648 387
rect 1684 335 1718 579
rect 1779 607 1845 649
rect 1779 573 1795 607
rect 1829 573 1845 607
rect 1779 514 1845 573
rect 1779 480 1795 514
rect 1829 480 1845 514
rect 1779 421 1845 480
rect 1779 387 1795 421
rect 1829 387 1845 421
rect 1779 371 1845 387
rect 1883 579 2057 613
rect 1684 319 1847 335
rect 1684 285 1803 319
rect 1837 285 1847 319
rect 1684 269 1847 285
rect 1287 241 1648 247
rect 1237 233 1648 241
rect 1883 233 1917 579
rect 1237 213 1917 233
rect 25 167 536 177
rect 25 143 486 167
rect 25 111 91 143
rect 459 133 486 143
rect 520 133 536 167
rect 683 145 800 179
rect 836 177 1154 211
rect 1570 199 1917 213
rect 1953 527 1987 543
rect 1953 413 1987 493
rect 2023 423 2057 579
rect 2093 600 2463 613
rect 2093 579 2413 600
rect 2093 510 2143 579
rect 2397 566 2413 579
rect 2447 566 2463 600
rect 2397 559 2463 566
rect 2499 600 2565 649
rect 2499 566 2515 600
rect 2549 566 2565 600
rect 2499 559 2565 566
rect 2628 577 2694 606
rect 2628 543 2644 577
rect 2678 543 2694 577
rect 2127 476 2143 510
rect 2186 531 2252 543
rect 2186 497 2202 531
rect 2236 519 2252 531
rect 2628 523 2694 543
rect 2786 590 2836 649
rect 2786 556 2802 590
rect 2786 540 2836 556
rect 2872 590 2938 606
rect 2872 556 2888 590
rect 2922 556 2938 590
rect 2872 540 2938 556
rect 2236 497 2392 519
rect 2186 485 2392 497
rect 2093 459 2143 476
rect 2272 433 2322 449
rect 2272 423 2288 433
rect 2023 399 2288 423
rect 2023 389 2322 399
rect 1953 353 1987 379
rect 2216 383 2322 389
rect 2358 383 2392 485
rect 2428 489 2694 523
rect 2733 498 2855 504
rect 2428 487 2483 489
rect 2428 453 2438 487
rect 2472 453 2483 487
rect 2733 470 2815 498
rect 2428 437 2483 453
rect 2519 419 2535 453
rect 2569 419 2680 453
rect 2733 436 2749 470
rect 2783 464 2815 470
rect 2849 464 2855 498
rect 2783 436 2855 464
rect 2733 420 2855 436
rect 2646 384 2680 419
rect 2904 384 2938 540
rect 1953 337 2180 353
rect 1953 303 2130 337
rect 2164 303 2180 337
rect 1953 287 2180 303
rect 1953 203 2019 287
rect 2216 251 2250 383
rect 1570 188 1648 199
rect 766 143 800 145
rect 1094 143 1228 177
rect 1262 143 1278 177
rect 1314 143 1534 177
rect 459 123 536 133
rect 25 77 41 111
rect 75 77 91 111
rect 25 53 91 77
rect 189 100 255 107
rect 189 66 205 100
rect 239 66 255 100
rect 189 17 255 66
rect 356 97 422 107
rect 356 63 372 97
rect 406 87 422 97
rect 601 87 647 134
rect 766 118 842 143
rect 406 63 647 87
rect 356 53 647 63
rect 696 93 730 111
rect 696 17 730 59
rect 766 84 794 118
rect 828 84 842 118
rect 766 53 842 84
rect 876 109 892 143
rect 926 109 942 143
rect 876 87 942 109
rect 1314 87 1348 143
rect 876 53 1348 87
rect 1399 91 1449 107
rect 1399 57 1415 91
rect 1399 17 1449 57
rect 1500 87 1534 143
rect 1570 154 1586 188
rect 1620 154 1648 188
rect 1953 169 1969 203
rect 2003 169 2019 203
rect 1953 163 2019 169
rect 1570 123 1648 154
rect 1684 129 2019 163
rect 1684 87 1718 129
rect 1953 103 2019 129
rect 2124 235 2250 251
rect 2124 201 2140 235
rect 2174 217 2250 235
rect 2358 349 2610 383
rect 2646 350 2938 384
rect 2984 597 3050 613
rect 2984 563 3000 597
rect 3034 563 3050 597
rect 2984 500 3050 563
rect 2984 466 3000 500
rect 3034 466 3050 500
rect 2984 403 3050 466
rect 2984 369 3000 403
rect 3034 369 3050 403
rect 3142 597 3208 649
rect 3142 563 3158 597
rect 3192 563 3208 597
rect 3142 519 3208 563
rect 3142 485 3158 519
rect 3192 485 3208 519
rect 3142 442 3208 485
rect 3142 408 3158 442
rect 3192 408 3208 442
rect 3142 392 3208 408
rect 3300 597 3366 613
rect 3300 563 3316 597
rect 3350 563 3366 597
rect 3300 500 3366 563
rect 3300 466 3316 500
rect 3350 466 3366 500
rect 3593 607 3659 649
rect 3593 573 3609 607
rect 3643 573 3659 607
rect 3593 510 3659 573
rect 3300 403 3366 466
rect 2174 201 2190 217
rect 2124 165 2190 201
rect 2358 181 2392 349
rect 2544 315 2560 349
rect 2594 315 2610 349
rect 2544 314 2610 315
rect 2984 314 3050 369
rect 3300 369 3316 403
rect 3350 369 3366 403
rect 2428 297 2494 313
rect 2428 263 2444 297
rect 2478 263 2494 297
rect 2544 298 2898 314
rect 2544 280 2827 298
rect 2428 244 2494 263
rect 2811 264 2827 280
rect 2861 264 2898 298
rect 2811 248 2898 264
rect 2937 298 3050 314
rect 2937 264 2953 298
rect 2987 264 3050 298
rect 2937 248 3050 264
rect 3086 309 3152 356
rect 3300 353 3366 369
rect 3086 275 3102 309
rect 3136 275 3152 309
rect 3086 259 3152 275
rect 3203 301 3269 317
rect 3203 267 3219 301
rect 3253 267 3269 301
rect 3203 251 3269 267
rect 2428 212 2572 244
rect 2864 212 2898 248
rect 3203 212 3237 251
rect 3332 215 3366 353
rect 2428 210 2828 212
rect 2124 131 2140 165
rect 2174 131 2190 165
rect 2124 115 2190 131
rect 2226 165 2392 181
rect 2538 191 2828 210
rect 2538 178 2794 191
rect 2226 131 2242 165
rect 2276 131 2392 165
rect 2226 115 2392 131
rect 2436 158 2502 174
rect 2436 124 2452 158
rect 2486 124 2502 158
rect 2778 157 2794 178
rect 2864 178 3237 212
rect 3289 199 3366 215
rect 2778 137 2828 157
rect 3289 165 3316 199
rect 3350 165 3366 199
rect 1500 53 1718 87
rect 1773 77 1839 93
rect 1773 43 1789 77
rect 1823 43 1839 77
rect 1953 69 1969 103
rect 2003 69 2019 103
rect 1953 53 2019 69
rect 1773 17 1839 43
rect 2436 17 2502 124
rect 2538 103 2604 119
rect 2538 69 2554 103
rect 2588 87 2604 103
rect 2900 114 3050 142
rect 2900 103 3000 114
rect 2900 87 2916 103
rect 2588 69 2916 87
rect 2950 80 3000 103
rect 3034 80 3050 114
rect 2950 69 3050 80
rect 2538 53 3050 69
rect 3142 109 3208 142
rect 3142 75 3158 109
rect 3192 75 3208 109
rect 3142 17 3208 75
rect 3289 103 3366 165
rect 3412 483 3478 499
rect 3412 449 3428 483
rect 3462 449 3478 483
rect 3412 413 3478 449
rect 3412 379 3428 413
rect 3462 379 3478 413
rect 3412 327 3478 379
rect 3593 476 3609 510
rect 3643 476 3659 510
rect 3593 413 3659 476
rect 3593 379 3609 413
rect 3643 379 3659 413
rect 3593 363 3659 379
rect 3751 597 3817 613
rect 3751 563 3767 597
rect 3801 563 3817 597
rect 3751 505 3817 563
rect 3751 471 3767 505
rect 3801 471 3817 505
rect 3751 413 3817 471
rect 3751 379 3767 413
rect 3801 379 3817 413
rect 3412 311 3715 327
rect 3412 277 3665 311
rect 3699 277 3715 311
rect 3412 261 3715 277
rect 3412 196 3478 261
rect 3412 162 3428 196
rect 3462 162 3478 196
rect 3412 133 3478 162
rect 3593 209 3659 225
rect 3593 175 3609 209
rect 3643 175 3659 209
rect 3289 69 3316 103
rect 3350 69 3366 103
rect 3289 53 3366 69
rect 3593 99 3659 175
rect 3593 65 3609 99
rect 3643 65 3659 99
rect 3593 17 3659 65
rect 3751 209 3817 379
rect 3751 175 3767 209
rect 3801 175 3817 209
rect 3751 103 3817 175
rect 3751 69 3767 103
rect 3801 69 3817 103
rect 3751 53 3817 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3840 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 3583 649 3617 683
rect 3679 649 3713 683
rect 3775 649 3809 683
rect 799 464 833 498
rect 1375 487 1409 498
rect 1375 464 1401 487
rect 1401 464 1409 487
rect 2815 464 2849 498
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
<< metal1 >>
rect 0 683 3840 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3775 683
rect 3809 649 3840 683
rect 0 617 3840 649
rect 787 498 845 504
rect 787 464 799 498
rect 833 495 845 498
rect 1363 498 1421 504
rect 1363 495 1375 498
rect 833 467 1375 495
rect 833 464 845 467
rect 787 458 845 464
rect 1363 464 1375 467
rect 1409 495 1421 498
rect 2803 498 2861 504
rect 2803 495 2815 498
rect 1409 467 2815 495
rect 1409 464 1421 467
rect 1363 458 1421 464
rect 2803 464 2815 467
rect 2849 464 2861 498
rect 2803 458 2861 464
rect 0 17 3840 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3840 17
rect 0 -49 3840 -17
<< labels >>
flabel pwell s 0 0 3840 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 3840 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel comment s 1073 36 1073 36 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfrbp_lp
flabel comment s 2957 175 2957 175 0 FreeSans 200 90 0 0 no_jumper_check
flabel comment s 2434 385 2434 385 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 799 464 833 498 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 3840 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 3840 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 3775 94 3809 128 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 168 3809 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 242 3809 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 316 3809 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 390 3809 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 464 3809 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3775 538 3809 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 3295 94 3329 128 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3295 168 3329 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 3103 316 3137 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3840 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry R90
string GDS_END 6481620
string GDS_START 6455860
<< end >>
