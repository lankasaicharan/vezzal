magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3026 1975
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 1 232 536 248
rect 829 232 939 275
rect 1 49 1727 232
rect 0 0 1728 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 273 368 309 592
rect 400 368 436 592
rect 501 392 537 592
rect 615 392 651 592
rect 788 392 824 592
rect 888 392 924 592
rect 1120 392 1156 592
rect 1214 392 1250 592
rect 1305 392 1341 592
rect 1419 392 1455 592
rect 1509 392 1545 592
rect 1603 392 1639 592
<< nmoslvt >>
rect 98 74 128 222
rect 184 74 214 222
rect 323 74 353 222
rect 423 74 453 222
rect 621 78 651 206
rect 810 78 840 206
rect 928 78 958 206
rect 1014 78 1044 206
rect 1120 78 1150 206
rect 1227 78 1257 206
rect 1314 78 1344 206
rect 1419 78 1449 206
rect 1525 78 1555 206
rect 1614 78 1644 206
<< ndiff >>
rect 27 188 98 222
rect 27 154 39 188
rect 73 154 98 188
rect 27 120 98 154
rect 27 86 53 120
rect 87 86 98 120
rect 27 74 98 86
rect 128 210 184 222
rect 128 176 139 210
rect 173 176 184 210
rect 128 120 184 176
rect 128 86 139 120
rect 173 86 184 120
rect 128 74 184 86
rect 214 120 323 222
rect 214 86 251 120
rect 285 86 323 120
rect 214 74 323 86
rect 353 194 423 222
rect 353 160 364 194
rect 398 160 423 194
rect 353 120 423 160
rect 353 86 364 120
rect 398 86 423 120
rect 353 74 423 86
rect 453 194 510 222
rect 855 237 913 249
rect 855 206 867 237
rect 453 160 464 194
rect 498 160 510 194
rect 571 181 621 206
rect 453 120 510 160
rect 453 86 464 120
rect 498 86 510 120
rect 453 74 510 86
rect 564 151 621 181
rect 564 117 576 151
rect 610 117 621 151
rect 564 78 621 117
rect 651 169 810 206
rect 651 135 676 169
rect 710 135 765 169
rect 799 135 810 169
rect 651 78 810 135
rect 840 203 867 206
rect 901 206 913 237
rect 901 203 928 206
rect 840 78 928 203
rect 958 172 1014 206
rect 958 138 969 172
rect 1003 138 1014 172
rect 958 78 1014 138
rect 1044 192 1120 206
rect 1044 158 1069 192
rect 1103 158 1120 192
rect 1044 124 1120 158
rect 1044 90 1069 124
rect 1103 90 1120 124
rect 1044 78 1120 90
rect 1150 124 1227 206
rect 1150 90 1169 124
rect 1203 90 1227 124
rect 1150 78 1227 90
rect 1257 194 1314 206
rect 1257 160 1269 194
rect 1303 160 1314 194
rect 1257 124 1314 160
rect 1257 90 1269 124
rect 1303 90 1314 124
rect 1257 78 1314 90
rect 1344 124 1419 206
rect 1344 90 1369 124
rect 1403 90 1419 124
rect 1344 78 1419 90
rect 1449 192 1525 206
rect 1449 158 1469 192
rect 1503 158 1525 192
rect 1449 120 1525 158
rect 1449 86 1469 120
rect 1503 86 1525 120
rect 1449 78 1525 86
rect 1555 124 1614 206
rect 1555 90 1569 124
rect 1603 90 1614 124
rect 1555 78 1614 90
rect 1644 192 1701 206
rect 1644 158 1655 192
rect 1689 158 1701 192
rect 1644 120 1701 158
rect 1644 86 1655 120
rect 1689 86 1701 120
rect 1644 78 1701 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 497 173 546
rect 119 463 129 497
rect 163 463 173 497
rect 119 414 173 463
rect 119 380 129 414
rect 163 380 173 414
rect 119 368 173 380
rect 209 582 273 592
rect 209 548 229 582
rect 263 548 273 582
rect 209 514 273 548
rect 209 480 229 514
rect 263 480 273 514
rect 209 446 273 480
rect 209 412 229 446
rect 263 412 273 446
rect 209 368 273 412
rect 309 580 400 592
rect 309 546 329 580
rect 363 546 400 580
rect 309 497 400 546
rect 309 463 329 497
rect 363 463 400 497
rect 309 414 400 463
rect 309 380 329 414
rect 363 380 400 414
rect 309 368 400 380
rect 436 582 501 592
rect 436 548 446 582
rect 480 548 501 582
rect 436 514 501 548
rect 436 480 446 514
rect 480 480 501 514
rect 436 446 501 480
rect 436 412 446 446
rect 480 412 501 446
rect 436 392 501 412
rect 537 580 615 592
rect 537 546 547 580
rect 581 546 615 580
rect 537 509 615 546
rect 537 475 547 509
rect 581 475 615 509
rect 537 438 615 475
rect 537 404 547 438
rect 581 404 615 438
rect 537 392 615 404
rect 651 580 788 592
rect 651 546 661 580
rect 695 546 744 580
rect 778 546 788 580
rect 651 508 788 546
rect 651 474 661 508
rect 695 474 744 508
rect 778 474 788 508
rect 651 392 788 474
rect 824 580 888 592
rect 824 546 834 580
rect 868 546 888 580
rect 824 509 888 546
rect 824 475 834 509
rect 868 475 888 509
rect 824 438 888 475
rect 824 404 834 438
rect 868 404 888 438
rect 824 392 888 404
rect 924 580 980 592
rect 924 546 934 580
rect 968 546 980 580
rect 924 512 980 546
rect 924 478 934 512
rect 968 478 980 512
rect 924 392 980 478
rect 1034 576 1120 592
rect 1034 542 1061 576
rect 1095 542 1120 576
rect 1034 392 1120 542
rect 1156 440 1214 592
rect 1156 406 1168 440
rect 1202 406 1214 440
rect 1156 392 1214 406
rect 1250 578 1305 592
rect 1250 544 1260 578
rect 1294 544 1305 578
rect 1250 392 1305 544
rect 1341 547 1419 592
rect 1341 513 1367 547
rect 1401 513 1419 547
rect 1341 392 1419 513
rect 1455 453 1509 592
rect 1455 419 1465 453
rect 1499 419 1509 453
rect 1455 392 1509 419
rect 1545 531 1603 592
rect 1545 497 1555 531
rect 1589 497 1603 531
rect 1545 444 1603 497
rect 1545 410 1555 444
rect 1589 410 1603 444
rect 1545 392 1603 410
rect 1639 580 1701 592
rect 1639 546 1655 580
rect 1689 546 1701 580
rect 1639 512 1701 546
rect 1639 478 1655 512
rect 1689 478 1701 512
rect 1639 444 1701 478
rect 1639 410 1655 444
rect 1689 410 1701 444
rect 1639 392 1701 410
rect 436 368 486 392
<< ndiffc >>
rect 39 154 73 188
rect 53 86 87 120
rect 139 176 173 210
rect 139 86 173 120
rect 251 86 285 120
rect 364 160 398 194
rect 364 86 398 120
rect 464 160 498 194
rect 464 86 498 120
rect 576 117 610 151
rect 676 135 710 169
rect 765 135 799 169
rect 867 203 901 237
rect 969 138 1003 172
rect 1069 158 1103 192
rect 1069 90 1103 124
rect 1169 90 1203 124
rect 1269 160 1303 194
rect 1269 90 1303 124
rect 1369 90 1403 124
rect 1469 158 1503 192
rect 1469 86 1503 120
rect 1569 90 1603 124
rect 1655 158 1689 192
rect 1655 86 1689 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 229 548 263 582
rect 229 480 263 514
rect 229 412 263 446
rect 329 546 363 580
rect 329 463 363 497
rect 329 380 363 414
rect 446 548 480 582
rect 446 480 480 514
rect 446 412 480 446
rect 547 546 581 580
rect 547 475 581 509
rect 547 404 581 438
rect 661 546 695 580
rect 744 546 778 580
rect 661 474 695 508
rect 744 474 778 508
rect 834 546 868 580
rect 834 475 868 509
rect 834 404 868 438
rect 934 546 968 580
rect 934 478 968 512
rect 1061 542 1095 576
rect 1168 406 1202 440
rect 1260 544 1294 578
rect 1367 513 1401 547
rect 1465 419 1499 453
rect 1555 497 1589 531
rect 1555 410 1589 444
rect 1655 546 1689 580
rect 1655 478 1689 512
rect 1655 410 1689 444
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 273 592 309 618
rect 400 592 436 618
rect 501 592 537 618
rect 615 592 651 618
rect 788 592 824 618
rect 888 592 924 618
rect 1120 592 1156 618
rect 1214 592 1250 618
rect 1305 592 1341 618
rect 1419 592 1455 618
rect 1509 592 1545 618
rect 1603 592 1639 618
rect 83 310 119 368
rect 173 310 209 368
rect 273 310 309 368
rect 400 310 436 368
rect 501 310 537 392
rect 615 353 651 392
rect 788 353 824 392
rect 888 372 924 392
rect 615 337 840 353
rect 888 344 1072 372
rect 888 342 1022 344
rect 615 323 715 337
rect 83 294 453 310
rect 83 260 267 294
rect 301 260 335 294
rect 369 260 403 294
rect 437 260 453 294
rect 83 244 453 260
rect 501 294 567 310
rect 501 260 517 294
rect 551 274 567 294
rect 699 303 715 323
rect 749 303 840 337
rect 699 294 840 303
rect 1006 310 1022 342
rect 1056 310 1072 344
rect 1006 294 1072 310
rect 1120 350 1156 392
rect 1214 350 1250 392
rect 1120 334 1250 350
rect 1120 300 1190 334
rect 1224 314 1250 334
rect 1224 300 1257 314
rect 551 260 651 274
rect 699 264 958 294
rect 501 244 651 260
rect 98 222 128 244
rect 184 222 214 244
rect 323 222 353 244
rect 423 222 453 244
rect 621 206 651 244
rect 810 206 840 264
rect 928 206 958 264
rect 1014 206 1044 294
rect 1120 284 1257 300
rect 1120 206 1150 284
rect 1227 206 1257 284
rect 1305 310 1341 392
rect 1419 360 1455 392
rect 1509 360 1545 392
rect 1419 344 1555 360
rect 1419 310 1437 344
rect 1471 310 1505 344
rect 1539 310 1555 344
rect 1305 294 1371 310
rect 1305 260 1321 294
rect 1355 260 1371 294
rect 1305 244 1371 260
rect 1419 294 1555 310
rect 1603 294 1639 392
rect 1314 206 1344 244
rect 1419 206 1449 294
rect 1525 206 1555 294
rect 1609 278 1707 294
rect 1609 244 1657 278
rect 1691 244 1707 278
rect 1609 228 1707 244
rect 1614 206 1644 228
rect 98 48 128 74
rect 184 48 214 74
rect 323 48 353 74
rect 423 48 453 74
rect 621 52 651 78
rect 810 52 840 78
rect 928 52 958 78
rect 1014 52 1044 78
rect 1120 52 1150 78
rect 1227 52 1257 78
rect 1314 52 1344 78
rect 1419 52 1449 78
rect 1525 52 1555 78
rect 1614 52 1644 78
<< polycont >>
rect 267 260 301 294
rect 335 260 369 294
rect 403 260 437 294
rect 517 260 551 294
rect 715 303 749 337
rect 1022 310 1056 344
rect 1190 300 1224 334
rect 1437 310 1471 344
rect 1505 310 1539 344
rect 1321 260 1355 294
rect 1657 244 1691 278
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 497 179 546
rect 113 463 129 497
rect 163 463 179 497
rect 113 414 179 463
rect 113 380 129 414
rect 163 380 179 414
rect 213 582 279 649
rect 213 548 229 582
rect 263 548 279 582
rect 213 514 279 548
rect 213 480 229 514
rect 263 480 279 514
rect 213 446 279 480
rect 213 412 229 446
rect 263 412 279 446
rect 313 580 379 596
rect 313 546 329 580
rect 363 546 379 580
rect 313 497 379 546
rect 313 463 329 497
rect 363 463 379 497
rect 313 414 379 463
rect 113 378 179 380
rect 313 380 329 414
rect 363 380 379 414
rect 430 582 496 649
rect 430 548 446 582
rect 480 548 496 582
rect 430 514 496 548
rect 430 480 446 514
rect 480 480 496 514
rect 430 446 496 480
rect 430 412 446 446
rect 480 412 496 446
rect 531 580 597 596
rect 531 546 547 580
rect 581 546 597 580
rect 531 509 597 546
rect 531 475 547 509
rect 581 475 597 509
rect 531 438 597 475
rect 645 580 784 649
rect 645 546 661 580
rect 695 546 744 580
rect 778 546 784 580
rect 645 508 784 546
rect 645 474 661 508
rect 695 474 744 508
rect 778 474 784 508
rect 645 458 784 474
rect 818 580 884 596
rect 818 546 834 580
rect 868 546 884 580
rect 818 509 884 546
rect 818 475 834 509
rect 868 475 884 509
rect 313 378 379 380
rect 531 404 547 438
rect 581 424 597 438
rect 818 438 884 475
rect 918 580 984 649
rect 1244 592 1705 615
rect 918 546 934 580
rect 968 546 984 580
rect 918 512 984 546
rect 1030 581 1705 592
rect 1030 578 1310 581
rect 1030 576 1260 578
rect 1030 542 1061 576
rect 1095 544 1260 576
rect 1294 544 1310 578
rect 1639 580 1705 581
rect 1095 542 1310 544
rect 1344 513 1367 547
rect 1401 531 1605 547
rect 1401 513 1555 531
rect 918 478 934 512
rect 968 508 984 512
rect 968 479 1310 508
rect 1589 497 1605 531
rect 968 478 1515 479
rect 918 474 1515 478
rect 918 462 984 474
rect 1276 453 1515 474
rect 818 424 834 438
rect 581 404 834 424
rect 868 428 884 438
rect 1150 428 1168 440
rect 868 406 1168 428
rect 1202 406 1220 440
rect 868 404 1220 406
rect 531 394 1220 404
rect 1276 419 1465 453
rect 1499 419 1515 453
rect 1276 394 1515 419
rect 1555 444 1605 497
rect 1589 410 1605 444
rect 1555 394 1605 410
rect 1639 546 1655 580
rect 1689 546 1705 580
rect 1639 512 1705 546
rect 1639 478 1655 512
rect 1689 478 1705 512
rect 1639 444 1705 478
rect 1639 410 1655 444
rect 1689 410 1705 444
rect 1639 394 1705 410
rect 531 390 884 394
rect 531 378 597 390
rect 818 388 884 390
rect 1106 390 1220 394
rect 113 344 379 378
rect 419 344 597 378
rect 113 330 179 344
rect 25 296 179 330
rect 419 310 453 344
rect 697 337 765 356
rect 25 262 71 296
rect 251 294 453 310
rect 25 228 189 262
rect 251 260 267 294
rect 301 260 335 294
rect 369 260 403 294
rect 437 260 453 294
rect 251 244 453 260
rect 501 294 582 310
rect 501 260 517 294
rect 551 260 582 294
rect 697 303 715 337
rect 749 303 765 337
rect 985 344 1072 360
rect 985 328 1022 344
rect 697 287 765 303
rect 799 310 1022 328
rect 1056 310 1072 344
rect 799 294 1072 310
rect 501 253 582 260
rect 799 253 833 294
rect 1106 260 1140 390
rect 1174 334 1240 356
rect 1174 300 1190 334
rect 1224 300 1240 334
rect 1421 344 1607 360
rect 1421 310 1437 344
rect 1471 310 1505 344
rect 1539 310 1607 344
rect 1174 284 1240 300
rect 1305 294 1387 310
rect 1421 294 1607 310
rect 501 244 833 253
rect 123 210 189 228
rect 548 219 833 244
rect 867 237 1140 260
rect 1305 260 1321 294
rect 1355 260 1387 294
rect 1641 278 1707 356
rect 1641 260 1657 278
rect 1305 244 1657 260
rect 1691 244 1707 278
rect 23 188 89 194
rect 23 154 39 188
rect 73 154 89 188
rect 23 120 89 154
rect 23 86 53 120
rect 87 86 89 120
rect 23 17 89 86
rect 123 176 139 210
rect 173 194 414 210
rect 173 176 364 194
rect 123 120 189 176
rect 348 160 364 176
rect 398 160 414 194
rect 123 86 139 120
rect 173 86 189 120
rect 123 70 189 86
rect 223 120 314 136
rect 223 86 251 120
rect 285 86 314 120
rect 223 17 314 86
rect 348 120 414 160
rect 348 86 364 120
rect 398 86 414 120
rect 348 70 414 86
rect 448 194 514 210
rect 448 160 464 194
rect 498 160 514 194
rect 901 226 1140 237
rect 1353 226 1707 244
rect 901 203 917 226
rect 867 187 917 203
rect 1253 194 1319 210
rect 1253 192 1269 194
rect 448 120 514 160
rect 448 86 464 120
rect 498 86 514 120
rect 448 17 514 86
rect 560 151 626 185
rect 560 117 576 151
rect 610 117 626 151
rect 660 169 815 185
rect 660 135 676 169
rect 710 135 765 169
rect 799 153 815 169
rect 953 172 1019 192
rect 953 153 969 172
rect 799 138 969 153
rect 1003 138 1019 172
rect 799 135 1019 138
rect 660 119 1019 135
rect 1053 158 1069 192
rect 1103 160 1269 192
rect 1303 192 1319 194
rect 1303 160 1469 192
rect 1103 158 1469 160
rect 1503 158 1655 192
rect 1689 158 1705 192
rect 1053 124 1119 158
rect 1253 124 1319 158
rect 560 85 626 117
rect 1053 90 1069 124
rect 1103 90 1119 124
rect 1053 85 1119 90
rect 560 51 1119 85
rect 1153 90 1169 124
rect 1203 90 1219 124
rect 1153 17 1219 90
rect 1253 90 1269 124
rect 1303 90 1319 124
rect 1253 74 1319 90
rect 1353 90 1369 124
rect 1403 90 1419 124
rect 1353 17 1419 90
rect 1453 120 1519 158
rect 1453 86 1469 120
rect 1503 86 1519 120
rect 1453 70 1519 86
rect 1553 90 1569 124
rect 1603 90 1619 124
rect 1553 17 1619 90
rect 1655 120 1705 158
rect 1689 86 1705 120
rect 1655 70 1705 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o311a_4
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 2371588
string GDS_START 2358390
<< end >>
