magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
rect 793 313 1603 331
<< pwell >>
rect 4 49 2052 241
rect 0 0 2112 49
<< scnmos >>
rect 83 47 113 215
rect 169 47 199 215
rect 255 47 285 215
rect 341 47 371 215
rect 427 47 457 215
rect 513 47 543 215
rect 599 47 629 215
rect 685 47 715 215
rect 793 47 823 215
rect 879 47 909 215
rect 979 47 1009 215
rect 1079 47 1109 215
rect 1258 47 1288 215
rect 1344 47 1374 215
rect 1430 47 1460 215
rect 1590 47 1620 215
rect 1685 47 1715 215
rect 1771 47 1801 215
rect 1857 47 1887 215
rect 1943 47 1973 215
<< scpmoshvt >>
rect 83 367 113 619
rect 169 367 199 619
rect 255 367 285 619
rect 341 367 371 619
rect 434 367 464 619
rect 520 367 550 619
rect 606 367 636 619
rect 692 367 722 619
rect 882 349 912 601
rect 968 349 998 601
rect 1054 349 1084 601
rect 1140 349 1170 601
rect 1226 349 1256 601
rect 1312 349 1342 601
rect 1398 349 1428 601
rect 1484 349 1514 601
rect 1685 367 1715 619
rect 1771 367 1801 619
rect 1857 367 1887 619
rect 1943 367 1973 619
<< ndiff >>
rect 30 203 83 215
rect 30 169 38 203
rect 72 169 83 203
rect 30 105 83 169
rect 30 71 38 105
rect 72 71 83 105
rect 30 47 83 71
rect 113 169 169 215
rect 113 135 124 169
rect 158 135 169 169
rect 113 47 169 135
rect 199 163 255 215
rect 199 129 210 163
rect 244 129 255 163
rect 199 93 255 129
rect 199 59 210 93
rect 244 59 255 93
rect 199 47 255 59
rect 285 169 341 215
rect 285 135 296 169
rect 330 135 341 169
rect 285 47 341 135
rect 371 163 427 215
rect 371 129 382 163
rect 416 129 427 163
rect 371 93 427 129
rect 371 59 382 93
rect 416 59 427 93
rect 371 47 427 59
rect 457 169 513 215
rect 457 135 468 169
rect 502 135 513 169
rect 457 47 513 135
rect 543 163 599 215
rect 543 129 554 163
rect 588 129 599 163
rect 543 93 599 129
rect 543 59 554 93
rect 588 59 599 93
rect 543 47 599 59
rect 629 173 685 215
rect 629 139 640 173
rect 674 139 685 173
rect 629 47 685 139
rect 715 163 793 215
rect 715 129 726 163
rect 760 129 793 163
rect 715 89 793 129
rect 715 55 726 89
rect 760 55 793 89
rect 715 47 793 55
rect 823 89 879 215
rect 823 55 834 89
rect 868 55 879 89
rect 823 47 879 55
rect 909 165 979 215
rect 909 131 920 165
rect 954 131 979 165
rect 909 92 979 131
rect 909 58 934 92
rect 968 58 979 92
rect 909 47 979 58
rect 1009 89 1079 215
rect 1009 55 1034 89
rect 1068 55 1079 89
rect 1009 47 1079 55
rect 1109 165 1258 215
rect 1109 131 1120 165
rect 1154 131 1258 165
rect 1109 127 1258 131
rect 1109 93 1202 127
rect 1236 93 1258 127
rect 1109 89 1258 93
rect 1109 55 1134 89
rect 1168 55 1258 89
rect 1109 47 1258 55
rect 1288 89 1344 215
rect 1288 55 1299 89
rect 1333 55 1344 89
rect 1288 47 1344 55
rect 1374 192 1430 215
rect 1374 158 1385 192
rect 1419 158 1430 192
rect 1374 101 1430 158
rect 1374 67 1385 101
rect 1419 67 1430 101
rect 1374 47 1430 67
rect 1460 124 1590 215
rect 1460 90 1471 124
rect 1505 90 1545 124
rect 1579 90 1590 124
rect 1460 47 1590 90
rect 1620 192 1685 215
rect 1620 158 1631 192
rect 1665 158 1685 192
rect 1620 101 1685 158
rect 1620 67 1631 101
rect 1665 67 1685 101
rect 1620 47 1685 67
rect 1715 124 1771 215
rect 1715 90 1726 124
rect 1760 90 1771 124
rect 1715 47 1771 90
rect 1801 192 1857 215
rect 1801 158 1812 192
rect 1846 158 1857 192
rect 1801 101 1857 158
rect 1801 67 1812 101
rect 1846 67 1857 101
rect 1801 47 1857 67
rect 1887 124 1943 215
rect 1887 90 1898 124
rect 1932 90 1943 124
rect 1887 47 1943 90
rect 1973 192 2026 215
rect 1973 158 1984 192
rect 2018 158 2026 192
rect 1973 101 2026 158
rect 1973 67 1984 101
rect 2018 67 2026 101
rect 1973 47 2026 67
<< pdiff >>
rect 30 599 83 619
rect 30 565 38 599
rect 72 565 83 599
rect 30 520 83 565
rect 30 486 38 520
rect 72 486 83 520
rect 30 438 83 486
rect 30 404 38 438
rect 72 404 83 438
rect 30 367 83 404
rect 113 538 169 619
rect 113 504 124 538
rect 158 504 169 538
rect 113 436 169 504
rect 113 402 124 436
rect 158 402 169 436
rect 113 367 169 402
rect 199 599 255 619
rect 199 565 210 599
rect 244 565 255 599
rect 199 504 255 565
rect 199 470 210 504
rect 244 470 255 504
rect 199 367 255 470
rect 285 538 341 619
rect 285 504 296 538
rect 330 504 341 538
rect 285 436 341 504
rect 285 402 296 436
rect 330 402 341 436
rect 285 367 341 402
rect 371 599 434 619
rect 371 565 389 599
rect 423 565 434 599
rect 371 504 434 565
rect 371 470 389 504
rect 423 470 434 504
rect 371 367 434 470
rect 464 568 520 619
rect 464 534 475 568
rect 509 534 520 568
rect 464 367 520 534
rect 550 599 606 619
rect 550 565 561 599
rect 595 565 606 599
rect 550 504 606 565
rect 550 470 561 504
rect 595 470 606 504
rect 550 367 606 470
rect 636 568 692 619
rect 636 534 647 568
rect 681 534 692 568
rect 636 367 692 534
rect 722 599 775 619
rect 1632 607 1685 619
rect 722 565 733 599
rect 767 565 775 599
rect 722 504 775 565
rect 722 470 733 504
rect 767 470 775 504
rect 722 367 775 470
rect 829 589 882 601
rect 829 555 837 589
rect 871 555 882 589
rect 829 504 882 555
rect 829 470 837 504
rect 871 470 882 504
rect 829 349 882 470
rect 912 531 968 601
rect 912 497 923 531
rect 957 497 968 531
rect 912 436 968 497
rect 912 402 923 436
rect 957 402 968 436
rect 912 349 968 402
rect 998 589 1054 601
rect 998 555 1009 589
rect 1043 555 1054 589
rect 998 504 1054 555
rect 998 470 1009 504
rect 1043 470 1054 504
rect 998 349 1054 470
rect 1084 531 1140 601
rect 1084 497 1095 531
rect 1129 497 1140 531
rect 1084 436 1140 497
rect 1084 402 1095 436
rect 1129 402 1140 436
rect 1084 349 1140 402
rect 1170 589 1226 601
rect 1170 555 1181 589
rect 1215 555 1226 589
rect 1170 504 1226 555
rect 1170 470 1181 504
rect 1215 470 1226 504
rect 1170 349 1226 470
rect 1256 529 1312 601
rect 1256 495 1267 529
rect 1301 495 1312 529
rect 1256 461 1312 495
rect 1256 427 1267 461
rect 1301 427 1312 461
rect 1256 391 1312 427
rect 1256 357 1267 391
rect 1301 357 1312 391
rect 1256 349 1312 357
rect 1342 589 1398 601
rect 1342 555 1353 589
rect 1387 555 1398 589
rect 1342 519 1398 555
rect 1342 485 1353 519
rect 1387 485 1398 519
rect 1342 451 1398 485
rect 1342 417 1353 451
rect 1387 417 1398 451
rect 1342 349 1398 417
rect 1428 531 1484 601
rect 1428 497 1439 531
rect 1473 497 1484 531
rect 1428 463 1484 497
rect 1428 429 1439 463
rect 1473 429 1484 463
rect 1428 391 1484 429
rect 1428 357 1439 391
rect 1473 357 1484 391
rect 1428 349 1484 357
rect 1514 589 1567 601
rect 1514 555 1525 589
rect 1559 555 1567 589
rect 1514 519 1567 555
rect 1514 485 1525 519
rect 1559 485 1567 519
rect 1514 451 1567 485
rect 1514 417 1525 451
rect 1559 417 1567 451
rect 1514 349 1567 417
rect 1632 573 1640 607
rect 1674 573 1685 607
rect 1632 518 1685 573
rect 1632 484 1640 518
rect 1674 484 1685 518
rect 1632 435 1685 484
rect 1632 401 1640 435
rect 1674 401 1685 435
rect 1632 367 1685 401
rect 1715 599 1771 619
rect 1715 565 1726 599
rect 1760 565 1771 599
rect 1715 506 1771 565
rect 1715 472 1726 506
rect 1760 472 1771 506
rect 1715 413 1771 472
rect 1715 379 1726 413
rect 1760 379 1771 413
rect 1715 367 1771 379
rect 1801 607 1857 619
rect 1801 573 1812 607
rect 1846 573 1857 607
rect 1801 518 1857 573
rect 1801 484 1812 518
rect 1846 484 1857 518
rect 1801 435 1857 484
rect 1801 401 1812 435
rect 1846 401 1857 435
rect 1801 367 1857 401
rect 1887 599 1943 619
rect 1887 565 1898 599
rect 1932 565 1943 599
rect 1887 506 1943 565
rect 1887 472 1898 506
rect 1932 472 1943 506
rect 1887 413 1943 472
rect 1887 379 1898 413
rect 1932 379 1943 413
rect 1887 367 1943 379
rect 1973 607 2026 619
rect 1973 573 1984 607
rect 2018 573 2026 607
rect 1973 504 2026 573
rect 1973 470 1984 504
rect 2018 470 2026 504
rect 1973 413 2026 470
rect 1973 379 1984 413
rect 2018 379 2026 413
rect 1973 367 2026 379
<< ndiffc >>
rect 38 169 72 203
rect 38 71 72 105
rect 124 135 158 169
rect 210 129 244 163
rect 210 59 244 93
rect 296 135 330 169
rect 382 129 416 163
rect 382 59 416 93
rect 468 135 502 169
rect 554 129 588 163
rect 554 59 588 93
rect 640 139 674 173
rect 726 129 760 163
rect 726 55 760 89
rect 834 55 868 89
rect 920 131 954 165
rect 934 58 968 92
rect 1034 55 1068 89
rect 1120 131 1154 165
rect 1202 93 1236 127
rect 1134 55 1168 89
rect 1299 55 1333 89
rect 1385 158 1419 192
rect 1385 67 1419 101
rect 1471 90 1505 124
rect 1545 90 1579 124
rect 1631 158 1665 192
rect 1631 67 1665 101
rect 1726 90 1760 124
rect 1812 158 1846 192
rect 1812 67 1846 101
rect 1898 90 1932 124
rect 1984 158 2018 192
rect 1984 67 2018 101
<< pdiffc >>
rect 38 565 72 599
rect 38 486 72 520
rect 38 404 72 438
rect 124 504 158 538
rect 124 402 158 436
rect 210 565 244 599
rect 210 470 244 504
rect 296 504 330 538
rect 296 402 330 436
rect 389 565 423 599
rect 389 470 423 504
rect 475 534 509 568
rect 561 565 595 599
rect 561 470 595 504
rect 647 534 681 568
rect 733 565 767 599
rect 733 470 767 504
rect 837 555 871 589
rect 837 470 871 504
rect 923 497 957 531
rect 923 402 957 436
rect 1009 555 1043 589
rect 1009 470 1043 504
rect 1095 497 1129 531
rect 1095 402 1129 436
rect 1181 555 1215 589
rect 1181 470 1215 504
rect 1267 495 1301 529
rect 1267 427 1301 461
rect 1267 357 1301 391
rect 1353 555 1387 589
rect 1353 485 1387 519
rect 1353 417 1387 451
rect 1439 497 1473 531
rect 1439 429 1473 463
rect 1439 357 1473 391
rect 1525 555 1559 589
rect 1525 485 1559 519
rect 1525 417 1559 451
rect 1640 573 1674 607
rect 1640 484 1674 518
rect 1640 401 1674 435
rect 1726 565 1760 599
rect 1726 472 1760 506
rect 1726 379 1760 413
rect 1812 573 1846 607
rect 1812 484 1846 518
rect 1812 401 1846 435
rect 1898 565 1932 599
rect 1898 472 1932 506
rect 1898 379 1932 413
rect 1984 573 2018 607
rect 1984 470 2018 504
rect 1984 379 2018 413
<< poly >>
rect 83 619 113 645
rect 169 619 199 645
rect 255 619 285 645
rect 341 619 371 645
rect 434 619 464 645
rect 520 619 550 645
rect 606 619 636 645
rect 692 619 722 645
rect 882 601 912 627
rect 968 601 998 627
rect 1054 601 1084 627
rect 1140 601 1170 627
rect 1226 601 1256 627
rect 1312 601 1342 627
rect 1398 601 1428 627
rect 1484 601 1514 627
rect 1685 619 1715 645
rect 1771 619 1801 645
rect 1857 619 1887 645
rect 1943 619 1973 645
rect 83 325 113 367
rect 169 325 199 367
rect 255 325 285 367
rect 341 325 371 367
rect 434 335 464 367
rect 520 335 550 367
rect 606 335 636 367
rect 692 335 722 367
rect 33 309 371 325
rect 33 275 49 309
rect 83 275 117 309
rect 151 275 185 309
rect 219 275 253 309
rect 287 275 321 309
rect 355 275 371 309
rect 33 259 371 275
rect 413 319 751 335
rect 413 285 429 319
rect 463 285 497 319
rect 531 285 565 319
rect 599 285 633 319
rect 667 285 701 319
rect 735 285 751 319
rect 882 317 912 349
rect 968 317 998 349
rect 1054 317 1084 349
rect 1140 317 1170 349
rect 413 269 751 285
rect 793 301 1170 317
rect 83 215 113 259
rect 169 215 199 259
rect 255 215 285 259
rect 341 215 371 259
rect 427 215 457 269
rect 513 215 543 269
rect 599 215 629 269
rect 685 215 715 269
rect 793 267 809 301
rect 843 267 877 301
rect 911 267 945 301
rect 979 267 1013 301
rect 1047 267 1081 301
rect 1115 267 1170 301
rect 793 251 1170 267
rect 1226 303 1256 349
rect 1312 303 1342 349
rect 1398 303 1428 349
rect 1484 303 1514 349
rect 1685 333 1715 367
rect 1771 333 1801 367
rect 1857 333 1887 367
rect 1943 333 1973 367
rect 1685 303 1973 333
rect 1226 287 1643 303
rect 1226 253 1253 287
rect 1287 253 1321 287
rect 1355 253 1389 287
rect 1423 253 1457 287
rect 1491 253 1525 287
rect 1559 253 1593 287
rect 1627 253 1643 287
rect 793 215 823 251
rect 879 215 909 251
rect 979 215 1009 251
rect 1079 215 1109 251
rect 1226 237 1643 253
rect 1685 287 2091 303
rect 1685 253 1701 287
rect 1735 253 1769 287
rect 1803 253 1837 287
rect 1871 253 1905 287
rect 1939 253 1973 287
rect 2007 253 2041 287
rect 2075 253 2091 287
rect 1685 237 2091 253
rect 1258 215 1288 237
rect 1344 215 1374 237
rect 1430 215 1460 237
rect 1590 215 1620 237
rect 1685 215 1715 237
rect 1771 215 1801 237
rect 1857 215 1887 237
rect 1943 215 1973 237
rect 83 21 113 47
rect 169 21 199 47
rect 255 21 285 47
rect 341 21 371 47
rect 427 21 457 47
rect 513 21 543 47
rect 599 21 629 47
rect 685 21 715 47
rect 793 21 823 47
rect 879 21 909 47
rect 979 21 1009 47
rect 1079 21 1109 47
rect 1258 21 1288 47
rect 1344 21 1374 47
rect 1430 21 1460 47
rect 1590 21 1620 47
rect 1685 21 1715 47
rect 1771 21 1801 47
rect 1857 21 1887 47
rect 1943 21 1973 47
<< polycont >>
rect 49 275 83 309
rect 117 275 151 309
rect 185 275 219 309
rect 253 275 287 309
rect 321 275 355 309
rect 429 285 463 319
rect 497 285 531 319
rect 565 285 599 319
rect 633 285 667 319
rect 701 285 735 319
rect 809 267 843 301
rect 877 267 911 301
rect 945 267 979 301
rect 1013 267 1047 301
rect 1081 267 1115 301
rect 1253 253 1287 287
rect 1321 253 1355 287
rect 1389 253 1423 287
rect 1457 253 1491 287
rect 1525 253 1559 287
rect 1593 253 1627 287
rect 1701 253 1735 287
rect 1769 253 1803 287
rect 1837 253 1871 287
rect 1905 253 1939 287
rect 1973 253 2007 287
rect 2041 253 2075 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 22 599 425 615
rect 22 565 38 599
rect 72 581 210 599
rect 72 565 74 581
rect 22 520 74 565
rect 208 565 210 581
rect 244 581 389 599
rect 244 565 246 581
rect 22 486 38 520
rect 72 486 74 520
rect 22 438 74 486
rect 22 404 38 438
rect 72 404 74 438
rect 22 388 74 404
rect 108 538 174 547
rect 108 504 124 538
rect 158 504 174 538
rect 108 436 174 504
rect 208 504 246 565
rect 387 565 389 581
rect 423 565 425 599
rect 208 470 210 504
rect 244 470 246 504
rect 208 454 246 470
rect 280 538 353 547
rect 280 504 296 538
rect 330 504 353 538
rect 108 402 124 436
rect 158 420 174 436
rect 280 436 353 504
rect 387 504 425 565
rect 459 568 525 649
rect 459 534 475 568
rect 509 534 525 568
rect 459 524 525 534
rect 559 599 597 615
rect 559 565 561 599
rect 595 565 597 599
rect 387 470 389 504
rect 423 490 425 504
rect 559 504 597 565
rect 631 568 697 649
rect 631 534 647 568
rect 681 534 697 568
rect 631 524 697 534
rect 731 599 783 615
rect 731 565 733 599
rect 767 565 783 599
rect 559 490 561 504
rect 423 470 561 490
rect 595 490 597 504
rect 731 504 783 565
rect 731 490 733 504
rect 595 470 733 490
rect 767 470 783 504
rect 387 454 783 470
rect 821 589 1575 615
rect 821 555 837 589
rect 871 581 1009 589
rect 871 555 875 581
rect 821 504 875 555
rect 998 555 1009 581
rect 1043 581 1181 589
rect 1043 555 1049 581
rect 821 470 837 504
rect 871 470 875 504
rect 821 454 875 470
rect 914 531 964 547
rect 914 497 923 531
rect 957 497 964 531
rect 280 420 296 436
rect 158 402 296 420
rect 330 420 353 436
rect 914 436 964 497
rect 998 504 1049 555
rect 1170 555 1181 581
rect 1215 581 1353 589
rect 1215 555 1224 581
rect 998 470 1009 504
rect 1043 470 1049 504
rect 998 454 1049 470
rect 1083 531 1136 547
rect 1083 497 1095 531
rect 1129 497 1136 531
rect 914 420 923 436
rect 330 402 923 420
rect 957 420 964 436
rect 1083 436 1136 497
rect 1170 504 1224 555
rect 1343 555 1353 581
rect 1387 581 1525 589
rect 1387 555 1395 581
rect 1170 470 1181 504
rect 1215 470 1224 504
rect 1170 454 1224 470
rect 1258 529 1309 547
rect 1258 495 1267 529
rect 1301 495 1309 529
rect 1258 461 1309 495
rect 1083 420 1095 436
rect 957 402 1095 420
rect 1129 420 1136 436
rect 1258 427 1267 461
rect 1301 427 1309 461
rect 1129 402 1201 420
rect 108 386 1201 402
rect 31 309 371 352
rect 31 275 49 309
rect 83 275 117 309
rect 151 275 185 309
rect 219 275 253 309
rect 287 275 321 309
rect 355 275 371 309
rect 413 319 751 352
rect 413 285 429 319
rect 463 285 497 319
rect 531 285 565 319
rect 599 285 633 319
rect 667 285 701 319
rect 735 285 751 319
rect 793 301 1131 352
rect 793 267 809 301
rect 843 267 877 301
rect 911 267 945 301
rect 979 267 1013 301
rect 1047 267 1081 301
rect 1115 267 1131 301
rect 114 233 682 235
rect 1167 233 1201 386
rect 1258 391 1309 427
rect 1343 519 1395 555
rect 1516 555 1525 581
rect 1559 555 1575 589
rect 1343 485 1353 519
rect 1387 485 1395 519
rect 1343 451 1395 485
rect 1343 417 1353 451
rect 1387 417 1395 451
rect 1343 401 1395 417
rect 1429 531 1482 547
rect 1429 497 1439 531
rect 1473 497 1482 531
rect 1429 463 1482 497
rect 1429 429 1439 463
rect 1473 429 1482 463
rect 1258 357 1267 391
rect 1301 367 1309 391
rect 1429 391 1482 429
rect 1516 519 1575 555
rect 1516 485 1525 519
rect 1559 485 1575 519
rect 1516 451 1575 485
rect 1516 417 1525 451
rect 1559 417 1575 451
rect 1516 401 1575 417
rect 1624 607 1690 649
rect 1624 573 1640 607
rect 1674 573 1690 607
rect 1624 518 1690 573
rect 1624 484 1640 518
rect 1674 484 1690 518
rect 1624 435 1690 484
rect 1624 401 1640 435
rect 1674 401 1690 435
rect 1724 599 1762 615
rect 1724 565 1726 599
rect 1760 565 1762 599
rect 1724 506 1762 565
rect 1724 472 1726 506
rect 1760 472 1762 506
rect 1724 413 1762 472
rect 1429 367 1439 391
rect 1301 357 1439 367
rect 1473 367 1482 391
rect 1724 379 1726 413
rect 1760 379 1762 413
rect 1796 607 1862 649
rect 1796 573 1812 607
rect 1846 573 1862 607
rect 1796 518 1862 573
rect 1796 484 1812 518
rect 1846 484 1862 518
rect 1796 435 1862 484
rect 1796 401 1812 435
rect 1846 401 1862 435
rect 1896 599 1942 615
rect 1896 565 1898 599
rect 1932 565 1942 599
rect 1896 506 1942 565
rect 1896 472 1898 506
rect 1932 472 1942 506
rect 1896 413 1942 472
rect 1724 367 1762 379
rect 1896 379 1898 413
rect 1932 379 1942 413
rect 1896 367 1942 379
rect 1473 357 1942 367
rect 1976 607 2034 649
rect 1976 573 1984 607
rect 2018 573 2034 607
rect 1976 504 2034 573
rect 1976 470 1984 504
rect 2018 470 2034 504
rect 1976 413 2034 470
rect 1976 379 1984 413
rect 2018 379 2034 413
rect 1976 363 2034 379
rect 1258 333 1942 357
rect 1237 287 1643 299
rect 1237 253 1253 287
rect 1287 253 1321 287
rect 1355 253 1389 287
rect 1423 253 1457 287
rect 1491 253 1525 287
rect 1559 253 1593 287
rect 1627 253 1643 287
rect 1237 242 1643 253
rect 1685 287 2091 299
rect 1685 253 1701 287
rect 1735 253 1769 287
rect 1803 253 1837 287
rect 1871 253 1905 287
rect 1939 253 1973 287
rect 2007 253 2041 287
rect 2075 253 2091 287
rect 1685 242 2091 253
rect 22 203 80 219
rect 22 169 38 203
rect 72 169 80 203
rect 22 105 80 169
rect 114 201 1201 233
rect 114 169 160 201
rect 114 135 124 169
rect 158 135 160 169
rect 294 169 332 201
rect 114 119 160 135
rect 194 163 260 167
rect 194 129 210 163
rect 244 129 260 163
rect 22 71 38 105
rect 72 85 80 105
rect 194 93 260 129
rect 294 135 296 169
rect 330 135 332 169
rect 466 169 504 201
rect 294 119 332 135
rect 366 163 432 167
rect 366 129 382 163
rect 416 129 432 163
rect 194 85 210 93
rect 72 71 210 85
rect 22 59 210 71
rect 244 85 260 93
rect 366 93 432 129
rect 466 135 468 169
rect 502 135 504 169
rect 638 199 1201 201
rect 638 173 676 199
rect 466 119 504 135
rect 538 163 604 167
rect 538 129 554 163
rect 588 129 604 163
rect 366 85 382 93
rect 244 59 382 85
rect 416 85 432 93
rect 538 93 604 129
rect 638 139 640 173
rect 674 139 676 173
rect 1235 192 2034 208
rect 1235 174 1385 192
rect 1235 165 1269 174
rect 638 123 676 139
rect 710 163 920 165
rect 710 129 726 163
rect 760 131 920 163
rect 954 131 1120 165
rect 1154 131 1269 165
rect 760 129 776 131
rect 538 85 554 93
rect 416 59 554 85
rect 588 89 604 93
rect 710 89 776 129
rect 588 59 726 89
rect 22 55 726 59
rect 760 55 776 89
rect 22 51 776 55
rect 818 89 884 97
rect 818 55 834 89
rect 868 55 884 89
rect 818 17 884 55
rect 918 92 984 131
rect 1118 129 1269 131
rect 1383 158 1385 174
rect 1419 174 1631 192
rect 1419 158 1428 174
rect 1118 127 1247 129
rect 918 58 934 92
rect 968 58 984 92
rect 918 51 984 58
rect 1018 89 1084 97
rect 1018 55 1034 89
rect 1068 55 1084 89
rect 1018 17 1084 55
rect 1118 93 1202 127
rect 1236 93 1247 127
rect 1383 101 1428 158
rect 1622 158 1631 174
rect 1665 174 1812 192
rect 1665 158 1676 174
rect 1118 89 1247 93
rect 1118 55 1134 89
rect 1168 55 1247 89
rect 1118 51 1247 55
rect 1281 89 1349 95
rect 1281 55 1299 89
rect 1333 55 1349 89
rect 1281 17 1349 55
rect 1383 67 1385 101
rect 1419 67 1428 101
rect 1383 51 1428 67
rect 1462 124 1588 140
rect 1462 90 1471 124
rect 1505 90 1545 124
rect 1579 90 1588 124
rect 1462 17 1588 90
rect 1622 101 1676 158
rect 1810 158 1812 174
rect 1846 174 1984 192
rect 1846 158 1848 174
rect 1622 67 1631 101
rect 1665 67 1676 101
rect 1622 51 1676 67
rect 1710 124 1776 140
rect 1710 90 1726 124
rect 1760 90 1776 124
rect 1710 17 1776 90
rect 1810 101 1848 158
rect 1982 158 1984 174
rect 2018 158 2034 192
rect 1810 67 1812 101
rect 1846 67 1848 101
rect 1810 51 1848 67
rect 1882 124 1948 140
rect 1882 90 1898 124
rect 1932 90 1948 124
rect 1882 17 1948 90
rect 1982 101 2034 158
rect 1982 67 1984 101
rect 2018 67 2034 101
rect 1982 51 2034 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o32ai_4
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1858158
string GDS_START 1839964
<< end >>
