magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 1 49 762 248
rect 0 0 768 49
<< scpmos >>
rect 88 368 118 592
rect 214 368 244 568
rect 304 368 334 568
rect 452 368 482 568
rect 542 368 572 568
rect 652 368 682 568
<< nmoslvt >>
rect 84 74 114 222
rect 229 94 259 222
rect 307 94 337 222
rect 415 94 445 222
rect 571 94 601 222
rect 649 94 679 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 126 229 222
rect 114 92 153 126
rect 187 94 229 126
rect 259 94 307 222
rect 337 94 415 222
rect 445 204 571 222
rect 445 170 456 204
rect 490 170 526 204
rect 560 170 571 204
rect 445 136 571 170
rect 445 102 456 136
rect 490 102 526 136
rect 560 102 571 136
rect 445 94 571 102
rect 601 94 649 222
rect 679 208 736 222
rect 679 174 690 208
rect 724 174 736 208
rect 679 140 736 174
rect 679 106 690 140
rect 724 106 736 140
rect 679 94 736 106
rect 187 92 214 94
rect 114 74 214 92
<< pdiff >>
rect 29 580 88 592
rect 29 546 41 580
rect 75 546 88 580
rect 29 497 88 546
rect 29 463 41 497
rect 75 463 88 497
rect 29 414 88 463
rect 29 380 41 414
rect 75 380 88 414
rect 29 368 88 380
rect 118 580 187 592
rect 118 546 141 580
rect 175 568 187 580
rect 175 546 214 568
rect 118 462 214 546
rect 118 428 153 462
rect 187 428 214 462
rect 118 368 214 428
rect 244 556 304 568
rect 244 522 257 556
rect 291 522 304 556
rect 244 453 304 522
rect 244 419 257 453
rect 291 419 304 453
rect 244 368 304 419
rect 334 530 452 568
rect 334 496 376 530
rect 410 496 452 530
rect 334 368 452 496
rect 482 556 542 568
rect 482 522 495 556
rect 529 522 542 556
rect 482 453 542 522
rect 482 419 495 453
rect 529 419 542 453
rect 482 368 542 419
rect 572 547 652 568
rect 572 513 595 547
rect 629 513 652 547
rect 572 479 652 513
rect 572 445 595 479
rect 629 445 652 479
rect 572 411 652 445
rect 572 377 595 411
rect 629 377 652 411
rect 572 368 652 377
rect 682 556 741 568
rect 682 522 695 556
rect 729 522 741 556
rect 682 485 741 522
rect 682 451 695 485
rect 729 451 741 485
rect 682 414 741 451
rect 682 380 695 414
rect 729 380 741 414
rect 682 368 741 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 153 92 187 126
rect 456 170 490 204
rect 526 170 560 204
rect 456 102 490 136
rect 526 102 560 136
rect 690 174 724 208
rect 690 106 724 140
<< pdiffc >>
rect 41 546 75 580
rect 41 463 75 497
rect 41 380 75 414
rect 141 546 175 580
rect 153 428 187 462
rect 257 522 291 556
rect 257 419 291 453
rect 376 496 410 530
rect 495 522 529 556
rect 495 419 529 453
rect 595 513 629 547
rect 595 445 629 479
rect 595 377 629 411
rect 695 522 729 556
rect 695 451 729 485
rect 695 380 729 414
<< poly >>
rect 88 592 118 618
rect 214 568 244 594
rect 304 568 334 594
rect 452 568 482 594
rect 542 568 572 594
rect 652 568 682 594
rect 88 353 118 368
rect 214 353 244 368
rect 304 353 334 368
rect 452 353 482 368
rect 542 353 572 368
rect 652 353 682 368
rect 85 326 121 353
rect 84 310 151 326
rect 211 310 247 353
rect 301 310 337 353
rect 449 310 485 353
rect 539 310 575 353
rect 649 310 685 353
rect 84 276 101 310
rect 135 276 151 310
rect 84 260 151 276
rect 193 294 259 310
rect 193 260 209 294
rect 243 260 259 294
rect 84 222 114 260
rect 193 244 259 260
rect 301 294 367 310
rect 301 260 317 294
rect 351 260 367 294
rect 301 244 367 260
rect 409 294 485 310
rect 409 260 425 294
rect 459 260 485 294
rect 409 244 485 260
rect 535 294 601 310
rect 535 260 551 294
rect 585 260 601 294
rect 535 244 601 260
rect 229 222 259 244
rect 307 222 337 244
rect 415 222 445 244
rect 571 222 601 244
rect 649 294 724 310
rect 649 260 674 294
rect 708 260 724 294
rect 649 244 724 260
rect 649 222 679 244
rect 84 48 114 74
rect 229 68 259 94
rect 307 68 337 94
rect 415 68 445 94
rect 571 68 601 94
rect 649 68 679 94
<< polycont >>
rect 101 276 135 310
rect 209 260 243 294
rect 317 260 351 294
rect 425 260 459 294
rect 551 260 585 294
rect 674 260 708 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 580 91 596
rect 17 546 41 580
rect 75 546 91 580
rect 17 497 91 546
rect 17 463 41 497
rect 75 463 91 497
rect 17 414 91 463
rect 17 380 41 414
rect 75 380 91 414
rect 125 580 203 649
rect 125 546 141 580
rect 175 546 203 580
rect 125 462 203 546
rect 125 428 153 462
rect 187 428 203 462
rect 125 412 203 428
rect 241 556 307 572
rect 241 522 257 556
rect 291 522 307 556
rect 241 453 307 522
rect 360 530 426 649
rect 360 496 376 530
rect 410 496 426 530
rect 360 480 426 496
rect 479 581 745 615
rect 479 556 545 581
rect 479 522 495 556
rect 529 522 545 556
rect 679 556 745 581
rect 241 419 257 453
rect 291 446 307 453
rect 479 453 545 522
rect 479 446 495 453
rect 291 419 495 446
rect 529 419 545 453
rect 241 412 545 419
rect 579 513 595 547
rect 629 513 645 547
rect 579 479 645 513
rect 579 445 595 479
rect 629 445 645 479
rect 17 364 91 380
rect 579 411 645 445
rect 579 378 595 411
rect 125 377 595 378
rect 629 377 645 411
rect 17 226 51 364
rect 125 344 645 377
rect 679 522 695 556
rect 729 522 745 556
rect 679 485 745 522
rect 679 451 695 485
rect 729 451 745 485
rect 679 414 745 451
rect 679 380 695 414
rect 729 380 745 414
rect 679 364 745 380
rect 125 326 159 344
rect 85 310 159 326
rect 85 276 101 310
rect 135 276 159 310
rect 85 260 159 276
rect 17 210 89 226
rect 17 176 39 210
rect 73 176 89 210
rect 17 120 89 176
rect 125 204 159 260
rect 193 294 263 310
rect 193 260 209 294
rect 243 260 263 294
rect 193 238 263 260
rect 301 294 367 310
rect 301 260 317 294
rect 351 260 367 294
rect 301 238 367 260
rect 409 294 475 310
rect 409 260 425 294
rect 459 260 475 294
rect 409 238 475 260
rect 509 294 601 310
rect 509 260 551 294
rect 585 260 601 294
rect 509 238 601 260
rect 658 294 743 310
rect 658 260 674 294
rect 708 260 743 294
rect 658 242 743 260
rect 125 170 456 204
rect 490 170 526 204
rect 560 170 576 204
rect 440 136 576 170
rect 17 86 39 120
rect 73 86 89 120
rect 17 70 89 86
rect 130 126 210 136
rect 130 92 153 126
rect 187 92 210 126
rect 130 17 210 92
rect 440 102 456 136
rect 490 102 526 136
rect 560 102 576 136
rect 440 86 576 102
rect 674 174 690 208
rect 724 174 740 208
rect 674 140 740 174
rect 674 106 690 140
rect 724 106 740 140
rect 674 17 740 106
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a32o_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 1041462
string GDS_START 1034424
<< end >>
