magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 21 49 2015 241
rect 0 0 2016 49
<< scnmos >>
rect 100 47 130 215
rect 186 47 216 215
rect 272 47 302 215
rect 358 47 388 215
rect 444 47 474 215
rect 530 47 560 215
rect 616 47 646 215
rect 702 47 732 215
rect 788 47 818 215
rect 874 47 904 215
rect 960 47 990 215
rect 1046 47 1076 215
rect 1132 47 1162 215
rect 1218 47 1248 215
rect 1304 47 1334 215
rect 1390 47 1420 215
rect 1476 47 1506 215
rect 1562 47 1592 215
rect 1648 47 1678 215
rect 1734 47 1764 215
rect 1820 47 1850 215
rect 1906 47 1936 215
<< scpmoshvt >>
rect 100 367 130 619
rect 186 367 216 619
rect 272 367 302 619
rect 358 367 388 619
rect 444 367 474 619
rect 530 367 560 619
rect 616 367 646 619
rect 702 367 732 619
rect 788 367 818 619
rect 874 367 904 619
rect 960 367 990 619
rect 1046 367 1076 619
rect 1132 367 1162 619
rect 1218 367 1248 619
rect 1304 367 1334 619
rect 1390 367 1420 619
rect 1476 367 1506 619
rect 1562 367 1592 619
rect 1648 367 1678 619
rect 1734 367 1764 619
rect 1820 367 1850 619
rect 1906 367 1936 619
<< ndiff >>
rect 47 192 100 215
rect 47 158 55 192
rect 89 158 100 192
rect 47 103 100 158
rect 47 69 55 103
rect 89 69 100 103
rect 47 47 100 69
rect 130 203 186 215
rect 130 169 141 203
rect 175 169 186 203
rect 130 135 186 169
rect 130 101 141 135
rect 175 101 186 135
rect 130 47 186 101
rect 216 159 272 215
rect 216 125 227 159
rect 261 125 272 159
rect 216 91 272 125
rect 216 57 227 91
rect 261 57 272 91
rect 216 47 272 57
rect 302 203 358 215
rect 302 169 313 203
rect 347 169 358 203
rect 302 135 358 169
rect 302 101 313 135
rect 347 101 358 135
rect 302 47 358 101
rect 388 129 444 215
rect 388 95 399 129
rect 433 95 444 129
rect 388 47 444 95
rect 474 203 530 215
rect 474 169 485 203
rect 519 169 530 203
rect 474 135 530 169
rect 474 101 485 135
rect 519 101 530 135
rect 474 47 530 101
rect 560 159 616 215
rect 560 125 571 159
rect 605 125 616 159
rect 560 91 616 125
rect 560 57 571 91
rect 605 57 616 91
rect 560 47 616 57
rect 646 185 702 215
rect 646 151 657 185
rect 691 151 702 185
rect 646 111 702 151
rect 646 77 657 111
rect 691 77 702 111
rect 646 47 702 77
rect 732 185 788 215
rect 732 151 743 185
rect 777 151 788 185
rect 732 111 788 151
rect 732 77 743 111
rect 777 77 788 111
rect 732 47 788 77
rect 818 185 874 215
rect 818 151 829 185
rect 863 151 874 185
rect 818 111 874 151
rect 818 77 829 111
rect 863 77 874 111
rect 818 47 874 77
rect 904 185 960 215
rect 904 151 915 185
rect 949 151 960 185
rect 904 111 960 151
rect 904 77 915 111
rect 949 77 960 111
rect 904 47 960 77
rect 990 185 1046 215
rect 990 151 1001 185
rect 1035 151 1046 185
rect 990 111 1046 151
rect 990 77 1001 111
rect 1035 77 1046 111
rect 990 47 1046 77
rect 1076 185 1132 215
rect 1076 151 1087 185
rect 1121 151 1132 185
rect 1076 111 1132 151
rect 1076 77 1087 111
rect 1121 77 1132 111
rect 1076 47 1132 77
rect 1162 185 1218 215
rect 1162 151 1173 185
rect 1207 151 1218 185
rect 1162 111 1218 151
rect 1162 77 1173 111
rect 1207 77 1218 111
rect 1162 47 1218 77
rect 1248 185 1304 215
rect 1248 151 1259 185
rect 1293 151 1304 185
rect 1248 111 1304 151
rect 1248 77 1259 111
rect 1293 77 1304 111
rect 1248 47 1304 77
rect 1334 185 1390 215
rect 1334 151 1345 185
rect 1379 151 1390 185
rect 1334 111 1390 151
rect 1334 77 1345 111
rect 1379 77 1390 111
rect 1334 47 1390 77
rect 1420 185 1476 215
rect 1420 151 1431 185
rect 1465 151 1476 185
rect 1420 111 1476 151
rect 1420 77 1431 111
rect 1465 77 1476 111
rect 1420 47 1476 77
rect 1506 185 1562 215
rect 1506 151 1517 185
rect 1551 151 1562 185
rect 1506 111 1562 151
rect 1506 77 1517 111
rect 1551 77 1562 111
rect 1506 47 1562 77
rect 1592 185 1648 215
rect 1592 151 1603 185
rect 1637 151 1648 185
rect 1592 111 1648 151
rect 1592 77 1603 111
rect 1637 77 1648 111
rect 1592 47 1648 77
rect 1678 185 1734 215
rect 1678 151 1689 185
rect 1723 151 1734 185
rect 1678 111 1734 151
rect 1678 77 1689 111
rect 1723 77 1734 111
rect 1678 47 1734 77
rect 1764 185 1820 215
rect 1764 151 1775 185
rect 1809 151 1820 185
rect 1764 111 1820 151
rect 1764 77 1775 111
rect 1809 77 1820 111
rect 1764 47 1820 77
rect 1850 185 1906 215
rect 1850 151 1861 185
rect 1895 151 1906 185
rect 1850 111 1906 151
rect 1850 77 1861 111
rect 1895 77 1906 111
rect 1850 47 1906 77
rect 1936 185 1989 215
rect 1936 151 1947 185
rect 1981 151 1989 185
rect 1936 111 1989 151
rect 1936 77 1947 111
rect 1981 77 1989 111
rect 1936 47 1989 77
<< pdiff >>
rect 47 590 100 619
rect 47 556 55 590
rect 89 556 100 590
rect 47 506 100 556
rect 47 472 55 506
rect 89 472 100 506
rect 47 422 100 472
rect 47 388 55 422
rect 89 388 100 422
rect 47 367 100 388
rect 130 590 186 619
rect 130 556 141 590
rect 175 556 186 590
rect 130 506 186 556
rect 130 472 141 506
rect 175 472 186 506
rect 130 422 186 472
rect 130 388 141 422
rect 175 388 186 422
rect 130 367 186 388
rect 216 605 272 619
rect 216 571 227 605
rect 261 571 272 605
rect 216 537 272 571
rect 216 503 227 537
rect 261 503 272 537
rect 216 469 272 503
rect 216 435 227 469
rect 261 435 272 469
rect 216 367 272 435
rect 302 590 358 619
rect 302 556 313 590
rect 347 556 358 590
rect 302 506 358 556
rect 302 472 313 506
rect 347 472 358 506
rect 302 422 358 472
rect 302 388 313 422
rect 347 388 358 422
rect 302 367 358 388
rect 388 605 444 619
rect 388 571 399 605
rect 433 571 444 605
rect 388 537 444 571
rect 388 503 399 537
rect 433 503 444 537
rect 388 469 444 503
rect 388 435 399 469
rect 433 435 444 469
rect 388 367 444 435
rect 474 590 530 619
rect 474 556 485 590
rect 519 556 530 590
rect 474 506 530 556
rect 474 472 485 506
rect 519 472 530 506
rect 474 422 530 472
rect 474 388 485 422
rect 519 388 530 422
rect 474 367 530 388
rect 560 605 616 619
rect 560 571 571 605
rect 605 571 616 605
rect 560 537 616 571
rect 560 503 571 537
rect 605 503 616 537
rect 560 469 616 503
rect 560 435 571 469
rect 605 435 616 469
rect 560 367 616 435
rect 646 590 702 619
rect 646 556 657 590
rect 691 556 702 590
rect 646 506 702 556
rect 646 472 657 506
rect 691 472 702 506
rect 646 422 702 472
rect 646 388 657 422
rect 691 388 702 422
rect 646 367 702 388
rect 732 595 788 619
rect 732 561 743 595
rect 777 561 788 595
rect 732 515 788 561
rect 732 481 743 515
rect 777 481 788 515
rect 732 434 788 481
rect 732 400 743 434
rect 777 400 788 434
rect 732 367 788 400
rect 818 590 874 619
rect 818 556 829 590
rect 863 556 874 590
rect 818 506 874 556
rect 818 472 829 506
rect 863 472 874 506
rect 818 422 874 472
rect 818 388 829 422
rect 863 388 874 422
rect 818 367 874 388
rect 904 595 960 619
rect 904 561 915 595
rect 949 561 960 595
rect 904 515 960 561
rect 904 481 915 515
rect 949 481 960 515
rect 904 434 960 481
rect 904 400 915 434
rect 949 400 960 434
rect 904 367 960 400
rect 990 590 1046 619
rect 990 556 1001 590
rect 1035 556 1046 590
rect 990 506 1046 556
rect 990 472 1001 506
rect 1035 472 1046 506
rect 990 422 1046 472
rect 990 388 1001 422
rect 1035 388 1046 422
rect 990 367 1046 388
rect 1076 595 1132 619
rect 1076 561 1087 595
rect 1121 561 1132 595
rect 1076 515 1132 561
rect 1076 481 1087 515
rect 1121 481 1132 515
rect 1076 434 1132 481
rect 1076 400 1087 434
rect 1121 400 1132 434
rect 1076 367 1132 400
rect 1162 590 1218 619
rect 1162 556 1173 590
rect 1207 556 1218 590
rect 1162 506 1218 556
rect 1162 472 1173 506
rect 1207 472 1218 506
rect 1162 422 1218 472
rect 1162 388 1173 422
rect 1207 388 1218 422
rect 1162 367 1218 388
rect 1248 595 1304 619
rect 1248 561 1259 595
rect 1293 561 1304 595
rect 1248 515 1304 561
rect 1248 481 1259 515
rect 1293 481 1304 515
rect 1248 434 1304 481
rect 1248 400 1259 434
rect 1293 400 1304 434
rect 1248 367 1304 400
rect 1334 590 1390 619
rect 1334 556 1345 590
rect 1379 556 1390 590
rect 1334 506 1390 556
rect 1334 472 1345 506
rect 1379 472 1390 506
rect 1334 422 1390 472
rect 1334 388 1345 422
rect 1379 388 1390 422
rect 1334 367 1390 388
rect 1420 595 1476 619
rect 1420 561 1431 595
rect 1465 561 1476 595
rect 1420 515 1476 561
rect 1420 481 1431 515
rect 1465 481 1476 515
rect 1420 434 1476 481
rect 1420 400 1431 434
rect 1465 400 1476 434
rect 1420 367 1476 400
rect 1506 590 1562 619
rect 1506 556 1517 590
rect 1551 556 1562 590
rect 1506 506 1562 556
rect 1506 472 1517 506
rect 1551 472 1562 506
rect 1506 422 1562 472
rect 1506 388 1517 422
rect 1551 388 1562 422
rect 1506 367 1562 388
rect 1592 595 1648 619
rect 1592 561 1603 595
rect 1637 561 1648 595
rect 1592 515 1648 561
rect 1592 481 1603 515
rect 1637 481 1648 515
rect 1592 434 1648 481
rect 1592 400 1603 434
rect 1637 400 1648 434
rect 1592 367 1648 400
rect 1678 590 1734 619
rect 1678 556 1689 590
rect 1723 556 1734 590
rect 1678 506 1734 556
rect 1678 472 1689 506
rect 1723 472 1734 506
rect 1678 422 1734 472
rect 1678 388 1689 422
rect 1723 388 1734 422
rect 1678 367 1734 388
rect 1764 595 1820 619
rect 1764 561 1775 595
rect 1809 561 1820 595
rect 1764 515 1820 561
rect 1764 481 1775 515
rect 1809 481 1820 515
rect 1764 434 1820 481
rect 1764 400 1775 434
rect 1809 400 1820 434
rect 1764 367 1820 400
rect 1850 590 1906 619
rect 1850 556 1861 590
rect 1895 556 1906 590
rect 1850 506 1906 556
rect 1850 472 1861 506
rect 1895 472 1906 506
rect 1850 422 1906 472
rect 1850 388 1861 422
rect 1895 388 1906 422
rect 1850 367 1906 388
rect 1936 595 1989 619
rect 1936 561 1947 595
rect 1981 561 1989 595
rect 1936 515 1989 561
rect 1936 481 1947 515
rect 1981 481 1989 515
rect 1936 434 1989 481
rect 1936 400 1947 434
rect 1981 400 1989 434
rect 1936 367 1989 400
<< ndiffc >>
rect 55 158 89 192
rect 55 69 89 103
rect 141 169 175 203
rect 141 101 175 135
rect 227 125 261 159
rect 227 57 261 91
rect 313 169 347 203
rect 313 101 347 135
rect 399 95 433 129
rect 485 169 519 203
rect 485 101 519 135
rect 571 125 605 159
rect 571 57 605 91
rect 657 151 691 185
rect 657 77 691 111
rect 743 151 777 185
rect 743 77 777 111
rect 829 151 863 185
rect 829 77 863 111
rect 915 151 949 185
rect 915 77 949 111
rect 1001 151 1035 185
rect 1001 77 1035 111
rect 1087 151 1121 185
rect 1087 77 1121 111
rect 1173 151 1207 185
rect 1173 77 1207 111
rect 1259 151 1293 185
rect 1259 77 1293 111
rect 1345 151 1379 185
rect 1345 77 1379 111
rect 1431 151 1465 185
rect 1431 77 1465 111
rect 1517 151 1551 185
rect 1517 77 1551 111
rect 1603 151 1637 185
rect 1603 77 1637 111
rect 1689 151 1723 185
rect 1689 77 1723 111
rect 1775 151 1809 185
rect 1775 77 1809 111
rect 1861 151 1895 185
rect 1861 77 1895 111
rect 1947 151 1981 185
rect 1947 77 1981 111
<< pdiffc >>
rect 55 556 89 590
rect 55 472 89 506
rect 55 388 89 422
rect 141 556 175 590
rect 141 472 175 506
rect 141 388 175 422
rect 227 571 261 605
rect 227 503 261 537
rect 227 435 261 469
rect 313 556 347 590
rect 313 472 347 506
rect 313 388 347 422
rect 399 571 433 605
rect 399 503 433 537
rect 399 435 433 469
rect 485 556 519 590
rect 485 472 519 506
rect 485 388 519 422
rect 571 571 605 605
rect 571 503 605 537
rect 571 435 605 469
rect 657 556 691 590
rect 657 472 691 506
rect 657 388 691 422
rect 743 561 777 595
rect 743 481 777 515
rect 743 400 777 434
rect 829 556 863 590
rect 829 472 863 506
rect 829 388 863 422
rect 915 561 949 595
rect 915 481 949 515
rect 915 400 949 434
rect 1001 556 1035 590
rect 1001 472 1035 506
rect 1001 388 1035 422
rect 1087 561 1121 595
rect 1087 481 1121 515
rect 1087 400 1121 434
rect 1173 556 1207 590
rect 1173 472 1207 506
rect 1173 388 1207 422
rect 1259 561 1293 595
rect 1259 481 1293 515
rect 1259 400 1293 434
rect 1345 556 1379 590
rect 1345 472 1379 506
rect 1345 388 1379 422
rect 1431 561 1465 595
rect 1431 481 1465 515
rect 1431 400 1465 434
rect 1517 556 1551 590
rect 1517 472 1551 506
rect 1517 388 1551 422
rect 1603 561 1637 595
rect 1603 481 1637 515
rect 1603 400 1637 434
rect 1689 556 1723 590
rect 1689 472 1723 506
rect 1689 388 1723 422
rect 1775 561 1809 595
rect 1775 481 1809 515
rect 1775 400 1809 434
rect 1861 556 1895 590
rect 1861 472 1895 506
rect 1861 388 1895 422
rect 1947 561 1981 595
rect 1947 481 1981 515
rect 1947 400 1981 434
<< poly >>
rect 100 619 130 645
rect 186 619 216 645
rect 272 619 302 645
rect 358 619 388 645
rect 444 619 474 645
rect 530 619 560 645
rect 616 619 646 645
rect 702 619 732 645
rect 788 619 818 645
rect 874 619 904 645
rect 960 619 990 645
rect 1046 619 1076 645
rect 1132 619 1162 645
rect 1218 619 1248 645
rect 1304 619 1334 645
rect 1390 619 1420 645
rect 1476 619 1506 645
rect 1562 619 1592 645
rect 1648 619 1678 645
rect 1734 619 1764 645
rect 1820 619 1850 645
rect 1906 619 1936 645
rect 100 329 130 367
rect 186 329 216 367
rect 272 329 302 367
rect 358 329 388 367
rect 444 329 474 367
rect 530 329 560 367
rect 73 313 560 329
rect 73 279 89 313
rect 123 279 157 313
rect 191 279 225 313
rect 259 279 293 313
rect 327 279 361 313
rect 395 279 429 313
rect 463 279 497 313
rect 531 279 560 313
rect 73 263 560 279
rect 100 215 130 263
rect 186 215 216 263
rect 272 215 302 263
rect 358 215 388 263
rect 444 215 474 263
rect 530 215 560 263
rect 616 345 646 367
rect 702 345 732 367
rect 616 331 732 345
rect 788 331 818 367
rect 874 331 904 367
rect 960 331 990 367
rect 1046 331 1076 367
rect 1132 331 1162 367
rect 1218 331 1248 367
rect 1304 331 1334 367
rect 1390 331 1420 367
rect 1476 331 1506 367
rect 1562 331 1592 367
rect 1648 331 1678 367
rect 1734 331 1764 367
rect 1820 331 1850 367
rect 1906 331 1936 367
rect 616 315 1936 331
rect 616 281 743 315
rect 777 281 915 315
rect 949 281 1087 315
rect 1121 281 1259 315
rect 1293 281 1431 315
rect 1465 281 1603 315
rect 1637 281 1775 315
rect 1809 281 1936 315
rect 616 267 1936 281
rect 616 215 646 267
rect 702 265 1936 267
rect 702 215 732 265
rect 788 215 818 265
rect 874 215 904 265
rect 960 215 990 265
rect 1046 215 1076 265
rect 1132 215 1162 265
rect 1218 215 1248 265
rect 1304 215 1334 265
rect 1390 215 1420 265
rect 1476 215 1506 265
rect 1562 215 1592 265
rect 1648 215 1678 265
rect 1734 215 1764 265
rect 1820 215 1850 265
rect 1906 215 1936 265
rect 100 21 130 47
rect 186 21 216 47
rect 272 21 302 47
rect 358 21 388 47
rect 444 21 474 47
rect 530 21 560 47
rect 616 21 646 47
rect 702 21 732 47
rect 788 21 818 47
rect 874 21 904 47
rect 960 21 990 47
rect 1046 21 1076 47
rect 1132 21 1162 47
rect 1218 21 1248 47
rect 1304 21 1334 47
rect 1390 21 1420 47
rect 1476 21 1506 47
rect 1562 21 1592 47
rect 1648 21 1678 47
rect 1734 21 1764 47
rect 1820 21 1850 47
rect 1906 21 1936 47
<< polycont >>
rect 89 279 123 313
rect 157 279 191 313
rect 225 279 259 313
rect 293 279 327 313
rect 361 279 395 313
rect 429 279 463 313
rect 497 279 531 313
rect 743 281 777 315
rect 915 281 949 315
rect 1087 281 1121 315
rect 1259 281 1293 315
rect 1431 281 1465 315
rect 1603 281 1637 315
rect 1775 281 1809 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 39 590 98 649
rect 39 556 55 590
rect 89 556 98 590
rect 39 506 98 556
rect 39 472 55 506
rect 89 472 98 506
rect 39 422 98 472
rect 39 388 55 422
rect 89 388 98 422
rect 39 363 98 388
rect 132 590 184 615
rect 132 556 141 590
rect 175 556 184 590
rect 132 506 184 556
rect 132 472 141 506
rect 175 472 184 506
rect 132 422 184 472
rect 132 388 141 422
rect 175 388 184 422
rect 218 605 270 649
rect 218 571 227 605
rect 261 571 270 605
rect 218 537 270 571
rect 218 503 227 537
rect 261 503 270 537
rect 218 469 270 503
rect 218 435 227 469
rect 261 435 270 469
rect 218 419 270 435
rect 304 590 356 615
rect 304 556 313 590
rect 347 556 356 590
rect 304 506 356 556
rect 304 472 313 506
rect 347 472 356 506
rect 304 422 356 472
rect 132 385 184 388
rect 304 388 313 422
rect 347 388 356 422
rect 390 605 442 649
rect 390 571 399 605
rect 433 571 442 605
rect 390 537 442 571
rect 390 503 399 537
rect 433 503 442 537
rect 390 469 442 503
rect 390 435 399 469
rect 433 435 442 469
rect 390 419 442 435
rect 476 590 528 615
rect 476 556 485 590
rect 519 556 528 590
rect 476 506 528 556
rect 476 472 485 506
rect 519 472 528 506
rect 476 422 528 472
rect 304 385 356 388
rect 476 388 485 422
rect 519 388 528 422
rect 562 605 619 649
rect 562 571 571 605
rect 605 571 619 605
rect 562 537 619 571
rect 562 503 571 537
rect 605 503 619 537
rect 562 469 619 503
rect 562 435 571 469
rect 605 435 619 469
rect 562 419 619 435
rect 653 590 700 615
rect 653 556 657 590
rect 691 556 700 590
rect 653 506 700 556
rect 653 472 657 506
rect 691 472 700 506
rect 653 424 700 472
rect 476 385 528 388
rect 653 388 657 424
rect 691 388 700 424
rect 132 351 619 385
rect 581 350 619 351
rect 73 313 547 317
rect 73 279 89 313
rect 123 279 157 313
rect 191 279 225 313
rect 259 279 293 313
rect 327 279 361 313
rect 395 279 429 313
rect 463 279 497 313
rect 531 279 547 313
rect 73 277 547 279
rect 581 316 583 350
rect 617 316 619 350
rect 39 192 98 215
rect 39 158 55 192
rect 89 158 98 192
rect 39 103 98 158
rect 39 69 55 103
rect 89 69 98 103
rect 132 209 347 243
rect 381 241 451 277
rect 581 243 619 316
rect 132 203 184 209
rect 132 169 141 203
rect 175 169 184 203
rect 306 207 347 209
rect 485 209 619 243
rect 485 207 528 209
rect 306 203 528 207
rect 132 135 184 169
rect 132 101 141 135
rect 175 101 184 135
rect 132 85 184 101
rect 218 159 272 175
rect 218 125 227 159
rect 261 125 272 159
rect 218 91 272 125
rect 39 17 98 69
rect 218 57 227 91
rect 261 57 272 91
rect 306 169 313 203
rect 347 173 485 203
rect 347 169 349 173
rect 306 135 349 169
rect 483 169 485 173
rect 519 169 528 203
rect 653 185 700 388
rect 734 595 786 649
rect 734 561 743 595
rect 777 561 786 595
rect 734 515 786 561
rect 734 481 743 515
rect 777 481 786 515
rect 734 434 786 481
rect 734 400 743 434
rect 777 400 786 434
rect 734 384 786 400
rect 820 590 872 615
rect 820 556 829 590
rect 863 556 872 590
rect 820 506 872 556
rect 820 472 829 506
rect 863 472 872 506
rect 820 424 872 472
rect 820 388 829 424
rect 863 388 872 424
rect 734 316 743 350
rect 777 316 786 350
rect 734 315 786 316
rect 734 281 743 315
rect 777 281 786 315
rect 734 265 786 281
rect 306 101 313 135
rect 347 101 349 135
rect 306 85 349 101
rect 383 129 449 139
rect 383 95 399 129
rect 433 95 449 129
rect 218 17 272 57
rect 383 17 449 95
rect 483 135 528 169
rect 483 101 485 135
rect 519 101 528 135
rect 483 85 528 101
rect 562 159 619 175
rect 562 125 571 159
rect 605 125 619 159
rect 562 91 619 125
rect 562 57 571 91
rect 605 57 619 91
rect 562 17 619 57
rect 653 151 657 185
rect 691 151 700 185
rect 653 111 700 151
rect 653 77 657 111
rect 691 77 700 111
rect 653 51 700 77
rect 734 185 786 215
rect 734 151 743 185
rect 777 151 786 185
rect 734 111 786 151
rect 734 77 743 111
rect 777 77 786 111
rect 734 17 786 77
rect 820 185 872 388
rect 906 595 958 649
rect 906 561 915 595
rect 949 561 958 595
rect 906 515 958 561
rect 906 481 915 515
rect 949 481 958 515
rect 906 434 958 481
rect 906 400 915 434
rect 949 400 958 434
rect 906 384 958 400
rect 992 590 1044 615
rect 992 556 1001 590
rect 1035 556 1044 590
rect 992 506 1044 556
rect 992 472 1001 506
rect 1035 472 1044 506
rect 992 424 1044 472
rect 992 388 1001 424
rect 1035 388 1044 424
rect 906 316 915 350
rect 949 316 958 350
rect 906 315 958 316
rect 906 281 915 315
rect 949 281 958 315
rect 906 265 958 281
rect 820 151 829 185
rect 863 151 872 185
rect 820 111 872 151
rect 820 77 829 111
rect 863 77 872 111
rect 820 51 872 77
rect 906 185 958 215
rect 906 151 915 185
rect 949 151 958 185
rect 906 111 958 151
rect 906 77 915 111
rect 949 77 958 111
rect 906 17 958 77
rect 992 185 1044 388
rect 1078 595 1130 649
rect 1078 561 1087 595
rect 1121 561 1130 595
rect 1078 515 1130 561
rect 1078 481 1087 515
rect 1121 481 1130 515
rect 1078 434 1130 481
rect 1078 400 1087 434
rect 1121 400 1130 434
rect 1078 384 1130 400
rect 1164 590 1216 615
rect 1164 556 1173 590
rect 1207 556 1216 590
rect 1164 506 1216 556
rect 1164 472 1173 506
rect 1207 472 1216 506
rect 1164 424 1216 472
rect 1164 388 1173 424
rect 1207 388 1216 424
rect 1078 316 1087 350
rect 1121 316 1130 350
rect 1078 315 1130 316
rect 1078 281 1087 315
rect 1121 281 1130 315
rect 1078 265 1130 281
rect 992 151 1001 185
rect 1035 151 1044 185
rect 992 111 1044 151
rect 992 77 1001 111
rect 1035 77 1044 111
rect 992 51 1044 77
rect 1078 185 1130 215
rect 1078 151 1087 185
rect 1121 151 1130 185
rect 1078 111 1130 151
rect 1078 77 1087 111
rect 1121 77 1130 111
rect 1078 17 1130 77
rect 1164 185 1216 388
rect 1250 595 1302 649
rect 1250 561 1259 595
rect 1293 561 1302 595
rect 1250 515 1302 561
rect 1250 481 1259 515
rect 1293 481 1302 515
rect 1250 434 1302 481
rect 1250 400 1259 434
rect 1293 400 1302 434
rect 1250 384 1302 400
rect 1336 590 1388 615
rect 1336 556 1345 590
rect 1379 556 1388 590
rect 1336 506 1388 556
rect 1336 472 1345 506
rect 1379 472 1388 506
rect 1336 424 1388 472
rect 1336 388 1345 424
rect 1379 388 1388 424
rect 1250 316 1259 350
rect 1293 316 1302 350
rect 1250 315 1302 316
rect 1250 281 1259 315
rect 1293 281 1302 315
rect 1250 265 1302 281
rect 1164 151 1173 185
rect 1207 151 1216 185
rect 1164 111 1216 151
rect 1164 77 1173 111
rect 1207 77 1216 111
rect 1164 51 1216 77
rect 1250 185 1302 215
rect 1250 151 1259 185
rect 1293 151 1302 185
rect 1250 111 1302 151
rect 1250 77 1259 111
rect 1293 77 1302 111
rect 1250 17 1302 77
rect 1336 185 1388 388
rect 1422 595 1474 649
rect 1422 561 1431 595
rect 1465 561 1474 595
rect 1422 515 1474 561
rect 1422 481 1431 515
rect 1465 481 1474 515
rect 1422 434 1474 481
rect 1422 400 1431 434
rect 1465 400 1474 434
rect 1422 384 1474 400
rect 1508 590 1560 615
rect 1508 556 1517 590
rect 1551 556 1560 590
rect 1508 506 1560 556
rect 1508 472 1517 506
rect 1551 472 1560 506
rect 1508 424 1560 472
rect 1508 388 1517 424
rect 1551 388 1560 424
rect 1422 316 1431 350
rect 1465 316 1474 350
rect 1422 315 1474 316
rect 1422 281 1431 315
rect 1465 281 1474 315
rect 1422 265 1474 281
rect 1336 151 1345 185
rect 1379 151 1388 185
rect 1336 111 1388 151
rect 1336 77 1345 111
rect 1379 77 1388 111
rect 1336 51 1388 77
rect 1422 185 1474 215
rect 1422 151 1431 185
rect 1465 151 1474 185
rect 1422 111 1474 151
rect 1422 77 1431 111
rect 1465 77 1474 111
rect 1422 17 1474 77
rect 1508 185 1560 388
rect 1594 595 1646 649
rect 1594 561 1603 595
rect 1637 561 1646 595
rect 1594 515 1646 561
rect 1594 481 1603 515
rect 1637 481 1646 515
rect 1594 434 1646 481
rect 1594 400 1603 434
rect 1637 400 1646 434
rect 1594 384 1646 400
rect 1680 590 1732 615
rect 1680 556 1689 590
rect 1723 556 1732 590
rect 1680 506 1732 556
rect 1680 472 1689 506
rect 1723 472 1732 506
rect 1680 424 1732 472
rect 1680 388 1689 424
rect 1723 388 1732 424
rect 1594 316 1603 350
rect 1637 316 1646 350
rect 1594 315 1646 316
rect 1594 281 1603 315
rect 1637 281 1646 315
rect 1594 265 1646 281
rect 1508 151 1517 185
rect 1551 151 1560 185
rect 1508 111 1560 151
rect 1508 77 1517 111
rect 1551 77 1560 111
rect 1508 51 1560 77
rect 1594 185 1646 215
rect 1594 151 1603 185
rect 1637 151 1646 185
rect 1594 111 1646 151
rect 1594 77 1603 111
rect 1637 77 1646 111
rect 1594 17 1646 77
rect 1680 185 1732 388
rect 1766 595 1818 649
rect 1766 561 1775 595
rect 1809 561 1818 595
rect 1766 515 1818 561
rect 1766 481 1775 515
rect 1809 481 1818 515
rect 1766 434 1818 481
rect 1766 400 1775 434
rect 1809 400 1818 434
rect 1766 384 1818 400
rect 1852 590 1904 615
rect 1852 556 1861 590
rect 1895 556 1904 590
rect 1852 506 1904 556
rect 1852 472 1861 506
rect 1895 472 1904 506
rect 1852 424 1904 472
rect 1852 388 1861 424
rect 1895 388 1904 424
rect 1766 316 1775 350
rect 1809 316 1818 350
rect 1766 315 1818 316
rect 1766 281 1775 315
rect 1809 281 1818 315
rect 1766 265 1818 281
rect 1680 151 1689 185
rect 1723 151 1732 185
rect 1680 111 1732 151
rect 1680 77 1689 111
rect 1723 77 1732 111
rect 1680 51 1732 77
rect 1766 185 1818 215
rect 1766 151 1775 185
rect 1809 151 1818 185
rect 1766 111 1818 151
rect 1766 77 1775 111
rect 1809 77 1818 111
rect 1766 17 1818 77
rect 1852 185 1904 388
rect 1938 595 1997 649
rect 1938 561 1947 595
rect 1981 561 1997 595
rect 1938 515 1997 561
rect 1938 481 1947 515
rect 1981 481 1997 515
rect 1938 434 1997 481
rect 1938 400 1947 434
rect 1981 400 1997 434
rect 1938 384 1997 400
rect 1852 151 1861 185
rect 1895 151 1904 185
rect 1852 111 1904 151
rect 1852 77 1861 111
rect 1895 77 1904 111
rect 1852 51 1904 77
rect 1938 185 1997 215
rect 1938 151 1947 185
rect 1981 151 1997 185
rect 1938 111 1997 151
rect 1938 77 1947 111
rect 1981 77 1997 111
rect 1938 17 1997 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 657 422 691 424
rect 657 390 691 422
rect 583 316 617 350
rect 829 422 863 424
rect 829 390 863 422
rect 743 316 777 350
rect 1001 422 1035 424
rect 1001 390 1035 422
rect 915 316 949 350
rect 1173 422 1207 424
rect 1173 390 1207 422
rect 1087 316 1121 350
rect 1345 422 1379 424
rect 1345 390 1379 422
rect 1259 316 1293 350
rect 1517 422 1551 424
rect 1517 390 1551 422
rect 1431 316 1465 350
rect 1689 422 1723 424
rect 1689 390 1723 422
rect 1603 316 1637 350
rect 1861 422 1895 424
rect 1861 390 1895 422
rect 1775 316 1809 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 645 424 1907 430
rect 645 390 657 424
rect 691 390 829 424
rect 863 390 1001 424
rect 1035 390 1173 424
rect 1207 390 1345 424
rect 1379 390 1517 424
rect 1551 390 1689 424
rect 1723 390 1861 424
rect 1895 390 1907 424
rect 645 384 1907 390
rect 571 350 1821 356
rect 571 316 583 350
rect 617 316 743 350
rect 777 316 915 350
rect 949 316 1087 350
rect 1121 316 1259 350
rect 1293 316 1431 350
rect 1465 316 1603 350
rect 1637 316 1775 350
rect 1809 316 1821 350
rect 571 310 1821 316
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 buf_16
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 645 384 1907 430 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5059460
string GDS_START 5042172
<< end >>
