magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 332 1478 704
<< pwell >>
rect 1 156 676 248
rect 848 156 1439 248
rect 1 49 1439 156
rect 0 0 1440 49
<< scpmos >>
rect 86 392 116 592
rect 176 392 206 592
rect 266 392 296 592
rect 366 392 396 592
rect 466 392 496 592
rect 566 392 596 592
rect 656 392 686 592
rect 746 392 776 592
rect 948 368 978 568
rect 1055 368 1085 592
rect 1145 368 1175 592
rect 1235 368 1265 592
rect 1325 368 1355 592
<< nmoslvt >>
rect 84 74 114 222
rect 198 74 228 222
rect 449 74 479 222
rect 563 74 593 222
rect 924 94 954 222
rect 1029 74 1059 222
rect 1140 74 1170 222
rect 1240 74 1270 222
rect 1326 74 1356 222
<< ndiff >>
rect 27 188 84 222
rect 27 154 39 188
rect 73 154 84 188
rect 27 120 84 154
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 120 198 222
rect 114 86 139 120
rect 173 86 198 120
rect 114 74 198 86
rect 228 188 449 222
rect 228 154 239 188
rect 273 154 314 188
rect 348 154 390 188
rect 424 154 449 188
rect 228 120 449 154
rect 228 86 239 120
rect 273 86 314 120
rect 348 86 390 120
rect 424 86 449 120
rect 228 74 449 86
rect 479 120 563 222
rect 479 86 492 120
rect 526 86 563 120
rect 479 74 563 86
rect 593 210 650 222
rect 593 176 604 210
rect 638 176 650 210
rect 593 120 650 176
rect 593 86 604 120
rect 638 86 650 120
rect 593 74 650 86
rect 874 130 924 222
rect 776 118 924 130
rect 776 84 788 118
rect 822 84 863 118
rect 897 94 924 118
rect 954 127 1029 222
rect 954 94 981 127
rect 897 84 909 94
rect 776 72 909 84
rect 969 93 981 94
rect 1015 93 1029 127
rect 969 74 1029 93
rect 1059 210 1140 222
rect 1059 176 1081 210
rect 1115 176 1140 210
rect 1059 120 1140 176
rect 1059 86 1081 120
rect 1115 86 1140 120
rect 1059 74 1140 86
rect 1170 133 1240 222
rect 1170 99 1181 133
rect 1215 99 1240 133
rect 1170 74 1240 99
rect 1270 210 1326 222
rect 1270 176 1281 210
rect 1315 176 1326 210
rect 1270 120 1326 176
rect 1270 86 1281 120
rect 1315 86 1326 120
rect 1270 74 1326 86
rect 1356 210 1413 222
rect 1356 176 1367 210
rect 1401 176 1413 210
rect 1356 120 1413 176
rect 1356 86 1367 120
rect 1401 86 1413 120
rect 1356 74 1413 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 509 86 546
rect 27 475 39 509
rect 73 475 86 509
rect 27 438 86 475
rect 27 404 39 438
rect 73 404 86 438
rect 27 392 86 404
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 508 176 546
rect 116 474 129 508
rect 163 474 176 508
rect 116 392 176 474
rect 206 578 266 592
rect 206 544 219 578
rect 253 544 266 578
rect 206 392 266 544
rect 296 580 366 592
rect 296 546 319 580
rect 353 546 366 580
rect 296 508 366 546
rect 296 474 319 508
rect 353 474 366 508
rect 296 392 366 474
rect 396 580 466 592
rect 396 546 419 580
rect 453 546 466 580
rect 396 510 466 546
rect 396 476 419 510
rect 453 476 466 510
rect 396 440 466 476
rect 396 406 419 440
rect 453 406 466 440
rect 396 392 466 406
rect 496 577 566 592
rect 496 543 519 577
rect 553 543 566 577
rect 496 392 566 543
rect 596 438 656 592
rect 596 404 609 438
rect 643 404 656 438
rect 596 392 656 404
rect 686 577 746 592
rect 686 543 699 577
rect 733 543 746 577
rect 686 392 746 543
rect 776 580 835 592
rect 776 546 789 580
rect 823 546 835 580
rect 996 580 1055 592
rect 996 568 1008 580
rect 776 462 835 546
rect 776 428 789 462
rect 823 428 835 462
rect 776 392 835 428
rect 889 556 948 568
rect 889 522 901 556
rect 935 522 948 556
rect 889 485 948 522
rect 889 451 901 485
rect 935 451 948 485
rect 889 414 948 451
rect 889 380 901 414
rect 935 380 948 414
rect 889 368 948 380
rect 978 546 1008 568
rect 1042 546 1055 580
rect 978 497 1055 546
rect 978 463 1008 497
rect 1042 463 1055 497
rect 978 414 1055 463
rect 978 380 1008 414
rect 1042 380 1055 414
rect 978 368 1055 380
rect 1085 580 1145 592
rect 1085 546 1098 580
rect 1132 546 1145 580
rect 1085 497 1145 546
rect 1085 463 1098 497
rect 1132 463 1145 497
rect 1085 414 1145 463
rect 1085 380 1098 414
rect 1132 380 1145 414
rect 1085 368 1145 380
rect 1175 580 1235 592
rect 1175 546 1188 580
rect 1222 546 1235 580
rect 1175 498 1235 546
rect 1175 464 1188 498
rect 1222 464 1235 498
rect 1175 368 1235 464
rect 1265 580 1325 592
rect 1265 546 1278 580
rect 1312 546 1325 580
rect 1265 497 1325 546
rect 1265 463 1278 497
rect 1312 463 1325 497
rect 1265 414 1325 463
rect 1265 380 1278 414
rect 1312 380 1325 414
rect 1265 368 1325 380
rect 1355 580 1413 592
rect 1355 546 1368 580
rect 1402 546 1413 580
rect 1355 498 1413 546
rect 1355 464 1368 498
rect 1402 464 1413 498
rect 1355 368 1413 464
<< ndiffc >>
rect 39 154 73 188
rect 39 86 73 120
rect 139 86 173 120
rect 239 154 273 188
rect 314 154 348 188
rect 390 154 424 188
rect 239 86 273 120
rect 314 86 348 120
rect 390 86 424 120
rect 492 86 526 120
rect 604 176 638 210
rect 604 86 638 120
rect 788 84 822 118
rect 863 84 897 118
rect 981 93 1015 127
rect 1081 176 1115 210
rect 1081 86 1115 120
rect 1181 99 1215 133
rect 1281 176 1315 210
rect 1281 86 1315 120
rect 1367 176 1401 210
rect 1367 86 1401 120
<< pdiffc >>
rect 39 546 73 580
rect 39 475 73 509
rect 39 404 73 438
rect 129 546 163 580
rect 129 474 163 508
rect 219 544 253 578
rect 319 546 353 580
rect 319 474 353 508
rect 419 546 453 580
rect 419 476 453 510
rect 419 406 453 440
rect 519 543 553 577
rect 609 404 643 438
rect 699 543 733 577
rect 789 546 823 580
rect 789 428 823 462
rect 901 522 935 556
rect 901 451 935 485
rect 901 380 935 414
rect 1008 546 1042 580
rect 1008 463 1042 497
rect 1008 380 1042 414
rect 1098 546 1132 580
rect 1098 463 1132 497
rect 1098 380 1132 414
rect 1188 546 1222 580
rect 1188 464 1222 498
rect 1278 546 1312 580
rect 1278 463 1312 497
rect 1278 380 1312 414
rect 1368 546 1402 580
rect 1368 464 1402 498
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 366 592 396 618
rect 466 592 496 618
rect 566 592 596 618
rect 656 592 686 618
rect 746 592 776 618
rect 948 568 978 594
rect 1055 592 1085 618
rect 1145 592 1175 618
rect 1235 592 1265 618
rect 1325 592 1355 618
rect 86 377 116 392
rect 176 377 206 392
rect 266 377 296 392
rect 366 377 396 392
rect 466 377 496 392
rect 566 377 596 392
rect 656 377 686 392
rect 746 377 776 392
rect 83 310 119 377
rect 53 294 119 310
rect 53 260 69 294
rect 103 260 119 294
rect 173 356 209 377
rect 263 356 299 377
rect 173 340 299 356
rect 173 306 217 340
rect 251 306 299 340
rect 363 310 399 377
rect 463 310 499 377
rect 563 360 599 377
rect 653 360 689 377
rect 563 344 701 360
rect 563 310 651 344
rect 685 310 701 344
rect 173 290 299 306
rect 341 294 407 310
rect 53 244 119 260
rect 84 222 114 244
rect 198 222 228 290
rect 341 260 357 294
rect 391 260 407 294
rect 341 244 407 260
rect 449 294 515 310
rect 449 260 465 294
rect 499 260 515 294
rect 449 244 515 260
rect 563 294 701 310
rect 743 302 779 377
rect 948 353 978 368
rect 1055 353 1085 368
rect 1145 353 1175 368
rect 1235 353 1265 368
rect 1325 353 1355 368
rect 945 310 981 353
rect 1052 330 1088 353
rect 1142 330 1178 353
rect 1232 330 1268 353
rect 449 222 479 244
rect 563 222 593 294
rect 665 134 695 294
rect 743 286 839 302
rect 743 252 789 286
rect 823 252 839 286
rect 743 236 839 252
rect 897 294 981 310
rect 897 260 913 294
rect 947 260 981 294
rect 897 244 981 260
rect 1029 327 1268 330
rect 1322 327 1358 353
rect 1029 314 1358 327
rect 1029 280 1045 314
rect 1079 280 1113 314
rect 1147 280 1181 314
rect 1215 294 1358 314
rect 1215 280 1356 294
rect 1029 264 1356 280
rect 924 222 954 244
rect 1029 222 1059 264
rect 1140 222 1170 264
rect 1240 222 1270 264
rect 1326 222 1356 264
rect 665 118 754 134
rect 665 84 704 118
rect 738 84 754 118
rect 84 48 114 74
rect 198 48 228 74
rect 449 48 479 74
rect 563 48 593 74
rect 665 68 754 84
rect 924 68 954 94
rect 1029 48 1059 74
rect 1140 48 1170 74
rect 1240 48 1270 74
rect 1326 48 1356 74
<< polycont >>
rect 69 260 103 294
rect 217 306 251 340
rect 651 310 685 344
rect 357 260 391 294
rect 465 260 499 294
rect 789 252 823 286
rect 913 260 947 294
rect 1045 280 1079 314
rect 1113 280 1147 314
rect 1181 280 1215 314
rect 704 84 738 118
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 509 89 546
rect 23 475 39 509
rect 73 475 89 509
rect 23 438 89 475
rect 129 580 163 596
rect 129 508 163 546
rect 203 578 269 649
rect 203 544 219 578
rect 253 544 269 578
rect 203 526 269 544
rect 303 580 369 596
rect 303 546 319 580
rect 353 546 369 580
rect 303 508 369 546
rect 303 492 319 508
rect 163 474 319 492
rect 353 474 369 508
rect 129 458 369 474
rect 403 580 469 596
rect 403 546 419 580
rect 453 546 469 580
rect 403 510 469 546
rect 503 577 749 596
rect 503 543 519 577
rect 553 543 699 577
rect 733 543 749 577
rect 503 540 749 543
rect 789 580 839 596
rect 823 546 839 580
rect 992 580 1042 649
rect 403 476 419 510
rect 453 506 469 510
rect 789 506 839 546
rect 453 476 839 506
rect 403 472 839 476
rect 23 404 39 438
rect 73 424 89 438
rect 403 440 469 472
rect 403 424 419 440
rect 73 406 419 424
rect 453 406 469 440
rect 789 462 839 472
rect 73 404 469 406
rect 23 390 469 404
rect 579 404 609 438
rect 643 404 659 438
rect 823 428 839 462
rect 789 412 839 428
rect 885 556 951 572
rect 885 522 901 556
rect 935 522 951 556
rect 885 485 951 522
rect 885 451 901 485
rect 935 451 951 485
rect 885 414 951 451
rect 23 388 89 390
rect 201 340 267 356
rect 25 294 167 310
rect 25 260 69 294
rect 103 260 167 294
rect 201 306 217 340
rect 251 306 267 340
rect 201 290 267 306
rect 341 294 407 310
rect 25 256 167 260
rect 341 260 357 294
rect 391 260 407 294
rect 341 256 407 260
rect 25 222 407 256
rect 449 294 545 356
rect 449 260 465 294
rect 499 276 545 294
rect 499 260 511 276
rect 449 242 511 260
rect 449 236 545 242
rect 579 226 613 404
rect 885 380 901 414
rect 935 380 951 414
rect 885 378 951 380
rect 693 360 951 378
rect 992 546 1008 580
rect 992 497 1042 546
rect 992 463 1008 497
rect 992 414 1042 463
rect 992 380 1008 414
rect 992 364 1042 380
rect 1082 580 1138 596
rect 1082 546 1098 580
rect 1132 546 1138 580
rect 1082 497 1138 546
rect 1082 463 1098 497
rect 1132 463 1138 497
rect 1172 580 1238 649
rect 1172 546 1188 580
rect 1222 546 1238 580
rect 1172 498 1238 546
rect 1172 464 1188 498
rect 1222 464 1238 498
rect 1272 580 1318 596
rect 1272 546 1278 580
rect 1312 546 1318 580
rect 1272 497 1318 546
rect 1082 430 1138 463
rect 1272 463 1278 497
rect 1312 463 1318 497
rect 1352 580 1418 649
rect 1352 546 1368 580
rect 1402 546 1418 580
rect 1352 498 1418 546
rect 1352 464 1368 498
rect 1402 464 1418 498
rect 1272 430 1318 463
rect 1082 414 1415 430
rect 1082 380 1098 414
rect 1132 380 1278 414
rect 1312 380 1415 414
rect 1082 364 1415 380
rect 647 344 951 360
rect 647 310 651 344
rect 685 310 727 344
rect 997 314 1231 330
rect 647 294 727 310
rect 773 286 839 302
rect 773 252 789 286
rect 823 276 839 286
rect 773 242 799 252
rect 833 242 839 276
rect 773 236 839 242
rect 889 294 963 310
rect 889 260 913 294
rect 947 260 963 294
rect 889 236 963 260
rect 997 280 1045 314
rect 1079 280 1113 314
rect 1147 280 1181 314
rect 1215 280 1231 314
rect 1273 294 1331 364
rect 997 264 1231 280
rect 579 210 654 226
rect 579 188 604 210
rect 23 154 39 188
rect 73 154 239 188
rect 273 154 314 188
rect 348 154 390 188
rect 424 176 604 188
rect 638 202 654 210
rect 997 202 1031 264
rect 1265 260 1331 294
rect 1265 230 1315 260
rect 638 176 1031 202
rect 424 168 1031 176
rect 1065 210 1315 230
rect 1065 176 1081 210
rect 1115 196 1281 210
rect 1115 176 1131 196
rect 424 154 654 168
rect 23 120 89 154
rect 223 120 440 154
rect 579 120 654 154
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 86 139 120
rect 173 86 189 120
rect 123 17 189 86
rect 223 86 239 120
rect 273 86 314 120
rect 348 86 390 120
rect 424 86 440 120
rect 223 70 440 86
rect 474 86 492 120
rect 526 86 545 120
rect 474 17 545 86
rect 579 86 604 120
rect 638 86 654 120
rect 579 70 654 86
rect 688 118 913 134
rect 688 84 704 118
rect 738 84 788 118
rect 822 84 863 118
rect 897 84 913 118
rect 688 68 913 84
rect 965 127 1031 134
rect 965 93 981 127
rect 1015 93 1031 127
rect 965 17 1031 93
rect 1065 120 1131 176
rect 1265 176 1281 196
rect 1065 86 1081 120
rect 1115 86 1131 120
rect 1065 70 1131 86
rect 1165 133 1231 162
rect 1165 99 1181 133
rect 1215 99 1231 133
rect 1165 17 1231 99
rect 1265 120 1315 176
rect 1265 86 1281 120
rect 1265 70 1315 86
rect 1351 210 1417 226
rect 1351 176 1367 210
rect 1401 176 1417 210
rect 1351 120 1417 176
rect 1351 86 1367 120
rect 1401 86 1417 120
rect 1351 17 1417 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 511 242 545 276
rect 799 252 823 276
rect 823 252 833 276
rect 799 242 833 252
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 499 276 557 282
rect 499 242 511 276
rect 545 273 557 276
rect 787 276 845 282
rect 787 273 799 276
rect 545 245 799 273
rect 545 242 557 245
rect 499 236 557 242
rect 787 242 799 245
rect 833 242 845 276
rect 787 236 845 242
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or4b_4
flabel comment s 680 282 680 282 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 511 242 545 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 1375 390 1409 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 1833084
string GDS_START 1820704
<< end >>
