magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4946 1975
<< nwell >>
rect -38 331 3686 704
rect 1498 275 1695 331
<< pwell >>
rect 3196 242 3645 247
rect 189 221 1051 226
rect 189 201 1651 221
rect 189 161 1974 201
rect 2567 161 2677 195
rect 189 158 2677 161
rect 2930 158 3645 242
rect 189 49 3645 158
rect 0 0 3648 49
<< scnmos >>
rect 319 116 349 200
rect 397 116 427 200
rect 560 116 590 200
rect 662 116 692 200
rect 817 116 847 200
rect 895 116 925 200
rect 1271 67 1301 195
rect 1343 67 1373 195
rect 1466 111 1496 195
rect 1538 111 1568 195
rect 1861 47 1891 175
rect 1970 51 2000 135
rect 2102 51 2132 135
rect 2463 51 2493 135
rect 2541 51 2571 135
rect 2795 48 2825 132
rect 2873 48 2903 132
rect 3006 48 3036 216
rect 3078 48 3108 216
rect 3279 137 3309 221
rect 3351 137 3381 221
rect 3460 53 3490 221
rect 3532 53 3562 221
<< scpmoshvt >>
rect 81 457 111 541
rect 167 457 197 541
rect 239 457 269 541
rect 346 494 376 578
rect 592 411 622 495
rect 678 411 708 495
rect 893 457 923 541
rect 1007 457 1037 541
rect 1079 457 1109 541
rect 1271 373 1301 541
rect 1343 373 1373 541
rect 1450 413 1480 541
rect 1522 413 1552 541
rect 1769 379 1799 463
rect 1876 379 1906 547
rect 2102 535 2132 619
rect 2608 510 2638 594
rect 2289 397 2319 481
rect 2421 397 2451 481
rect 2493 397 2523 481
rect 2801 367 2831 495
rect 2873 367 2903 495
rect 3006 367 3036 619
rect 3078 367 3108 619
rect 3279 367 3309 495
rect 3351 367 3381 495
rect 3460 367 3490 619
rect 3532 367 3562 619
<< ndiff >>
rect 215 172 319 200
rect 215 138 227 172
rect 261 138 319 172
rect 215 116 319 138
rect 349 116 397 200
rect 427 175 560 200
rect 427 141 515 175
rect 549 141 560 175
rect 427 116 560 141
rect 590 175 662 200
rect 590 141 617 175
rect 651 141 662 175
rect 590 116 662 141
rect 692 116 817 200
rect 847 116 895 200
rect 925 116 1025 200
rect 940 98 1025 116
rect 940 64 959 98
rect 993 64 1025 98
rect 1214 170 1271 195
rect 1214 136 1226 170
rect 1260 136 1271 170
rect 1214 67 1271 136
rect 1301 67 1343 195
rect 1373 183 1466 195
rect 1373 149 1398 183
rect 1432 149 1466 183
rect 1373 113 1466 149
rect 1373 79 1398 113
rect 1432 111 1466 113
rect 1496 111 1538 195
rect 1568 170 1625 195
rect 1568 136 1579 170
rect 1613 136 1625 170
rect 1568 111 1625 136
rect 1788 133 1861 175
rect 1432 79 1444 111
rect 1788 99 1800 133
rect 1834 99 1861 133
rect 1373 67 1444 79
rect 940 52 1025 64
rect 1788 47 1861 99
rect 1891 135 1948 175
rect 2593 157 2651 169
rect 2593 135 2605 157
rect 1891 133 1970 135
rect 1891 99 1902 133
rect 1936 99 1970 133
rect 1891 51 1970 99
rect 2000 51 2102 135
rect 2132 97 2463 135
rect 2132 63 2143 97
rect 2177 63 2463 97
rect 2132 51 2463 63
rect 2493 51 2541 135
rect 2571 123 2605 135
rect 2639 123 2651 157
rect 2956 132 3006 216
rect 2571 51 2651 123
rect 2738 111 2795 132
rect 2738 77 2750 111
rect 2784 77 2795 111
rect 1891 47 1948 51
rect 2738 48 2795 77
rect 2825 48 2873 132
rect 2903 94 3006 132
rect 2903 60 2914 94
rect 2948 60 3006 94
rect 2903 48 3006 60
rect 3036 48 3078 216
rect 3108 204 3165 216
rect 3108 170 3119 204
rect 3153 170 3165 204
rect 3108 103 3165 170
rect 3222 196 3279 221
rect 3222 162 3234 196
rect 3268 162 3279 196
rect 3222 137 3279 162
rect 3309 137 3351 221
rect 3381 209 3460 221
rect 3381 175 3415 209
rect 3449 175 3460 209
rect 3381 137 3460 175
rect 3108 69 3119 103
rect 3153 69 3165 103
rect 3108 48 3165 69
rect 3403 99 3460 137
rect 3403 65 3415 99
rect 3449 65 3460 99
rect 3403 53 3460 65
rect 3490 53 3532 221
rect 3562 209 3619 221
rect 3562 175 3573 209
rect 3607 175 3619 209
rect 3562 103 3619 175
rect 3562 69 3573 103
rect 3607 69 3619 103
rect 3562 53 3619 69
<< pdiff >>
rect 291 566 346 578
rect 291 541 301 566
rect 27 516 81 541
rect 27 482 36 516
rect 70 482 81 516
rect 27 457 81 482
rect 111 515 167 541
rect 111 481 122 515
rect 156 481 167 515
rect 111 457 167 481
rect 197 457 239 541
rect 269 532 301 541
rect 335 532 346 566
rect 269 494 346 532
rect 376 553 430 578
rect 376 519 387 553
rect 421 519 430 553
rect 376 494 430 519
rect 484 512 543 524
rect 269 457 319 494
rect 484 478 493 512
rect 527 495 543 512
rect 817 582 871 594
rect 817 548 827 582
rect 861 548 871 582
rect 938 582 992 594
rect 817 541 871 548
rect 938 548 948 582
rect 982 548 992 582
rect 938 541 992 548
rect 2045 589 2102 619
rect 2045 555 2057 589
rect 2091 555 2102 589
rect 527 478 592 495
rect 484 411 592 478
rect 622 457 678 495
rect 622 423 633 457
rect 667 423 678 457
rect 622 411 678 423
rect 708 470 763 495
rect 708 436 719 470
rect 753 436 763 470
rect 817 457 893 541
rect 923 457 1007 541
rect 1037 457 1079 541
rect 1109 520 1163 541
rect 1109 486 1120 520
rect 1154 486 1163 520
rect 1109 457 1163 486
rect 1217 529 1271 541
rect 1217 495 1226 529
rect 1260 495 1271 529
rect 708 411 763 436
rect 1217 419 1271 495
rect 1217 385 1226 419
rect 1260 385 1271 419
rect 1217 373 1271 385
rect 1301 373 1343 541
rect 1373 529 1450 541
rect 1373 495 1384 529
rect 1418 495 1450 529
rect 1373 413 1450 495
rect 1480 413 1522 541
rect 1552 413 1630 541
rect 1821 527 1876 547
rect 1821 493 1831 527
rect 1865 493 1876 527
rect 1821 463 1876 493
rect 1373 373 1428 413
rect 1574 357 1630 413
rect 1712 438 1769 463
rect 1712 404 1724 438
rect 1758 404 1769 438
rect 1712 379 1769 404
rect 1799 379 1876 463
rect 1906 425 1963 547
rect 2045 535 2102 555
rect 2132 594 2189 619
rect 2947 607 3006 619
rect 2132 560 2143 594
rect 2177 560 2189 594
rect 2132 535 2189 560
rect 2545 582 2608 594
rect 2545 548 2563 582
rect 2597 548 2608 582
rect 1906 391 1917 425
rect 1951 391 1963 425
rect 1906 379 1963 391
rect 1574 323 1584 357
rect 1618 323 1630 357
rect 1574 311 1630 323
rect 2545 510 2608 548
rect 2638 569 2692 594
rect 2638 535 2649 569
rect 2683 535 2692 569
rect 2638 510 2692 535
rect 2947 573 2959 607
rect 2993 573 3006 607
rect 2545 481 2593 510
rect 2185 456 2289 481
rect 2185 422 2197 456
rect 2231 422 2289 456
rect 2185 397 2289 422
rect 2319 450 2421 481
rect 2319 416 2353 450
rect 2387 416 2421 450
rect 2319 397 2421 416
rect 2451 397 2493 481
rect 2523 445 2593 481
rect 2523 397 2575 445
rect 2947 508 3006 573
rect 2947 495 2959 508
rect 2746 460 2801 495
rect 2746 426 2756 460
rect 2790 426 2801 460
rect 2746 367 2801 426
rect 2831 367 2873 495
rect 2903 474 2959 495
rect 2993 474 3006 508
rect 2903 367 3006 474
rect 3036 367 3078 619
rect 3108 597 3165 619
rect 3108 563 3119 597
rect 3153 563 3165 597
rect 3108 505 3165 563
rect 3403 607 3460 619
rect 3403 573 3415 607
rect 3449 573 3460 607
rect 3108 471 3119 505
rect 3153 471 3165 505
rect 3403 510 3460 573
rect 3403 495 3415 510
rect 3108 413 3165 471
rect 3108 379 3119 413
rect 3153 379 3165 413
rect 3108 367 3165 379
rect 3222 483 3279 495
rect 3222 449 3234 483
rect 3268 449 3279 483
rect 3222 413 3279 449
rect 3222 379 3234 413
rect 3268 379 3279 413
rect 3222 367 3279 379
rect 3309 367 3351 495
rect 3381 476 3415 495
rect 3449 476 3460 510
rect 3381 413 3460 476
rect 3381 379 3415 413
rect 3449 379 3460 413
rect 3381 367 3460 379
rect 3490 367 3532 619
rect 3562 597 3619 619
rect 3562 563 3573 597
rect 3607 563 3619 597
rect 3562 505 3619 563
rect 3562 471 3573 505
rect 3607 471 3619 505
rect 3562 413 3619 471
rect 3562 379 3573 413
rect 3607 379 3619 413
rect 3562 367 3619 379
<< ndiffc >>
rect 227 138 261 172
rect 515 141 549 175
rect 617 141 651 175
rect 959 64 993 98
rect 1226 136 1260 170
rect 1398 149 1432 183
rect 1398 79 1432 113
rect 1579 136 1613 170
rect 1800 99 1834 133
rect 1902 99 1936 133
rect 2143 63 2177 97
rect 2605 123 2639 157
rect 2750 77 2784 111
rect 2914 60 2948 94
rect 3119 170 3153 204
rect 3234 162 3268 196
rect 3415 175 3449 209
rect 3119 69 3153 103
rect 3415 65 3449 99
rect 3573 175 3607 209
rect 3573 69 3607 103
<< pdiffc >>
rect 36 482 70 516
rect 122 481 156 515
rect 301 532 335 566
rect 387 519 421 553
rect 493 478 527 512
rect 827 548 861 582
rect 948 548 982 582
rect 2057 555 2091 589
rect 633 423 667 457
rect 719 436 753 470
rect 1120 486 1154 520
rect 1226 495 1260 529
rect 1226 385 1260 419
rect 1384 495 1418 529
rect 1831 493 1865 527
rect 1724 404 1758 438
rect 2143 560 2177 594
rect 2563 548 2597 582
rect 1917 391 1951 425
rect 1584 323 1618 357
rect 2649 535 2683 569
rect 2959 573 2993 607
rect 2197 422 2231 456
rect 2353 416 2387 450
rect 2756 426 2790 460
rect 2959 474 2993 508
rect 3119 563 3153 597
rect 3415 573 3449 607
rect 3119 471 3153 505
rect 3119 379 3153 413
rect 3234 449 3268 483
rect 3234 379 3268 413
rect 3415 476 3449 510
rect 3415 379 3449 413
rect 3573 563 3607 597
rect 3573 471 3607 505
rect 3573 379 3607 413
<< poly >>
rect 81 615 376 645
rect 81 541 111 615
rect 346 578 376 615
rect 592 615 1480 645
rect 2102 619 2132 645
rect 167 541 197 567
rect 239 541 269 567
rect 81 431 111 457
rect 167 356 197 457
rect 239 356 269 457
rect 167 340 269 356
rect 167 306 213 340
rect 247 306 269 340
rect 167 272 269 306
rect 346 324 376 494
rect 592 495 622 615
rect 1450 599 1480 615
rect 893 541 923 567
rect 1450 569 1906 599
rect 1007 541 1037 567
rect 1079 541 1109 567
rect 1271 541 1301 567
rect 1343 541 1373 567
rect 1450 541 1480 569
rect 1522 541 1552 569
rect 1876 547 1906 569
rect 678 495 708 521
rect 893 425 923 457
rect 1007 432 1037 457
rect 1079 432 1109 457
rect 592 389 622 411
rect 560 359 622 389
rect 346 294 463 324
rect 167 238 213 272
rect 247 252 269 272
rect 397 276 463 294
rect 247 238 349 252
rect 167 222 349 238
rect 319 200 349 222
rect 397 242 413 276
rect 447 242 463 276
rect 397 215 463 242
rect 397 200 427 215
rect 560 200 590 359
rect 678 292 708 411
rect 875 409 941 425
rect 875 375 891 409
rect 925 375 941 409
rect 1007 402 1109 432
rect 875 341 941 375
rect 875 321 891 341
rect 817 307 891 321
rect 925 307 941 341
rect 662 276 769 292
rect 662 242 719 276
rect 753 242 769 276
rect 662 215 769 242
rect 817 291 941 307
rect 989 340 1055 402
rect 1769 463 1799 489
rect 989 306 1005 340
rect 1039 306 1055 340
rect 662 200 692 215
rect 817 200 847 291
rect 989 290 1055 306
rect 1108 338 1174 354
rect 1108 304 1124 338
rect 1158 304 1174 338
rect 989 245 1019 290
rect 895 215 1019 245
rect 1108 270 1174 304
rect 1108 236 1124 270
rect 1158 250 1174 270
rect 1271 250 1301 373
rect 1343 250 1373 373
rect 1450 296 1480 413
rect 1522 296 1552 413
rect 2608 594 2638 620
rect 3006 619 3036 645
rect 3078 619 3108 645
rect 3460 619 3490 645
rect 3532 619 3562 645
rect 1450 266 1568 296
rect 1769 269 1799 379
rect 1876 305 1906 379
rect 1876 275 2054 305
rect 1158 236 1373 250
rect 1108 220 1373 236
rect 895 200 925 215
rect 1271 195 1301 220
rect 1343 195 1373 220
rect 1466 195 1496 266
rect 1538 195 1568 266
rect 1682 253 1799 269
rect 1682 219 1698 253
rect 1732 227 1799 253
rect 1970 253 2054 275
rect 1732 219 1891 227
rect 1682 197 1891 219
rect 319 48 349 116
rect 397 90 427 116
rect 560 90 590 116
rect 662 90 692 116
rect 817 90 847 116
rect 895 48 925 116
rect 1682 185 1748 197
rect 1682 151 1698 185
rect 1732 151 1748 185
rect 1861 175 1891 197
rect 1970 219 2004 253
rect 2038 219 2054 253
rect 1970 203 2054 219
rect 2102 269 2132 535
rect 2289 481 2319 507
rect 2421 481 2451 507
rect 2493 481 2523 507
rect 2289 339 2319 397
rect 2243 323 2319 339
rect 2243 289 2259 323
rect 2293 289 2319 323
rect 2243 273 2319 289
rect 2421 356 2451 397
rect 2493 356 2523 397
rect 2421 340 2523 356
rect 2421 306 2441 340
rect 2475 326 2523 340
rect 2608 384 2638 510
rect 2801 495 2831 521
rect 2873 495 2903 521
rect 2608 368 2674 384
rect 2608 334 2624 368
rect 2658 334 2674 368
rect 3279 495 3309 521
rect 3351 495 3381 521
rect 2475 306 2493 326
rect 2421 272 2493 306
rect 2102 253 2168 269
rect 2102 219 2118 253
rect 2152 219 2168 253
rect 2421 238 2441 272
rect 2475 238 2493 272
rect 2421 222 2493 238
rect 2102 203 2168 219
rect 1682 135 1748 151
rect 1466 85 1496 111
rect 1538 85 1568 111
rect 319 18 925 48
rect 1271 41 1301 67
rect 1343 41 1373 67
rect 1970 135 2000 203
rect 2102 135 2132 203
rect 2463 135 2493 222
rect 2608 318 2674 334
rect 2608 214 2638 318
rect 2801 282 2831 367
rect 2765 266 2831 282
rect 2765 232 2781 266
rect 2815 246 2831 266
rect 2873 246 2903 367
rect 3006 335 3036 367
rect 2945 319 3036 335
rect 2945 285 2961 319
rect 2995 299 3036 319
rect 3078 299 3108 367
rect 3279 299 3309 367
rect 3351 299 3381 367
rect 3460 327 3490 367
rect 3532 327 3562 367
rect 2995 285 3381 299
rect 2945 269 3381 285
rect 2815 232 2903 246
rect 2765 216 2903 232
rect 3006 216 3036 269
rect 3078 216 3108 269
rect 3279 221 3309 269
rect 3351 221 3381 269
rect 3455 311 3562 327
rect 3455 277 3471 311
rect 3505 277 3562 311
rect 3455 261 3562 277
rect 3460 221 3490 261
rect 3532 221 3562 261
rect 2541 184 2638 214
rect 2541 135 2571 184
rect 2795 132 2825 216
rect 2873 132 2903 216
rect 1861 21 1891 47
rect 1970 25 2000 51
rect 2102 25 2132 51
rect 2463 25 2493 51
rect 2541 25 2571 51
rect 3279 111 3309 137
rect 3351 111 3381 137
rect 2795 22 2825 48
rect 2873 22 2903 48
rect 3006 22 3036 48
rect 3078 22 3108 48
rect 3460 27 3490 53
rect 3532 27 3562 53
<< polycont >>
rect 213 306 247 340
rect 213 238 247 272
rect 413 242 447 276
rect 891 375 925 409
rect 891 307 925 341
rect 719 242 753 276
rect 1005 306 1039 340
rect 1124 304 1158 338
rect 1124 236 1158 270
rect 1698 219 1732 253
rect 1698 151 1732 185
rect 2004 219 2038 253
rect 2259 289 2293 323
rect 2441 306 2475 340
rect 2624 334 2658 368
rect 2118 219 2152 253
rect 2441 238 2475 272
rect 2781 232 2815 266
rect 2961 285 2995 319
rect 3471 277 3505 311
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3648 683
rect 20 579 242 613
rect 20 516 70 579
rect 20 482 36 516
rect 20 453 70 482
rect 106 515 172 543
rect 106 481 122 515
rect 156 481 172 515
rect 106 426 172 481
rect 208 496 242 579
rect 285 566 351 649
rect 477 582 877 613
rect 285 532 301 566
rect 335 532 351 566
rect 387 553 437 582
rect 421 519 437 553
rect 387 496 437 519
rect 208 462 437 496
rect 477 579 827 582
rect 477 512 527 579
rect 811 548 827 579
rect 861 548 877 582
rect 477 478 493 512
rect 477 462 527 478
rect 563 509 769 543
rect 811 532 877 548
rect 932 582 998 649
rect 932 548 948 582
rect 982 548 998 582
rect 932 532 998 548
rect 563 426 597 509
rect 106 392 597 426
rect 633 457 667 473
rect 197 350 263 356
rect 197 340 223 350
rect 197 306 213 340
rect 257 316 263 350
rect 247 306 263 316
rect 197 272 263 306
rect 197 238 213 272
rect 247 238 263 272
rect 197 222 263 238
rect 313 276 463 292
rect 313 242 413 276
rect 447 242 463 276
rect 211 172 263 188
rect 211 138 227 172
rect 261 140 263 172
rect 261 138 277 140
rect 211 17 277 138
rect 313 88 463 242
rect 499 175 565 392
rect 633 371 667 423
rect 703 470 769 509
rect 1104 520 1170 545
rect 1104 496 1120 520
rect 703 436 719 470
rect 753 436 769 470
rect 703 407 769 436
rect 805 486 1120 496
rect 1154 486 1170 520
rect 805 462 1170 486
rect 1210 529 1276 545
rect 1210 495 1226 529
rect 1260 495 1276 529
rect 805 371 839 462
rect 1210 443 1276 495
rect 1368 529 1434 649
rect 1368 495 1384 529
rect 1418 495 1434 529
rect 1368 479 1434 495
rect 1724 589 2091 613
rect 1724 579 2057 589
rect 1210 426 1688 443
rect 633 337 839 371
rect 633 200 667 337
rect 499 141 515 175
rect 549 141 565 175
rect 499 116 565 141
rect 601 175 667 200
rect 601 141 617 175
rect 651 141 667 175
rect 703 276 769 292
rect 703 242 719 276
rect 753 242 769 276
rect 703 184 769 242
rect 805 254 839 337
rect 875 419 1688 426
rect 875 409 1226 419
rect 875 375 891 409
rect 925 392 1226 409
rect 925 375 941 392
rect 875 341 941 375
rect 1210 385 1226 392
rect 1260 409 1688 419
rect 1260 385 1276 409
rect 875 307 891 341
rect 925 307 941 341
rect 875 291 941 307
rect 985 350 1055 356
rect 985 316 991 350
rect 1025 340 1055 350
rect 985 306 1005 316
rect 1039 306 1055 340
rect 985 290 1055 306
rect 1108 338 1174 354
rect 1108 304 1124 338
rect 1158 304 1174 338
rect 1108 270 1174 304
rect 1108 254 1124 270
rect 805 236 1124 254
rect 1158 236 1174 270
rect 805 220 1174 236
rect 703 150 1079 184
rect 601 116 667 141
rect 943 98 1009 114
rect 943 64 959 98
rect 993 64 1009 98
rect 943 17 1009 64
rect 1045 87 1079 150
rect 1210 170 1276 385
rect 1563 357 1618 373
rect 1563 323 1584 357
rect 1563 269 1618 323
rect 1654 339 1688 409
rect 1724 438 1774 579
rect 1815 527 2021 543
rect 2057 531 2091 555
rect 2127 594 2177 649
rect 2127 560 2143 594
rect 2127 531 2177 560
rect 2213 579 2527 613
rect 1815 493 1831 527
rect 1865 493 2021 527
rect 1815 477 2021 493
rect 2213 485 2247 579
rect 1758 404 1774 438
rect 1724 375 1774 404
rect 1816 425 1951 441
rect 1816 391 1917 425
rect 1816 375 1951 391
rect 1816 339 1850 375
rect 1987 339 2021 477
rect 2181 456 2247 485
rect 2181 422 2197 456
rect 2231 422 2247 456
rect 2181 393 2247 422
rect 2283 509 2457 543
rect 2283 339 2317 509
rect 1654 305 1850 339
rect 1210 136 1226 170
rect 1260 136 1276 170
rect 1210 123 1276 136
rect 1312 253 1748 269
rect 1312 235 1698 253
rect 1312 87 1346 235
rect 1045 53 1346 87
rect 1382 183 1448 199
rect 1382 149 1398 183
rect 1432 149 1448 183
rect 1382 113 1448 149
rect 1382 79 1398 113
rect 1432 79 1448 113
rect 1563 170 1629 235
rect 1563 136 1579 170
rect 1613 136 1629 170
rect 1563 107 1629 136
rect 1682 219 1698 235
rect 1732 219 1748 253
rect 1682 185 1748 219
rect 1682 151 1698 185
rect 1732 151 1748 185
rect 1682 135 1748 151
rect 1784 133 1850 305
rect 1382 17 1448 79
rect 1784 99 1800 133
rect 1834 99 1850 133
rect 1784 53 1850 99
rect 1886 323 2317 339
rect 1886 305 2259 323
rect 1886 133 1952 305
rect 2243 289 2259 305
rect 2293 289 2317 323
rect 2243 273 2317 289
rect 2353 450 2387 473
rect 1988 253 2054 269
rect 1988 219 2004 253
rect 2038 219 2054 253
rect 1988 167 2054 219
rect 2102 253 2168 269
rect 2102 219 2118 253
rect 2152 237 2168 253
rect 2353 237 2387 416
rect 2423 426 2457 509
rect 2493 496 2527 579
rect 2563 582 2597 649
rect 2943 607 3009 649
rect 2563 532 2597 548
rect 2633 569 2699 598
rect 2633 535 2649 569
rect 2683 535 2699 569
rect 2633 496 2699 535
rect 2943 573 2959 607
rect 2993 573 3009 607
rect 2943 508 3009 573
rect 2493 462 2699 496
rect 2740 460 2806 499
rect 2740 426 2756 460
rect 2790 426 2806 460
rect 2943 474 2959 508
rect 2993 474 3009 508
rect 2943 458 3009 474
rect 3103 597 3169 613
rect 3103 563 3119 597
rect 3153 563 3169 597
rect 3103 505 3169 563
rect 3103 471 3119 505
rect 3153 471 3169 505
rect 3399 607 3465 649
rect 3399 573 3415 607
rect 3449 573 3465 607
rect 3399 510 3465 573
rect 2423 392 2674 426
rect 2608 368 2674 392
rect 2740 422 2806 426
rect 2740 388 3067 422
rect 2152 219 2387 237
rect 2425 350 2491 356
rect 2425 316 2431 350
rect 2465 340 2491 350
rect 2425 306 2441 316
rect 2475 306 2491 340
rect 2608 334 2624 368
rect 2658 352 2674 368
rect 2658 334 2997 352
rect 2608 319 2997 334
rect 2608 318 2961 319
rect 2425 272 2491 306
rect 2945 285 2961 318
rect 2995 285 2997 319
rect 2425 238 2441 272
rect 2475 238 2491 272
rect 2425 222 2491 238
rect 2713 266 2855 282
rect 2945 269 2997 285
rect 2713 232 2781 266
rect 2815 232 2855 266
rect 2102 203 2387 219
rect 2713 216 2855 232
rect 2353 173 2387 203
rect 3033 180 3067 388
rect 1988 133 2263 167
rect 1886 99 1902 133
rect 1936 99 1952 133
rect 1886 53 1952 99
rect 2127 63 2143 97
rect 2177 63 2193 97
rect 2127 17 2193 63
rect 2229 87 2263 133
rect 2353 157 2655 173
rect 2353 123 2605 157
rect 2639 123 2655 157
rect 2734 146 3067 180
rect 3103 413 3169 471
rect 3103 379 3119 413
rect 3153 379 3169 413
rect 3103 204 3169 379
rect 3103 170 3119 204
rect 3153 170 3169 204
rect 2734 111 2800 146
rect 2734 87 2750 111
rect 2229 77 2750 87
rect 2784 77 2800 111
rect 2229 53 2800 77
rect 2898 94 2964 110
rect 2898 60 2914 94
rect 2948 60 2964 94
rect 2898 17 2964 60
rect 3103 103 3169 170
rect 3218 483 3284 499
rect 3218 449 3234 483
rect 3268 449 3284 483
rect 3218 413 3284 449
rect 3218 379 3234 413
rect 3268 379 3284 413
rect 3218 327 3284 379
rect 3399 476 3415 510
rect 3449 476 3465 510
rect 3399 413 3465 476
rect 3399 379 3415 413
rect 3449 379 3465 413
rect 3399 363 3465 379
rect 3557 597 3623 613
rect 3557 563 3573 597
rect 3607 563 3623 597
rect 3557 505 3623 563
rect 3557 471 3573 505
rect 3607 471 3623 505
rect 3557 413 3623 471
rect 3557 379 3573 413
rect 3607 379 3623 413
rect 3218 311 3521 327
rect 3218 277 3471 311
rect 3505 277 3521 311
rect 3218 261 3521 277
rect 3218 196 3284 261
rect 3218 162 3234 196
rect 3268 162 3284 196
rect 3218 133 3284 162
rect 3399 209 3465 225
rect 3399 175 3415 209
rect 3449 175 3465 209
rect 3103 69 3119 103
rect 3153 69 3169 103
rect 3103 53 3169 69
rect 3399 99 3465 175
rect 3399 65 3415 99
rect 3449 65 3465 99
rect 3399 17 3465 65
rect 3557 209 3623 379
rect 3557 175 3573 209
rect 3607 175 3623 209
rect 3557 103 3623 175
rect 3557 69 3573 103
rect 3607 69 3623 103
rect 3557 53 3623 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3648 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 3583 649 3617 683
rect 223 340 257 350
rect 223 316 247 340
rect 247 316 257 340
rect 991 340 1025 350
rect 991 316 1005 340
rect 1005 316 1025 340
rect 2431 340 2465 350
rect 2431 316 2441 340
rect 2441 316 2465 340
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
<< metal1 >>
rect 0 683 3648 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3648 683
rect 0 617 3648 649
rect 211 350 269 356
rect 211 316 223 350
rect 257 347 269 350
rect 979 350 1037 356
rect 979 347 991 350
rect 257 319 991 347
rect 257 316 269 319
rect 211 310 269 316
rect 979 316 991 319
rect 1025 347 1037 350
rect 2419 350 2477 356
rect 2419 347 2431 350
rect 1025 319 2431 347
rect 1025 316 1037 319
rect 979 310 1037 316
rect 2419 316 2431 319
rect 2465 316 2477 350
rect 2419 310 2477 316
rect 0 17 3648 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3648 17
rect 0 -49 3648 -17
<< labels >>
flabel pwell s 0 0 3648 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 3648 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfrbp_lp
flabel metal1 s 2431 316 2465 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 3648 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 3648 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 2719 242 2753 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2815 242 2849 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 3583 94 3617 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3583 168 3617 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3583 242 3617 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3583 316 3617 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3583 390 3617 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3583 464 3617 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3583 538 3617 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3103 94 3137 128 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3103 168 3137 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3103 242 3137 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3103 316 3137 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3103 390 3137 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3103 464 3137 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3103 538 3137 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3648 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry R90
string GDS_END 4569760
string GDS_START 4547784
<< end >>
