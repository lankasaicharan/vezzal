magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 106 162 623 278
rect 1 49 728 162
rect 0 0 768 49
<< scnmos >>
rect 80 52 110 136
rect 232 52 282 252
rect 447 52 497 252
rect 619 52 649 136
<< scpmoshvt >>
rect 80 367 110 619
rect 232 419 282 619
rect 447 419 497 619
rect 619 367 649 619
<< ndiff >>
rect 132 136 232 252
rect 27 111 80 136
rect 27 77 35 111
rect 69 77 80 111
rect 27 52 80 77
rect 110 111 232 136
rect 110 77 132 111
rect 166 77 232 111
rect 110 52 232 77
rect 282 240 335 252
rect 282 206 293 240
rect 327 206 335 240
rect 282 172 335 206
rect 282 138 293 172
rect 327 138 335 172
rect 282 104 335 138
rect 282 70 293 104
rect 327 70 335 104
rect 282 52 335 70
rect 394 227 447 252
rect 394 193 402 227
rect 436 193 447 227
rect 394 104 447 193
rect 394 70 402 104
rect 436 70 447 104
rect 394 52 447 70
rect 497 136 597 252
rect 497 118 619 136
rect 497 84 558 118
rect 592 84 619 118
rect 497 52 619 84
rect 649 112 702 136
rect 649 78 660 112
rect 694 78 702 112
rect 649 52 702 78
<< pdiff >>
rect 27 600 80 619
rect 27 566 35 600
rect 69 566 80 600
rect 27 532 80 566
rect 27 498 35 532
rect 69 498 80 532
rect 27 456 80 498
rect 27 422 35 456
rect 69 422 80 456
rect 27 367 80 422
rect 110 594 232 619
rect 110 560 135 594
rect 169 560 232 594
rect 110 515 232 560
rect 110 481 135 515
rect 169 481 232 515
rect 110 419 232 481
rect 282 606 335 619
rect 282 572 293 606
rect 327 572 335 606
rect 282 538 335 572
rect 282 504 293 538
rect 327 504 335 538
rect 282 470 335 504
rect 282 436 293 470
rect 327 436 335 470
rect 282 419 335 436
rect 394 599 447 619
rect 394 565 402 599
rect 436 565 447 599
rect 394 466 447 565
rect 394 432 402 466
rect 436 432 447 466
rect 394 419 447 432
rect 497 607 619 619
rect 497 573 558 607
rect 592 573 619 607
rect 497 539 619 573
rect 497 505 558 539
rect 592 505 619 539
rect 497 471 619 505
rect 497 437 558 471
rect 592 437 619 471
rect 497 419 619 437
rect 110 367 160 419
rect 569 367 619 419
rect 649 599 702 619
rect 649 565 660 599
rect 694 565 702 599
rect 649 510 702 565
rect 649 476 660 510
rect 694 476 702 510
rect 649 413 702 476
rect 649 379 660 413
rect 694 379 702 413
rect 649 367 702 379
<< ndiffc >>
rect 35 77 69 111
rect 132 77 166 111
rect 293 206 327 240
rect 293 138 327 172
rect 293 70 327 104
rect 402 193 436 227
rect 402 70 436 104
rect 558 84 592 118
rect 660 78 694 112
<< pdiffc >>
rect 35 566 69 600
rect 35 498 69 532
rect 35 422 69 456
rect 135 560 169 594
rect 135 481 169 515
rect 293 572 327 606
rect 293 504 327 538
rect 293 436 327 470
rect 402 565 436 599
rect 402 432 436 466
rect 558 573 592 607
rect 558 505 592 539
rect 558 437 592 471
rect 660 565 694 599
rect 660 476 694 510
rect 660 379 694 413
<< poly >>
rect 80 619 110 645
rect 232 619 282 645
rect 447 619 497 645
rect 619 619 649 645
rect 232 386 282 419
rect 182 370 316 386
rect 80 333 110 367
rect 44 317 110 333
rect 44 283 60 317
rect 94 283 110 317
rect 44 267 110 283
rect 182 336 266 370
rect 300 336 316 370
rect 447 340 497 419
rect 182 324 316 336
rect 182 290 200 324
rect 234 320 316 324
rect 403 324 547 340
rect 234 290 282 320
rect 182 274 282 290
rect 403 290 419 324
rect 453 290 487 324
rect 521 290 547 324
rect 403 274 547 290
rect 619 325 649 367
rect 619 309 685 325
rect 619 275 635 309
rect 669 275 685 309
rect 80 136 110 267
rect 232 252 282 274
rect 447 252 497 274
rect 619 259 685 275
rect 619 136 649 259
rect 80 26 110 52
rect 232 26 282 52
rect 447 26 497 52
rect 619 26 649 52
<< polycont >>
rect 60 283 94 317
rect 266 336 300 370
rect 200 290 234 324
rect 419 290 453 324
rect 487 290 521 324
rect 635 275 669 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 19 600 85 615
rect 19 566 35 600
rect 69 566 85 600
rect 19 532 85 566
rect 19 498 35 532
rect 69 498 85 532
rect 19 456 85 498
rect 119 594 185 615
rect 119 545 135 594
rect 169 545 185 594
rect 119 515 185 545
rect 119 481 135 515
rect 169 481 185 515
rect 119 476 185 481
rect 277 606 368 615
rect 277 572 293 606
rect 327 572 368 606
rect 277 538 368 572
rect 277 504 293 538
rect 327 504 368 538
rect 277 479 368 504
rect 19 422 35 456
rect 69 441 85 456
rect 289 470 368 479
rect 69 422 253 441
rect 19 406 253 422
rect 289 436 293 470
rect 327 436 368 470
rect 289 420 368 436
rect 182 386 253 406
rect 20 317 110 372
rect 20 283 60 317
rect 94 283 110 317
rect 20 238 110 283
rect 182 370 300 386
rect 182 336 266 370
rect 182 324 300 336
rect 182 290 200 324
rect 234 320 300 324
rect 334 331 368 420
rect 402 599 452 615
rect 436 565 452 599
rect 402 466 452 565
rect 436 450 452 466
rect 542 607 608 615
rect 542 545 558 607
rect 592 545 608 607
rect 542 539 608 545
rect 542 505 558 539
rect 592 505 608 539
rect 542 471 608 505
rect 436 432 508 450
rect 542 437 558 471
rect 592 437 608 471
rect 542 433 608 437
rect 646 599 750 615
rect 646 565 660 599
rect 694 565 750 599
rect 646 510 750 565
rect 646 476 660 510
rect 694 476 750 510
rect 402 416 508 432
rect 474 399 508 416
rect 646 413 750 476
rect 474 365 605 399
rect 334 324 537 331
rect 234 290 253 320
rect 182 204 253 290
rect 334 290 419 324
rect 453 290 487 324
rect 521 290 537 324
rect 334 277 537 290
rect 571 325 605 365
rect 646 379 660 413
rect 694 379 750 413
rect 646 363 750 379
rect 571 309 669 325
rect 334 256 368 277
rect 19 164 253 204
rect 287 240 368 256
rect 571 275 635 309
rect 571 259 669 275
rect 571 243 605 259
rect 287 206 293 240
rect 327 206 368 240
rect 287 172 368 206
rect 19 111 82 164
rect 287 138 293 172
rect 327 138 368 172
rect 19 77 35 111
rect 69 77 82 111
rect 19 61 82 77
rect 116 111 182 130
rect 116 77 132 111
rect 166 77 182 111
rect 116 17 182 77
rect 287 104 368 138
rect 287 70 293 104
rect 327 70 368 104
rect 287 54 368 70
rect 402 227 605 243
rect 436 196 605 227
rect 436 193 452 196
rect 402 104 452 193
rect 436 70 452 104
rect 402 54 452 70
rect 542 118 608 134
rect 703 128 750 363
rect 542 84 558 118
rect 592 84 608 118
rect 542 17 608 84
rect 642 112 750 128
rect 642 78 660 112
rect 694 78 750 112
rect 642 62 750 78
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 135 560 169 579
rect 135 545 169 560
rect 558 573 592 579
rect 558 545 592 573
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 14 579 754 589
rect 14 545 135 579
rect 169 545 558 579
rect 592 545 754 579
rect 14 535 754 545
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlybuf4s25kapwr_1
flabel metal1 s 14 535 754 589 0 FreeSans 200 0 0 0 KAPWR
port 2 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 464 737 498 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 703 94 737 128 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y
string GDS_END 3557414
string GDS_START 3549934
<< end >>
