magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 24 157 212 241
rect 24 49 749 157
rect 0 0 768 49
<< scnmos >>
rect 103 47 133 215
rect 241 47 271 131
rect 338 47 368 131
rect 455 47 485 131
rect 541 47 571 131
rect 619 47 649 131
<< scpmoshvt >>
rect 122 367 152 619
rect 475 529 505 613
rect 561 529 591 613
rect 647 529 677 613
rect 241 367 271 451
rect 319 367 349 451
<< ndiff >>
rect 50 203 103 215
rect 50 169 58 203
rect 92 169 103 203
rect 50 101 103 169
rect 50 67 58 101
rect 92 67 103 101
rect 50 47 103 67
rect 133 203 186 215
rect 133 169 144 203
rect 178 169 186 203
rect 133 131 186 169
rect 133 93 241 131
rect 133 59 144 93
rect 178 59 241 93
rect 133 47 241 59
rect 271 106 338 131
rect 271 72 293 106
rect 327 72 338 106
rect 271 47 338 72
rect 368 96 455 131
rect 368 62 394 96
rect 428 62 455 96
rect 368 47 455 62
rect 485 106 541 131
rect 485 72 496 106
rect 530 72 541 106
rect 485 47 541 72
rect 571 47 619 131
rect 649 106 723 131
rect 649 72 681 106
rect 715 72 723 106
rect 649 47 723 72
<< pdiff >>
rect 69 599 122 619
rect 69 565 77 599
rect 111 565 122 599
rect 69 506 122 565
rect 69 472 77 506
rect 111 472 122 506
rect 69 413 122 472
rect 69 379 77 413
rect 111 379 122 413
rect 69 367 122 379
rect 152 575 205 619
rect 152 541 163 575
rect 197 541 205 575
rect 152 451 205 541
rect 422 588 475 613
rect 422 554 430 588
rect 464 554 475 588
rect 422 529 475 554
rect 505 588 561 613
rect 505 554 516 588
rect 550 554 561 588
rect 505 529 561 554
rect 591 588 647 613
rect 591 554 602 588
rect 636 554 647 588
rect 591 529 647 554
rect 677 588 730 613
rect 677 554 688 588
rect 722 554 730 588
rect 677 529 730 554
rect 152 367 241 451
rect 271 367 319 451
rect 349 413 402 451
rect 349 379 360 413
rect 394 379 402 413
rect 349 367 402 379
<< ndiffc >>
rect 58 169 92 203
rect 58 67 92 101
rect 144 169 178 203
rect 144 59 178 93
rect 293 72 327 106
rect 394 62 428 96
rect 496 72 530 106
rect 681 72 715 106
<< pdiffc >>
rect 77 565 111 599
rect 77 472 111 506
rect 77 379 111 413
rect 163 541 197 575
rect 430 554 464 588
rect 516 554 550 588
rect 602 554 636 588
rect 688 554 722 588
rect 360 379 394 413
<< poly >>
rect 122 619 152 645
rect 475 613 505 639
rect 561 613 591 639
rect 647 613 677 639
rect 241 451 271 477
rect 319 451 349 477
rect 475 458 505 529
rect 463 428 505 458
rect 122 335 152 367
rect 241 335 271 367
rect 91 319 157 335
rect 91 285 107 319
rect 141 285 157 319
rect 91 269 157 285
rect 205 319 274 335
rect 205 285 221 319
rect 255 285 274 319
rect 103 215 133 269
rect 205 251 274 285
rect 205 217 224 251
rect 258 217 274 251
rect 205 201 274 217
rect 319 321 349 367
rect 463 335 493 428
rect 561 380 591 529
rect 647 452 677 529
rect 647 422 711 452
rect 319 305 385 321
rect 319 271 335 305
rect 369 271 385 305
rect 319 237 385 271
rect 319 203 335 237
rect 369 203 385 237
rect 241 131 271 201
rect 319 187 385 203
rect 427 319 493 335
rect 427 285 443 319
rect 477 285 493 319
rect 427 251 493 285
rect 427 217 443 251
rect 477 217 493 251
rect 427 201 493 217
rect 541 364 633 380
rect 541 330 583 364
rect 617 330 633 364
rect 541 296 633 330
rect 541 262 583 296
rect 617 262 633 296
rect 541 246 633 262
rect 681 302 711 422
rect 681 286 747 302
rect 681 252 697 286
rect 731 252 747 286
rect 338 131 368 187
rect 455 131 485 201
rect 541 131 571 246
rect 681 218 747 252
rect 681 198 697 218
rect 619 184 697 198
rect 731 184 747 218
rect 619 168 747 184
rect 619 131 649 168
rect 103 21 133 47
rect 241 21 271 47
rect 338 21 368 47
rect 455 21 485 47
rect 541 21 571 47
rect 619 21 649 47
<< polycont >>
rect 107 285 141 319
rect 221 285 255 319
rect 224 217 258 251
rect 335 271 369 305
rect 335 203 369 237
rect 443 285 477 319
rect 443 217 477 251
rect 583 330 617 364
rect 583 262 617 296
rect 697 252 731 286
rect 697 184 731 218
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 21 599 113 615
rect 21 565 77 599
rect 111 565 113 599
rect 21 506 113 565
rect 147 575 213 649
rect 147 541 163 575
rect 197 541 213 575
rect 147 533 213 541
rect 414 588 473 604
rect 414 554 430 588
rect 464 554 473 588
rect 21 472 77 506
rect 111 472 113 506
rect 414 499 473 554
rect 21 413 113 472
rect 21 379 77 413
rect 111 379 113 413
rect 21 363 113 379
rect 151 465 473 499
rect 507 588 552 604
rect 507 554 516 588
rect 550 554 552 588
rect 507 513 552 554
rect 586 588 652 649
rect 586 554 602 588
rect 636 554 652 588
rect 586 547 652 554
rect 686 588 738 604
rect 686 554 688 588
rect 722 554 738 588
rect 686 513 738 554
rect 507 479 738 513
rect 21 219 57 363
rect 151 329 185 465
rect 434 445 473 465
rect 91 319 185 329
rect 91 285 107 319
rect 141 285 185 319
rect 91 269 185 285
rect 221 319 259 431
rect 356 413 398 429
rect 356 379 360 413
rect 394 379 398 413
rect 434 411 547 445
rect 356 375 398 379
rect 356 341 477 375
rect 255 285 259 319
rect 422 319 477 341
rect 221 251 259 285
rect 21 203 101 219
rect 21 169 58 203
rect 92 169 101 203
rect 21 101 101 169
rect 21 67 58 101
rect 92 67 101 101
rect 21 51 101 67
rect 135 203 187 219
rect 135 169 144 203
rect 178 169 187 203
rect 135 93 187 169
rect 135 59 144 93
rect 178 59 187 93
rect 221 217 224 251
rect 258 217 259 251
rect 221 74 259 217
rect 293 271 335 305
rect 369 271 385 305
rect 293 237 385 271
rect 293 203 335 237
rect 369 203 385 237
rect 422 285 443 319
rect 422 251 477 285
rect 422 217 443 251
rect 422 201 477 217
rect 422 167 456 201
rect 293 133 456 167
rect 513 135 547 411
rect 293 106 343 133
rect 135 17 187 59
rect 327 72 343 106
rect 490 106 547 135
rect 293 56 343 72
rect 378 96 444 99
rect 378 62 394 96
rect 428 62 444 96
rect 378 17 444 62
rect 490 72 496 106
rect 530 72 547 106
rect 490 56 547 72
rect 583 364 643 445
rect 617 330 643 364
rect 583 296 643 330
rect 617 262 643 296
rect 583 56 643 262
rect 677 286 751 445
rect 677 252 697 286
rect 731 252 751 286
rect 677 218 751 252
rect 677 184 697 218
rect 731 184 751 218
rect 677 168 751 184
rect 677 106 731 122
rect 677 72 681 106
rect 715 72 731 106
rect 677 17 731 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2bb2o_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5903388
string GDS_START 5895012
<< end >>
