magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 11 49 671 167
rect 0 0 672 49
<< scnmos >>
rect 110 57 140 141
rect 202 57 232 141
rect 314 57 344 141
rect 400 57 430 141
rect 486 57 516 141
rect 558 57 588 141
<< scpmoshvt >>
rect 100 410 150 610
rect 206 410 256 610
rect 310 410 360 610
rect 418 410 468 610
rect 524 410 574 610
<< ndiff >>
rect 37 116 110 141
rect 37 82 49 116
rect 83 82 110 116
rect 37 57 110 82
rect 140 116 202 141
rect 140 82 151 116
rect 185 82 202 116
rect 140 57 202 82
rect 232 103 314 141
rect 232 69 253 103
rect 287 69 314 103
rect 232 57 314 69
rect 344 116 400 141
rect 344 82 355 116
rect 389 82 400 116
rect 344 57 400 82
rect 430 116 486 141
rect 430 82 441 116
rect 475 82 486 116
rect 430 57 486 82
rect 516 57 558 141
rect 588 116 645 141
rect 588 82 599 116
rect 633 82 645 116
rect 588 57 645 82
<< pdiff >>
rect 43 598 100 610
rect 43 564 55 598
rect 89 564 100 598
rect 43 515 100 564
rect 43 481 55 515
rect 89 481 100 515
rect 43 410 100 481
rect 150 597 206 610
rect 150 563 161 597
rect 195 563 206 597
rect 150 526 206 563
rect 150 492 161 526
rect 195 492 206 526
rect 150 456 206 492
rect 150 422 161 456
rect 195 422 206 456
rect 150 410 206 422
rect 256 410 310 610
rect 360 410 418 610
rect 468 598 524 610
rect 468 564 479 598
rect 513 564 524 598
rect 468 524 524 564
rect 468 490 479 524
rect 513 490 524 524
rect 468 410 524 490
rect 574 597 631 610
rect 574 563 585 597
rect 619 563 631 597
rect 574 526 631 563
rect 574 492 585 526
rect 619 492 631 526
rect 574 456 631 492
rect 574 422 585 456
rect 619 422 631 456
rect 574 410 631 422
<< ndiffc >>
rect 49 82 83 116
rect 151 82 185 116
rect 253 69 287 103
rect 355 82 389 116
rect 441 82 475 116
rect 599 82 633 116
<< pdiffc >>
rect 55 564 89 598
rect 55 481 89 515
rect 161 563 195 597
rect 161 492 195 526
rect 161 422 195 456
rect 479 564 513 598
rect 479 490 513 524
rect 585 563 619 597
rect 585 492 619 526
rect 585 422 619 456
<< poly >>
rect 100 610 150 636
rect 206 610 256 636
rect 310 610 360 636
rect 418 610 468 636
rect 524 610 574 636
rect 100 359 150 410
rect 206 359 256 410
rect 310 368 360 410
rect 418 368 468 410
rect 88 343 154 359
rect 88 309 104 343
rect 138 309 154 343
rect 88 275 154 309
rect 88 241 104 275
rect 138 241 154 275
rect 88 225 154 241
rect 196 343 262 359
rect 196 309 212 343
rect 246 309 262 343
rect 196 275 262 309
rect 196 241 212 275
rect 246 241 262 275
rect 196 225 262 241
rect 304 352 370 368
rect 304 318 320 352
rect 354 318 370 352
rect 304 284 370 318
rect 304 250 320 284
rect 354 250 370 284
rect 304 234 370 250
rect 412 352 478 368
rect 412 318 428 352
rect 462 318 478 352
rect 524 320 574 410
rect 412 284 478 318
rect 412 250 428 284
rect 462 250 478 284
rect 412 234 478 250
rect 520 304 588 320
rect 520 270 536 304
rect 570 270 588 304
rect 520 236 588 270
rect 110 141 140 225
rect 202 141 232 225
rect 314 141 344 234
rect 412 186 442 234
rect 520 202 536 236
rect 570 202 588 236
rect 520 186 588 202
rect 400 156 442 186
rect 486 156 588 186
rect 400 141 430 156
rect 486 141 516 156
rect 558 141 588 156
rect 110 31 140 57
rect 202 31 232 57
rect 314 31 344 57
rect 400 31 430 57
rect 486 31 516 57
rect 558 31 588 57
<< polycont >>
rect 104 309 138 343
rect 104 241 138 275
rect 212 309 246 343
rect 212 241 246 275
rect 320 318 354 352
rect 320 250 354 284
rect 428 318 462 352
rect 428 250 462 284
rect 536 270 570 304
rect 536 202 570 236
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 39 598 105 649
rect 39 564 55 598
rect 89 564 105 598
rect 39 515 105 564
rect 39 481 55 515
rect 89 481 105 515
rect 39 465 105 481
rect 145 597 211 613
rect 145 563 161 597
rect 195 563 211 597
rect 145 526 211 563
rect 145 492 161 526
rect 195 492 211 526
rect 145 456 211 492
rect 463 598 529 649
rect 463 564 479 598
rect 513 564 529 598
rect 463 524 529 564
rect 463 490 479 524
rect 513 490 529 524
rect 463 474 529 490
rect 585 597 654 613
rect 619 563 654 597
rect 585 526 654 563
rect 619 492 654 526
rect 145 429 161 456
rect 18 422 161 429
rect 195 438 211 456
rect 585 456 654 492
rect 195 422 549 438
rect 18 404 549 422
rect 18 395 211 404
rect 18 145 52 395
rect 88 343 161 359
rect 88 309 104 343
rect 138 309 161 343
rect 88 275 161 309
rect 88 241 104 275
rect 138 241 161 275
rect 88 225 161 241
rect 197 343 263 359
rect 197 309 212 343
rect 246 309 263 343
rect 197 275 263 309
rect 197 241 212 275
rect 246 241 263 275
rect 197 225 263 241
rect 304 352 370 368
rect 304 318 320 352
rect 354 318 370 352
rect 304 284 370 318
rect 304 250 320 284
rect 354 250 370 284
rect 304 234 370 250
rect 409 352 478 368
rect 409 318 428 352
rect 462 318 478 352
rect 409 284 478 318
rect 409 250 428 284
rect 462 250 478 284
rect 409 234 478 250
rect 515 320 549 404
rect 619 422 654 456
rect 585 384 654 422
rect 515 304 584 320
rect 515 270 536 304
rect 570 270 584 304
rect 515 236 584 270
rect 515 202 536 236
rect 570 202 584 236
rect 135 155 389 189
rect 515 186 584 202
rect 18 116 99 145
rect 18 82 49 116
rect 83 82 99 116
rect 18 53 99 82
rect 135 116 201 155
rect 135 82 151 116
rect 185 82 201 116
rect 135 53 201 82
rect 237 103 303 119
rect 237 69 253 103
rect 287 69 303 103
rect 237 17 303 69
rect 339 116 389 155
rect 620 145 654 384
rect 339 82 355 116
rect 339 53 389 82
rect 425 116 491 145
rect 425 82 441 116
rect 475 82 491 116
rect 425 17 491 82
rect 583 116 654 145
rect 583 82 599 116
rect 633 82 654 116
rect 583 53 654 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o31a_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1236880
string GDS_START 1229896
<< end >>
