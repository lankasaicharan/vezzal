magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
rect 465 319 907 331
<< pwell >>
rect 1072 241 1533 263
rect 2 49 1533 241
rect 0 0 1536 49
<< scnmos >>
rect 81 47 111 215
rect 167 47 197 215
rect 261 47 291 215
rect 347 47 377 215
rect 435 47 465 215
rect 521 47 551 215
rect 607 47 637 215
rect 693 47 723 215
rect 847 47 877 215
rect 933 47 963 215
rect 1151 69 1181 237
rect 1252 69 1282 237
rect 1338 69 1368 237
rect 1424 69 1454 237
<< scpmoshvt >>
rect 81 367 111 619
rect 167 367 197 619
rect 253 367 283 619
rect 347 367 377 619
rect 573 355 603 607
rect 659 355 689 607
rect 769 355 799 607
rect 893 367 923 619
rect 979 367 1009 619
rect 1065 367 1095 619
rect 1151 367 1181 619
rect 1237 367 1267 619
rect 1338 367 1368 619
rect 1424 367 1454 619
<< ndiff >>
rect 28 203 81 215
rect 28 169 36 203
rect 70 169 81 203
rect 28 93 81 169
rect 28 59 36 93
rect 70 59 81 93
rect 28 47 81 59
rect 111 197 167 215
rect 111 163 122 197
rect 156 163 167 197
rect 111 101 167 163
rect 111 67 122 101
rect 156 67 167 101
rect 111 47 167 67
rect 197 181 261 215
rect 197 147 211 181
rect 245 147 261 181
rect 197 89 261 147
rect 197 55 211 89
rect 245 55 261 89
rect 197 47 261 55
rect 291 203 347 215
rect 291 169 302 203
rect 336 169 347 203
rect 291 101 347 169
rect 291 67 302 101
rect 336 67 347 101
rect 291 47 347 67
rect 377 181 435 215
rect 377 147 388 181
rect 422 147 435 181
rect 377 93 435 147
rect 377 59 388 93
rect 422 59 435 93
rect 377 47 435 59
rect 465 203 521 215
rect 465 169 476 203
rect 510 169 521 203
rect 465 101 521 169
rect 465 67 476 101
rect 510 67 521 101
rect 465 47 521 67
rect 551 171 607 215
rect 551 137 562 171
rect 596 137 607 171
rect 551 93 607 137
rect 551 59 562 93
rect 596 59 607 93
rect 551 47 607 59
rect 637 203 693 215
rect 637 169 648 203
rect 682 169 693 203
rect 637 101 693 169
rect 637 67 648 101
rect 682 67 693 101
rect 637 47 693 67
rect 723 171 847 215
rect 723 137 734 171
rect 768 137 802 171
rect 836 137 847 171
rect 723 93 847 137
rect 723 59 734 93
rect 768 59 802 93
rect 836 59 847 93
rect 723 47 847 59
rect 877 203 933 215
rect 877 169 888 203
rect 922 169 933 203
rect 877 101 933 169
rect 877 67 888 101
rect 922 67 933 101
rect 877 47 933 67
rect 963 169 1030 215
rect 963 135 974 169
rect 1008 135 1030 169
rect 963 93 1030 135
rect 963 59 974 93
rect 1008 59 1030 93
rect 1098 151 1151 237
rect 1098 117 1106 151
rect 1140 117 1151 151
rect 1098 69 1151 117
rect 1181 229 1252 237
rect 1181 195 1199 229
rect 1233 195 1252 229
rect 1181 153 1252 195
rect 1181 119 1199 153
rect 1233 119 1252 153
rect 1181 69 1252 119
rect 1282 219 1338 237
rect 1282 185 1293 219
rect 1327 185 1338 219
rect 1282 115 1338 185
rect 1282 81 1293 115
rect 1327 81 1338 115
rect 1282 69 1338 81
rect 1368 229 1424 237
rect 1368 195 1379 229
rect 1413 195 1424 229
rect 1368 153 1424 195
rect 1368 119 1379 153
rect 1413 119 1424 153
rect 1368 69 1424 119
rect 1454 192 1507 237
rect 1454 158 1465 192
rect 1499 158 1507 192
rect 1454 115 1507 158
rect 1454 81 1465 115
rect 1499 81 1507 115
rect 1454 69 1507 81
rect 963 47 1030 59
<< pdiff >>
rect 28 599 81 619
rect 28 565 36 599
rect 70 565 81 599
rect 28 507 81 565
rect 28 473 36 507
rect 70 473 81 507
rect 28 418 81 473
rect 28 384 36 418
rect 70 384 81 418
rect 28 367 81 384
rect 111 531 167 619
rect 111 497 122 531
rect 156 497 167 531
rect 111 436 167 497
rect 111 402 122 436
rect 156 402 167 436
rect 111 367 167 402
rect 197 599 253 619
rect 197 565 208 599
rect 242 565 253 599
rect 197 507 253 565
rect 197 473 208 507
rect 242 473 253 507
rect 197 418 253 473
rect 197 384 208 418
rect 242 384 253 418
rect 197 367 253 384
rect 283 531 347 619
rect 283 497 298 531
rect 332 497 347 531
rect 283 434 347 497
rect 283 400 298 434
rect 332 400 347 434
rect 283 367 347 400
rect 377 599 430 619
rect 377 565 388 599
rect 422 565 430 599
rect 377 502 430 565
rect 377 468 388 502
rect 422 468 430 502
rect 377 367 430 468
rect 501 607 551 619
rect 704 611 754 623
rect 704 607 712 611
rect 501 573 509 607
rect 543 573 573 607
rect 501 355 573 573
rect 603 397 659 607
rect 603 363 614 397
rect 648 363 659 397
rect 603 355 659 363
rect 689 577 712 607
rect 746 607 754 611
rect 821 607 893 619
rect 746 577 769 607
rect 689 355 769 577
rect 799 401 893 607
rect 799 367 829 401
rect 863 367 893 401
rect 923 611 979 619
rect 923 577 934 611
rect 968 577 979 611
rect 923 367 979 577
rect 1009 599 1065 619
rect 1009 565 1020 599
rect 1054 565 1065 599
rect 1009 486 1065 565
rect 1009 452 1020 486
rect 1054 452 1065 486
rect 1009 367 1065 452
rect 1095 562 1151 619
rect 1095 528 1106 562
rect 1140 528 1151 562
rect 1095 367 1151 528
rect 1181 599 1237 619
rect 1181 565 1192 599
rect 1226 565 1237 599
rect 1181 486 1237 565
rect 1181 452 1192 486
rect 1226 452 1237 486
rect 1181 367 1237 452
rect 1267 562 1338 619
rect 1267 528 1285 562
rect 1319 528 1338 562
rect 1267 367 1338 528
rect 1368 599 1424 619
rect 1368 565 1379 599
rect 1413 565 1424 599
rect 1368 507 1424 565
rect 1368 473 1379 507
rect 1413 473 1424 507
rect 1368 413 1424 473
rect 1368 379 1379 413
rect 1413 379 1424 413
rect 1368 367 1424 379
rect 1454 607 1507 619
rect 1454 573 1465 607
rect 1499 573 1507 607
rect 1454 513 1507 573
rect 1454 479 1465 513
rect 1499 479 1507 513
rect 1454 418 1507 479
rect 1454 384 1465 418
rect 1499 384 1507 418
rect 1454 367 1507 384
rect 799 355 871 367
<< ndiffc >>
rect 36 169 70 203
rect 36 59 70 93
rect 122 163 156 197
rect 122 67 156 101
rect 211 147 245 181
rect 211 55 245 89
rect 302 169 336 203
rect 302 67 336 101
rect 388 147 422 181
rect 388 59 422 93
rect 476 169 510 203
rect 476 67 510 101
rect 562 137 596 171
rect 562 59 596 93
rect 648 169 682 203
rect 648 67 682 101
rect 734 137 768 171
rect 802 137 836 171
rect 734 59 768 93
rect 802 59 836 93
rect 888 169 922 203
rect 888 67 922 101
rect 974 135 1008 169
rect 974 59 1008 93
rect 1106 117 1140 151
rect 1199 195 1233 229
rect 1199 119 1233 153
rect 1293 185 1327 219
rect 1293 81 1327 115
rect 1379 195 1413 229
rect 1379 119 1413 153
rect 1465 158 1499 192
rect 1465 81 1499 115
<< pdiffc >>
rect 36 565 70 599
rect 36 473 70 507
rect 36 384 70 418
rect 122 497 156 531
rect 122 402 156 436
rect 208 565 242 599
rect 208 473 242 507
rect 208 384 242 418
rect 298 497 332 531
rect 298 400 332 434
rect 388 565 422 599
rect 388 468 422 502
rect 509 573 543 607
rect 614 363 648 397
rect 712 577 746 611
rect 829 367 863 401
rect 934 577 968 611
rect 1020 565 1054 599
rect 1020 452 1054 486
rect 1106 528 1140 562
rect 1192 565 1226 599
rect 1192 452 1226 486
rect 1285 528 1319 562
rect 1379 565 1413 599
rect 1379 473 1413 507
rect 1379 379 1413 413
rect 1465 573 1499 607
rect 1465 479 1499 513
rect 1465 384 1499 418
<< poly >>
rect 81 619 111 645
rect 167 619 197 645
rect 253 619 283 645
rect 347 619 377 645
rect 573 607 603 633
rect 659 607 689 633
rect 81 308 111 367
rect 167 308 197 367
rect 253 333 283 367
rect 347 333 377 367
rect 769 607 799 633
rect 893 619 923 645
rect 979 619 1009 645
rect 1065 619 1095 645
rect 1151 619 1181 645
rect 1237 619 1267 645
rect 1338 619 1368 645
rect 1424 619 1454 645
rect 32 292 197 308
rect 32 258 48 292
rect 82 258 197 292
rect 239 317 377 333
rect 573 323 603 355
rect 659 323 689 355
rect 769 340 799 355
rect 893 340 923 367
rect 769 323 923 340
rect 239 283 255 317
rect 289 283 323 317
rect 357 283 377 317
rect 239 258 377 283
rect 32 242 197 258
rect 81 215 111 242
rect 167 215 197 242
rect 261 215 291 258
rect 347 215 377 258
rect 435 310 923 323
rect 979 333 1009 367
rect 1065 333 1095 367
rect 979 317 1095 333
rect 435 307 799 310
rect 435 273 451 307
rect 485 273 519 307
rect 553 273 587 307
rect 621 273 655 307
rect 689 273 723 307
rect 757 293 799 307
rect 757 273 773 293
rect 435 257 773 273
rect 979 283 1020 317
rect 1054 283 1095 317
rect 979 268 1095 283
rect 871 267 1095 268
rect 1151 335 1181 367
rect 1237 335 1267 367
rect 1151 319 1289 335
rect 1151 285 1171 319
rect 1205 285 1239 319
rect 1273 285 1289 319
rect 1151 269 1289 285
rect 1338 325 1368 367
rect 1424 325 1454 367
rect 1338 309 1515 325
rect 1338 275 1465 309
rect 1499 275 1515 309
rect 435 215 465 257
rect 521 215 551 257
rect 607 215 637 257
rect 693 215 723 257
rect 847 238 1055 267
rect 847 232 963 238
rect 1151 237 1181 269
rect 1252 237 1282 269
rect 1338 259 1515 275
rect 1338 237 1368 259
rect 1424 237 1454 259
rect 847 215 877 232
rect 933 215 963 232
rect 81 21 111 47
rect 167 21 197 47
rect 261 21 291 47
rect 347 21 377 47
rect 435 21 465 47
rect 521 21 551 47
rect 607 21 637 47
rect 693 21 723 47
rect 847 21 877 47
rect 933 21 963 47
rect 1151 43 1181 69
rect 1252 43 1282 69
rect 1338 43 1368 69
rect 1424 43 1454 69
<< polycont >>
rect 48 258 82 292
rect 255 283 289 317
rect 323 283 357 317
rect 451 273 485 307
rect 519 273 553 307
rect 587 273 621 307
rect 655 273 689 307
rect 723 273 757 307
rect 1020 283 1054 317
rect 1171 285 1205 319
rect 1239 285 1273 319
rect 1465 275 1499 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 20 599 424 615
rect 20 565 36 599
rect 70 581 208 599
rect 70 565 86 581
rect 20 507 86 565
rect 192 565 208 581
rect 242 581 388 599
rect 242 565 258 581
rect 20 473 36 507
rect 70 473 86 507
rect 20 418 86 473
rect 20 384 36 418
rect 70 384 86 418
rect 120 531 158 547
rect 120 497 122 531
rect 156 497 158 531
rect 120 436 158 497
rect 120 402 122 436
rect 156 402 158 436
rect 17 292 86 350
rect 17 258 48 292
rect 82 258 86 292
rect 17 242 86 258
rect 120 249 158 402
rect 192 507 258 565
rect 372 565 388 581
rect 422 565 424 599
rect 493 607 559 649
rect 493 573 509 607
rect 543 573 559 607
rect 696 611 762 649
rect 696 577 712 611
rect 746 577 762 611
rect 696 573 762 577
rect 918 611 984 649
rect 918 577 934 611
rect 968 577 984 611
rect 918 573 984 577
rect 1018 599 1056 615
rect 192 473 208 507
rect 242 473 258 507
rect 192 418 258 473
rect 192 384 208 418
rect 242 384 258 418
rect 292 531 338 547
rect 292 497 298 531
rect 332 497 338 531
rect 292 434 338 497
rect 372 502 424 565
rect 1018 565 1020 599
rect 1054 565 1056 599
rect 1018 539 1056 565
rect 372 468 388 502
rect 422 468 424 502
rect 372 452 424 468
rect 458 505 1056 539
rect 1090 562 1156 649
rect 1090 528 1106 562
rect 1140 528 1156 562
rect 1090 520 1156 528
rect 1190 599 1232 615
rect 1190 565 1192 599
rect 1226 565 1232 599
rect 292 400 298 434
rect 332 418 338 434
rect 458 418 492 505
rect 1004 486 1056 505
rect 1190 486 1232 565
rect 1269 562 1335 649
rect 1269 528 1285 562
rect 1319 528 1335 562
rect 1269 520 1335 528
rect 1369 599 1415 615
rect 1369 565 1379 599
rect 1413 565 1415 599
rect 1369 507 1415 565
rect 1369 486 1379 507
rect 332 400 492 418
rect 292 384 492 400
rect 528 437 947 471
rect 1004 452 1020 486
rect 1054 452 1192 486
rect 1226 473 1379 486
rect 1413 473 1415 507
rect 1226 452 1415 473
rect 194 317 373 350
rect 528 317 562 437
rect 913 418 947 437
rect 598 401 879 403
rect 598 397 829 401
rect 598 363 614 397
rect 648 367 829 397
rect 863 367 879 401
rect 913 384 1343 418
rect 648 363 879 367
rect 598 350 879 363
rect 194 283 255 317
rect 289 283 323 317
rect 357 283 373 317
rect 407 307 562 317
rect 407 273 451 307
rect 485 273 519 307
rect 553 273 587 307
rect 621 273 655 307
rect 689 273 723 307
rect 757 273 773 307
rect 812 281 945 350
rect 979 317 1121 350
rect 979 283 1020 317
rect 1054 283 1121 317
rect 1155 319 1275 350
rect 1155 285 1171 319
rect 1205 285 1239 319
rect 1273 285 1275 319
rect 407 249 441 273
rect 120 215 441 249
rect 812 239 846 281
rect 1155 269 1275 285
rect 1309 329 1343 384
rect 1377 413 1415 452
rect 1377 379 1379 413
rect 1413 379 1415 413
rect 1449 607 1515 649
rect 1449 573 1465 607
rect 1499 573 1515 607
rect 1449 513 1515 573
rect 1449 479 1465 513
rect 1499 479 1515 513
rect 1449 418 1515 479
rect 1449 384 1465 418
rect 1499 384 1515 418
rect 1377 363 1415 379
rect 1309 269 1429 329
rect 20 203 86 208
rect 20 169 36 203
rect 70 169 86 203
rect 20 93 86 169
rect 20 59 36 93
rect 70 59 86 93
rect 20 17 86 59
rect 120 197 161 215
rect 120 163 122 197
rect 156 163 161 197
rect 295 203 338 215
rect 120 101 161 163
rect 120 67 122 101
rect 156 67 161 101
rect 120 51 161 67
rect 195 147 211 181
rect 245 147 261 181
rect 195 89 261 147
rect 195 55 211 89
rect 245 55 261 89
rect 195 17 261 55
rect 295 169 302 203
rect 336 169 338 203
rect 475 205 846 239
rect 886 235 1076 247
rect 886 229 1249 235
rect 886 213 1199 229
rect 475 203 512 205
rect 295 101 338 169
rect 295 67 302 101
rect 336 67 338 101
rect 295 51 338 67
rect 372 147 388 181
rect 422 147 438 181
rect 372 93 438 147
rect 372 59 388 93
rect 422 59 438 93
rect 372 17 438 59
rect 475 169 476 203
rect 510 169 512 203
rect 646 203 684 205
rect 475 101 512 169
rect 475 67 476 101
rect 510 67 512 101
rect 475 51 512 67
rect 546 137 562 171
rect 596 137 612 171
rect 546 93 612 137
rect 546 59 562 93
rect 596 59 612 93
rect 546 17 612 59
rect 646 169 648 203
rect 682 169 684 203
rect 886 203 924 213
rect 646 101 684 169
rect 646 67 648 101
rect 682 67 684 101
rect 646 51 684 67
rect 718 137 734 171
rect 768 137 802 171
rect 836 137 852 171
rect 718 93 852 137
rect 718 59 734 93
rect 768 59 802 93
rect 836 59 852 93
rect 718 17 852 59
rect 886 169 888 203
rect 922 169 924 203
rect 1042 201 1199 213
rect 1183 195 1199 201
rect 1233 195 1249 229
rect 886 101 924 169
rect 886 67 888 101
rect 922 67 924 101
rect 886 51 924 67
rect 958 135 974 169
rect 1008 135 1024 169
rect 958 93 1024 135
rect 958 59 974 93
rect 1008 59 1024 93
rect 958 17 1024 59
rect 1090 151 1149 167
rect 1090 117 1106 151
rect 1140 117 1149 151
rect 1183 153 1249 195
rect 1183 119 1199 153
rect 1233 119 1249 153
rect 1283 219 1329 235
rect 1283 185 1293 219
rect 1327 185 1329 219
rect 1090 85 1149 117
rect 1283 115 1329 185
rect 1363 229 1429 269
rect 1463 309 1519 350
rect 1463 275 1465 309
rect 1499 275 1519 309
rect 1463 242 1519 275
rect 1363 195 1379 229
rect 1413 195 1429 229
rect 1363 153 1429 195
rect 1363 119 1379 153
rect 1413 119 1429 153
rect 1463 192 1515 208
rect 1463 158 1465 192
rect 1499 158 1515 192
rect 1283 85 1293 115
rect 1090 81 1293 85
rect 1327 85 1329 115
rect 1463 115 1515 158
rect 1463 85 1465 115
rect 1327 81 1465 85
rect 1499 81 1515 115
rect 1090 51 1515 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a311o_4
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2826362
string GDS_START 2813456
<< end >>
