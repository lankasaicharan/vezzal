magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 3 241 297 267
rect 579 241 767 263
rect 3 49 767 241
rect 0 0 768 49
<< scnmos >>
rect 86 73 116 241
rect 182 73 212 241
rect 378 47 408 215
rect 464 47 494 215
rect 658 69 688 237
<< scpmoshvt >>
rect 110 367 140 619
rect 206 367 236 619
rect 304 367 334 619
rect 428 367 458 619
rect 650 367 680 619
<< ndiff >>
rect 29 219 86 241
rect 29 185 37 219
rect 71 185 86 219
rect 29 119 86 185
rect 29 85 37 119
rect 71 85 86 119
rect 29 73 86 85
rect 116 229 182 241
rect 116 195 127 229
rect 161 195 182 229
rect 116 153 182 195
rect 116 119 127 153
rect 161 119 182 153
rect 116 73 182 119
rect 212 229 271 241
rect 212 195 227 229
rect 261 195 271 229
rect 212 153 271 195
rect 212 119 227 153
rect 261 119 271 153
rect 212 73 271 119
rect 325 181 378 215
rect 325 147 333 181
rect 367 147 378 181
rect 325 93 378 147
rect 325 59 333 93
rect 367 59 378 93
rect 325 47 378 59
rect 408 165 464 215
rect 408 131 419 165
rect 453 131 464 165
rect 408 93 464 131
rect 408 59 419 93
rect 453 59 464 93
rect 408 47 464 59
rect 494 203 547 215
rect 494 169 505 203
rect 539 169 547 203
rect 494 101 547 169
rect 494 67 505 101
rect 539 67 547 101
rect 605 203 658 237
rect 605 169 613 203
rect 647 169 658 203
rect 605 122 658 169
rect 605 88 613 122
rect 647 88 658 122
rect 605 69 658 88
rect 688 208 741 237
rect 688 174 699 208
rect 733 174 741 208
rect 688 115 741 174
rect 688 81 699 115
rect 733 81 741 115
rect 688 69 741 81
rect 494 47 547 67
<< pdiff >>
rect 52 599 110 619
rect 52 565 65 599
rect 99 565 110 599
rect 52 515 110 565
rect 52 481 65 515
rect 99 481 110 515
rect 52 436 110 481
rect 52 402 60 436
rect 94 402 110 436
rect 52 367 110 402
rect 140 424 206 619
rect 140 390 151 424
rect 185 390 206 424
rect 140 367 206 390
rect 236 367 304 619
rect 334 607 428 619
rect 334 573 375 607
rect 409 573 428 607
rect 334 536 428 573
rect 334 502 375 536
rect 409 502 428 536
rect 334 465 428 502
rect 334 431 375 465
rect 409 431 428 465
rect 334 367 428 431
rect 458 599 511 619
rect 458 565 469 599
rect 503 565 511 599
rect 458 508 511 565
rect 458 474 469 508
rect 503 474 511 508
rect 458 413 511 474
rect 458 379 469 413
rect 503 379 511 413
rect 458 367 511 379
rect 597 599 650 619
rect 597 565 605 599
rect 639 565 650 599
rect 597 517 650 565
rect 597 483 605 517
rect 639 483 650 517
rect 597 426 650 483
rect 597 392 605 426
rect 639 392 650 426
rect 597 367 650 392
rect 680 607 733 619
rect 680 573 691 607
rect 725 573 733 607
rect 680 514 733 573
rect 680 480 691 514
rect 725 480 733 514
rect 680 418 733 480
rect 680 384 691 418
rect 725 384 733 418
rect 680 367 733 384
<< ndiffc >>
rect 37 185 71 219
rect 37 85 71 119
rect 127 195 161 229
rect 127 119 161 153
rect 227 195 261 229
rect 227 119 261 153
rect 333 147 367 181
rect 333 59 367 93
rect 419 131 453 165
rect 419 59 453 93
rect 505 169 539 203
rect 505 67 539 101
rect 613 169 647 203
rect 613 88 647 122
rect 699 174 733 208
rect 699 81 733 115
<< pdiffc >>
rect 65 565 99 599
rect 65 481 99 515
rect 60 402 94 436
rect 151 390 185 424
rect 375 573 409 607
rect 375 502 409 536
rect 375 431 409 465
rect 469 565 503 599
rect 469 474 503 508
rect 469 379 503 413
rect 605 565 639 599
rect 605 483 639 517
rect 605 392 639 426
rect 691 573 725 607
rect 691 480 725 514
rect 691 384 725 418
<< poly >>
rect 110 619 140 645
rect 206 619 236 645
rect 304 619 334 645
rect 428 619 458 645
rect 650 619 680 645
rect 110 335 140 367
rect 206 335 236 367
rect 44 319 140 335
rect 44 285 60 319
rect 94 305 140 319
rect 182 319 262 335
rect 94 285 116 305
rect 44 269 116 285
rect 86 241 116 269
rect 182 285 212 319
rect 246 285 262 319
rect 182 269 262 285
rect 304 333 334 367
rect 428 345 458 367
rect 650 345 680 367
rect 304 317 380 333
rect 304 283 320 317
rect 354 283 380 317
rect 428 315 729 345
rect 182 241 212 269
rect 304 267 380 283
rect 304 237 408 267
rect 378 215 408 237
rect 464 215 494 315
rect 650 309 729 315
rect 650 275 679 309
rect 713 275 729 309
rect 650 259 729 275
rect 658 237 688 259
rect 86 47 116 73
rect 182 47 212 73
rect 378 21 408 47
rect 464 21 494 47
rect 658 43 688 69
<< polycont >>
rect 60 285 94 319
rect 212 285 246 319
rect 320 283 354 317
rect 679 275 713 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 40 599 106 615
rect 40 565 65 599
rect 99 565 106 599
rect 40 515 106 565
rect 40 481 65 515
rect 99 510 106 515
rect 359 607 425 649
rect 359 573 375 607
rect 409 573 425 607
rect 359 536 425 573
rect 99 481 325 510
rect 40 462 325 481
rect 40 436 94 462
rect 40 402 60 436
rect 40 386 94 402
rect 128 424 257 428
rect 128 390 151 424
rect 185 390 257 424
rect 128 386 257 390
rect 291 397 325 462
rect 359 502 375 536
rect 409 502 425 536
rect 359 465 425 502
rect 359 431 375 465
rect 409 431 425 465
rect 459 599 519 615
rect 459 565 469 599
rect 503 565 519 599
rect 459 508 519 565
rect 459 474 469 508
rect 503 474 519 508
rect 459 413 519 474
rect 459 397 469 413
rect 17 319 94 352
rect 17 285 60 319
rect 17 269 94 285
rect 128 235 162 386
rect 291 379 469 397
rect 503 379 519 413
rect 291 368 519 379
rect 294 363 519 368
rect 589 599 641 615
rect 589 565 605 599
rect 639 565 641 599
rect 589 517 641 565
rect 589 483 605 517
rect 639 483 641 517
rect 589 426 641 483
rect 589 392 605 426
rect 639 392 641 426
rect 196 319 262 350
rect 196 285 212 319
rect 246 285 262 319
rect 589 317 641 392
rect 675 607 741 649
rect 675 573 691 607
rect 725 573 741 607
rect 675 514 741 573
rect 675 480 691 514
rect 725 480 741 514
rect 675 418 741 480
rect 675 384 691 418
rect 725 384 741 418
rect 304 283 320 317
rect 354 283 641 317
rect 21 219 77 235
rect 21 185 37 219
rect 71 185 77 219
rect 21 119 77 185
rect 111 233 162 235
rect 111 229 177 233
rect 111 195 127 229
rect 161 195 177 229
rect 111 153 177 195
rect 111 119 127 153
rect 161 119 177 153
rect 211 229 555 249
rect 211 195 227 229
rect 261 215 555 229
rect 261 195 277 215
rect 211 153 277 195
rect 498 203 555 215
rect 211 119 227 153
rect 261 119 277 153
rect 317 147 333 181
rect 367 147 383 181
rect 21 85 37 119
rect 71 85 77 119
rect 317 93 383 147
rect 317 85 333 93
rect 21 59 333 85
rect 367 59 383 93
rect 21 51 383 59
rect 417 165 461 181
rect 417 131 419 165
rect 453 131 461 165
rect 417 93 461 131
rect 417 59 419 93
rect 453 59 461 93
rect 417 17 461 59
rect 498 169 505 203
rect 539 169 555 203
rect 498 101 555 169
rect 498 67 505 101
rect 539 67 555 101
rect 597 219 641 283
rect 675 309 751 350
rect 675 275 679 309
rect 713 275 751 309
rect 675 242 751 275
rect 597 203 649 219
rect 597 169 613 203
rect 647 169 649 203
rect 597 122 649 169
rect 597 88 613 122
rect 647 88 649 122
rect 597 72 649 88
rect 683 174 699 208
rect 733 174 749 208
rect 683 115 749 174
rect 683 81 699 115
rect 733 81 749 115
rect 498 51 555 67
rect 683 17 749 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2i_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3839984
string GDS_START 3832892
<< end >>
