magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 70 49 954 241
rect 0 0 960 49
<< scnmos >>
rect 149 47 179 215
rect 235 47 265 215
rect 353 47 383 215
rect 439 47 469 215
rect 565 47 595 215
rect 673 47 703 215
rect 759 47 789 215
rect 845 47 875 215
<< scpmoshvt >>
rect 102 367 132 619
rect 231 367 261 619
rect 317 367 347 619
rect 493 367 523 619
rect 579 367 609 619
rect 673 367 703 619
rect 759 367 789 619
rect 845 367 875 619
<< ndiff >>
rect 96 203 149 215
rect 96 169 104 203
rect 138 169 149 203
rect 96 101 149 169
rect 96 67 104 101
rect 138 67 149 101
rect 96 47 149 67
rect 179 159 235 215
rect 179 125 190 159
rect 224 125 235 159
rect 179 91 235 125
rect 179 57 190 91
rect 224 57 235 91
rect 179 47 235 57
rect 265 89 353 215
rect 265 55 292 89
rect 326 55 353 89
rect 265 47 353 55
rect 383 159 439 215
rect 383 125 394 159
rect 428 125 439 159
rect 383 91 439 125
rect 383 57 394 91
rect 428 57 439 91
rect 383 47 439 57
rect 469 203 565 215
rect 469 169 498 203
rect 532 169 565 203
rect 469 99 565 169
rect 469 65 498 99
rect 532 65 565 99
rect 469 47 565 65
rect 595 159 673 215
rect 595 125 612 159
rect 646 125 673 159
rect 595 91 673 125
rect 595 57 612 91
rect 646 57 673 91
rect 595 47 673 57
rect 703 96 759 215
rect 703 62 714 96
rect 748 62 759 96
rect 703 47 759 62
rect 789 151 845 215
rect 789 117 800 151
rect 834 117 845 151
rect 789 47 845 117
rect 875 203 928 215
rect 875 169 886 203
rect 920 169 928 203
rect 875 101 928 169
rect 875 67 886 101
rect 920 67 928 101
rect 875 47 928 67
<< pdiff >>
rect 420 630 478 638
rect 420 619 432 630
rect 49 599 102 619
rect 49 565 57 599
rect 91 565 102 599
rect 49 508 102 565
rect 49 474 57 508
rect 91 474 102 508
rect 49 421 102 474
rect 49 387 57 421
rect 91 387 102 421
rect 49 367 102 387
rect 132 568 231 619
rect 132 534 166 568
rect 200 534 231 568
rect 132 367 231 534
rect 261 599 317 619
rect 261 565 272 599
rect 306 565 317 599
rect 261 492 317 565
rect 261 458 272 492
rect 306 458 317 492
rect 261 367 317 458
rect 347 596 432 619
rect 466 619 478 630
rect 466 596 493 619
rect 347 568 493 596
rect 347 534 358 568
rect 392 534 493 568
rect 347 367 493 534
rect 523 571 579 619
rect 523 537 534 571
rect 568 537 579 571
rect 523 367 579 537
rect 609 487 673 619
rect 609 453 628 487
rect 662 453 673 487
rect 609 367 673 453
rect 703 596 759 619
rect 703 562 714 596
rect 748 562 759 596
rect 703 367 759 562
rect 789 503 845 619
rect 789 469 800 503
rect 834 469 845 503
rect 789 367 845 469
rect 875 599 928 619
rect 875 565 886 599
rect 920 565 928 599
rect 875 516 928 565
rect 875 482 886 516
rect 920 482 928 516
rect 875 448 928 482
rect 875 414 886 448
rect 920 414 928 448
rect 875 367 928 414
<< ndiffc >>
rect 104 169 138 203
rect 104 67 138 101
rect 190 125 224 159
rect 190 57 224 91
rect 292 55 326 89
rect 394 125 428 159
rect 394 57 428 91
rect 498 169 532 203
rect 498 65 532 99
rect 612 125 646 159
rect 612 57 646 91
rect 714 62 748 96
rect 800 117 834 151
rect 886 169 920 203
rect 886 67 920 101
<< pdiffc >>
rect 57 565 91 599
rect 57 474 91 508
rect 57 387 91 421
rect 166 534 200 568
rect 272 565 306 599
rect 272 458 306 492
rect 432 596 466 630
rect 358 534 392 568
rect 534 537 568 571
rect 628 453 662 487
rect 714 562 748 596
rect 800 469 834 503
rect 886 565 920 599
rect 886 482 920 516
rect 886 414 920 448
<< poly >>
rect 102 619 132 645
rect 231 619 261 645
rect 317 619 347 645
rect 493 619 523 645
rect 579 619 609 645
rect 673 619 703 645
rect 759 619 789 645
rect 845 619 875 645
rect 102 335 132 367
rect 102 319 179 335
rect 102 285 127 319
rect 161 285 179 319
rect 102 269 179 285
rect 231 299 261 367
rect 317 335 347 367
rect 493 335 523 367
rect 579 335 609 367
rect 673 335 703 367
rect 759 335 789 367
rect 317 319 383 335
rect 317 299 333 319
rect 231 285 333 299
rect 367 285 383 319
rect 231 269 383 285
rect 425 319 523 335
rect 425 285 441 319
rect 475 305 523 319
rect 565 319 631 335
rect 475 285 493 305
rect 425 269 493 285
rect 565 285 581 319
rect 615 285 631 319
rect 565 269 631 285
rect 673 319 789 335
rect 673 285 729 319
rect 763 285 789 319
rect 673 269 789 285
rect 149 215 179 269
rect 235 215 265 269
rect 353 215 383 269
rect 439 215 469 269
rect 565 215 595 269
rect 673 215 703 269
rect 759 215 789 269
rect 845 335 875 367
rect 845 319 911 335
rect 845 285 861 319
rect 895 285 911 319
rect 845 269 911 285
rect 845 215 875 269
rect 149 21 179 47
rect 235 21 265 47
rect 353 21 383 47
rect 439 21 469 47
rect 565 21 595 47
rect 673 21 703 47
rect 759 21 789 47
rect 845 21 875 47
<< polycont >>
rect 127 285 161 319
rect 333 285 367 319
rect 441 285 475 319
rect 581 285 615 319
rect 729 285 763 319
rect 861 285 895 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 41 599 107 615
rect 41 565 57 599
rect 91 565 107 599
rect 41 508 107 565
rect 150 568 216 649
rect 342 630 482 649
rect 150 534 166 568
rect 200 534 216 568
rect 150 526 216 534
rect 256 599 308 615
rect 256 565 272 599
rect 306 565 308 599
rect 41 474 57 508
rect 91 492 107 508
rect 256 492 308 565
rect 342 596 432 630
rect 466 596 482 630
rect 342 589 482 596
rect 518 599 936 615
rect 518 596 886 599
rect 342 568 408 589
rect 342 534 358 568
rect 392 534 408 568
rect 518 571 714 596
rect 518 555 534 571
rect 342 526 408 534
rect 442 537 534 555
rect 568 562 714 571
rect 748 565 886 596
rect 920 565 936 599
rect 748 562 936 565
rect 568 553 936 562
rect 568 537 745 553
rect 442 521 745 537
rect 442 492 476 521
rect 91 474 272 492
rect 41 458 272 474
rect 306 458 476 492
rect 784 503 848 519
rect 784 487 800 503
rect 41 421 91 458
rect 510 453 628 487
rect 662 469 800 487
rect 834 469 848 503
rect 662 453 848 469
rect 882 516 936 553
rect 882 482 886 516
rect 920 482 936 516
rect 41 387 57 421
rect 41 371 91 387
rect 125 390 475 424
rect 125 319 177 390
rect 125 285 127 319
rect 161 285 177 319
rect 125 269 177 285
rect 211 319 383 356
rect 211 285 333 319
rect 367 285 383 319
rect 211 269 383 285
rect 425 319 475 390
rect 425 285 441 319
rect 425 269 475 285
rect 510 235 547 453
rect 882 448 936 482
rect 581 385 833 419
rect 882 414 886 448
rect 920 414 936 448
rect 882 398 936 414
rect 581 319 631 385
rect 797 350 833 385
rect 615 285 631 319
rect 581 269 631 285
rect 673 319 763 350
rect 673 285 729 319
rect 673 269 763 285
rect 797 319 911 350
rect 797 285 861 319
rect 895 285 911 319
rect 797 269 911 285
rect 510 233 936 235
rect 88 203 936 233
rect 88 169 104 203
rect 138 199 498 203
rect 88 101 138 169
rect 482 169 498 199
rect 532 201 886 203
rect 532 169 548 201
rect 88 67 104 101
rect 88 51 138 67
rect 174 159 444 165
rect 174 125 190 159
rect 224 131 394 159
rect 224 125 240 131
rect 174 91 240 125
rect 378 125 394 131
rect 428 125 444 159
rect 174 57 190 91
rect 224 57 240 91
rect 174 53 240 57
rect 276 89 342 97
rect 276 55 292 89
rect 326 55 342 89
rect 276 17 342 55
rect 378 91 444 125
rect 378 57 394 91
rect 428 57 444 91
rect 378 53 444 57
rect 482 99 548 169
rect 880 169 886 201
rect 920 169 936 203
rect 482 65 498 99
rect 532 65 548 99
rect 482 51 548 65
rect 596 159 846 167
rect 596 125 612 159
rect 646 151 846 159
rect 646 133 800 151
rect 646 125 664 133
rect 596 91 664 125
rect 798 117 800 133
rect 834 117 846 151
rect 798 101 846 117
rect 880 101 936 169
rect 596 57 612 91
rect 646 57 664 91
rect 596 51 664 57
rect 698 96 764 99
rect 698 62 714 96
rect 748 62 764 96
rect 698 17 764 62
rect 880 67 886 101
rect 920 67 936 101
rect 880 51 936 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a22oi_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 383438
string GDS_START 375300
<< end >>
