magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 17 241 473 263
rect 17 49 1114 241
rect 0 0 1152 49
<< scnmos >>
rect 96 69 126 237
rect 182 69 212 237
rect 268 69 298 237
rect 354 69 384 237
rect 575 47 605 215
rect 661 47 691 215
rect 747 47 777 215
rect 833 47 863 215
rect 919 47 949 215
rect 1005 47 1035 215
<< scpmoshvt >>
rect 96 367 126 619
rect 182 367 212 619
rect 268 367 298 619
rect 354 367 384 619
rect 440 367 470 619
rect 526 367 556 619
rect 747 367 777 619
rect 833 367 863 619
rect 919 367 949 619
rect 1005 367 1035 619
<< ndiff >>
rect 43 192 96 237
rect 43 158 51 192
rect 85 158 96 192
rect 43 115 96 158
rect 43 81 51 115
rect 85 81 96 115
rect 43 69 96 81
rect 126 229 182 237
rect 126 195 137 229
rect 171 195 182 229
rect 126 153 182 195
rect 126 119 137 153
rect 171 119 182 153
rect 126 69 182 119
rect 212 192 268 237
rect 212 158 223 192
rect 257 158 268 192
rect 212 115 268 158
rect 212 81 223 115
rect 257 81 268 115
rect 212 69 268 81
rect 298 124 354 237
rect 298 90 309 124
rect 343 90 354 124
rect 298 69 354 90
rect 384 225 447 237
rect 384 191 405 225
rect 439 191 447 225
rect 384 153 447 191
rect 384 119 405 153
rect 439 119 447 153
rect 384 69 447 119
rect 522 193 575 215
rect 522 159 530 193
rect 564 159 575 193
rect 522 47 575 159
rect 605 113 661 215
rect 605 79 616 113
rect 650 79 661 113
rect 605 47 661 79
rect 691 203 747 215
rect 691 169 702 203
rect 736 169 747 203
rect 691 101 747 169
rect 691 67 702 101
rect 736 67 747 101
rect 691 47 747 67
rect 777 127 833 215
rect 777 93 788 127
rect 822 93 833 127
rect 777 47 833 93
rect 863 203 919 215
rect 863 169 874 203
rect 908 169 919 203
rect 863 101 919 169
rect 863 67 874 101
rect 908 67 919 101
rect 863 47 919 67
rect 949 127 1005 215
rect 949 93 960 127
rect 994 93 1005 127
rect 949 47 1005 93
rect 1035 203 1088 215
rect 1035 169 1046 203
rect 1080 169 1088 203
rect 1035 101 1088 169
rect 1035 67 1046 101
rect 1080 67 1088 101
rect 1035 47 1088 67
<< pdiff >>
rect 43 607 96 619
rect 43 573 51 607
rect 85 573 96 607
rect 43 518 96 573
rect 43 484 51 518
rect 85 484 96 518
rect 43 435 96 484
rect 43 401 51 435
rect 85 401 96 435
rect 43 367 96 401
rect 126 599 182 619
rect 126 565 137 599
rect 171 565 182 599
rect 126 506 182 565
rect 126 472 137 506
rect 171 472 182 506
rect 126 413 182 472
rect 126 379 137 413
rect 171 379 182 413
rect 126 367 182 379
rect 212 607 268 619
rect 212 573 223 607
rect 257 573 268 607
rect 212 531 268 573
rect 212 497 223 531
rect 257 497 268 531
rect 212 453 268 497
rect 212 419 223 453
rect 257 419 268 453
rect 212 367 268 419
rect 298 599 354 619
rect 298 565 309 599
rect 343 565 354 599
rect 298 508 354 565
rect 298 474 309 508
rect 343 474 354 508
rect 298 413 354 474
rect 298 379 309 413
rect 343 379 354 413
rect 298 367 354 379
rect 384 607 440 619
rect 384 573 395 607
rect 429 573 440 607
rect 384 531 440 573
rect 384 497 395 531
rect 429 497 440 531
rect 384 453 440 497
rect 384 419 395 453
rect 429 419 440 453
rect 384 367 440 419
rect 470 599 526 619
rect 470 565 481 599
rect 515 565 526 599
rect 470 508 526 565
rect 470 474 481 508
rect 515 474 526 508
rect 470 413 526 474
rect 470 379 481 413
rect 515 379 526 413
rect 470 367 526 379
rect 556 607 609 619
rect 556 573 567 607
rect 601 573 609 607
rect 556 527 609 573
rect 556 493 567 527
rect 601 493 609 527
rect 556 439 609 493
rect 556 405 567 439
rect 601 405 609 439
rect 556 367 609 405
rect 694 599 747 619
rect 694 565 702 599
rect 736 565 747 599
rect 694 529 747 565
rect 694 495 702 529
rect 736 495 747 529
rect 694 455 747 495
rect 694 421 702 455
rect 736 421 747 455
rect 694 367 747 421
rect 777 547 833 619
rect 777 513 788 547
rect 822 513 833 547
rect 777 479 833 513
rect 777 445 788 479
rect 822 445 833 479
rect 777 411 833 445
rect 777 377 788 411
rect 822 377 833 411
rect 777 367 833 377
rect 863 599 919 619
rect 863 565 874 599
rect 908 565 919 599
rect 863 502 919 565
rect 863 468 874 502
rect 908 468 919 502
rect 863 413 919 468
rect 863 379 874 413
rect 908 379 919 413
rect 863 367 919 379
rect 949 607 1005 619
rect 949 573 960 607
rect 994 573 1005 607
rect 949 514 1005 573
rect 949 480 960 514
rect 994 480 1005 514
rect 949 423 1005 480
rect 949 389 960 423
rect 994 389 1005 423
rect 949 367 1005 389
rect 1035 599 1088 619
rect 1035 565 1046 599
rect 1080 565 1088 599
rect 1035 502 1088 565
rect 1035 468 1046 502
rect 1080 468 1088 502
rect 1035 413 1088 468
rect 1035 379 1046 413
rect 1080 379 1088 413
rect 1035 367 1088 379
<< ndiffc >>
rect 51 158 85 192
rect 51 81 85 115
rect 137 195 171 229
rect 137 119 171 153
rect 223 158 257 192
rect 223 81 257 115
rect 309 90 343 124
rect 405 191 439 225
rect 405 119 439 153
rect 530 159 564 193
rect 616 79 650 113
rect 702 169 736 203
rect 702 67 736 101
rect 788 93 822 127
rect 874 169 908 203
rect 874 67 908 101
rect 960 93 994 127
rect 1046 169 1080 203
rect 1046 67 1080 101
<< pdiffc >>
rect 51 573 85 607
rect 51 484 85 518
rect 51 401 85 435
rect 137 565 171 599
rect 137 472 171 506
rect 137 379 171 413
rect 223 573 257 607
rect 223 497 257 531
rect 223 419 257 453
rect 309 565 343 599
rect 309 474 343 508
rect 309 379 343 413
rect 395 573 429 607
rect 395 497 429 531
rect 395 419 429 453
rect 481 565 515 599
rect 481 474 515 508
rect 481 379 515 413
rect 567 573 601 607
rect 567 493 601 527
rect 567 405 601 439
rect 702 565 736 599
rect 702 495 736 529
rect 702 421 736 455
rect 788 513 822 547
rect 788 445 822 479
rect 788 377 822 411
rect 874 565 908 599
rect 874 468 908 502
rect 874 379 908 413
rect 960 573 994 607
rect 960 480 994 514
rect 960 389 994 423
rect 1046 565 1080 599
rect 1046 468 1080 502
rect 1046 379 1080 413
<< poly >>
rect 96 619 126 645
rect 182 619 212 645
rect 268 619 298 645
rect 354 619 384 645
rect 440 619 470 645
rect 526 619 556 645
rect 747 619 777 645
rect 833 619 863 645
rect 919 619 949 645
rect 1005 619 1035 645
rect 96 325 126 367
rect 182 325 212 367
rect 268 325 298 367
rect 354 325 384 367
rect 35 309 212 325
rect 35 275 51 309
rect 85 275 212 309
rect 35 259 212 275
rect 254 309 398 325
rect 254 275 270 309
rect 304 275 348 309
rect 382 275 398 309
rect 254 259 398 275
rect 440 303 470 367
rect 526 303 556 367
rect 747 303 777 367
rect 833 303 863 367
rect 440 287 691 303
rect 440 273 505 287
rect 96 237 126 259
rect 182 237 212 259
rect 268 237 298 259
rect 354 237 384 259
rect 474 253 505 273
rect 539 253 573 287
rect 607 253 641 287
rect 675 253 691 287
rect 474 237 691 253
rect 575 215 605 237
rect 661 215 691 237
rect 747 287 863 303
rect 747 253 789 287
rect 823 253 863 287
rect 747 237 863 253
rect 747 215 777 237
rect 833 215 863 237
rect 919 303 949 367
rect 1005 303 1035 367
rect 919 287 1035 303
rect 919 253 985 287
rect 1019 253 1035 287
rect 919 237 1035 253
rect 919 215 949 237
rect 1005 215 1035 237
rect 96 43 126 69
rect 182 43 212 69
rect 268 43 298 69
rect 354 43 384 69
rect 575 21 605 47
rect 661 21 691 47
rect 747 21 777 47
rect 833 21 863 47
rect 919 21 949 47
rect 1005 21 1035 47
<< polycont >>
rect 51 275 85 309
rect 270 275 304 309
rect 348 275 382 309
rect 505 253 539 287
rect 573 253 607 287
rect 641 253 675 287
rect 789 253 823 287
rect 985 253 1019 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 35 607 85 649
rect 35 573 51 607
rect 35 518 85 573
rect 35 484 51 518
rect 35 435 85 484
rect 35 401 51 435
rect 35 385 85 401
rect 119 599 173 615
rect 119 565 137 599
rect 171 565 173 599
rect 119 506 173 565
rect 119 472 137 506
rect 171 472 173 506
rect 119 413 173 472
rect 207 607 273 649
rect 207 573 223 607
rect 257 573 273 607
rect 207 531 273 573
rect 207 497 223 531
rect 257 497 273 531
rect 207 453 273 497
rect 207 419 223 453
rect 257 419 273 453
rect 307 599 345 615
rect 307 565 309 599
rect 343 565 345 599
rect 307 508 345 565
rect 307 474 309 508
rect 343 474 345 508
rect 119 379 137 413
rect 171 385 173 413
rect 307 413 345 474
rect 379 607 445 649
rect 379 573 395 607
rect 429 573 445 607
rect 379 531 445 573
rect 379 497 395 531
rect 429 497 445 531
rect 379 453 445 497
rect 379 419 395 453
rect 429 419 445 453
rect 479 599 515 615
rect 479 565 481 599
rect 479 508 515 565
rect 479 474 481 508
rect 307 385 309 413
rect 171 379 309 385
rect 343 385 345 413
rect 479 413 515 474
rect 479 385 481 413
rect 343 379 481 385
rect 551 607 617 649
rect 551 573 567 607
rect 601 573 617 607
rect 551 527 617 573
rect 551 493 567 527
rect 601 493 617 527
rect 551 439 617 493
rect 551 405 567 439
rect 601 405 617 439
rect 686 599 910 615
rect 686 565 702 599
rect 736 581 874 599
rect 736 565 738 581
rect 686 529 738 565
rect 872 565 874 581
rect 908 565 910 599
rect 686 495 702 529
rect 736 495 738 529
rect 686 455 738 495
rect 686 421 702 455
rect 736 421 738 455
rect 686 405 738 421
rect 772 513 788 547
rect 822 513 838 547
rect 772 479 838 513
rect 772 445 788 479
rect 822 445 838 479
rect 772 411 838 445
rect 119 371 515 379
rect 772 377 788 411
rect 822 377 838 411
rect 772 371 838 377
rect 119 351 838 371
rect 17 309 85 350
rect 17 275 51 309
rect 17 242 85 275
rect 119 233 187 351
rect 477 337 838 351
rect 872 502 910 565
rect 872 468 874 502
rect 908 468 910 502
rect 872 413 910 468
rect 872 379 874 413
rect 908 379 910 413
rect 944 607 1010 649
rect 944 573 960 607
rect 994 573 1010 607
rect 944 514 1010 573
rect 944 480 960 514
rect 994 480 1010 514
rect 944 423 1010 480
rect 944 389 960 423
rect 994 389 1010 423
rect 1044 599 1096 615
rect 1044 565 1046 599
rect 1080 565 1096 599
rect 1044 502 1096 565
rect 1044 468 1046 502
rect 1080 468 1096 502
rect 1044 413 1096 468
rect 872 355 910 379
rect 1044 379 1046 413
rect 1080 379 1096 413
rect 1044 355 1096 379
rect 872 321 1096 355
rect 221 275 270 309
rect 304 275 348 309
rect 382 275 398 309
rect 489 287 739 303
rect 221 242 355 275
rect 489 253 505 287
rect 539 253 573 287
rect 607 253 641 287
rect 675 253 739 287
rect 121 229 187 233
rect 35 192 87 208
rect 35 158 51 192
rect 85 158 87 192
rect 35 115 87 158
rect 121 195 137 229
rect 171 195 187 229
rect 389 225 455 241
rect 489 237 739 253
rect 773 253 789 287
rect 823 253 935 287
rect 773 237 935 253
rect 969 253 985 287
rect 1019 253 1135 287
rect 969 237 1135 253
rect 389 208 405 225
rect 121 153 187 195
rect 121 119 137 153
rect 171 119 187 153
rect 223 192 405 208
rect 257 191 405 192
rect 439 191 455 225
rect 257 174 455 191
rect 257 158 267 174
rect 35 81 51 115
rect 85 85 87 115
rect 223 115 267 158
rect 389 153 455 174
rect 514 193 702 203
rect 514 159 530 193
rect 564 169 702 193
rect 736 169 874 203
rect 908 169 1046 203
rect 1080 169 1096 203
rect 564 159 738 169
rect 514 155 738 159
rect 85 81 223 85
rect 257 81 267 115
rect 35 51 267 81
rect 301 124 355 140
rect 301 90 309 124
rect 343 90 355 124
rect 389 119 405 153
rect 439 119 455 153
rect 301 85 355 90
rect 600 113 666 121
rect 600 85 616 113
rect 301 79 616 85
rect 650 79 666 113
rect 301 51 666 79
rect 700 101 738 155
rect 700 67 702 101
rect 736 67 738 101
rect 700 51 738 67
rect 772 127 838 135
rect 772 93 788 127
rect 822 93 838 127
rect 772 17 838 93
rect 872 101 910 169
rect 872 67 874 101
rect 908 67 910 101
rect 872 51 910 67
rect 944 127 1010 135
rect 944 93 960 127
rect 994 93 1010 127
rect 944 17 1010 93
rect 1044 101 1096 169
rect 1044 67 1046 101
rect 1080 67 1096 101
rect 1044 51 1096 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2111ai_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4758838
string GDS_START 4747920
<< end >>
