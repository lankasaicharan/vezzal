magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 1 49 1531 259
rect 0 0 1536 49
<< scnmos >>
rect 80 65 110 233
rect 166 65 196 233
rect 252 65 282 233
rect 338 65 368 233
rect 424 65 454 233
rect 510 65 540 233
rect 596 65 626 233
rect 682 65 712 233
rect 768 65 798 233
rect 854 65 884 233
rect 954 65 984 233
rect 1054 65 1084 233
rect 1154 65 1184 233
rect 1246 65 1276 233
rect 1332 65 1362 233
rect 1418 65 1448 233
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 252 367 282 619
rect 338 367 368 619
rect 424 367 454 619
rect 510 367 540 619
rect 596 367 626 619
rect 682 367 712 619
rect 768 367 798 619
rect 854 367 884 619
rect 954 367 984 619
rect 1054 367 1084 619
rect 1154 367 1184 619
rect 1246 367 1276 619
rect 1332 367 1362 619
rect 1418 367 1448 619
<< ndiff >>
rect 27 221 80 233
rect 27 187 35 221
rect 69 187 80 221
rect 27 111 80 187
rect 27 77 35 111
rect 69 77 80 111
rect 27 65 80 77
rect 110 181 166 233
rect 110 147 121 181
rect 155 147 166 181
rect 110 111 166 147
rect 110 77 121 111
rect 155 77 166 111
rect 110 65 166 77
rect 196 221 252 233
rect 196 187 207 221
rect 241 187 252 221
rect 196 111 252 187
rect 196 77 207 111
rect 241 77 252 111
rect 196 65 252 77
rect 282 181 338 233
rect 282 147 293 181
rect 327 147 338 181
rect 282 107 338 147
rect 282 73 293 107
rect 327 73 338 107
rect 282 65 338 73
rect 368 221 424 233
rect 368 187 379 221
rect 413 187 424 221
rect 368 111 424 187
rect 368 77 379 111
rect 413 77 424 111
rect 368 65 424 77
rect 454 181 510 233
rect 454 147 465 181
rect 499 147 510 181
rect 454 107 510 147
rect 454 73 465 107
rect 499 73 510 107
rect 454 65 510 73
rect 540 221 596 233
rect 540 187 551 221
rect 585 187 596 221
rect 540 111 596 187
rect 540 77 551 111
rect 585 77 596 111
rect 540 65 596 77
rect 626 181 682 233
rect 626 147 637 181
rect 671 147 682 181
rect 626 107 682 147
rect 626 73 637 107
rect 671 73 682 107
rect 626 65 682 73
rect 712 221 768 233
rect 712 187 723 221
rect 757 187 768 221
rect 712 111 768 187
rect 712 77 723 111
rect 757 77 768 111
rect 712 65 768 77
rect 798 225 854 233
rect 798 191 809 225
rect 843 191 854 225
rect 798 157 854 191
rect 798 123 809 157
rect 843 123 854 157
rect 798 65 854 123
rect 884 183 954 233
rect 884 149 909 183
rect 943 149 954 183
rect 884 107 954 149
rect 884 73 909 107
rect 943 73 954 107
rect 884 65 954 73
rect 984 225 1054 233
rect 984 191 1009 225
rect 1043 191 1054 225
rect 984 157 1054 191
rect 984 123 1009 157
rect 1043 123 1054 157
rect 984 65 1054 123
rect 1084 181 1154 233
rect 1084 147 1109 181
rect 1143 147 1154 181
rect 1084 107 1154 147
rect 1084 73 1109 107
rect 1143 73 1154 107
rect 1084 65 1154 73
rect 1184 178 1246 233
rect 1184 144 1201 178
rect 1235 144 1246 178
rect 1184 65 1246 144
rect 1276 181 1332 233
rect 1276 147 1287 181
rect 1321 147 1332 181
rect 1276 107 1332 147
rect 1276 73 1287 107
rect 1321 73 1332 107
rect 1276 65 1332 73
rect 1362 225 1418 233
rect 1362 191 1373 225
rect 1407 191 1418 225
rect 1362 157 1418 191
rect 1362 123 1373 157
rect 1407 123 1418 157
rect 1362 65 1418 123
rect 1448 221 1505 233
rect 1448 187 1459 221
rect 1493 187 1505 221
rect 1448 111 1505 187
rect 1448 77 1459 111
rect 1493 77 1505 111
rect 1448 65 1505 77
<< pdiff >>
rect 27 607 80 619
rect 27 573 35 607
rect 69 573 80 607
rect 27 509 80 573
rect 27 475 35 509
rect 69 475 80 509
rect 27 414 80 475
rect 27 380 35 414
rect 69 380 80 414
rect 27 367 80 380
rect 110 599 166 619
rect 110 565 121 599
rect 155 565 166 599
rect 110 509 166 565
rect 110 475 121 509
rect 155 475 166 509
rect 110 413 166 475
rect 110 379 121 413
rect 155 379 166 413
rect 110 367 166 379
rect 196 607 252 619
rect 196 573 207 607
rect 241 573 252 607
rect 196 533 252 573
rect 196 499 207 533
rect 241 499 252 533
rect 196 455 252 499
rect 196 421 207 455
rect 241 421 252 455
rect 196 367 252 421
rect 282 599 338 619
rect 282 565 293 599
rect 327 565 338 599
rect 282 509 338 565
rect 282 475 293 509
rect 327 475 338 509
rect 282 413 338 475
rect 282 379 293 413
rect 327 379 338 413
rect 282 367 338 379
rect 368 607 424 619
rect 368 573 379 607
rect 413 573 424 607
rect 368 488 424 573
rect 368 454 379 488
rect 413 454 424 488
rect 368 367 424 454
rect 454 599 510 619
rect 454 565 465 599
rect 499 565 510 599
rect 454 517 510 565
rect 454 483 465 517
rect 499 483 510 517
rect 454 436 510 483
rect 454 402 465 436
rect 499 402 510 436
rect 454 367 510 402
rect 540 607 596 619
rect 540 573 551 607
rect 585 573 596 607
rect 540 488 596 573
rect 540 454 551 488
rect 585 454 596 488
rect 540 367 596 454
rect 626 599 682 619
rect 626 565 637 599
rect 671 565 682 599
rect 626 509 682 565
rect 626 475 637 509
rect 671 475 682 509
rect 626 413 682 475
rect 626 379 637 413
rect 671 379 682 413
rect 626 367 682 379
rect 712 611 768 619
rect 712 577 723 611
rect 757 577 768 611
rect 712 543 768 577
rect 712 509 723 543
rect 757 509 768 543
rect 712 457 768 509
rect 712 423 723 457
rect 757 423 768 457
rect 712 367 768 423
rect 798 599 854 619
rect 798 565 809 599
rect 843 565 854 599
rect 798 509 854 565
rect 798 475 809 509
rect 843 475 854 509
rect 798 413 854 475
rect 798 379 809 413
rect 843 379 854 413
rect 798 367 854 379
rect 884 607 954 619
rect 884 573 902 607
rect 936 573 954 607
rect 884 488 954 573
rect 884 454 902 488
rect 936 454 954 488
rect 884 367 954 454
rect 984 599 1054 619
rect 984 565 1002 599
rect 1036 565 1054 599
rect 984 519 1054 565
rect 984 485 1002 519
rect 1036 485 1054 519
rect 984 436 1054 485
rect 984 402 1002 436
rect 1036 402 1054 436
rect 984 367 1054 402
rect 1084 607 1154 619
rect 1084 573 1102 607
rect 1136 573 1154 607
rect 1084 488 1154 573
rect 1084 454 1102 488
rect 1136 454 1154 488
rect 1084 367 1154 454
rect 1184 599 1246 619
rect 1184 565 1201 599
rect 1235 565 1246 599
rect 1184 508 1246 565
rect 1184 474 1201 508
rect 1235 474 1246 508
rect 1184 413 1246 474
rect 1184 379 1201 413
rect 1235 379 1246 413
rect 1184 367 1246 379
rect 1276 607 1332 619
rect 1276 573 1287 607
rect 1321 573 1332 607
rect 1276 537 1332 573
rect 1276 503 1287 537
rect 1321 503 1332 537
rect 1276 453 1332 503
rect 1276 419 1287 453
rect 1321 419 1332 453
rect 1276 367 1332 419
rect 1362 599 1418 619
rect 1362 565 1373 599
rect 1407 565 1418 599
rect 1362 508 1418 565
rect 1362 474 1373 508
rect 1407 474 1418 508
rect 1362 413 1418 474
rect 1362 379 1373 413
rect 1407 379 1418 413
rect 1362 367 1418 379
rect 1448 607 1501 619
rect 1448 573 1459 607
rect 1493 573 1501 607
rect 1448 508 1501 573
rect 1448 474 1459 508
rect 1493 474 1501 508
rect 1448 413 1501 474
rect 1448 379 1459 413
rect 1493 379 1501 413
rect 1448 367 1501 379
<< ndiffc >>
rect 35 187 69 221
rect 35 77 69 111
rect 121 147 155 181
rect 121 77 155 111
rect 207 187 241 221
rect 207 77 241 111
rect 293 147 327 181
rect 293 73 327 107
rect 379 187 413 221
rect 379 77 413 111
rect 465 147 499 181
rect 465 73 499 107
rect 551 187 585 221
rect 551 77 585 111
rect 637 147 671 181
rect 637 73 671 107
rect 723 187 757 221
rect 723 77 757 111
rect 809 191 843 225
rect 809 123 843 157
rect 909 149 943 183
rect 909 73 943 107
rect 1009 191 1043 225
rect 1009 123 1043 157
rect 1109 147 1143 181
rect 1109 73 1143 107
rect 1201 144 1235 178
rect 1287 147 1321 181
rect 1287 73 1321 107
rect 1373 191 1407 225
rect 1373 123 1407 157
rect 1459 187 1493 221
rect 1459 77 1493 111
<< pdiffc >>
rect 35 573 69 607
rect 35 475 69 509
rect 35 380 69 414
rect 121 565 155 599
rect 121 475 155 509
rect 121 379 155 413
rect 207 573 241 607
rect 207 499 241 533
rect 207 421 241 455
rect 293 565 327 599
rect 293 475 327 509
rect 293 379 327 413
rect 379 573 413 607
rect 379 454 413 488
rect 465 565 499 599
rect 465 483 499 517
rect 465 402 499 436
rect 551 573 585 607
rect 551 454 585 488
rect 637 565 671 599
rect 637 475 671 509
rect 637 379 671 413
rect 723 577 757 611
rect 723 509 757 543
rect 723 423 757 457
rect 809 565 843 599
rect 809 475 843 509
rect 809 379 843 413
rect 902 573 936 607
rect 902 454 936 488
rect 1002 565 1036 599
rect 1002 485 1036 519
rect 1002 402 1036 436
rect 1102 573 1136 607
rect 1102 454 1136 488
rect 1201 565 1235 599
rect 1201 474 1235 508
rect 1201 379 1235 413
rect 1287 573 1321 607
rect 1287 503 1321 537
rect 1287 419 1321 453
rect 1373 565 1407 599
rect 1373 474 1407 508
rect 1373 379 1407 413
rect 1459 573 1493 607
rect 1459 474 1493 508
rect 1459 379 1493 413
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 252 619 282 645
rect 338 619 368 645
rect 424 619 454 645
rect 510 619 540 645
rect 596 619 626 645
rect 682 619 712 645
rect 768 619 798 645
rect 854 619 884 645
rect 954 619 984 645
rect 1054 619 1084 645
rect 1154 619 1184 645
rect 1246 619 1276 645
rect 1332 619 1362 645
rect 1418 619 1448 645
rect 80 335 110 367
rect 166 335 196 367
rect 252 335 282 367
rect 338 335 368 367
rect 424 335 454 367
rect 510 335 540 367
rect 596 335 626 367
rect 682 335 712 367
rect 80 319 712 335
rect 80 285 107 319
rect 141 285 175 319
rect 209 285 243 319
rect 277 285 311 319
rect 345 285 379 319
rect 413 285 447 319
rect 481 285 515 319
rect 549 285 583 319
rect 617 285 651 319
rect 685 285 712 319
rect 80 269 712 285
rect 80 233 110 269
rect 166 233 196 269
rect 252 233 282 269
rect 338 233 368 269
rect 424 233 454 269
rect 510 233 540 269
rect 596 233 626 269
rect 682 233 712 269
rect 768 335 798 367
rect 854 335 884 367
rect 954 335 984 367
rect 1054 335 1084 367
rect 1154 335 1184 367
rect 1246 335 1276 367
rect 1332 335 1362 367
rect 1418 335 1448 367
rect 768 319 1448 335
rect 768 285 902 319
rect 936 285 970 319
rect 1004 285 1038 319
rect 1072 285 1106 319
rect 1140 285 1448 319
rect 768 269 1448 285
rect 768 233 798 269
rect 854 233 884 269
rect 954 233 984 269
rect 1054 233 1084 269
rect 1154 233 1184 269
rect 1246 233 1276 269
rect 1332 233 1362 269
rect 1418 233 1448 269
rect 80 39 110 65
rect 166 39 196 65
rect 252 39 282 65
rect 338 39 368 65
rect 424 39 454 65
rect 510 39 540 65
rect 596 39 626 65
rect 682 39 712 65
rect 768 39 798 65
rect 854 39 884 65
rect 954 39 984 65
rect 1054 39 1084 65
rect 1154 39 1184 65
rect 1246 39 1276 65
rect 1332 39 1362 65
rect 1418 39 1448 65
<< polycont >>
rect 107 285 141 319
rect 175 285 209 319
rect 243 285 277 319
rect 311 285 345 319
rect 379 285 413 319
rect 447 285 481 319
rect 515 285 549 319
rect 583 285 617 319
rect 651 285 685 319
rect 902 285 936 319
rect 970 285 1004 319
rect 1038 285 1072 319
rect 1106 285 1140 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 19 607 85 649
rect 19 573 35 607
rect 69 573 85 607
rect 19 509 85 573
rect 19 475 35 509
rect 69 475 85 509
rect 19 414 85 475
rect 19 380 35 414
rect 69 380 85 414
rect 19 364 85 380
rect 119 599 157 615
rect 119 565 121 599
rect 155 565 157 599
rect 119 509 157 565
rect 119 475 121 509
rect 155 475 157 509
rect 119 413 157 475
rect 191 607 257 649
rect 191 573 207 607
rect 241 573 257 607
rect 191 533 257 573
rect 191 499 207 533
rect 241 499 257 533
rect 191 455 257 499
rect 191 421 207 455
rect 241 421 257 455
rect 291 599 329 615
rect 291 565 293 599
rect 327 565 329 599
rect 291 509 329 565
rect 291 475 293 509
rect 327 475 329 509
rect 119 379 121 413
rect 155 387 157 413
rect 291 420 329 475
rect 363 607 429 649
rect 363 573 379 607
rect 413 573 429 607
rect 363 488 429 573
rect 363 454 379 488
rect 413 454 429 488
rect 463 599 501 615
rect 463 565 465 599
rect 499 565 501 599
rect 463 517 501 565
rect 463 483 465 517
rect 499 483 501 517
rect 463 436 501 483
rect 535 607 601 649
rect 535 573 551 607
rect 585 573 601 607
rect 535 488 601 573
rect 535 454 551 488
rect 585 454 601 488
rect 635 599 673 615
rect 635 565 637 599
rect 671 565 673 599
rect 635 509 673 565
rect 635 475 637 509
rect 671 475 673 509
rect 463 420 465 436
rect 291 413 465 420
rect 291 387 293 413
rect 155 379 293 387
rect 327 402 465 413
rect 499 420 501 436
rect 635 420 673 475
rect 707 611 773 649
rect 707 577 723 611
rect 757 577 773 611
rect 707 543 773 577
rect 707 509 723 543
rect 757 509 773 543
rect 707 457 773 509
rect 707 423 723 457
rect 757 423 773 457
rect 807 599 852 615
rect 807 565 809 599
rect 843 565 852 599
rect 807 509 852 565
rect 807 475 809 509
rect 843 475 852 509
rect 499 413 673 420
rect 499 402 637 413
rect 327 386 637 402
rect 119 353 327 379
rect 625 379 637 386
rect 671 389 673 413
rect 807 420 852 475
rect 886 607 952 649
rect 886 573 902 607
rect 936 573 952 607
rect 886 488 952 573
rect 886 454 902 488
rect 936 454 952 488
rect 986 599 1052 615
rect 986 565 1002 599
rect 1036 565 1052 599
rect 986 519 1052 565
rect 986 485 1002 519
rect 1036 485 1052 519
rect 986 436 1052 485
rect 1086 607 1152 649
rect 1086 573 1102 607
rect 1136 573 1152 607
rect 1086 488 1152 573
rect 1086 454 1102 488
rect 1136 454 1152 488
rect 1190 599 1237 615
rect 1190 565 1201 599
rect 1235 565 1237 599
rect 1190 508 1237 565
rect 1190 474 1201 508
rect 1235 474 1237 508
rect 986 420 1002 436
rect 807 413 1002 420
rect 807 389 809 413
rect 671 379 809 389
rect 843 402 1002 413
rect 1036 420 1052 436
rect 1190 420 1237 474
rect 1036 413 1237 420
rect 1271 607 1337 649
rect 1271 573 1287 607
rect 1321 573 1337 607
rect 1271 537 1337 573
rect 1271 503 1287 537
rect 1321 503 1337 537
rect 1271 453 1337 503
rect 1271 419 1287 453
rect 1321 419 1337 453
rect 1371 599 1411 615
rect 1371 565 1373 599
rect 1407 565 1411 599
rect 1371 508 1411 565
rect 1371 474 1373 508
rect 1407 474 1411 508
rect 1036 402 1201 413
rect 843 386 1201 402
rect 843 379 852 386
rect 625 355 852 379
rect 363 321 565 352
rect 363 319 701 321
rect 91 285 107 319
rect 141 285 175 319
rect 209 285 243 319
rect 277 285 311 319
rect 345 285 379 319
rect 413 285 447 319
rect 481 285 515 319
rect 549 285 583 319
rect 617 285 651 319
rect 685 285 701 319
rect 91 283 701 285
rect 793 251 852 355
rect 1190 379 1201 386
rect 1235 385 1237 413
rect 1371 413 1411 474
rect 1371 385 1373 413
rect 1235 379 1373 385
rect 1407 379 1411 413
rect 886 319 1156 352
rect 886 285 902 319
rect 936 285 970 319
rect 1004 285 1038 319
rect 1072 285 1106 319
rect 1140 285 1156 319
rect 1190 300 1411 379
rect 1455 607 1497 649
rect 1455 573 1459 607
rect 1493 573 1497 607
rect 1455 508 1497 573
rect 1455 474 1459 508
rect 1493 474 1497 508
rect 1455 413 1497 474
rect 1455 379 1459 413
rect 1493 379 1497 413
rect 1455 363 1497 379
rect 1190 251 1423 300
rect 19 221 759 249
rect 19 187 35 221
rect 69 215 207 221
rect 69 187 71 215
rect 19 111 71 187
rect 205 187 207 215
rect 241 215 379 221
rect 19 77 35 111
rect 69 77 71 111
rect 19 61 71 77
rect 105 147 121 181
rect 155 147 171 181
rect 105 111 171 147
rect 105 77 121 111
rect 155 77 171 111
rect 105 17 171 77
rect 205 111 241 187
rect 377 187 379 215
rect 413 215 551 221
rect 413 187 415 215
rect 205 77 207 111
rect 205 61 241 77
rect 277 147 293 181
rect 327 147 343 181
rect 277 107 343 147
rect 277 73 293 107
rect 327 73 343 107
rect 277 17 343 73
rect 377 111 415 187
rect 549 187 551 215
rect 585 215 723 221
rect 585 187 587 215
rect 377 77 379 111
rect 413 77 415 111
rect 377 61 415 77
rect 449 147 465 181
rect 499 147 515 181
rect 449 107 515 147
rect 449 73 465 107
rect 499 73 515 107
rect 449 17 515 73
rect 549 111 587 187
rect 721 187 723 215
rect 757 187 759 221
rect 549 77 551 111
rect 585 77 587 111
rect 549 61 587 77
rect 621 147 637 181
rect 671 147 687 181
rect 621 107 687 147
rect 621 73 637 107
rect 671 73 687 107
rect 621 17 687 73
rect 721 111 759 187
rect 793 231 1423 251
rect 793 225 1244 231
rect 793 191 809 225
rect 843 217 1009 225
rect 843 191 859 217
rect 793 157 859 191
rect 993 191 1009 217
rect 1043 215 1244 225
rect 1043 191 1059 215
rect 793 123 809 157
rect 843 123 859 157
rect 793 119 859 123
rect 893 149 909 183
rect 943 149 959 183
rect 721 77 723 111
rect 757 85 759 111
rect 893 107 959 149
rect 993 157 1059 191
rect 993 123 1009 157
rect 1043 123 1059 157
rect 993 119 1059 123
rect 1093 147 1109 181
rect 1143 147 1159 181
rect 893 85 909 107
rect 757 77 909 85
rect 721 73 909 77
rect 943 85 959 107
rect 1093 107 1159 147
rect 1193 178 1244 215
rect 1357 225 1423 231
rect 1193 144 1201 178
rect 1235 144 1244 178
rect 1193 121 1244 144
rect 1278 181 1323 197
rect 1278 147 1287 181
rect 1321 147 1323 181
rect 1093 85 1109 107
rect 943 73 1109 85
rect 1143 87 1159 107
rect 1278 107 1323 147
rect 1357 191 1373 225
rect 1407 191 1423 225
rect 1357 157 1423 191
rect 1357 123 1373 157
rect 1407 123 1423 157
rect 1357 121 1423 123
rect 1457 221 1509 238
rect 1457 187 1459 221
rect 1493 187 1509 221
rect 1278 87 1287 107
rect 1143 73 1287 87
rect 1321 87 1323 107
rect 1457 111 1509 187
rect 1457 87 1459 111
rect 1321 77 1459 87
rect 1493 77 1509 111
rect 1321 73 1509 77
rect 721 51 1509 73
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2_8
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5807526
string GDS_START 5794664
<< end >>
