magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3230 1852
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 34 201 1523 203
rect 34 23 1926 201
rect 34 21 257 23
rect 784 21 996 23
rect 1438 21 1926 23
rect 34 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 116 47 146 177
rect 246 93 276 177
rect 488 49 518 177
rect 608 49 638 177
rect 890 47 920 177
rect 1086 49 1116 177
rect 1248 49 1278 133
rect 1407 49 1437 177
rect 1546 47 1576 167
rect 1657 47 1687 175
rect 1813 47 1843 175
<< scpmoshvt >>
rect 118 297 154 497
rect 248 297 284 425
rect 472 325 508 493
rect 588 325 624 493
rect 839 297 875 497
rect 1078 297 1114 465
rect 1240 297 1276 425
rect 1425 329 1461 457
rect 1538 329 1574 497
rect 1649 297 1685 497
rect 1805 297 1841 497
<< ndiff >>
rect 60 129 116 177
rect 60 95 68 129
rect 102 95 116 129
rect 60 47 116 95
rect 146 93 246 177
rect 276 169 370 177
rect 276 135 324 169
rect 358 135 370 169
rect 276 93 370 135
rect 424 165 488 177
rect 424 131 434 165
rect 468 131 488 165
rect 146 89 231 93
rect 146 55 178 89
rect 212 55 231 89
rect 146 47 231 55
rect 424 49 488 131
rect 518 91 608 177
rect 518 57 528 91
rect 562 57 608 91
rect 518 49 608 57
rect 638 169 737 177
rect 638 135 690 169
rect 724 135 737 169
rect 638 49 737 135
rect 810 157 890 177
rect 810 123 826 157
rect 860 123 890 157
rect 810 89 890 123
rect 810 55 826 89
rect 860 55 890 89
rect 810 47 890 55
rect 920 161 972 177
rect 920 127 930 161
rect 964 127 972 161
rect 920 121 972 127
rect 920 47 970 121
rect 1026 105 1086 177
rect 1024 97 1086 105
rect 1024 63 1032 97
rect 1066 63 1086 97
rect 1024 49 1086 63
rect 1116 133 1217 177
rect 1303 169 1407 177
rect 1303 135 1349 169
rect 1383 135 1407 169
rect 1303 133 1407 135
rect 1116 126 1248 133
rect 1116 92 1126 126
rect 1160 92 1248 126
rect 1116 49 1248 92
rect 1278 49 1407 133
rect 1437 167 1497 177
rect 1597 167 1657 175
rect 1437 93 1546 167
rect 1437 59 1459 93
rect 1493 59 1546 93
rect 1437 49 1546 59
rect 1464 47 1546 49
rect 1576 142 1657 167
rect 1576 108 1603 142
rect 1637 108 1657 142
rect 1576 47 1657 108
rect 1687 97 1813 175
rect 1687 63 1726 97
rect 1760 63 1813 97
rect 1687 47 1813 63
rect 1843 101 1900 175
rect 1843 67 1853 101
rect 1887 67 1900 101
rect 1843 47 1900 67
<< pdiff >>
rect 60 477 118 497
rect 60 443 72 477
rect 106 443 118 477
rect 60 409 118 443
rect 60 375 72 409
rect 106 375 118 409
rect 60 341 118 375
rect 60 307 72 341
rect 106 307 118 341
rect 60 297 118 307
rect 154 477 231 497
rect 154 443 183 477
rect 217 443 231 477
rect 154 425 231 443
rect 154 297 248 425
rect 284 341 342 425
rect 284 307 296 341
rect 330 307 342 341
rect 406 413 472 493
rect 406 379 426 413
rect 460 379 472 413
rect 406 325 472 379
rect 508 481 588 493
rect 508 447 529 481
rect 563 447 588 481
rect 508 325 588 447
rect 624 481 731 493
rect 624 447 686 481
rect 720 447 731 481
rect 624 325 731 447
rect 785 481 839 497
rect 785 447 793 481
rect 827 447 839 481
rect 284 297 342 307
rect 785 297 839 447
rect 875 349 937 497
rect 1478 489 1538 497
rect 991 405 1078 465
rect 991 371 999 405
rect 1033 371 1078 405
rect 991 365 1078 371
rect 875 343 939 349
rect 875 309 887 343
rect 921 309 939 343
rect 875 297 939 309
rect 993 297 1078 365
rect 1114 425 1216 465
rect 1478 457 1490 489
rect 1338 425 1425 457
rect 1114 409 1240 425
rect 1114 375 1167 409
rect 1201 375 1240 409
rect 1114 341 1240 375
rect 1114 307 1167 341
rect 1201 307 1240 341
rect 1114 297 1240 307
rect 1276 421 1425 425
rect 1276 387 1379 421
rect 1413 387 1425 421
rect 1276 329 1425 387
rect 1461 455 1490 457
rect 1524 455 1538 489
rect 1461 329 1538 455
rect 1574 341 1649 497
rect 1574 329 1603 341
rect 1276 297 1373 329
rect 1591 307 1603 329
rect 1637 307 1649 341
rect 1591 297 1649 307
rect 1685 489 1805 497
rect 1685 455 1728 489
rect 1762 455 1805 489
rect 1685 297 1805 455
rect 1841 477 1900 497
rect 1841 443 1854 477
rect 1888 443 1900 477
rect 1841 409 1900 443
rect 1841 375 1854 409
rect 1888 375 1900 409
rect 1841 297 1900 375
<< ndiffc >>
rect 68 95 102 129
rect 324 135 358 169
rect 434 131 468 165
rect 178 55 212 89
rect 528 57 562 91
rect 690 135 724 169
rect 826 123 860 157
rect 826 55 860 89
rect 930 127 964 161
rect 1032 63 1066 97
rect 1349 135 1383 169
rect 1126 92 1160 126
rect 1459 59 1493 93
rect 1603 108 1637 142
rect 1726 63 1760 97
rect 1853 67 1887 101
<< pdiffc >>
rect 72 443 106 477
rect 72 375 106 409
rect 72 307 106 341
rect 183 443 217 477
rect 296 307 330 341
rect 426 379 460 413
rect 529 447 563 481
rect 686 447 720 481
rect 793 447 827 481
rect 999 371 1033 405
rect 887 309 921 343
rect 1167 375 1201 409
rect 1167 307 1201 341
rect 1379 387 1413 421
rect 1490 455 1524 489
rect 1603 307 1637 341
rect 1728 455 1762 489
rect 1854 443 1888 477
rect 1854 375 1888 409
<< poly >>
rect 118 497 154 523
rect 472 493 508 519
rect 588 493 624 519
rect 839 497 875 523
rect 246 451 286 483
rect 248 425 284 451
rect 472 310 508 325
rect 588 310 624 325
rect 118 282 154 297
rect 248 282 284 297
rect 116 265 156 282
rect 246 265 286 282
rect 470 271 510 310
rect 470 265 519 271
rect 586 265 626 310
rect 1076 493 1463 523
rect 1538 497 1574 523
rect 1649 497 1685 523
rect 1805 497 1841 523
rect 1076 491 1116 493
rect 1078 465 1114 491
rect 1423 483 1463 493
rect 1425 457 1461 483
rect 1240 425 1276 451
rect 1425 314 1461 329
rect 1538 314 1574 329
rect 839 282 875 297
rect 1078 282 1114 297
rect 1240 282 1276 297
rect 116 249 204 265
rect 116 215 160 249
rect 194 215 204 249
rect 116 199 204 215
rect 246 249 519 265
rect 246 215 397 249
rect 431 215 465 249
rect 499 215 519 249
rect 246 199 519 215
rect 574 249 638 265
rect 574 215 584 249
rect 618 215 638 249
rect 837 247 877 282
rect 1076 247 1116 282
rect 1238 265 1278 282
rect 1423 265 1463 314
rect 837 217 1116 247
rect 574 199 638 215
rect 116 177 146 199
rect 246 177 276 199
rect 488 197 519 199
rect 488 177 518 197
rect 608 177 638 199
rect 890 177 920 217
rect 1086 177 1116 217
rect 1158 249 1278 265
rect 1158 215 1168 249
rect 1202 215 1278 249
rect 1158 199 1278 215
rect 246 67 276 93
rect 116 21 146 47
rect 488 21 518 49
rect 608 21 638 49
rect 1248 133 1278 199
rect 1407 249 1471 265
rect 1536 255 1576 314
rect 1649 282 1685 297
rect 1805 282 1841 297
rect 1647 265 1687 282
rect 1803 265 1843 282
rect 1407 215 1417 249
rect 1451 215 1471 249
rect 1407 199 1471 215
rect 1513 239 1576 255
rect 1513 205 1523 239
rect 1557 205 1576 239
rect 1407 177 1437 199
rect 1513 189 1576 205
rect 1619 249 1687 265
rect 1619 215 1629 249
rect 1663 215 1687 249
rect 1619 199 1687 215
rect 1791 249 1855 265
rect 1791 215 1801 249
rect 1835 215 1855 249
rect 1791 199 1855 215
rect 1546 167 1576 189
rect 1657 175 1687 199
rect 1813 175 1843 199
rect 890 21 920 47
rect 1086 21 1116 49
rect 1248 23 1278 49
rect 1407 21 1437 49
rect 1546 21 1576 47
rect 1657 21 1687 47
rect 1813 21 1843 47
<< polycont >>
rect 160 215 194 249
rect 397 215 431 249
rect 465 215 499 249
rect 584 215 618 249
rect 1168 215 1202 249
rect 1417 215 1451 249
rect 1523 205 1557 239
rect 1629 215 1663 249
rect 1801 215 1835 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 17 477 122 493
rect 17 443 72 477
rect 106 443 122 477
rect 166 477 233 527
rect 777 481 843 527
rect 1671 489 1810 527
rect 166 443 183 477
rect 217 443 233 477
rect 270 447 529 481
rect 563 447 609 481
rect 662 447 686 481
rect 720 447 743 481
rect 777 447 793 481
rect 827 447 843 481
rect 930 455 1490 489
rect 1524 455 1589 489
rect 1671 455 1728 489
rect 1762 455 1810 489
rect 1854 477 1913 493
rect 17 409 122 443
rect 270 409 314 447
rect 709 413 743 447
rect 930 413 964 455
rect 17 375 72 409
rect 106 375 122 409
rect 17 341 122 375
rect 17 307 72 341
rect 106 307 122 341
rect 17 288 122 307
rect 160 375 314 409
rect 394 379 426 413
rect 460 379 675 413
rect 709 379 964 413
rect 999 405 1033 421
rect 17 185 80 288
rect 160 249 200 375
rect 247 307 296 341
rect 330 307 597 341
rect 194 215 200 249
rect 17 129 118 185
rect 160 173 200 215
rect 160 139 290 173
rect 17 95 68 129
rect 102 95 118 129
rect 17 70 118 95
rect 162 89 212 105
rect 162 55 178 89
rect 162 17 212 55
rect 246 85 290 139
rect 324 169 358 307
rect 563 265 597 307
rect 641 339 675 379
rect 641 323 747 339
rect 641 305 713 323
rect 690 289 713 305
rect 690 275 747 289
rect 392 249 529 265
rect 392 215 397 249
rect 431 215 465 249
rect 499 215 529 249
rect 392 199 529 215
rect 563 249 628 265
rect 563 215 584 249
rect 618 215 628 249
rect 563 199 628 215
rect 690 169 724 275
rect 781 241 815 379
rect 861 309 887 343
rect 921 309 964 343
rect 861 289 964 309
rect 324 119 358 135
rect 414 131 434 165
rect 468 131 656 165
rect 498 85 528 91
rect 246 57 528 85
rect 562 57 578 91
rect 246 51 578 57
rect 612 85 656 131
rect 690 119 724 135
rect 758 207 815 241
rect 758 85 792 207
rect 906 187 964 289
rect 612 51 792 85
rect 826 157 860 173
rect 826 89 860 123
rect 906 153 907 187
rect 941 161 964 187
rect 906 127 930 153
rect 906 83 964 127
rect 999 119 1033 371
rect 1067 178 1101 455
rect 1888 443 1913 477
rect 1854 421 1913 443
rect 1149 375 1167 409
rect 1201 375 1232 409
rect 1149 341 1232 375
rect 1149 307 1167 341
rect 1201 323 1232 341
rect 1349 387 1379 421
rect 1413 409 1913 421
rect 1413 387 1854 409
rect 1201 307 1203 323
rect 1149 289 1203 307
rect 1237 289 1315 323
rect 1152 249 1237 254
rect 1152 215 1168 249
rect 1202 215 1237 249
rect 1152 199 1237 215
rect 1194 187 1237 199
rect 1067 165 1121 178
rect 1067 144 1160 165
rect 1077 131 1160 144
rect 1126 126 1160 131
rect 1194 153 1203 187
rect 1194 126 1237 153
rect 999 85 1009 119
rect 826 17 860 55
rect 999 63 1032 85
rect 1066 63 1082 97
rect 1126 64 1160 92
rect 1281 85 1315 289
rect 1349 169 1383 387
rect 1806 375 1854 387
rect 1888 375 1913 409
rect 1417 289 1543 345
rect 1587 307 1603 341
rect 1637 307 1823 341
rect 1587 299 1823 307
rect 1417 249 1461 289
rect 1789 265 1823 299
rect 1451 215 1461 249
rect 1417 199 1461 215
rect 1495 239 1557 255
rect 1495 205 1523 239
rect 1601 249 1739 265
rect 1601 215 1629 249
rect 1663 215 1739 249
rect 1789 249 1845 265
rect 1789 215 1801 249
rect 1835 215 1845 249
rect 1495 189 1557 205
rect 1789 199 1845 215
rect 1495 187 1536 189
rect 1495 153 1499 187
rect 1533 153 1536 187
rect 1789 181 1823 199
rect 1495 146 1536 153
rect 1603 150 1823 181
rect 1595 147 1823 150
rect 1349 119 1383 135
rect 1595 142 1653 147
rect 1595 119 1603 142
rect 1417 85 1459 93
rect 999 53 1082 63
rect 1281 59 1459 85
rect 1493 59 1520 93
rect 1595 85 1601 119
rect 1637 108 1653 142
rect 1879 117 1913 375
rect 1635 85 1653 108
rect 1595 59 1653 85
rect 1697 97 1787 113
rect 1697 63 1726 97
rect 1760 63 1787 97
rect 1281 51 1520 59
rect 1697 17 1787 63
rect 1853 101 1913 117
rect 1887 67 1913 101
rect 1853 51 1913 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 713 289 747 323
rect 907 161 941 187
rect 907 153 930 161
rect 930 153 941 161
rect 1203 289 1237 323
rect 1203 153 1237 187
rect 1009 97 1043 119
rect 1009 85 1032 97
rect 1032 85 1043 97
rect 1499 153 1533 187
rect 1601 108 1603 119
rect 1603 108 1635 119
rect 1601 85 1635 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 701 323 759 329
rect 701 289 713 323
rect 747 320 759 323
rect 1191 323 1249 329
rect 1191 320 1203 323
rect 747 292 1203 320
rect 747 289 759 292
rect 701 283 759 289
rect 1191 289 1203 292
rect 1237 289 1249 323
rect 1191 283 1249 289
rect 895 187 953 193
rect 895 153 907 187
rect 941 184 953 187
rect 1191 187 1249 193
rect 1191 184 1203 187
rect 941 156 1203 184
rect 941 153 953 156
rect 895 147 953 153
rect 1191 153 1203 156
rect 1237 184 1249 187
rect 1487 187 1545 193
rect 1487 184 1499 187
rect 1237 156 1499 184
rect 1237 153 1249 156
rect 1191 147 1249 153
rect 1487 153 1499 156
rect 1533 153 1545 187
rect 1487 147 1545 153
rect 997 119 1055 125
rect 997 85 1009 119
rect 1043 116 1055 119
rect 1589 119 1647 125
rect 1589 116 1601 119
rect 1043 88 1601 116
rect 1043 85 1055 88
rect 997 79 1055 85
rect 1589 85 1601 88
rect 1635 85 1647 119
rect 1589 79 1647 85
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 29 357 63 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 404 221 438 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1417 289 1543 345 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1685 221 1719 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xor3_1
rlabel locali s 1417 199 1461 289 1 B
port 2 nsew signal input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2972232
string GDS_START 2959748
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
