magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
rect 475 313 988 331
<< pwell >>
rect 51 49 1606 241
rect 0 0 1632 49
<< scnmos >>
rect 130 47 160 215
rect 216 47 246 215
rect 302 47 332 215
rect 404 47 434 215
rect 490 47 520 215
rect 697 47 727 215
rect 783 47 813 215
rect 869 47 899 215
rect 1067 47 1097 215
rect 1153 47 1183 215
rect 1239 47 1269 215
rect 1325 47 1355 215
rect 1411 47 1441 215
rect 1497 47 1527 215
<< scpmoshvt >>
rect 116 367 146 619
rect 202 367 232 619
rect 288 367 318 619
rect 374 367 404 619
rect 564 349 594 601
rect 650 349 680 601
rect 783 349 813 601
rect 869 349 899 601
rect 1067 367 1097 619
rect 1153 367 1183 619
rect 1239 367 1269 619
rect 1325 367 1355 619
rect 1411 367 1441 619
rect 1497 367 1527 619
<< ndiff >>
rect 77 203 130 215
rect 77 169 85 203
rect 119 169 130 203
rect 77 101 130 169
rect 77 67 85 101
rect 119 67 130 101
rect 77 47 130 67
rect 160 177 216 215
rect 160 143 171 177
rect 205 143 216 177
rect 160 93 216 143
rect 160 59 171 93
rect 205 59 216 93
rect 160 47 216 59
rect 246 203 302 215
rect 246 169 257 203
rect 291 169 302 203
rect 246 101 302 169
rect 246 67 257 101
rect 291 67 302 101
rect 246 47 302 67
rect 332 163 404 215
rect 332 129 351 163
rect 385 129 404 163
rect 332 89 404 129
rect 332 55 351 89
rect 385 55 404 89
rect 332 47 404 55
rect 434 203 490 215
rect 434 169 445 203
rect 479 169 490 203
rect 434 101 490 169
rect 434 67 445 101
rect 479 67 490 101
rect 434 47 490 67
rect 520 163 697 215
rect 520 129 531 163
rect 565 129 652 163
rect 686 129 697 163
rect 520 89 697 129
rect 520 55 531 89
rect 565 55 652 89
rect 686 55 697 89
rect 520 47 697 55
rect 727 203 783 215
rect 727 169 738 203
rect 772 169 783 203
rect 727 101 783 169
rect 727 67 738 101
rect 772 67 783 101
rect 727 47 783 67
rect 813 161 869 215
rect 813 127 824 161
rect 858 127 869 161
rect 813 47 869 127
rect 899 91 956 215
rect 899 57 910 91
rect 944 57 956 91
rect 899 47 956 57
rect 1010 110 1067 215
rect 1010 76 1022 110
rect 1056 76 1067 110
rect 1010 47 1067 76
rect 1097 192 1153 215
rect 1097 158 1108 192
rect 1142 158 1153 192
rect 1097 101 1153 158
rect 1097 67 1108 101
rect 1142 67 1153 101
rect 1097 47 1153 67
rect 1183 203 1239 215
rect 1183 169 1194 203
rect 1228 169 1239 203
rect 1183 89 1239 169
rect 1183 55 1194 89
rect 1228 55 1239 89
rect 1183 47 1239 55
rect 1269 203 1325 215
rect 1269 169 1280 203
rect 1314 169 1325 203
rect 1269 101 1325 169
rect 1269 67 1280 101
rect 1314 67 1325 101
rect 1269 47 1325 67
rect 1355 179 1411 215
rect 1355 145 1366 179
rect 1400 145 1411 179
rect 1355 89 1411 145
rect 1355 55 1366 89
rect 1400 55 1411 89
rect 1355 47 1411 55
rect 1441 203 1497 215
rect 1441 169 1452 203
rect 1486 169 1497 203
rect 1441 101 1497 169
rect 1441 67 1452 101
rect 1486 67 1497 101
rect 1441 47 1497 67
rect 1527 179 1580 215
rect 1527 145 1538 179
rect 1572 145 1580 179
rect 1527 93 1580 145
rect 1527 59 1538 93
rect 1572 59 1580 93
rect 1527 47 1580 59
<< pdiff >>
rect 63 599 116 619
rect 63 565 71 599
rect 105 565 116 599
rect 63 512 116 565
rect 63 478 71 512
rect 105 478 116 512
rect 63 434 116 478
rect 63 400 71 434
rect 105 400 116 434
rect 63 367 116 400
rect 146 541 202 619
rect 146 507 157 541
rect 191 507 202 541
rect 146 423 202 507
rect 146 389 157 423
rect 191 389 202 423
rect 146 367 202 389
rect 232 599 288 619
rect 232 565 243 599
rect 277 565 288 599
rect 232 512 288 565
rect 232 478 243 512
rect 277 478 288 512
rect 232 438 288 478
rect 232 404 243 438
rect 277 404 288 438
rect 232 367 288 404
rect 318 541 374 619
rect 318 507 329 541
rect 363 507 374 541
rect 318 426 374 507
rect 318 392 329 426
rect 363 392 374 426
rect 318 367 374 392
rect 404 599 457 619
rect 1014 607 1067 619
rect 404 565 415 599
rect 449 565 457 599
rect 404 506 457 565
rect 404 472 415 506
rect 449 472 457 506
rect 404 367 457 472
rect 511 589 564 601
rect 511 555 519 589
rect 553 555 564 589
rect 511 494 564 555
rect 511 460 519 494
rect 553 460 564 494
rect 511 349 564 460
rect 594 531 650 601
rect 594 497 605 531
rect 639 497 650 531
rect 594 459 650 497
rect 594 425 605 459
rect 639 425 650 459
rect 594 391 650 425
rect 594 357 605 391
rect 639 357 650 391
rect 594 349 650 357
rect 680 587 783 601
rect 680 553 715 587
rect 749 553 783 587
rect 680 506 783 553
rect 680 472 715 506
rect 749 472 783 506
rect 680 425 783 472
rect 680 391 715 425
rect 749 391 783 425
rect 680 349 783 391
rect 813 589 869 601
rect 813 555 824 589
rect 858 555 869 589
rect 813 501 869 555
rect 813 467 824 501
rect 858 467 869 501
rect 813 349 869 467
rect 899 589 952 601
rect 899 555 910 589
rect 944 555 952 589
rect 899 509 952 555
rect 899 475 910 509
rect 944 475 952 509
rect 899 425 952 475
rect 899 391 910 425
rect 944 391 952 425
rect 899 349 952 391
rect 1014 573 1022 607
rect 1056 573 1067 607
rect 1014 501 1067 573
rect 1014 467 1022 501
rect 1056 467 1067 501
rect 1014 367 1067 467
rect 1097 587 1153 619
rect 1097 553 1108 587
rect 1142 553 1153 587
rect 1097 519 1153 553
rect 1097 485 1108 519
rect 1142 485 1153 519
rect 1097 451 1153 485
rect 1097 417 1108 451
rect 1142 417 1153 451
rect 1097 367 1153 417
rect 1183 607 1239 619
rect 1183 573 1194 607
rect 1228 573 1239 607
rect 1183 516 1239 573
rect 1183 482 1194 516
rect 1228 482 1239 516
rect 1183 425 1239 482
rect 1183 391 1194 425
rect 1228 391 1239 425
rect 1183 367 1239 391
rect 1269 599 1325 619
rect 1269 565 1280 599
rect 1314 565 1325 599
rect 1269 506 1325 565
rect 1269 472 1280 506
rect 1314 472 1325 506
rect 1269 413 1325 472
rect 1269 379 1280 413
rect 1314 379 1325 413
rect 1269 367 1325 379
rect 1355 607 1411 619
rect 1355 573 1366 607
rect 1400 573 1411 607
rect 1355 533 1411 573
rect 1355 499 1366 533
rect 1400 499 1411 533
rect 1355 453 1411 499
rect 1355 419 1366 453
rect 1400 419 1411 453
rect 1355 367 1411 419
rect 1441 599 1497 619
rect 1441 565 1452 599
rect 1486 565 1497 599
rect 1441 506 1497 565
rect 1441 472 1452 506
rect 1486 472 1497 506
rect 1441 413 1497 472
rect 1441 379 1452 413
rect 1486 379 1497 413
rect 1441 367 1497 379
rect 1527 607 1580 619
rect 1527 573 1538 607
rect 1572 573 1580 607
rect 1527 533 1580 573
rect 1527 499 1538 533
rect 1572 499 1580 533
rect 1527 455 1580 499
rect 1527 421 1538 455
rect 1572 421 1580 455
rect 1527 367 1580 421
<< ndiffc >>
rect 85 169 119 203
rect 85 67 119 101
rect 171 143 205 177
rect 171 59 205 93
rect 257 169 291 203
rect 257 67 291 101
rect 351 129 385 163
rect 351 55 385 89
rect 445 169 479 203
rect 445 67 479 101
rect 531 129 565 163
rect 652 129 686 163
rect 531 55 565 89
rect 652 55 686 89
rect 738 169 772 203
rect 738 67 772 101
rect 824 127 858 161
rect 910 57 944 91
rect 1022 76 1056 110
rect 1108 158 1142 192
rect 1108 67 1142 101
rect 1194 169 1228 203
rect 1194 55 1228 89
rect 1280 169 1314 203
rect 1280 67 1314 101
rect 1366 145 1400 179
rect 1366 55 1400 89
rect 1452 169 1486 203
rect 1452 67 1486 101
rect 1538 145 1572 179
rect 1538 59 1572 93
<< pdiffc >>
rect 71 565 105 599
rect 71 478 105 512
rect 71 400 105 434
rect 157 507 191 541
rect 157 389 191 423
rect 243 565 277 599
rect 243 478 277 512
rect 243 404 277 438
rect 329 507 363 541
rect 329 392 363 426
rect 415 565 449 599
rect 415 472 449 506
rect 519 555 553 589
rect 519 460 553 494
rect 605 497 639 531
rect 605 425 639 459
rect 605 357 639 391
rect 715 553 749 587
rect 715 472 749 506
rect 715 391 749 425
rect 824 555 858 589
rect 824 467 858 501
rect 910 555 944 589
rect 910 475 944 509
rect 910 391 944 425
rect 1022 573 1056 607
rect 1022 467 1056 501
rect 1108 553 1142 587
rect 1108 485 1142 519
rect 1108 417 1142 451
rect 1194 573 1228 607
rect 1194 482 1228 516
rect 1194 391 1228 425
rect 1280 565 1314 599
rect 1280 472 1314 506
rect 1280 379 1314 413
rect 1366 573 1400 607
rect 1366 499 1400 533
rect 1366 419 1400 453
rect 1452 565 1486 599
rect 1452 472 1486 506
rect 1452 379 1486 413
rect 1538 573 1572 607
rect 1538 499 1572 533
rect 1538 421 1572 455
<< poly >>
rect 116 619 146 645
rect 202 619 232 645
rect 288 619 318 645
rect 374 619 404 645
rect 564 601 594 627
rect 650 601 680 627
rect 783 601 813 627
rect 869 601 899 627
rect 1067 619 1097 645
rect 1153 619 1183 645
rect 1239 619 1269 645
rect 1325 619 1355 645
rect 1411 619 1441 645
rect 1497 619 1527 645
rect 116 335 146 367
rect 41 319 160 335
rect 41 285 57 319
rect 91 299 160 319
rect 202 299 232 367
rect 288 335 318 367
rect 374 335 404 367
rect 288 319 434 335
rect 91 285 246 299
rect 41 269 246 285
rect 288 285 304 319
rect 338 285 384 319
rect 418 285 434 319
rect 288 269 434 285
rect 564 317 594 349
rect 650 317 680 349
rect 564 301 741 317
rect 564 281 609 301
rect 130 215 160 269
rect 216 215 246 269
rect 302 215 332 269
rect 404 215 434 269
rect 490 267 609 281
rect 643 267 691 301
rect 725 267 741 301
rect 490 251 741 267
rect 783 267 813 349
rect 869 303 899 349
rect 1067 303 1097 367
rect 1153 303 1183 367
rect 869 287 1005 303
rect 869 267 955 287
rect 783 253 955 267
rect 989 253 1005 287
rect 490 215 520 251
rect 697 215 727 251
rect 783 237 1005 253
rect 1067 287 1183 303
rect 1067 253 1120 287
rect 1154 253 1183 287
rect 1067 237 1183 253
rect 783 215 813 237
rect 869 215 899 237
rect 1067 215 1097 237
rect 1153 215 1183 237
rect 1239 331 1269 367
rect 1325 331 1355 367
rect 1411 331 1441 367
rect 1497 331 1527 367
rect 1239 315 1527 331
rect 1239 281 1255 315
rect 1289 281 1323 315
rect 1357 281 1391 315
rect 1425 281 1459 315
rect 1493 281 1527 315
rect 1239 265 1527 281
rect 1239 215 1269 265
rect 1325 215 1355 265
rect 1411 215 1441 265
rect 1497 215 1527 265
rect 130 21 160 47
rect 216 21 246 47
rect 302 21 332 47
rect 404 21 434 47
rect 490 21 520 47
rect 697 21 727 47
rect 783 21 813 47
rect 869 21 899 47
rect 1067 21 1097 47
rect 1153 21 1183 47
rect 1239 21 1269 47
rect 1325 21 1355 47
rect 1411 21 1441 47
rect 1497 21 1527 47
<< polycont >>
rect 57 285 91 319
rect 304 285 338 319
rect 384 285 418 319
rect 609 267 643 301
rect 691 267 725 301
rect 955 253 989 287
rect 1120 253 1154 287
rect 1255 281 1289 315
rect 1323 281 1357 315
rect 1391 281 1425 315
rect 1459 281 1493 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 55 599 465 615
rect 55 565 71 599
rect 105 581 243 599
rect 105 565 107 581
rect 55 512 107 565
rect 241 565 243 581
rect 277 581 415 599
rect 277 565 279 581
rect 55 478 71 512
rect 105 478 107 512
rect 55 434 107 478
rect 55 400 71 434
rect 105 400 107 434
rect 55 384 107 400
rect 141 541 207 547
rect 141 507 157 541
rect 191 507 207 541
rect 141 423 207 507
rect 141 389 157 423
rect 191 389 207 423
rect 141 386 207 389
rect 241 512 279 565
rect 413 565 415 581
rect 449 565 465 599
rect 241 478 243 512
rect 277 478 279 512
rect 241 438 279 478
rect 241 404 243 438
rect 277 404 279 438
rect 241 388 279 404
rect 313 541 379 547
rect 313 507 329 541
rect 363 507 379 541
rect 313 426 379 507
rect 413 506 465 565
rect 413 472 415 506
rect 449 472 465 506
rect 413 456 465 472
rect 503 589 765 615
rect 503 555 519 589
rect 553 587 765 589
rect 553 581 715 587
rect 553 555 569 581
rect 503 494 569 555
rect 699 553 715 581
rect 749 553 765 587
rect 503 460 519 494
rect 553 460 569 494
rect 503 456 569 460
rect 603 531 641 547
rect 603 497 605 531
rect 639 497 641 531
rect 603 459 641 497
rect 313 392 329 426
rect 363 422 379 426
rect 603 425 605 459
rect 639 425 641 459
rect 603 422 641 425
rect 363 392 641 422
rect 313 391 641 392
rect 699 506 765 553
rect 699 472 715 506
rect 749 472 765 506
rect 699 425 765 472
rect 808 589 874 649
rect 1006 607 1072 649
rect 808 555 824 589
rect 858 555 874 589
rect 808 501 874 555
rect 808 467 824 501
rect 858 467 874 501
rect 808 459 874 467
rect 908 589 960 605
rect 908 555 910 589
rect 944 555 960 589
rect 908 509 960 555
rect 908 475 910 509
rect 944 475 960 509
rect 908 425 960 475
rect 1006 573 1022 607
rect 1056 573 1072 607
rect 1006 501 1072 573
rect 1006 467 1022 501
rect 1056 467 1072 501
rect 1006 459 1072 467
rect 1106 587 1144 615
rect 1106 553 1108 587
rect 1142 553 1144 587
rect 1106 519 1144 553
rect 1106 485 1108 519
rect 1142 485 1144 519
rect 1106 451 1144 485
rect 1106 425 1108 451
rect 699 391 715 425
rect 749 391 910 425
rect 944 417 1108 425
rect 1142 417 1144 451
rect 944 391 1144 417
rect 1178 607 1244 649
rect 1178 573 1194 607
rect 1228 573 1244 607
rect 1178 516 1244 573
rect 1178 482 1194 516
rect 1228 482 1244 516
rect 1178 425 1244 482
rect 1178 391 1194 425
rect 1228 391 1244 425
rect 1278 599 1316 615
rect 1278 565 1280 599
rect 1314 565 1316 599
rect 1278 506 1316 565
rect 1278 472 1280 506
rect 1314 472 1316 506
rect 1278 413 1316 472
rect 1350 607 1416 649
rect 1350 573 1366 607
rect 1400 573 1416 607
rect 1350 533 1416 573
rect 1350 499 1366 533
rect 1400 499 1416 533
rect 1350 453 1416 499
rect 1350 419 1366 453
rect 1400 419 1416 453
rect 1450 599 1488 615
rect 1450 565 1452 599
rect 1486 565 1488 599
rect 1450 506 1488 565
rect 1450 472 1452 506
rect 1486 472 1488 506
rect 313 388 605 391
rect 17 319 107 350
rect 17 285 57 319
rect 91 285 107 319
rect 141 247 187 386
rect 593 357 605 388
rect 639 357 641 391
rect 1278 379 1280 413
rect 1314 385 1316 413
rect 1450 413 1488 472
rect 1522 607 1588 649
rect 1522 573 1538 607
rect 1572 573 1588 607
rect 1522 533 1588 573
rect 1522 499 1538 533
rect 1572 499 1588 533
rect 1522 455 1588 499
rect 1522 421 1538 455
rect 1572 421 1588 455
rect 1450 385 1452 413
rect 1314 379 1452 385
rect 1486 385 1488 413
rect 1486 379 1615 385
rect 221 319 559 354
rect 593 341 641 357
rect 221 285 304 319
rect 338 285 384 319
rect 418 285 559 319
rect 675 307 833 357
rect 593 301 833 307
rect 593 267 609 301
rect 643 267 691 301
rect 725 267 833 301
rect 869 323 1240 357
rect 1278 349 1615 379
rect 69 231 291 247
rect 869 231 903 323
rect 1204 315 1240 323
rect 939 287 1034 289
rect 939 253 955 287
rect 989 253 1034 287
rect 939 242 1034 253
rect 1068 287 1170 289
rect 1068 253 1120 287
rect 1154 253 1170 287
rect 1204 281 1255 315
rect 1289 281 1323 315
rect 1357 281 1391 315
rect 1425 281 1459 315
rect 1493 281 1509 315
rect 1068 242 1170 253
rect 1543 247 1615 349
rect 69 213 903 231
rect 69 203 121 213
rect 69 169 85 203
rect 119 169 121 203
rect 255 203 903 213
rect 1278 213 1615 247
rect 69 101 121 169
rect 69 67 85 101
rect 119 67 121 101
rect 69 51 121 67
rect 155 143 171 177
rect 205 143 221 177
rect 155 93 221 143
rect 155 59 171 93
rect 205 59 221 93
rect 155 17 221 59
rect 255 169 257 203
rect 291 197 445 203
rect 291 169 301 197
rect 255 101 301 169
rect 435 169 445 197
rect 479 197 738 203
rect 479 169 481 197
rect 255 67 257 101
rect 291 67 301 101
rect 255 51 301 67
rect 335 129 351 163
rect 385 129 401 163
rect 335 89 401 129
rect 335 55 351 89
rect 385 55 401 89
rect 335 17 401 55
rect 435 101 481 169
rect 736 169 738 197
rect 772 197 903 203
rect 772 169 774 197
rect 435 67 445 101
rect 479 67 481 101
rect 435 51 481 67
rect 515 129 531 163
rect 565 129 652 163
rect 686 129 702 163
rect 515 89 702 129
rect 515 55 531 89
rect 565 55 652 89
rect 686 55 702 89
rect 515 17 702 55
rect 736 101 774 169
rect 937 192 1144 208
rect 937 163 1108 192
rect 808 161 1108 163
rect 808 127 824 161
rect 858 158 1108 161
rect 1142 158 1144 192
rect 858 152 1144 158
rect 858 127 972 152
rect 736 67 738 101
rect 772 93 774 101
rect 1006 110 1072 118
rect 772 91 960 93
rect 772 67 910 91
rect 736 57 910 67
rect 944 57 960 91
rect 736 51 960 57
rect 1006 76 1022 110
rect 1056 76 1072 110
rect 1006 17 1072 76
rect 1106 101 1144 152
rect 1106 67 1108 101
rect 1142 67 1144 101
rect 1106 51 1144 67
rect 1178 203 1244 208
rect 1178 169 1194 203
rect 1228 169 1244 203
rect 1178 89 1244 169
rect 1178 55 1194 89
rect 1228 55 1244 89
rect 1178 17 1244 55
rect 1278 203 1316 213
rect 1278 169 1280 203
rect 1314 169 1316 203
rect 1450 203 1488 213
rect 1278 101 1316 169
rect 1278 67 1280 101
rect 1314 67 1316 101
rect 1278 51 1316 67
rect 1350 145 1366 179
rect 1400 145 1416 179
rect 1350 89 1416 145
rect 1350 55 1366 89
rect 1400 55 1416 89
rect 1350 17 1416 55
rect 1450 169 1452 203
rect 1486 169 1488 203
rect 1450 101 1488 169
rect 1450 67 1452 101
rect 1486 67 1488 101
rect 1450 51 1488 67
rect 1522 145 1538 179
rect 1572 145 1588 179
rect 1522 93 1588 145
rect 1522 59 1538 93
rect 1572 59 1588 93
rect 1522 17 1588 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2111o_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1077716
string GDS_START 1063836
<< end >>
