magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 12 49 1055 241
rect 0 0 1056 49
<< scnmos >>
rect 91 131 121 215
rect 282 47 312 215
rect 368 47 398 215
rect 454 47 484 215
rect 540 47 570 215
rect 688 47 718 215
rect 774 47 804 215
rect 860 47 890 215
rect 946 47 976 215
<< scpmoshvt >>
rect 80 535 110 619
rect 282 367 312 619
rect 368 367 398 619
rect 454 367 484 619
rect 540 367 570 619
rect 642 367 672 619
rect 774 367 804 619
rect 860 367 890 619
rect 946 367 976 619
<< ndiff >>
rect 38 197 91 215
rect 38 163 46 197
rect 80 163 91 197
rect 38 131 91 163
rect 121 183 282 215
rect 121 149 189 183
rect 223 149 282 183
rect 121 131 282 149
rect 213 93 282 131
rect 213 59 221 93
rect 255 59 282 93
rect 213 47 282 59
rect 312 183 368 215
rect 312 149 323 183
rect 357 149 368 183
rect 312 101 368 149
rect 312 67 323 101
rect 357 67 368 101
rect 312 47 368 67
rect 398 107 454 215
rect 398 73 409 107
rect 443 73 454 107
rect 398 47 454 73
rect 484 183 540 215
rect 484 149 495 183
rect 529 149 540 183
rect 484 101 540 149
rect 484 67 495 101
rect 529 67 540 101
rect 484 47 540 67
rect 570 107 688 215
rect 570 73 613 107
rect 647 73 688 107
rect 570 47 688 73
rect 718 192 774 215
rect 718 158 729 192
rect 763 158 774 192
rect 718 101 774 158
rect 718 67 729 101
rect 763 67 774 101
rect 718 47 774 67
rect 804 132 860 215
rect 804 98 815 132
rect 849 98 860 132
rect 804 47 860 98
rect 890 192 946 215
rect 890 158 901 192
rect 935 158 946 192
rect 890 103 946 158
rect 890 69 901 103
rect 935 69 946 103
rect 890 47 946 69
rect 976 203 1029 215
rect 976 169 987 203
rect 1021 169 1029 203
rect 976 93 1029 169
rect 976 59 987 93
rect 1021 59 1029 93
rect 976 47 1029 59
<< pdiff >>
rect 27 594 80 619
rect 27 560 35 594
rect 69 560 80 594
rect 27 535 80 560
rect 110 594 163 619
rect 110 560 121 594
rect 155 560 163 594
rect 110 535 163 560
rect 229 599 282 619
rect 229 565 237 599
rect 271 565 282 599
rect 229 527 282 565
rect 229 493 237 527
rect 271 493 282 527
rect 229 457 282 493
rect 229 423 237 457
rect 271 423 282 457
rect 229 367 282 423
rect 312 581 368 619
rect 312 547 323 581
rect 357 547 368 581
rect 312 367 368 547
rect 398 413 454 619
rect 398 379 409 413
rect 443 379 454 413
rect 398 367 454 379
rect 484 581 540 619
rect 484 547 495 581
rect 529 547 540 581
rect 484 367 540 547
rect 570 607 642 619
rect 570 573 597 607
rect 631 573 642 607
rect 570 537 642 573
rect 570 503 597 537
rect 631 503 642 537
rect 570 463 642 503
rect 570 429 597 463
rect 631 429 642 463
rect 570 367 642 429
rect 672 607 774 619
rect 672 573 704 607
rect 738 573 774 607
rect 672 531 774 573
rect 672 497 704 531
rect 738 497 774 531
rect 672 367 774 497
rect 804 529 860 619
rect 804 495 815 529
rect 849 495 860 529
rect 804 367 860 495
rect 890 607 946 619
rect 890 573 901 607
rect 935 573 946 607
rect 890 367 946 573
rect 976 451 1029 619
rect 976 417 987 451
rect 1021 417 1029 451
rect 976 367 1029 417
<< ndiffc >>
rect 46 163 80 197
rect 189 149 223 183
rect 221 59 255 93
rect 323 149 357 183
rect 323 67 357 101
rect 409 73 443 107
rect 495 149 529 183
rect 495 67 529 101
rect 613 73 647 107
rect 729 158 763 192
rect 729 67 763 101
rect 815 98 849 132
rect 901 158 935 192
rect 901 69 935 103
rect 987 169 1021 203
rect 987 59 1021 93
<< pdiffc >>
rect 35 560 69 594
rect 121 560 155 594
rect 237 565 271 599
rect 237 493 271 527
rect 237 423 271 457
rect 323 547 357 581
rect 409 379 443 413
rect 495 547 529 581
rect 597 573 631 607
rect 597 503 631 537
rect 597 429 631 463
rect 704 573 738 607
rect 704 497 738 531
rect 815 495 849 529
rect 901 573 935 607
rect 987 417 1021 451
<< poly >>
rect 80 619 110 645
rect 282 619 312 645
rect 368 619 398 645
rect 454 619 484 645
rect 540 619 570 645
rect 642 619 672 645
rect 774 619 804 645
rect 860 619 890 645
rect 946 619 976 645
rect 80 303 110 535
rect 282 303 312 367
rect 21 287 110 303
rect 21 253 37 287
rect 71 267 110 287
rect 163 287 312 303
rect 71 253 121 267
rect 21 237 121 253
rect 163 253 179 287
rect 213 253 312 287
rect 163 237 312 253
rect 91 215 121 237
rect 282 215 312 237
rect 368 335 398 367
rect 454 335 484 367
rect 368 319 484 335
rect 368 285 414 319
rect 448 285 484 319
rect 540 303 570 367
rect 642 335 672 367
rect 642 319 732 335
rect 368 269 484 285
rect 368 215 398 269
rect 454 215 484 269
rect 526 287 592 303
rect 526 253 542 287
rect 576 253 592 287
rect 642 285 682 319
rect 716 285 732 319
rect 642 269 732 285
rect 774 303 804 367
rect 860 303 890 367
rect 774 287 890 303
rect 526 237 592 253
rect 540 215 570 237
rect 688 215 718 269
rect 774 253 840 287
rect 874 253 890 287
rect 774 237 890 253
rect 774 215 804 237
rect 860 215 890 237
rect 946 303 976 367
rect 946 287 1029 303
rect 946 253 979 287
rect 1013 253 1029 287
rect 946 237 1029 253
rect 946 215 976 237
rect 91 105 121 131
rect 282 21 312 47
rect 368 21 398 47
rect 454 21 484 47
rect 540 21 570 47
rect 688 21 718 47
rect 774 21 804 47
rect 860 21 890 47
rect 946 21 976 47
<< polycont >>
rect 37 253 71 287
rect 179 253 213 287
rect 414 285 448 319
rect 542 253 576 287
rect 682 285 716 319
rect 840 253 874 287
rect 979 253 1013 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 19 594 71 610
rect 19 560 35 594
rect 69 560 71 594
rect 19 373 71 560
rect 105 594 171 649
rect 105 560 121 594
rect 155 560 171 594
rect 105 544 171 560
rect 221 599 282 615
rect 581 607 647 615
rect 221 565 237 599
rect 271 565 282 599
rect 221 527 282 565
rect 316 581 547 602
rect 316 547 323 581
rect 357 547 495 581
rect 529 547 547 581
rect 316 531 547 547
rect 581 573 597 607
rect 631 573 647 607
rect 581 537 647 573
rect 221 493 237 527
rect 271 497 282 527
rect 581 503 597 537
rect 631 503 647 537
rect 581 497 647 503
rect 688 607 951 615
rect 688 573 704 607
rect 738 573 901 607
rect 935 573 951 607
rect 688 567 951 573
rect 688 531 754 567
rect 987 533 1039 649
rect 688 497 704 531
rect 738 497 754 531
rect 799 529 1039 533
rect 271 493 647 497
rect 221 463 647 493
rect 799 495 815 529
rect 849 495 1039 529
rect 799 491 1039 495
rect 221 457 283 463
rect 221 423 237 457
rect 271 423 283 457
rect 581 429 597 463
rect 631 457 763 463
rect 631 451 1037 457
rect 631 429 987 451
rect 221 407 283 423
rect 317 413 547 429
rect 317 379 409 413
rect 443 395 547 413
rect 729 417 987 429
rect 1021 417 1037 451
rect 729 401 1037 417
rect 443 379 646 395
rect 19 339 283 373
rect 317 361 646 379
rect 17 287 71 303
rect 17 253 37 287
rect 17 237 71 253
rect 105 201 139 339
rect 249 327 283 339
rect 249 319 464 327
rect 173 287 213 303
rect 173 253 179 287
rect 249 285 414 319
rect 448 285 464 319
rect 498 287 576 303
rect 173 251 213 253
rect 498 253 542 287
rect 498 251 576 253
rect 173 217 576 251
rect 612 235 646 361
rect 680 323 1039 357
rect 680 319 732 323
rect 680 285 682 319
rect 716 285 732 319
rect 680 269 732 285
rect 774 287 929 289
rect 774 253 840 287
rect 874 253 929 287
rect 774 242 929 253
rect 963 287 1039 323
rect 963 253 979 287
rect 1013 253 1039 287
rect 963 237 1039 253
rect 30 197 139 201
rect 30 163 46 197
rect 80 163 139 197
rect 612 208 740 235
rect 612 192 937 208
rect 612 183 729 192
rect 30 159 139 163
rect 173 149 189 183
rect 223 149 273 183
rect 173 93 273 149
rect 173 59 221 93
rect 255 59 273 93
rect 173 17 273 59
rect 307 149 323 183
rect 357 149 495 183
rect 529 158 729 183
rect 763 174 901 192
rect 763 158 765 174
rect 529 149 765 158
rect 307 101 359 149
rect 307 67 323 101
rect 357 67 359 101
rect 307 51 359 67
rect 393 107 459 115
rect 393 73 409 107
rect 443 73 459 107
rect 393 17 459 73
rect 493 101 545 149
rect 493 67 495 101
rect 529 67 545 101
rect 493 51 545 67
rect 597 107 663 115
rect 597 73 613 107
rect 647 73 663 107
rect 597 17 663 73
rect 713 101 765 149
rect 899 158 901 174
rect 935 158 937 192
rect 713 67 729 101
rect 763 67 765 101
rect 713 51 765 67
rect 799 132 865 140
rect 799 98 815 132
rect 849 98 865 132
rect 799 17 865 98
rect 899 103 937 158
rect 899 69 901 103
rect 935 69 937 103
rect 899 53 937 69
rect 971 169 987 203
rect 1021 169 1037 203
rect 971 93 1037 169
rect 971 59 987 93
rect 1021 59 1037 93
rect 971 17 1037 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4b_2
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1793290
string GDS_START 1784524
<< end >>
