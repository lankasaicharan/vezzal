magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 41 178 504 235
rect 41 49 863 178
rect 0 0 864 49
<< scnmos >>
rect 124 125 154 209
rect 202 125 232 209
rect 320 125 350 209
rect 398 125 428 209
rect 500 68 530 152
rect 592 68 622 152
rect 678 68 708 152
rect 750 68 780 152
<< scpmoshvt >>
rect 102 419 152 619
rect 194 419 244 619
rect 300 419 350 619
rect 392 419 442 619
rect 498 419 548 619
rect 598 419 648 619
rect 706 419 756 619
<< ndiff >>
rect 67 182 124 209
rect 67 148 79 182
rect 113 148 124 182
rect 67 125 124 148
rect 154 125 202 209
rect 232 125 320 209
rect 350 125 398 209
rect 428 152 478 209
rect 428 127 500 152
rect 428 125 455 127
rect 247 114 305 125
rect 247 80 259 114
rect 293 80 305 114
rect 247 68 305 80
rect 443 93 455 125
rect 489 93 500 127
rect 443 68 500 93
rect 530 68 592 152
rect 622 120 678 152
rect 622 86 633 120
rect 667 86 678 120
rect 622 68 678 86
rect 708 68 750 152
rect 780 127 837 152
rect 780 93 791 127
rect 825 93 837 127
rect 780 68 837 93
<< pdiff >>
rect 29 597 102 619
rect 29 563 41 597
rect 75 563 102 597
rect 29 465 102 563
rect 29 431 41 465
rect 75 431 102 465
rect 29 419 102 431
rect 152 419 194 619
rect 244 596 300 619
rect 244 562 255 596
rect 289 562 300 596
rect 244 419 300 562
rect 350 419 392 619
rect 442 597 498 619
rect 442 563 453 597
rect 487 563 498 597
rect 442 469 498 563
rect 442 435 453 469
rect 487 435 498 469
rect 442 419 498 435
rect 548 419 598 619
rect 648 607 706 619
rect 648 573 659 607
rect 693 573 706 607
rect 648 538 706 573
rect 648 504 659 538
rect 693 504 706 538
rect 648 469 706 504
rect 648 435 659 469
rect 693 435 706 469
rect 648 419 706 435
rect 756 597 813 619
rect 756 563 767 597
rect 801 563 813 597
rect 756 465 813 563
rect 756 431 767 465
rect 801 431 813 465
rect 756 419 813 431
<< ndiffc >>
rect 79 148 113 182
rect 259 80 293 114
rect 455 93 489 127
rect 633 86 667 120
rect 791 93 825 127
<< pdiffc >>
rect 41 563 75 597
rect 41 431 75 465
rect 255 562 289 596
rect 453 563 487 597
rect 453 435 487 469
rect 659 573 693 607
rect 659 504 693 538
rect 659 435 693 469
rect 767 563 801 597
rect 767 431 801 465
<< poly >>
rect 102 619 152 645
rect 194 619 244 645
rect 300 619 350 645
rect 392 619 442 645
rect 498 619 548 645
rect 598 619 648 645
rect 706 619 756 645
rect 102 379 152 419
rect 86 363 152 379
rect 86 329 102 363
rect 136 329 152 363
rect 86 295 152 329
rect 194 387 244 419
rect 300 387 350 419
rect 194 371 350 387
rect 194 337 300 371
rect 334 337 350 371
rect 194 323 350 337
rect 86 261 102 295
rect 136 275 152 295
rect 202 321 350 323
rect 136 261 154 275
rect 86 245 154 261
rect 124 209 154 245
rect 202 209 232 321
rect 320 209 350 321
rect 392 275 442 419
rect 498 383 548 419
rect 598 383 648 419
rect 484 367 550 383
rect 484 333 500 367
rect 534 333 550 367
rect 484 317 550 333
rect 592 367 658 383
rect 592 333 608 367
rect 642 333 658 367
rect 592 299 658 333
rect 592 275 608 299
rect 392 265 608 275
rect 642 265 658 299
rect 392 245 658 265
rect 706 331 756 419
rect 706 315 772 331
rect 706 281 722 315
rect 756 281 772 315
rect 706 247 772 281
rect 398 209 428 245
rect 500 152 530 178
rect 592 152 622 245
rect 706 213 722 247
rect 756 213 772 247
rect 706 197 772 213
rect 678 167 780 197
rect 678 152 708 167
rect 750 152 780 167
rect 124 51 154 125
rect 202 99 232 125
rect 320 99 350 125
rect 398 99 428 125
rect 500 51 530 68
rect 124 21 530 51
rect 592 42 622 68
rect 678 42 708 68
rect 750 42 780 68
<< polycont >>
rect 102 329 136 363
rect 300 337 334 371
rect 102 261 136 295
rect 500 333 534 367
rect 608 333 642 367
rect 608 265 642 299
rect 722 281 756 315
rect 722 213 756 247
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 18 597 91 613
rect 18 563 41 597
rect 75 563 91 597
rect 18 500 91 563
rect 239 596 305 649
rect 239 562 255 596
rect 289 562 305 596
rect 239 536 305 562
rect 437 597 503 613
rect 437 563 453 597
rect 487 563 503 597
rect 437 500 503 563
rect 18 469 503 500
rect 18 466 453 469
rect 18 465 91 466
rect 18 431 41 465
rect 75 431 91 465
rect 18 415 91 431
rect 437 435 453 466
rect 487 435 503 469
rect 18 209 52 415
rect 88 363 152 379
rect 88 329 102 363
rect 136 329 152 363
rect 88 295 152 329
rect 217 371 359 430
rect 437 419 503 435
rect 643 607 709 649
rect 643 573 659 607
rect 693 573 709 607
rect 643 538 709 573
rect 643 504 659 538
rect 693 504 709 538
rect 643 469 709 504
rect 643 435 659 469
rect 693 435 709 469
rect 643 419 709 435
rect 751 597 842 613
rect 751 563 767 597
rect 801 563 842 597
rect 751 465 842 563
rect 751 431 767 465
rect 801 431 842 465
rect 751 384 842 431
rect 217 337 300 371
rect 334 337 359 371
rect 217 321 359 337
rect 484 367 550 383
rect 484 333 500 367
rect 534 333 550 367
rect 88 261 102 295
rect 136 283 152 295
rect 484 283 550 333
rect 136 261 550 283
rect 88 249 550 261
rect 592 367 658 383
rect 592 333 608 367
rect 642 333 658 367
rect 592 299 658 333
rect 592 265 608 299
rect 642 265 658 299
rect 592 249 658 265
rect 705 315 772 331
rect 705 281 722 315
rect 756 281 772 315
rect 88 245 263 249
rect 217 236 263 245
rect 705 247 772 281
rect 705 213 722 247
rect 756 213 772 247
rect 18 200 129 209
rect 299 200 772 213
rect 18 197 772 200
rect 18 182 739 197
rect 18 175 79 182
rect 63 148 79 175
rect 113 179 739 182
rect 113 166 333 179
rect 113 148 129 166
rect 63 121 129 148
rect 243 114 309 130
rect 243 80 259 114
rect 293 80 309 114
rect 243 17 309 80
rect 439 127 505 179
rect 808 156 842 384
rect 439 93 455 127
rect 489 93 505 127
rect 439 64 505 93
rect 617 120 683 143
rect 617 86 633 120
rect 667 86 683 120
rect 617 17 683 86
rect 775 127 842 156
rect 775 93 791 127
rect 825 93 842 127
rect 775 64 842 93
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 maj3_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6751622
string GDS_START 6744790
<< end >>
