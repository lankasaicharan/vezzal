magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3794 1975
<< nwell >>
rect -38 331 2534 704
rect 1763 299 1971 331
<< pwell >>
rect 367 209 803 229
rect 4 157 803 209
rect 1066 157 1733 201
rect 4 49 1733 157
rect 1963 49 2495 243
rect 0 0 2496 49
<< scnmos >>
rect 83 99 113 183
rect 242 99 272 183
rect 446 119 476 203
rect 532 119 562 203
rect 618 119 648 203
rect 690 119 720 203
rect 884 47 914 131
rect 956 47 986 131
rect 1145 47 1175 175
rect 1217 47 1247 175
rect 1326 91 1356 175
rect 1398 91 1428 175
rect 1470 91 1500 175
rect 1624 91 1654 175
rect 2042 49 2072 217
rect 2128 49 2158 217
rect 2214 49 2244 217
rect 2300 49 2330 217
rect 2386 49 2416 217
<< scpmoshvt >>
rect 114 465 144 593
rect 200 465 230 593
rect 488 463 518 547
rect 574 463 604 547
rect 660 463 690 547
rect 732 463 762 547
rect 841 463 871 547
rect 927 463 957 547
rect 1064 379 1094 547
rect 1254 407 1284 491
rect 1359 407 1389 575
rect 1574 457 1604 541
rect 1660 457 1690 541
rect 1852 335 1882 419
rect 2042 367 2072 619
rect 2128 367 2158 619
rect 2214 367 2244 619
rect 2300 367 2330 619
rect 2386 367 2416 619
<< ndiff >>
rect 30 158 83 183
rect 30 124 38 158
rect 72 124 83 158
rect 30 99 83 124
rect 113 158 242 183
rect 113 124 197 158
rect 231 124 242 158
rect 113 99 242 124
rect 272 158 325 183
rect 272 124 283 158
rect 317 124 325 158
rect 272 99 325 124
rect 393 178 446 203
rect 393 144 401 178
rect 435 144 446 178
rect 393 119 446 144
rect 476 178 532 203
rect 476 144 487 178
rect 521 144 532 178
rect 476 119 532 144
rect 562 167 618 203
rect 562 133 573 167
rect 607 133 618 167
rect 562 119 618 133
rect 648 119 690 203
rect 720 161 777 203
rect 720 127 731 161
rect 765 127 777 161
rect 1092 161 1145 175
rect 1092 131 1100 161
rect 720 119 777 127
rect 831 107 884 131
rect 831 73 839 107
rect 873 73 884 107
rect 831 47 884 73
rect 914 47 956 131
rect 986 127 1100 131
rect 1134 127 1145 161
rect 986 106 1145 127
rect 986 72 997 106
rect 1031 93 1145 106
rect 1031 72 1100 93
rect 986 59 1100 72
rect 1134 59 1145 93
rect 986 47 1145 59
rect 1175 47 1217 175
rect 1247 163 1326 175
rect 1247 129 1281 163
rect 1315 129 1326 163
rect 1247 95 1326 129
rect 1247 61 1258 95
rect 1292 91 1326 95
rect 1356 91 1398 175
rect 1428 91 1470 175
rect 1500 148 1624 175
rect 1500 114 1511 148
rect 1545 114 1579 148
rect 1613 114 1624 148
rect 1500 91 1624 114
rect 1654 141 1707 175
rect 1654 107 1665 141
rect 1699 107 1707 141
rect 1654 91 1707 107
rect 1989 205 2042 217
rect 1989 171 1997 205
rect 2031 171 2042 205
rect 1292 61 1300 91
rect 1247 47 1300 61
rect 1989 101 2042 171
rect 1989 67 1997 101
rect 2031 67 2042 101
rect 1989 49 2042 67
rect 2072 205 2128 217
rect 2072 171 2083 205
rect 2117 171 2128 205
rect 2072 95 2128 171
rect 2072 61 2083 95
rect 2117 61 2128 95
rect 2072 49 2128 61
rect 2158 205 2214 217
rect 2158 171 2169 205
rect 2203 171 2214 205
rect 2158 101 2214 171
rect 2158 67 2169 101
rect 2203 67 2214 101
rect 2158 49 2214 67
rect 2244 181 2300 217
rect 2244 147 2255 181
rect 2289 147 2300 181
rect 2244 95 2300 147
rect 2244 61 2255 95
rect 2289 61 2300 95
rect 2244 49 2300 61
rect 2330 205 2386 217
rect 2330 171 2341 205
rect 2375 171 2386 205
rect 2330 101 2386 171
rect 2330 67 2341 101
rect 2375 67 2386 101
rect 2330 49 2386 67
rect 2416 181 2469 217
rect 2416 147 2427 181
rect 2461 147 2469 181
rect 2416 95 2469 147
rect 2416 61 2427 95
rect 2461 61 2469 95
rect 2416 49 2469 61
<< pdiff >>
rect 57 579 114 593
rect 57 545 65 579
rect 99 545 114 579
rect 57 511 114 545
rect 57 477 65 511
rect 99 477 114 511
rect 57 465 114 477
rect 144 570 200 593
rect 144 536 155 570
rect 189 536 200 570
rect 144 465 200 536
rect 230 578 283 593
rect 230 544 241 578
rect 275 544 283 578
rect 1411 609 1461 621
rect 1411 575 1419 609
rect 1453 575 1461 609
rect 230 465 283 544
rect 435 527 488 547
rect 435 493 443 527
rect 477 493 488 527
rect 435 481 488 493
rect 438 463 488 481
rect 518 522 574 547
rect 518 488 529 522
rect 563 488 574 522
rect 518 463 574 488
rect 604 522 660 547
rect 604 488 615 522
rect 649 488 660 522
rect 604 463 660 488
rect 690 463 732 547
rect 762 522 841 547
rect 762 488 777 522
rect 811 488 841 522
rect 762 463 841 488
rect 871 522 927 547
rect 871 488 882 522
rect 916 488 927 522
rect 871 463 927 488
rect 957 539 1064 547
rect 957 505 1019 539
rect 1053 505 1064 539
rect 957 471 1064 505
rect 957 463 1019 471
rect 1011 437 1019 463
rect 1053 437 1064 471
rect 1011 379 1064 437
rect 1094 535 1147 547
rect 1094 501 1105 535
rect 1139 501 1147 535
rect 1094 467 1147 501
rect 1306 491 1359 575
rect 1094 433 1105 467
rect 1139 433 1147 467
rect 1094 379 1147 433
rect 1201 466 1254 491
rect 1201 432 1209 466
rect 1243 432 1254 466
rect 1201 407 1254 432
rect 1284 455 1359 491
rect 1284 421 1309 455
rect 1343 421 1359 455
rect 1284 407 1359 421
rect 1389 407 1461 575
rect 1521 521 1574 541
rect 1521 487 1529 521
rect 1563 487 1574 521
rect 1521 457 1574 487
rect 1604 516 1660 541
rect 1604 482 1615 516
rect 1649 482 1660 516
rect 1604 457 1660 482
rect 1690 516 1743 541
rect 1690 482 1701 516
rect 1735 482 1743 516
rect 1989 599 2042 619
rect 1989 565 1997 599
rect 2031 565 2042 599
rect 1989 505 2042 565
rect 1690 457 1743 482
rect 1989 471 1997 505
rect 2031 471 2042 505
rect 1799 394 1852 419
rect 1799 360 1807 394
rect 1841 360 1852 394
rect 1799 335 1852 360
rect 1882 394 1935 419
rect 1882 360 1893 394
rect 1927 360 1935 394
rect 1989 413 2042 471
rect 1989 379 1997 413
rect 2031 379 2042 413
rect 1989 367 2042 379
rect 2072 607 2128 619
rect 2072 573 2083 607
rect 2117 573 2128 607
rect 2072 507 2128 573
rect 2072 473 2083 507
rect 2117 473 2128 507
rect 2072 409 2128 473
rect 2072 375 2083 409
rect 2117 375 2128 409
rect 2072 367 2128 375
rect 2158 599 2214 619
rect 2158 565 2169 599
rect 2203 565 2214 599
rect 2158 505 2214 565
rect 2158 471 2169 505
rect 2203 471 2214 505
rect 2158 413 2214 471
rect 2158 379 2169 413
rect 2203 379 2214 413
rect 2158 367 2214 379
rect 2244 611 2300 619
rect 2244 577 2255 611
rect 2289 577 2300 611
rect 2244 533 2300 577
rect 2244 499 2255 533
rect 2289 499 2300 533
rect 2244 455 2300 499
rect 2244 421 2255 455
rect 2289 421 2300 455
rect 2244 367 2300 421
rect 2330 599 2386 619
rect 2330 565 2341 599
rect 2375 565 2386 599
rect 2330 505 2386 565
rect 2330 471 2341 505
rect 2375 471 2386 505
rect 2330 413 2386 471
rect 2330 379 2341 413
rect 2375 379 2386 413
rect 2330 367 2386 379
rect 2416 607 2469 619
rect 2416 573 2427 607
rect 2461 573 2469 607
rect 2416 533 2469 573
rect 2416 499 2427 533
rect 2461 499 2469 533
rect 2416 455 2469 499
rect 2416 421 2427 455
rect 2461 421 2469 455
rect 2416 367 2469 421
rect 1882 335 1935 360
<< ndiffc >>
rect 38 124 72 158
rect 197 124 231 158
rect 283 124 317 158
rect 401 144 435 178
rect 487 144 521 178
rect 573 133 607 167
rect 731 127 765 161
rect 839 73 873 107
rect 1100 127 1134 161
rect 997 72 1031 106
rect 1100 59 1134 93
rect 1281 129 1315 163
rect 1258 61 1292 95
rect 1511 114 1545 148
rect 1579 114 1613 148
rect 1665 107 1699 141
rect 1997 171 2031 205
rect 1997 67 2031 101
rect 2083 171 2117 205
rect 2083 61 2117 95
rect 2169 171 2203 205
rect 2169 67 2203 101
rect 2255 147 2289 181
rect 2255 61 2289 95
rect 2341 171 2375 205
rect 2341 67 2375 101
rect 2427 147 2461 181
rect 2427 61 2461 95
<< pdiffc >>
rect 65 545 99 579
rect 65 477 99 511
rect 155 536 189 570
rect 241 544 275 578
rect 1419 575 1453 609
rect 443 493 477 527
rect 529 488 563 522
rect 615 488 649 522
rect 777 488 811 522
rect 882 488 916 522
rect 1019 505 1053 539
rect 1019 437 1053 471
rect 1105 501 1139 535
rect 1105 433 1139 467
rect 1209 432 1243 466
rect 1309 421 1343 455
rect 1529 487 1563 521
rect 1615 482 1649 516
rect 1701 482 1735 516
rect 1997 565 2031 599
rect 1997 471 2031 505
rect 1807 360 1841 394
rect 1893 360 1927 394
rect 1997 379 2031 413
rect 2083 573 2117 607
rect 2083 473 2117 507
rect 2083 375 2117 409
rect 2169 565 2203 599
rect 2169 471 2203 505
rect 2169 379 2203 413
rect 2255 577 2289 611
rect 2255 499 2289 533
rect 2255 421 2289 455
rect 2341 565 2375 599
rect 2341 471 2375 505
rect 2341 379 2375 413
rect 2427 573 2461 607
rect 2427 499 2461 533
rect 2427 421 2461 455
<< poly >>
rect 114 593 144 619
rect 200 615 1389 645
rect 200 593 230 615
rect 488 547 518 573
rect 574 547 604 573
rect 660 547 690 615
rect 1359 575 1389 615
rect 732 547 762 573
rect 841 547 871 573
rect 927 547 957 573
rect 1064 547 1094 573
rect 114 339 144 465
rect 200 433 230 465
rect 340 441 406 449
rect 488 441 518 463
rect 340 433 518 441
rect 200 417 272 433
rect 200 383 216 417
rect 250 383 272 417
rect 340 399 356 433
rect 390 411 518 433
rect 390 399 406 411
rect 340 383 406 399
rect 200 349 272 383
rect 83 323 158 339
rect 83 289 108 323
rect 142 289 158 323
rect 200 315 216 349
rect 250 315 272 349
rect 200 299 272 315
rect 83 255 158 289
rect 83 221 108 255
rect 142 221 158 255
rect 83 205 158 221
rect 83 183 113 205
rect 242 183 272 299
rect 376 255 406 383
rect 454 347 520 363
rect 454 313 470 347
rect 504 327 520 347
rect 574 327 604 463
rect 660 437 690 463
rect 732 431 762 463
rect 732 415 798 431
rect 732 381 748 415
rect 782 381 798 415
rect 732 365 798 381
rect 504 313 648 327
rect 454 297 648 313
rect 376 225 476 255
rect 446 203 476 225
rect 532 203 562 229
rect 618 203 648 297
rect 732 291 762 365
rect 841 317 871 463
rect 927 431 957 463
rect 913 415 979 431
rect 913 381 929 415
rect 963 381 979 415
rect 913 365 979 381
rect 1254 491 1284 517
rect 1476 615 1955 645
rect 2042 619 2072 645
rect 2128 619 2158 645
rect 2214 619 2244 645
rect 2300 619 2330 645
rect 2386 619 2416 645
rect 1064 317 1094 379
rect 690 275 762 291
rect 690 241 712 275
rect 746 241 762 275
rect 827 301 1094 317
rect 827 267 843 301
rect 877 287 1094 301
rect 877 267 914 287
rect 827 251 914 267
rect 690 225 762 241
rect 690 203 720 225
rect 884 131 914 251
rect 1064 227 1094 287
rect 1136 319 1202 335
rect 1136 285 1152 319
rect 1186 305 1202 319
rect 1254 305 1284 407
rect 1359 385 1389 407
rect 1186 285 1284 305
rect 1136 275 1284 285
rect 1326 355 1389 385
rect 1136 269 1247 275
rect 956 205 1022 221
rect 956 171 972 205
rect 1006 171 1022 205
rect 1064 197 1175 227
rect 1145 175 1175 197
rect 1217 175 1247 269
rect 1326 175 1356 355
rect 1476 307 1506 615
rect 1574 541 1604 615
rect 1889 605 1955 615
rect 1889 571 1905 605
rect 1939 571 1955 605
rect 1660 541 1690 567
rect 1889 537 1955 571
rect 1889 503 1905 537
rect 1939 503 1955 537
rect 1889 487 1955 503
rect 1574 431 1604 457
rect 1660 383 1690 457
rect 1852 419 1882 445
rect 1398 277 1506 307
rect 1548 367 1690 383
rect 1548 333 1564 367
rect 1598 333 1690 367
rect 1548 299 1690 333
rect 1398 175 1428 277
rect 1548 265 1564 299
rect 1598 265 1690 299
rect 1548 249 1690 265
rect 1852 313 1882 335
rect 2042 313 2072 367
rect 2128 335 2158 367
rect 2214 335 2244 367
rect 2300 335 2330 367
rect 2386 335 2416 367
rect 1852 283 2072 313
rect 1548 227 1578 249
rect 1852 241 1882 283
rect 1470 197 1578 227
rect 1787 225 1882 241
rect 1470 175 1500 197
rect 1624 175 1654 201
rect 1787 191 1803 225
rect 1837 191 1882 225
rect 2042 217 2072 283
rect 2125 319 2416 335
rect 2125 285 2141 319
rect 2175 285 2209 319
rect 2243 285 2277 319
rect 2311 285 2345 319
rect 2379 285 2416 319
rect 2125 269 2416 285
rect 2128 217 2158 269
rect 2214 217 2244 269
rect 2300 217 2330 269
rect 2386 217 2416 269
rect 956 155 1022 171
rect 956 131 986 155
rect 83 73 113 99
rect 242 51 272 99
rect 446 93 476 119
rect 532 51 562 119
rect 618 93 648 119
rect 690 93 720 119
rect 242 21 562 51
rect 1787 157 1882 191
rect 1787 123 1803 157
rect 1837 123 1882 157
rect 1787 107 1882 123
rect 1326 65 1356 91
rect 1398 65 1428 91
rect 1470 65 1500 91
rect 1624 69 1654 91
rect 1787 69 1817 107
rect 884 21 914 47
rect 956 21 986 47
rect 1145 21 1175 47
rect 1217 21 1247 47
rect 1624 39 1817 69
rect 2042 23 2072 49
rect 2128 23 2158 49
rect 2214 23 2244 49
rect 2300 23 2330 49
rect 2386 23 2416 49
<< polycont >>
rect 216 383 250 417
rect 356 399 390 433
rect 108 289 142 323
rect 216 315 250 349
rect 108 221 142 255
rect 470 313 504 347
rect 748 381 782 415
rect 929 381 963 415
rect 712 241 746 275
rect 843 267 877 301
rect 1152 285 1186 319
rect 972 171 1006 205
rect 1905 571 1939 605
rect 1905 503 1939 537
rect 1564 333 1598 367
rect 1564 265 1598 299
rect 1803 191 1837 225
rect 2141 285 2175 319
rect 2209 285 2243 319
rect 2277 285 2311 319
rect 2345 285 2379 319
rect 1803 123 1837 157
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 34 579 105 595
rect 34 545 65 579
rect 99 545 105 579
rect 34 511 105 545
rect 139 570 205 649
rect 139 536 155 570
rect 189 536 205 570
rect 139 528 205 536
rect 239 578 320 594
rect 239 544 241 578
rect 275 544 320 578
rect 239 528 320 544
rect 34 477 65 511
rect 99 494 105 511
rect 99 477 252 494
rect 34 460 252 477
rect 34 158 72 460
rect 34 124 38 158
rect 34 108 72 124
rect 106 323 163 426
rect 106 289 108 323
rect 142 289 163 323
rect 200 417 252 460
rect 200 383 216 417
rect 250 383 252 417
rect 200 349 252 383
rect 200 315 216 349
rect 250 315 252 349
rect 200 299 252 315
rect 286 349 320 528
rect 427 527 493 649
rect 427 493 443 527
rect 477 493 493 527
rect 427 483 493 493
rect 527 522 573 538
rect 527 488 529 522
rect 563 488 573 522
rect 354 433 468 449
rect 354 399 356 433
rect 390 399 468 433
rect 354 383 468 399
rect 527 417 573 488
rect 607 522 660 538
rect 607 488 615 522
rect 649 488 660 522
rect 607 459 660 488
rect 761 522 827 649
rect 1003 539 1055 649
rect 761 488 777 522
rect 811 488 827 522
rect 761 472 827 488
rect 861 522 932 538
rect 861 488 882 522
rect 916 488 932 522
rect 527 383 590 417
rect 286 347 520 349
rect 286 313 470 347
rect 504 313 520 347
rect 106 255 163 289
rect 106 221 108 255
rect 142 221 163 255
rect 106 76 163 221
rect 286 297 520 313
rect 286 276 363 297
rect 286 242 319 276
rect 353 242 363 276
rect 556 251 590 383
rect 286 187 363 242
rect 479 217 590 251
rect 626 345 660 459
rect 861 465 932 488
rect 1003 505 1019 539
rect 1053 505 1055 539
rect 1003 471 1055 505
rect 861 431 895 465
rect 1003 437 1019 471
rect 1053 437 1055 471
rect 732 415 895 431
rect 732 381 748 415
rect 782 381 895 415
rect 732 379 895 381
rect 929 415 969 431
rect 1003 421 1055 437
rect 1089 609 1469 613
rect 1089 575 1419 609
rect 1453 575 1469 609
rect 1089 573 1469 575
rect 1089 535 1155 573
rect 1089 501 1105 535
rect 1139 501 1155 535
rect 1089 467 1155 501
rect 1089 433 1105 467
rect 1139 433 1155 467
rect 1089 421 1155 433
rect 1193 521 1565 539
rect 1193 505 1529 521
rect 1193 466 1259 505
rect 1513 487 1529 505
rect 1563 487 1565 521
rect 1513 471 1565 487
rect 1599 516 1665 649
rect 1599 482 1615 516
rect 1649 482 1665 516
rect 1599 471 1665 482
rect 1699 516 1767 532
rect 1699 482 1701 516
rect 1735 482 1767 516
rect 1193 432 1209 466
rect 1243 432 1259 466
rect 1193 421 1259 432
rect 1304 455 1359 471
rect 1304 421 1309 455
rect 1343 437 1359 455
rect 1699 437 1767 482
rect 1343 421 1767 437
rect 963 387 969 415
rect 1304 403 1767 421
rect 963 381 1270 387
rect 929 367 1270 381
rect 929 353 1564 367
rect 626 311 893 345
rect 197 158 241 174
rect 231 124 241 158
rect 197 17 241 124
rect 275 158 363 187
rect 275 124 283 158
rect 317 124 363 158
rect 275 108 363 124
rect 397 178 445 194
rect 397 144 401 178
rect 435 144 445 178
rect 397 17 445 144
rect 479 178 530 217
rect 626 183 660 311
rect 827 301 893 311
rect 696 275 762 277
rect 696 241 712 275
rect 746 241 762 275
rect 827 267 843 301
rect 877 267 893 301
rect 827 265 893 267
rect 696 231 762 241
rect 696 197 889 231
rect 479 144 487 178
rect 521 144 530 178
rect 479 128 530 144
rect 564 167 660 183
rect 564 133 573 167
rect 607 133 660 167
rect 564 117 660 133
rect 715 161 781 163
rect 715 127 731 161
rect 765 127 781 161
rect 715 17 781 127
rect 823 107 889 197
rect 929 205 1022 353
rect 1236 333 1564 353
rect 1598 333 1697 367
rect 1074 285 1152 319
rect 1186 285 1202 319
rect 1074 276 1202 285
rect 1074 242 1087 276
rect 1121 242 1202 276
rect 1236 299 1697 333
rect 1236 265 1564 299
rect 1598 265 1697 299
rect 1074 230 1202 242
rect 1731 241 1767 403
rect 1801 394 1853 649
rect 1801 360 1807 394
rect 1841 360 1853 394
rect 1801 344 1853 360
rect 1887 605 1955 615
rect 1887 571 1905 605
rect 1939 571 1955 605
rect 1887 537 1955 571
rect 1887 503 1905 537
rect 1939 503 1955 537
rect 1887 394 1955 503
rect 1887 360 1893 394
rect 1927 360 1955 394
rect 1731 225 1853 241
rect 929 171 972 205
rect 1006 171 1022 205
rect 1242 191 1803 225
rect 1837 191 1853 225
rect 929 156 1022 171
rect 1084 161 1150 177
rect 1084 127 1100 161
rect 1134 127 1150 161
rect 1084 122 1150 127
rect 823 73 839 107
rect 873 73 889 107
rect 823 57 889 73
rect 981 106 1150 122
rect 981 72 997 106
rect 1031 93 1150 106
rect 1031 72 1100 93
rect 981 59 1100 72
rect 1134 59 1150 93
rect 981 17 1150 59
rect 1242 163 1341 191
rect 1242 129 1281 163
rect 1315 129 1341 163
rect 1787 157 1853 191
rect 1242 95 1341 129
rect 1242 61 1258 95
rect 1292 61 1341 95
rect 1242 51 1341 61
rect 1495 148 1629 157
rect 1495 114 1511 148
rect 1545 114 1579 148
rect 1613 114 1629 148
rect 1495 17 1629 114
rect 1663 141 1715 157
rect 1663 107 1665 141
rect 1699 107 1715 141
rect 1787 123 1803 157
rect 1837 123 1853 157
rect 1787 121 1853 123
rect 1663 87 1715 107
rect 1887 87 1955 360
rect 1663 53 1955 87
rect 1989 599 2041 615
rect 1989 565 1997 599
rect 2031 565 2041 599
rect 1989 505 2041 565
rect 1989 471 1997 505
rect 2031 471 2041 505
rect 1989 413 2041 471
rect 1989 379 1997 413
rect 2031 379 2041 413
rect 1989 319 2041 379
rect 2075 607 2126 649
rect 2075 573 2083 607
rect 2117 573 2126 607
rect 2075 507 2126 573
rect 2075 473 2083 507
rect 2117 473 2126 507
rect 2075 409 2126 473
rect 2075 375 2083 409
rect 2117 375 2126 409
rect 2075 359 2126 375
rect 2160 599 2205 615
rect 2160 565 2169 599
rect 2203 565 2205 599
rect 2160 505 2205 565
rect 2160 471 2169 505
rect 2203 471 2205 505
rect 2160 413 2205 471
rect 2239 611 2305 649
rect 2239 577 2255 611
rect 2289 577 2305 611
rect 2239 533 2305 577
rect 2239 499 2255 533
rect 2289 499 2305 533
rect 2239 455 2305 499
rect 2239 421 2255 455
rect 2289 421 2305 455
rect 2339 599 2377 615
rect 2339 565 2341 599
rect 2375 565 2377 599
rect 2339 505 2377 565
rect 2339 471 2341 505
rect 2375 471 2377 505
rect 2160 379 2169 413
rect 2203 387 2205 413
rect 2339 413 2377 471
rect 2411 607 2477 649
rect 2411 573 2427 607
rect 2461 573 2477 607
rect 2411 533 2477 573
rect 2411 499 2427 533
rect 2461 499 2477 533
rect 2411 455 2477 499
rect 2411 421 2427 455
rect 2461 421 2477 455
rect 2339 387 2341 413
rect 2203 379 2341 387
rect 2375 387 2377 413
rect 2375 379 2478 387
rect 2160 353 2478 379
rect 1989 285 2141 319
rect 2175 285 2209 319
rect 2243 285 2277 319
rect 2311 285 2345 319
rect 2379 285 2395 319
rect 1989 205 2040 285
rect 2429 249 2478 353
rect 1989 171 1997 205
rect 2031 171 2040 205
rect 1989 101 2040 171
rect 1989 67 1997 101
rect 2031 67 2040 101
rect 1989 51 2040 67
rect 2074 205 2126 221
rect 2074 171 2083 205
rect 2117 171 2126 205
rect 2074 95 2126 171
rect 2074 61 2083 95
rect 2117 61 2126 95
rect 2074 17 2126 61
rect 2160 215 2478 249
rect 2160 205 2205 215
rect 2160 171 2169 205
rect 2203 171 2205 205
rect 2339 205 2377 215
rect 2160 101 2205 171
rect 2160 67 2169 101
rect 2203 67 2205 101
rect 2160 51 2205 67
rect 2239 147 2255 181
rect 2289 147 2305 181
rect 2239 95 2305 147
rect 2239 61 2255 95
rect 2289 61 2305 95
rect 2239 17 2305 61
rect 2339 171 2341 205
rect 2375 171 2377 205
rect 2339 101 2377 171
rect 2339 67 2341 101
rect 2375 67 2377 101
rect 2339 51 2377 67
rect 2411 147 2427 181
rect 2461 147 2477 181
rect 2411 95 2477 147
rect 2411 61 2427 95
rect 2461 61 2477 95
rect 2411 17 2477 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 319 242 353 276
rect 1087 242 1121 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 683 2496 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 0 617 2496 649
rect 307 276 365 282
rect 307 242 319 276
rect 353 273 365 276
rect 1075 276 1133 282
rect 1075 273 1087 276
rect 353 245 1087 273
rect 353 242 365 245
rect 307 236 365 242
rect 1075 242 1087 245
rect 1121 242 1133 276
rect 1075 236 1133 242
rect 0 17 2496 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
rect 0 -49 2496 -17
<< labels >>
flabel pwell s 0 0 2496 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2496 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel comment s 745 332 745 332 0 FreeSans 200 90 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfstp_4
flabel metal1 s 0 617 2496 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2496 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2431 242 2465 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2496 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 55838
string GDS_START 37570
<< end >>
