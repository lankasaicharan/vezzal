magic
tech sky130A
magscale 1 2
timestamp 1627202622
<< checkpaint >>
rect -1326 -1303 5358 2157
<< nwell >>
rect -66 377 4098 897
rect 3281 344 3619 377
<< pwell >>
rect 39 217 305 241
rect 2292 236 2703 283
rect 947 217 2703 236
rect 3327 251 3585 283
rect 3768 251 4026 317
rect 3327 217 4026 251
rect 39 43 4026 217
rect -26 -43 4058 43
<< mvnmos >>
rect 122 131 222 215
rect 418 107 518 191
rect 560 107 660 191
rect 716 107 816 191
rect 858 107 958 191
rect 1034 126 1134 210
rect 1190 126 1290 210
rect 1469 126 1569 210
rect 1743 126 1843 210
rect 1899 126 1999 210
rect 2041 126 2141 210
rect 2183 126 2283 210
rect 2368 107 2468 257
rect 2524 107 2624 257
rect 2699 107 2799 191
rect 2841 107 2941 191
rect 2998 107 3098 191
rect 3140 107 3240 191
rect 3406 107 3506 257
rect 3672 141 3772 225
rect 3847 141 3947 291
<< mvpmos >>
rect 122 649 222 733
rect 396 655 496 739
rect 538 655 638 739
rect 694 655 794 739
rect 836 655 936 739
rect 1000 655 1100 739
rect 1190 593 1290 743
rect 1716 659 1816 743
rect 1872 659 1972 743
rect 2014 659 2114 743
rect 2170 659 2270 743
rect 1486 449 1586 599
rect 2436 543 2536 743
rect 2592 543 2692 743
rect 2771 543 2871 627
rect 2913 543 3013 627
rect 3069 543 3169 627
rect 3225 543 3325 627
rect 3400 410 3500 710
rect 3666 443 3766 593
rect 3845 443 3945 743
<< mvndiff >>
rect 65 190 122 215
rect 65 156 77 190
rect 111 156 122 190
rect 65 131 122 156
rect 222 190 279 215
rect 2318 210 2368 257
rect 973 191 1034 210
rect 222 156 233 190
rect 267 156 279 190
rect 222 131 279 156
rect 361 166 418 191
rect 361 132 373 166
rect 407 132 418 166
rect 361 107 418 132
rect 518 107 560 191
rect 660 170 716 191
rect 660 136 671 170
rect 705 136 716 170
rect 660 107 716 136
rect 816 107 858 191
rect 958 151 1034 191
rect 958 117 969 151
rect 1003 126 1034 151
rect 1134 183 1190 210
rect 1134 149 1145 183
rect 1179 149 1190 183
rect 1134 126 1190 149
rect 1290 183 1347 210
rect 1290 149 1301 183
rect 1335 149 1347 183
rect 1290 126 1347 149
rect 1412 183 1469 210
rect 1412 149 1424 183
rect 1458 149 1469 183
rect 1412 126 1469 149
rect 1569 183 1626 210
rect 1569 149 1580 183
rect 1614 149 1626 183
rect 1569 126 1626 149
rect 1686 187 1743 210
rect 1686 153 1698 187
rect 1732 153 1743 187
rect 1686 126 1743 153
rect 1843 187 1899 210
rect 1843 153 1854 187
rect 1888 153 1899 187
rect 1843 126 1899 153
rect 1999 126 2041 210
rect 2141 126 2183 210
rect 2283 149 2368 210
rect 2283 126 2311 149
rect 1003 117 1019 126
rect 958 107 1019 117
rect 2298 115 2311 126
rect 2345 115 2368 149
rect 2298 107 2368 115
rect 2468 249 2524 257
rect 2468 215 2479 249
rect 2513 215 2524 249
rect 2468 157 2524 215
rect 2468 123 2479 157
rect 2513 123 2524 157
rect 2468 107 2524 123
rect 2624 243 2677 257
rect 2624 209 2635 243
rect 2669 209 2677 243
rect 2624 191 2677 209
rect 3353 245 3406 257
rect 3353 211 3361 245
rect 3395 211 3406 245
rect 2624 173 2699 191
rect 2624 139 2635 173
rect 2669 139 2699 173
rect 2624 107 2699 139
rect 2799 107 2841 191
rect 2941 164 2998 191
rect 2941 130 2952 164
rect 2986 130 2998 164
rect 2941 107 2998 130
rect 3098 107 3140 191
rect 3240 166 3293 191
rect 3240 132 3251 166
rect 3285 132 3293 166
rect 3240 107 3293 132
rect 3353 153 3406 211
rect 3353 119 3361 153
rect 3395 119 3406 153
rect 3353 107 3406 119
rect 3506 245 3559 257
rect 3506 211 3517 245
rect 3551 211 3559 245
rect 3794 279 3847 291
rect 3794 245 3802 279
rect 3836 245 3847 279
rect 3794 225 3847 245
rect 3506 153 3559 211
rect 3506 119 3517 153
rect 3551 119 3559 153
rect 3619 200 3672 225
rect 3619 166 3627 200
rect 3661 166 3672 200
rect 3619 141 3672 166
rect 3772 187 3847 225
rect 3772 153 3802 187
rect 3836 153 3847 187
rect 3772 141 3847 153
rect 3947 279 4000 291
rect 3947 245 3958 279
rect 3992 245 4000 279
rect 3947 187 4000 245
rect 3947 153 3958 187
rect 3992 153 4000 187
rect 3947 141 4000 153
rect 3506 107 3559 119
<< mvpdiff >>
rect 1133 739 1190 743
rect 65 708 122 733
rect 65 674 77 708
rect 111 674 122 708
rect 65 649 122 674
rect 222 708 279 733
rect 222 674 233 708
rect 267 674 279 708
rect 222 649 279 674
rect 339 714 396 739
rect 339 680 351 714
rect 385 680 396 714
rect 339 655 396 680
rect 496 655 538 739
rect 638 719 694 739
rect 638 685 649 719
rect 683 685 694 719
rect 638 655 694 685
rect 794 655 836 739
rect 936 714 1000 739
rect 936 680 947 714
rect 981 680 1000 714
rect 936 655 1000 680
rect 1100 721 1190 739
rect 1100 687 1145 721
rect 1179 687 1190 721
rect 1100 655 1190 687
rect 1133 593 1190 655
rect 1290 655 1347 743
rect 1659 718 1716 743
rect 1659 684 1671 718
rect 1705 684 1716 718
rect 1659 659 1716 684
rect 1816 718 1872 743
rect 1816 684 1827 718
rect 1861 684 1872 718
rect 1816 659 1872 684
rect 1972 659 2014 743
rect 2114 718 2170 743
rect 2114 684 2125 718
rect 2159 684 2170 718
rect 2114 659 2170 684
rect 2270 718 2323 743
rect 2270 684 2281 718
rect 2315 684 2323 718
rect 2270 659 2323 684
rect 2383 731 2436 743
rect 2383 697 2391 731
rect 2425 697 2436 731
rect 1290 621 1301 655
rect 1335 621 1347 655
rect 1290 593 1347 621
rect 1429 591 1486 599
rect 1429 557 1441 591
rect 1475 557 1486 591
rect 1429 491 1486 557
rect 1429 457 1441 491
rect 1475 457 1486 491
rect 1429 449 1486 457
rect 1586 587 1639 599
rect 1586 553 1597 587
rect 1631 553 1639 587
rect 1586 495 1639 553
rect 1586 461 1597 495
rect 1631 461 1639 495
rect 1586 449 1639 461
rect 2383 653 2436 697
rect 2383 619 2391 653
rect 2425 619 2436 653
rect 2383 543 2436 619
rect 2536 735 2592 743
rect 2536 701 2547 735
rect 2581 701 2592 735
rect 2536 660 2592 701
rect 2536 626 2547 660
rect 2581 626 2592 660
rect 2536 585 2592 626
rect 2536 551 2547 585
rect 2581 551 2592 585
rect 2536 543 2592 551
rect 2692 735 2749 743
rect 2692 701 2703 735
rect 2737 701 2749 735
rect 3788 735 3845 743
rect 2692 627 2749 701
rect 3347 698 3400 710
rect 3347 664 3355 698
rect 3389 664 3400 698
rect 3347 627 3400 664
rect 2692 609 2771 627
rect 2692 575 2703 609
rect 2737 575 2771 609
rect 2692 543 2771 575
rect 2871 543 2913 627
rect 3013 602 3069 627
rect 3013 568 3024 602
rect 3058 568 3069 602
rect 3013 543 3069 568
rect 3169 602 3225 627
rect 3169 568 3180 602
rect 3214 568 3225 602
rect 3169 543 3225 568
rect 3325 623 3400 627
rect 3325 589 3355 623
rect 3389 589 3400 623
rect 3325 546 3400 589
rect 3325 543 3355 546
rect 3347 512 3355 543
rect 3389 512 3400 546
rect 3347 471 3400 512
rect 3347 437 3355 471
rect 3389 437 3400 471
rect 3347 410 3400 437
rect 3500 698 3553 710
rect 3500 664 3511 698
rect 3545 664 3553 698
rect 3500 618 3553 664
rect 3788 701 3800 735
rect 3834 701 3845 735
rect 3788 652 3845 701
rect 3500 584 3511 618
rect 3545 584 3553 618
rect 3788 618 3800 652
rect 3834 618 3845 652
rect 3788 593 3845 618
rect 3500 536 3553 584
rect 3500 502 3511 536
rect 3545 502 3553 536
rect 3500 456 3553 502
rect 3500 422 3511 456
rect 3545 422 3553 456
rect 3613 581 3666 593
rect 3613 547 3621 581
rect 3655 547 3666 581
rect 3613 489 3666 547
rect 3613 455 3621 489
rect 3655 455 3666 489
rect 3613 443 3666 455
rect 3766 568 3845 593
rect 3766 534 3800 568
rect 3834 534 3845 568
rect 3766 485 3845 534
rect 3766 451 3800 485
rect 3834 451 3845 485
rect 3766 443 3845 451
rect 3945 735 4002 743
rect 3945 701 3956 735
rect 3990 701 4002 735
rect 3945 652 4002 701
rect 3945 618 3956 652
rect 3990 618 4002 652
rect 3945 568 4002 618
rect 3945 534 3956 568
rect 3990 534 4002 568
rect 3945 485 4002 534
rect 3945 451 3956 485
rect 3990 451 4002 485
rect 3945 443 4002 451
rect 3500 410 3553 422
<< mvndiffc >>
rect 77 156 111 190
rect 233 156 267 190
rect 373 132 407 166
rect 671 136 705 170
rect 969 117 1003 151
rect 1145 149 1179 183
rect 1301 149 1335 183
rect 1424 149 1458 183
rect 1580 149 1614 183
rect 1698 153 1732 187
rect 1854 153 1888 187
rect 2311 115 2345 149
rect 2479 215 2513 249
rect 2479 123 2513 157
rect 2635 209 2669 243
rect 3361 211 3395 245
rect 2635 139 2669 173
rect 2952 130 2986 164
rect 3251 132 3285 166
rect 3361 119 3395 153
rect 3517 211 3551 245
rect 3802 245 3836 279
rect 3517 119 3551 153
rect 3627 166 3661 200
rect 3802 153 3836 187
rect 3958 245 3992 279
rect 3958 153 3992 187
<< mvpdiffc >>
rect 77 674 111 708
rect 233 674 267 708
rect 351 680 385 714
rect 649 685 683 719
rect 947 680 981 714
rect 1145 687 1179 721
rect 1671 684 1705 718
rect 1827 684 1861 718
rect 2125 684 2159 718
rect 2281 684 2315 718
rect 2391 697 2425 731
rect 1301 621 1335 655
rect 1441 557 1475 591
rect 1441 457 1475 491
rect 1597 553 1631 587
rect 1597 461 1631 495
rect 2391 619 2425 653
rect 2547 701 2581 735
rect 2547 626 2581 660
rect 2547 551 2581 585
rect 2703 701 2737 735
rect 3355 664 3389 698
rect 2703 575 2737 609
rect 3024 568 3058 602
rect 3180 568 3214 602
rect 3355 589 3389 623
rect 3355 512 3389 546
rect 3355 437 3389 471
rect 3511 664 3545 698
rect 3800 701 3834 735
rect 3511 584 3545 618
rect 3800 618 3834 652
rect 3511 502 3545 536
rect 3511 422 3545 456
rect 3621 547 3655 581
rect 3621 455 3655 489
rect 3800 534 3834 568
rect 3800 451 3834 485
rect 3956 701 3990 735
rect 3956 618 3990 652
rect 3956 534 3990 568
rect 3956 451 3990 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4032 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4032 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
rect 3967 797 4001 831
<< poly >>
rect 122 733 222 759
rect 396 739 496 765
rect 538 739 638 765
rect 694 739 794 765
rect 836 739 936 765
rect 1000 739 1100 765
rect 1190 743 1290 769
rect 1716 743 1816 769
rect 1872 743 1972 769
rect 2014 743 2114 769
rect 2170 743 2270 769
rect 2436 743 2536 769
rect 2592 743 2692 769
rect 3845 743 3945 769
rect 122 623 222 649
rect 122 583 354 623
rect 122 549 303 583
rect 337 549 354 583
rect 122 523 354 549
rect 122 377 222 523
rect 122 343 147 377
rect 181 343 222 377
rect 122 309 222 343
rect 122 275 147 309
rect 181 275 222 309
rect 396 427 496 655
rect 538 567 638 655
rect 694 603 794 655
rect 538 533 558 567
rect 592 561 638 567
rect 592 533 700 561
rect 538 513 700 533
rect 396 393 416 427
rect 450 393 496 427
rect 396 359 496 393
rect 396 325 416 359
rect 450 325 496 359
rect 546 443 612 463
rect 546 409 562 443
rect 596 409 612 443
rect 546 375 612 409
rect 546 341 562 375
rect 596 341 612 375
rect 546 325 612 341
rect 654 378 700 513
rect 742 512 794 603
rect 836 567 936 655
rect 836 554 886 567
rect 870 533 886 554
rect 920 533 936 567
rect 1000 633 1100 655
rect 1000 533 1117 633
rect 1716 637 1816 659
rect 1486 599 1586 625
rect 1654 599 1816 637
rect 742 480 808 512
rect 742 446 758 480
rect 792 446 808 480
rect 870 499 936 533
rect 870 465 886 499
rect 920 465 936 499
rect 870 449 936 465
rect 742 426 808 446
rect 654 358 816 378
rect 654 326 736 358
rect 396 305 496 325
rect 122 215 222 275
rect 418 283 496 305
rect 560 284 612 325
rect 710 324 736 326
rect 770 324 816 358
rect 710 290 816 324
rect 418 191 518 283
rect 560 191 660 284
rect 710 256 736 290
rect 770 256 816 290
rect 710 225 816 256
rect 716 191 816 225
rect 858 377 958 397
rect 858 343 891 377
rect 925 343 958 377
rect 858 309 958 343
rect 858 275 891 309
rect 925 275 958 309
rect 858 191 958 275
rect 1014 377 1117 533
rect 1190 508 1290 593
rect 1014 343 1063 377
rect 1097 343 1117 377
rect 1170 488 1290 508
rect 1170 454 1190 488
rect 1224 454 1290 488
rect 1170 420 1290 454
rect 1654 565 1687 599
rect 1721 565 1816 599
rect 1654 538 1816 565
rect 1654 531 1741 538
rect 1654 497 1687 531
rect 1721 497 1741 531
rect 1654 477 1741 497
rect 1872 519 1972 659
rect 2014 637 2114 659
rect 2014 537 2128 637
rect 1872 496 1918 519
rect 1783 485 1918 496
rect 1952 485 1972 519
rect 1783 451 1972 485
rect 1170 386 1190 420
rect 1224 386 1290 420
rect 1170 353 1290 386
rect 1486 355 1586 449
rect 1014 311 1117 343
rect 1014 309 1134 311
rect 1014 275 1063 309
rect 1097 275 1134 309
rect 1014 237 1134 275
rect 1034 210 1134 237
rect 1190 210 1290 353
rect 1469 319 1586 355
rect 1469 285 1489 319
rect 1523 313 1586 319
rect 1783 417 1918 451
rect 1952 417 1972 451
rect 1783 397 1972 417
rect 1783 313 1857 397
rect 2041 393 2128 537
rect 2170 633 2270 659
rect 2170 533 2283 633
rect 3400 710 3500 736
rect 2771 627 2871 653
rect 2913 627 3013 653
rect 3069 627 3169 653
rect 3225 627 3325 653
rect 2183 427 2283 533
rect 2436 517 2536 543
rect 2592 517 2692 543
rect 2183 393 2199 427
rect 2233 393 2283 427
rect 2335 495 2536 517
rect 2335 461 2355 495
rect 2389 461 2536 495
rect 2335 417 2536 461
rect 2578 469 2722 517
rect 2578 435 2594 469
rect 2628 435 2722 469
rect 2771 495 2871 543
rect 2771 461 2820 495
rect 2854 461 2871 495
rect 2771 441 2871 461
rect 2913 521 3013 543
rect 3069 521 3169 543
rect 2913 495 3026 521
rect 2913 461 2976 495
rect 3010 461 3026 495
rect 2913 445 3026 461
rect 2041 373 2141 393
rect 1523 285 1857 313
rect 1469 225 1857 285
rect 1899 305 1999 355
rect 1899 271 1945 305
rect 1979 271 1999 305
rect 1469 210 1569 225
rect 1743 210 1843 225
rect 1899 210 1999 271
rect 2041 339 2061 373
rect 2095 339 2141 373
rect 2041 305 2141 339
rect 2041 271 2061 305
rect 2095 271 2141 305
rect 2041 210 2141 271
rect 2183 359 2283 393
rect 2183 325 2199 359
rect 2233 325 2283 359
rect 2183 210 2283 325
rect 2368 257 2468 417
rect 2578 399 2722 435
rect 2524 329 2635 357
rect 2677 347 2799 399
rect 2524 295 2581 329
rect 2615 295 2635 329
rect 2524 279 2635 295
rect 2524 257 2624 279
rect 122 105 222 131
rect 418 81 518 107
rect 560 81 660 107
rect 716 81 816 107
rect 858 81 958 107
rect 1034 58 1134 126
rect 1190 100 1290 126
rect 1469 100 1569 126
rect 1743 100 1843 126
rect 1899 100 1999 126
rect 2041 100 2141 126
rect 2183 58 2283 126
rect 2692 217 2799 347
rect 2913 313 2956 445
rect 3068 421 3169 521
rect 3068 403 3098 421
rect 2699 191 2799 217
rect 2841 213 2956 313
rect 2998 387 3098 403
rect 2998 353 3018 387
rect 3052 353 3098 387
rect 3225 384 3325 543
rect 3666 593 3766 619
rect 3666 417 3766 443
rect 3845 417 3945 443
rect 3400 384 3500 410
rect 3666 384 3772 417
rect 3225 379 3772 384
rect 2998 319 3098 353
rect 2998 285 3018 319
rect 3052 285 3098 319
rect 2841 191 2941 213
rect 2998 191 3098 285
rect 3140 331 3772 379
rect 3140 297 3189 331
rect 3223 297 3772 331
rect 3834 381 3947 417
rect 3834 347 3854 381
rect 3888 347 3947 381
rect 3834 317 3947 347
rect 3140 279 3772 297
rect 3847 291 3947 317
rect 3140 263 3243 279
rect 3140 229 3189 263
rect 3223 229 3243 263
rect 3406 257 3506 279
rect 3140 213 3243 229
rect 3140 191 3240 213
rect 3672 225 3772 279
rect 3672 115 3772 141
rect 3847 115 3947 141
rect 2368 81 2468 107
rect 2524 81 2624 107
rect 2699 81 2799 107
rect 2841 81 2941 107
rect 2998 81 3098 107
rect 3140 81 3240 107
rect 3406 81 3506 107
rect 1034 28 2283 58
<< polycont >>
rect 303 549 337 583
rect 147 343 181 377
rect 147 275 181 309
rect 558 533 592 567
rect 416 393 450 427
rect 416 325 450 359
rect 562 409 596 443
rect 562 341 596 375
rect 886 533 920 567
rect 758 446 792 480
rect 886 465 920 499
rect 736 324 770 358
rect 736 256 770 290
rect 891 343 925 377
rect 891 275 925 309
rect 1063 343 1097 377
rect 1190 454 1224 488
rect 1687 565 1721 599
rect 1687 497 1721 531
rect 1918 485 1952 519
rect 1190 386 1224 420
rect 1063 275 1097 309
rect 1489 285 1523 319
rect 1918 417 1952 451
rect 2199 393 2233 427
rect 2355 461 2389 495
rect 2594 435 2628 469
rect 2820 461 2854 495
rect 2976 461 3010 495
rect 1945 271 1979 305
rect 2061 339 2095 373
rect 2061 271 2095 305
rect 2199 325 2233 359
rect 2581 295 2615 329
rect 3018 353 3052 387
rect 3018 285 3052 319
rect 3189 297 3223 331
rect 3854 347 3888 381
rect 3189 229 3223 263
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4032 831
rect 18 735 197 741
rect 18 701 19 735
rect 53 708 91 735
rect 53 701 77 708
rect 125 701 163 735
rect 18 674 77 701
rect 111 674 197 701
rect 18 641 197 674
rect 233 708 283 741
rect 267 674 283 708
rect 233 641 283 674
rect 335 714 423 747
rect 335 680 351 714
rect 385 680 423 714
rect 335 647 423 680
rect 509 735 699 747
rect 509 701 515 735
rect 549 701 587 735
rect 621 719 659 735
rect 621 701 649 719
rect 693 701 699 735
rect 509 685 649 701
rect 683 685 699 701
rect 509 673 699 685
rect 931 714 981 747
rect 931 680 947 714
rect 233 497 267 641
rect 389 637 423 647
rect 931 637 981 680
rect 1017 735 1195 751
rect 1051 701 1089 735
rect 1123 721 1161 735
rect 1123 701 1145 721
rect 1017 687 1145 701
rect 1179 687 1195 701
rect 1017 673 1195 687
rect 1231 727 1405 761
rect 1231 637 1265 727
rect 389 603 1265 637
rect 1301 655 1335 691
rect 303 583 353 599
rect 337 567 353 583
rect 337 549 558 567
rect 303 533 558 549
rect 592 533 608 567
rect 654 533 886 567
rect 920 533 936 567
rect 654 497 688 533
rect 233 463 688 497
rect 870 499 936 533
rect 742 480 808 496
rect 131 377 197 393
rect 131 343 147 377
rect 181 343 197 377
rect 131 309 197 343
rect 131 275 147 309
rect 181 275 197 309
rect 131 259 197 275
rect 18 190 127 223
rect 18 156 77 190
rect 111 156 127 190
rect 18 113 127 156
rect 18 79 19 113
rect 53 79 91 113
rect 125 79 127 113
rect 18 73 127 79
rect 163 87 197 259
rect 233 190 267 463
rect 546 443 612 463
rect 313 393 416 427
rect 450 393 466 427
rect 313 359 466 393
rect 313 325 416 359
rect 450 325 466 359
rect 546 409 562 443
rect 596 409 612 443
rect 546 375 612 409
rect 742 446 758 480
rect 792 446 808 480
rect 870 465 886 499
rect 920 465 936 499
rect 742 431 808 446
rect 742 395 941 431
rect 546 341 562 375
rect 596 341 612 375
rect 875 377 941 395
rect 546 325 612 341
rect 697 358 839 359
rect 697 324 736 358
rect 770 324 839 358
rect 697 290 839 324
rect 697 289 736 290
rect 233 123 267 156
rect 303 256 736 289
rect 770 256 839 290
rect 875 343 891 377
rect 925 343 941 377
rect 875 309 941 343
rect 875 275 891 309
rect 925 275 941 309
rect 875 259 941 275
rect 303 255 839 256
rect 303 87 337 255
rect 977 219 1011 603
rect 1174 488 1240 504
rect 1174 454 1190 488
rect 1224 454 1240 488
rect 1047 424 1127 430
rect 1047 390 1087 424
rect 1121 390 1127 424
rect 1047 377 1127 390
rect 1047 343 1063 377
rect 1097 343 1127 377
rect 1174 420 1240 454
rect 1174 386 1190 420
rect 1224 386 1240 420
rect 1174 370 1240 386
rect 1047 309 1127 343
rect 1047 275 1063 309
rect 1097 275 1127 309
rect 1047 259 1127 275
rect 1301 335 1335 621
rect 1371 405 1405 727
rect 1441 735 1475 741
rect 1441 591 1475 701
rect 1655 718 1721 751
rect 1655 685 1671 718
rect 1441 491 1475 557
rect 1441 441 1475 457
rect 1511 684 1671 685
rect 1705 685 1721 718
rect 1827 718 1877 751
rect 1705 684 1791 685
rect 1511 651 1791 684
rect 1511 405 1545 651
rect 1671 603 1721 615
rect 1371 371 1545 405
rect 1581 599 1721 603
rect 1581 587 1687 599
rect 1581 553 1597 587
rect 1631 565 1687 587
rect 1631 553 1721 565
rect 1581 531 1721 553
rect 1581 497 1687 531
rect 1581 495 1721 497
rect 1581 461 1597 495
rect 1631 461 1721 495
rect 1581 445 1721 461
rect 1301 319 1539 335
rect 1301 301 1489 319
rect 163 53 337 87
rect 373 166 423 199
rect 407 132 423 166
rect 373 87 423 132
rect 655 185 1011 219
rect 655 170 721 185
rect 655 136 671 170
rect 705 136 721 170
rect 1055 183 1245 199
rect 655 123 721 136
rect 953 117 969 151
rect 1003 117 1019 151
rect 953 87 1019 117
rect 373 53 1019 87
rect 1055 149 1145 183
rect 1179 149 1245 183
rect 1055 113 1245 149
rect 1055 79 1061 113
rect 1095 79 1133 113
rect 1167 79 1205 113
rect 1239 79 1245 113
rect 1301 183 1335 301
rect 1473 285 1489 301
rect 1523 285 1539 319
rect 1473 269 1539 285
rect 1581 199 1630 445
rect 1757 199 1791 651
rect 1580 183 1630 199
rect 1301 99 1335 149
rect 1374 149 1424 183
rect 1458 149 1544 183
rect 1374 113 1544 149
rect 1055 73 1245 79
rect 1374 79 1390 113
rect 1424 79 1494 113
rect 1528 79 1544 113
rect 1374 73 1544 79
rect 1614 149 1630 183
rect 1580 87 1630 149
rect 1682 187 1791 199
rect 1682 153 1698 187
rect 1732 153 1791 187
rect 1682 123 1791 153
rect 1861 684 1877 718
rect 1827 615 1877 684
rect 1985 735 2175 751
rect 1985 701 1991 735
rect 2025 701 2063 735
rect 2097 718 2135 735
rect 2097 701 2125 718
rect 2169 701 2175 735
rect 1985 684 2125 701
rect 2159 684 2175 701
rect 1985 651 2175 684
rect 2265 718 2355 747
rect 2265 684 2281 718
rect 2315 684 2355 718
rect 2265 615 2355 684
rect 1827 581 2355 615
rect 2391 735 2509 747
rect 2391 731 2397 735
rect 2431 701 2469 735
rect 2503 701 2509 735
rect 2425 697 2509 701
rect 2391 653 2509 697
rect 2425 619 2509 653
rect 2391 603 2509 619
rect 2547 735 2597 751
rect 2581 701 2597 735
rect 2547 660 2597 701
rect 2581 626 2597 660
rect 1827 199 1861 581
rect 2265 567 2355 581
rect 2547 585 2597 626
rect 1902 519 1968 535
rect 2265 533 2389 567
rect 1902 485 1918 519
rect 1952 497 1968 519
rect 1952 485 2319 497
rect 1902 463 2319 485
rect 1902 451 1968 463
rect 1902 417 1918 451
rect 1952 417 1968 451
rect 1902 401 1968 417
rect 2137 424 2199 427
rect 2137 390 2143 424
rect 2177 393 2199 424
rect 2233 393 2249 427
rect 2177 390 2249 393
rect 2045 373 2101 389
rect 1940 305 1995 351
rect 1940 271 1945 305
rect 1979 271 1995 305
rect 1940 219 1995 271
rect 2045 339 2061 373
rect 2095 339 2101 373
rect 2045 305 2101 339
rect 2137 359 2249 390
rect 2285 409 2319 463
rect 2355 495 2389 533
rect 2581 551 2597 585
rect 2687 735 2753 751
rect 2687 701 2703 735
rect 2737 701 2753 735
rect 2687 609 2753 701
rect 2960 735 3144 741
rect 2960 701 2963 735
rect 2997 701 3035 735
rect 3069 701 3107 735
rect 3141 701 3144 735
rect 2687 575 2703 609
rect 2737 575 2924 609
rect 2547 539 2597 551
rect 2547 505 2714 539
rect 2355 445 2389 461
rect 2425 435 2594 469
rect 2628 435 2644 469
rect 2425 409 2459 435
rect 2285 375 2459 409
rect 2680 399 2714 505
rect 2137 325 2199 359
rect 2233 325 2249 359
rect 2495 365 2714 399
rect 2045 271 2061 305
rect 2095 289 2101 305
rect 2495 289 2529 365
rect 2095 271 2529 289
rect 2045 255 2529 271
rect 2463 249 2529 255
rect 1827 187 1904 199
rect 1827 153 1854 187
rect 1888 153 1904 187
rect 1827 123 1904 153
rect 1940 185 2429 219
rect 1940 87 1995 185
rect 1580 53 1995 87
rect 2154 115 2311 149
rect 2345 115 2361 149
rect 2154 113 2361 115
rect 2154 79 2160 113
rect 2194 79 2232 113
rect 2266 79 2304 113
rect 2338 79 2361 113
rect 2154 73 2361 79
rect 2395 87 2429 185
rect 2463 215 2479 249
rect 2513 215 2529 249
rect 2463 157 2529 215
rect 2463 123 2479 157
rect 2513 123 2529 157
rect 2565 295 2581 329
rect 2615 295 2631 329
rect 2565 87 2599 295
rect 2750 259 2784 575
rect 2635 243 2784 259
rect 2669 225 2784 243
rect 2820 495 2854 511
rect 2669 209 2685 225
rect 2635 173 2685 209
rect 2669 139 2685 173
rect 2635 123 2685 139
rect 2820 87 2854 461
rect 2890 249 2924 575
rect 2960 602 3144 701
rect 3266 735 3451 741
rect 3266 701 3269 735
rect 3303 701 3341 735
rect 3375 701 3413 735
rect 3447 701 3451 735
rect 3707 735 3897 751
rect 3266 698 3451 701
rect 3266 664 3355 698
rect 3389 664 3451 698
rect 2960 568 3024 602
rect 3058 568 3144 602
rect 2960 535 3144 568
rect 3180 602 3230 635
rect 3214 568 3230 602
rect 3180 499 3230 568
rect 2960 495 3230 499
rect 2960 461 2976 495
rect 3010 461 3230 495
rect 2960 460 3230 461
rect 3001 390 3007 424
rect 3041 390 3137 424
rect 3001 387 3137 390
rect 3001 353 3018 387
rect 3052 353 3137 387
rect 3196 401 3230 460
rect 3266 623 3451 664
rect 3266 589 3355 623
rect 3389 589 3451 623
rect 3266 546 3451 589
rect 3266 512 3355 546
rect 3389 512 3451 546
rect 3266 471 3451 512
rect 3266 437 3355 471
rect 3389 437 3451 471
rect 3487 698 3567 714
rect 3487 664 3511 698
rect 3545 664 3567 698
rect 3487 618 3567 664
rect 3487 584 3511 618
rect 3545 584 3567 618
rect 3707 701 3713 735
rect 3747 701 3785 735
rect 3834 701 3857 735
rect 3891 701 3897 735
rect 3707 652 3897 701
rect 3707 618 3800 652
rect 3834 618 3897 652
rect 3487 536 3567 584
rect 3487 502 3511 536
rect 3545 502 3567 536
rect 3487 456 3567 502
rect 3487 422 3511 456
rect 3545 422 3567 456
rect 3196 367 3309 401
rect 3001 319 3137 353
rect 3001 285 3018 319
rect 3052 285 3137 319
rect 3173 297 3189 331
rect 3223 297 3239 331
rect 3173 263 3239 297
rect 3173 249 3189 263
rect 2890 229 3189 249
rect 3223 229 3239 263
rect 2890 215 3239 229
rect 3275 179 3309 367
rect 2395 53 2854 87
rect 2890 164 3080 179
rect 2890 130 2952 164
rect 2986 130 3080 164
rect 2890 113 3080 130
rect 2890 79 2896 113
rect 2930 79 2968 113
rect 3002 79 3040 113
rect 3074 79 3080 113
rect 3235 166 3309 179
rect 3235 132 3251 166
rect 3285 132 3309 166
rect 3235 103 3309 132
rect 3345 245 3451 261
rect 3345 211 3361 245
rect 3395 211 3451 245
rect 3345 153 3451 211
rect 3345 119 3361 153
rect 3395 119 3451 153
rect 3345 113 3451 119
rect 2890 73 3080 79
rect 3379 79 3417 113
rect 3487 245 3567 422
rect 3487 211 3517 245
rect 3551 211 3567 245
rect 3487 153 3567 211
rect 3487 119 3517 153
rect 3551 119 3567 153
rect 3605 581 3671 597
rect 3605 547 3621 581
rect 3655 547 3671 581
rect 3605 489 3671 547
rect 3605 455 3621 489
rect 3655 455 3671 489
rect 3605 397 3671 455
rect 3707 568 3897 618
rect 3707 534 3800 568
rect 3834 534 3897 568
rect 3707 485 3897 534
rect 3707 451 3800 485
rect 3834 451 3897 485
rect 3707 435 3897 451
rect 3940 735 4008 751
rect 3940 701 3956 735
rect 3990 701 4008 735
rect 3940 652 4008 701
rect 3940 618 3956 652
rect 3990 618 4008 652
rect 3940 568 4008 618
rect 3940 534 3956 568
rect 3990 534 4008 568
rect 3940 485 4008 534
rect 3940 451 3956 485
rect 3990 451 4008 485
rect 3605 381 3904 397
rect 3605 347 3854 381
rect 3888 347 3904 381
rect 3605 331 3904 347
rect 3605 200 3677 331
rect 3605 166 3627 200
rect 3661 166 3677 200
rect 3605 137 3677 166
rect 3713 279 3903 295
rect 3713 245 3802 279
rect 3836 245 3903 279
rect 3713 187 3903 245
rect 3713 153 3802 187
rect 3836 153 3903 187
rect 3487 103 3567 119
rect 3713 113 3903 153
rect 3940 279 4008 451
rect 3940 245 3958 279
rect 3992 245 4008 279
rect 3940 187 4008 245
rect 3940 153 3958 187
rect 3992 153 4008 187
rect 3940 137 4008 153
rect 3345 73 3451 79
rect 3713 79 3719 113
rect 3753 79 3791 113
rect 3825 79 3863 113
rect 3897 79 3903 113
rect 3713 73 3903 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4032 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
rect 3967 797 4001 831
rect 19 701 53 735
rect 91 708 125 735
rect 91 701 111 708
rect 111 701 125 708
rect 163 701 197 735
rect 515 701 549 735
rect 587 701 621 735
rect 659 719 693 735
rect 659 701 683 719
rect 683 701 693 719
rect 1017 701 1051 735
rect 1089 701 1123 735
rect 1161 721 1195 735
rect 1161 701 1179 721
rect 1179 701 1195 721
rect 19 79 53 113
rect 91 79 125 113
rect 1087 390 1121 424
rect 1441 701 1475 735
rect 1061 79 1095 113
rect 1133 79 1167 113
rect 1205 79 1239 113
rect 1390 79 1424 113
rect 1494 79 1528 113
rect 1991 701 2025 735
rect 2063 701 2097 735
rect 2135 718 2169 735
rect 2135 701 2159 718
rect 2159 701 2169 718
rect 2397 731 2431 735
rect 2397 701 2425 731
rect 2425 701 2431 731
rect 2469 701 2503 735
rect 2143 390 2177 424
rect 2963 701 2997 735
rect 3035 701 3069 735
rect 3107 701 3141 735
rect 2160 79 2194 113
rect 2232 79 2266 113
rect 2304 79 2338 113
rect 3269 701 3303 735
rect 3341 701 3375 735
rect 3413 701 3447 735
rect 3007 390 3041 424
rect 3713 701 3747 735
rect 3785 701 3800 735
rect 3800 701 3819 735
rect 3857 701 3891 735
rect 2896 79 2930 113
rect 2968 79 3002 113
rect 3040 79 3074 113
rect 3345 79 3379 113
rect 3417 79 3451 113
rect 3719 79 3753 113
rect 3791 79 3825 113
rect 3863 79 3897 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
<< metal1 >>
rect 0 831 4032 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4032 831
rect 0 791 4032 797
rect 0 735 4032 763
rect 0 701 19 735
rect 53 701 91 735
rect 125 701 163 735
rect 197 701 515 735
rect 549 701 587 735
rect 621 701 659 735
rect 693 701 1017 735
rect 1051 701 1089 735
rect 1123 701 1161 735
rect 1195 701 1441 735
rect 1475 701 1991 735
rect 2025 701 2063 735
rect 2097 701 2135 735
rect 2169 701 2397 735
rect 2431 701 2469 735
rect 2503 701 2963 735
rect 2997 701 3035 735
rect 3069 701 3107 735
rect 3141 701 3269 735
rect 3303 701 3341 735
rect 3375 701 3413 735
rect 3447 701 3713 735
rect 3747 701 3785 735
rect 3819 701 3857 735
rect 3891 701 4032 735
rect 0 689 4032 701
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1121 393 2143 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 2131 390 2143 393
rect 2177 421 2189 424
rect 2995 424 3053 430
rect 2995 421 3007 424
rect 2177 393 3007 421
rect 2177 390 2189 393
rect 2131 384 2189 390
rect 2995 390 3007 393
rect 3041 390 3053 424
rect 2995 384 3053 390
rect 0 113 4032 125
rect 0 79 19 113
rect 53 79 91 113
rect 125 79 1061 113
rect 1095 79 1133 113
rect 1167 79 1205 113
rect 1239 79 1390 113
rect 1424 79 1494 113
rect 1528 79 2160 113
rect 2194 79 2232 113
rect 2266 79 2304 113
rect 2338 79 2896 113
rect 2930 79 2968 113
rect 3002 79 3040 113
rect 3074 79 3345 113
rect 3379 79 3417 113
rect 3451 79 3719 113
rect 3753 79 3791 113
rect 3825 79 3863 113
rect 3897 79 4032 113
rect 0 51 4032 79
rect 0 17 4032 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4032 17
rect 0 -23 4032 -17
<< labels >>
flabel comment s 678 453 678 453 0 FreeSans 200 90 0 0 no_jumper_check
flabel comment s 182 498 182 498 0 FreeSans 200 90 0 0 no_jumper_check
flabel comment s 1700 286 1700 286 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfrbp_1
flabel comment s 1623 43 1623 43 0 FreeSans 300 0 0 0 no_jumper_check
flabel metal1 s 0 51 4032 125 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 0 0 4032 23 0 FreeSans 340 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 0 689 4032 763 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 791 4032 814 0 FreeSans 340 0 0 0 VPB
port 8 nsew power bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 3007 390 3041 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 3103 390 3137 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 1183 464 1217 498 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 3967 168 4001 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 242 4001 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 316 4001 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 390 4001 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 464 4001 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 538 4001 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3967 612 4001 646 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 3487 168 3521 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 242 3521 276 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 316 3521 350 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 390 3521 424 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 464 3521 498 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 538 3521 572 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3487 612 3521 646 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
rlabel viali s 3007 390 3041 424 1 RESET_B
port 3 nsew signal input
rlabel locali s 3001 285 3137 424 1 RESET_B
port 3 nsew signal input
rlabel metal1 s 2995 421 3053 430 1 RESET_B
port 3 nsew signal input
rlabel metal1 s 2995 384 3053 393 1 RESET_B
port 3 nsew signal input
rlabel metal1 s 2131 421 2189 430 1 RESET_B
port 3 nsew signal input
rlabel metal1 s 2131 384 2189 393 1 RESET_B
port 3 nsew signal input
rlabel metal1 s 1075 421 1133 430 1 RESET_B
port 3 nsew signal input
rlabel metal1 s 1075 393 3053 421 1 RESET_B
port 3 nsew signal input
rlabel metal1 s 1075 384 1133 393 1 RESET_B
port 3 nsew signal input
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 4032 814
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string LEFsymmetry X Y
string GDS_END 1105218
string GDS_START 1071124
<< end >>
