magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 80 49 556 192
rect 0 0 576 49
<< scnmos >>
rect 159 82 189 166
rect 231 82 261 166
rect 303 82 333 166
rect 447 82 477 166
<< scpmoshvt >>
rect 139 500 169 584
rect 225 500 255 584
rect 311 500 341 584
rect 397 500 427 584
<< ndiff >>
rect 106 128 159 166
rect 106 94 114 128
rect 148 94 159 128
rect 106 82 159 94
rect 189 82 231 166
rect 261 82 303 166
rect 333 154 447 166
rect 333 120 398 154
rect 432 120 447 154
rect 333 82 447 120
rect 477 128 530 166
rect 477 94 488 128
rect 522 94 530 128
rect 477 82 530 94
<< pdiff >>
rect 86 572 139 584
rect 86 538 94 572
rect 128 538 139 572
rect 86 500 139 538
rect 169 542 225 584
rect 169 508 180 542
rect 214 508 225 542
rect 169 500 225 508
rect 255 576 311 584
rect 255 542 266 576
rect 300 542 311 576
rect 255 500 311 542
rect 341 542 397 584
rect 341 508 352 542
rect 386 508 397 542
rect 341 500 397 508
rect 427 546 480 584
rect 427 512 438 546
rect 472 512 480 546
rect 427 500 480 512
<< ndiffc >>
rect 114 94 148 128
rect 398 120 432 154
rect 488 94 522 128
<< pdiffc >>
rect 94 538 128 572
rect 180 508 214 542
rect 266 542 300 576
rect 352 508 386 542
rect 438 512 472 546
<< poly >>
rect 139 584 169 610
rect 225 584 255 610
rect 311 584 341 610
rect 397 584 427 610
rect 139 478 169 500
rect 57 448 169 478
rect 57 322 87 448
rect 225 400 255 500
rect 311 400 341 500
rect 397 478 427 500
rect 397 448 447 478
rect 21 306 87 322
rect 21 272 37 306
rect 71 272 87 306
rect 21 238 87 272
rect 195 384 261 400
rect 195 350 211 384
rect 245 350 261 384
rect 195 316 261 350
rect 195 282 211 316
rect 245 282 261 316
rect 195 266 261 282
rect 21 204 37 238
rect 71 218 87 238
rect 71 204 189 218
rect 21 188 189 204
rect 159 166 189 188
rect 231 166 261 266
rect 303 384 369 400
rect 303 350 319 384
rect 353 350 369 384
rect 417 376 447 448
rect 303 316 369 350
rect 303 282 319 316
rect 353 282 369 316
rect 303 266 369 282
rect 411 360 477 376
rect 411 326 427 360
rect 461 326 477 360
rect 411 292 477 326
rect 303 166 333 266
rect 411 258 427 292
rect 461 258 477 292
rect 411 242 477 258
rect 447 166 477 242
rect 159 56 189 82
rect 231 56 261 82
rect 303 56 333 82
rect 447 56 477 82
<< polycont >>
rect 37 272 71 306
rect 211 350 245 384
rect 211 282 245 316
rect 37 204 71 238
rect 319 350 353 384
rect 319 282 353 316
rect 427 326 461 360
rect 427 258 461 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 78 572 144 649
rect 78 538 94 572
rect 128 538 144 572
rect 250 576 316 649
rect 78 534 144 538
rect 180 542 214 558
rect 250 542 266 576
rect 300 542 316 576
rect 250 538 316 542
rect 352 542 390 558
rect 180 502 214 508
rect 386 508 390 542
rect 352 502 390 508
rect 31 306 71 498
rect 180 468 390 502
rect 434 546 545 562
rect 434 512 438 546
rect 472 512 545 546
rect 434 496 545 512
rect 31 272 37 306
rect 31 238 71 272
rect 31 204 37 238
rect 31 168 71 204
rect 211 384 257 424
rect 245 350 257 384
rect 211 316 257 350
rect 245 282 257 316
rect 98 128 164 132
rect 98 94 114 128
rect 148 94 164 128
rect 211 94 257 282
rect 319 384 353 424
rect 319 316 353 350
rect 319 94 353 282
rect 415 376 449 424
rect 415 360 461 376
rect 415 326 427 360
rect 415 292 461 326
rect 415 258 427 292
rect 415 242 461 258
rect 511 202 545 496
rect 394 168 545 202
rect 394 154 436 168
rect 394 120 398 154
rect 432 120 436 154
rect 394 104 436 120
rect 472 128 538 132
rect 472 94 488 128
rect 522 94 538 128
rect 98 17 164 94
rect 472 17 538 94
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a31oi_m
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3462606
string GDS_START 3455702
<< end >>
