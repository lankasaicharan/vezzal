magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 1 49 1999 241
rect 0 0 2016 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 252 47 282 215
rect 338 47 368 215
rect 424 47 454 215
rect 510 47 540 215
rect 596 47 626 215
rect 682 47 712 215
rect 872 47 902 215
rect 958 47 988 215
rect 1044 47 1074 215
rect 1130 47 1160 215
rect 1216 47 1246 215
rect 1302 47 1332 215
rect 1388 47 1418 215
rect 1474 47 1504 215
rect 1632 47 1662 215
rect 1718 47 1748 215
rect 1804 47 1834 215
rect 1890 47 1920 215
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 252 367 282 619
rect 338 367 368 619
rect 424 367 454 619
rect 510 367 540 619
rect 596 367 626 619
rect 682 367 712 619
rect 836 367 866 619
rect 922 367 952 619
rect 1008 367 1038 619
rect 1094 367 1124 619
rect 1180 367 1210 619
rect 1266 367 1296 619
rect 1352 367 1382 619
rect 1438 367 1468 619
rect 1628 367 1658 619
rect 1714 367 1744 619
rect 1800 367 1830 619
rect 1886 367 1916 619
<< ndiff >>
rect 27 163 80 215
rect 27 129 35 163
rect 69 129 80 163
rect 27 93 80 129
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 190 166 215
rect 110 156 121 190
rect 155 156 166 190
rect 110 47 166 156
rect 196 97 252 215
rect 196 63 207 97
rect 241 63 252 97
rect 196 47 252 63
rect 282 190 338 215
rect 282 156 293 190
rect 327 156 338 190
rect 282 47 338 156
rect 368 199 424 215
rect 368 165 379 199
rect 413 165 424 199
rect 368 101 424 165
rect 368 67 379 101
rect 413 67 424 101
rect 368 47 424 67
rect 454 163 510 215
rect 454 129 465 163
rect 499 129 510 163
rect 454 93 510 129
rect 454 59 465 93
rect 499 59 510 93
rect 454 47 510 59
rect 540 181 596 215
rect 540 147 551 181
rect 585 147 596 181
rect 540 47 596 147
rect 626 93 682 215
rect 626 59 637 93
rect 671 59 682 93
rect 626 47 682 59
rect 712 181 765 215
rect 712 147 723 181
rect 757 147 765 181
rect 712 47 765 147
rect 819 181 872 215
rect 819 147 827 181
rect 861 147 872 181
rect 819 47 872 147
rect 902 169 958 215
rect 902 135 913 169
rect 947 135 958 169
rect 902 93 958 135
rect 902 59 913 93
rect 947 59 958 93
rect 902 47 958 59
rect 988 169 1044 215
rect 988 135 999 169
rect 1033 135 1044 169
rect 988 47 1044 135
rect 1074 169 1130 215
rect 1074 135 1085 169
rect 1119 135 1130 169
rect 1074 93 1130 135
rect 1074 59 1085 93
rect 1119 59 1130 93
rect 1074 47 1130 59
rect 1160 203 1216 215
rect 1160 169 1171 203
rect 1205 169 1216 203
rect 1160 101 1216 169
rect 1160 67 1171 101
rect 1205 67 1216 101
rect 1160 47 1216 67
rect 1246 169 1302 215
rect 1246 135 1257 169
rect 1291 135 1302 169
rect 1246 93 1302 135
rect 1246 59 1257 93
rect 1291 59 1302 93
rect 1246 47 1302 59
rect 1332 203 1388 215
rect 1332 169 1343 203
rect 1377 169 1388 203
rect 1332 101 1388 169
rect 1332 67 1343 101
rect 1377 67 1388 101
rect 1332 47 1388 67
rect 1418 132 1474 215
rect 1418 98 1429 132
rect 1463 98 1474 132
rect 1418 47 1474 98
rect 1504 207 1632 215
rect 1504 173 1515 207
rect 1549 203 1632 207
rect 1549 173 1587 203
rect 1504 169 1587 173
rect 1621 169 1632 203
rect 1504 101 1632 169
rect 1504 67 1515 101
rect 1549 67 1587 101
rect 1621 67 1632 101
rect 1504 47 1632 67
rect 1662 167 1718 215
rect 1662 133 1673 167
rect 1707 133 1718 167
rect 1662 93 1718 133
rect 1662 59 1673 93
rect 1707 59 1718 93
rect 1662 47 1718 59
rect 1748 203 1804 215
rect 1748 169 1759 203
rect 1793 169 1804 203
rect 1748 101 1804 169
rect 1748 67 1759 101
rect 1793 67 1804 101
rect 1748 47 1804 67
rect 1834 167 1890 215
rect 1834 133 1845 167
rect 1879 133 1890 167
rect 1834 93 1890 133
rect 1834 59 1845 93
rect 1879 59 1890 93
rect 1834 47 1890 59
rect 1920 203 1973 215
rect 1920 169 1931 203
rect 1965 169 1973 203
rect 1920 101 1973 169
rect 1920 67 1931 101
rect 1965 67 1973 101
rect 1920 47 1973 67
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 504 80 565
rect 27 470 35 504
rect 69 470 80 504
rect 27 413 80 470
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 607 166 619
rect 110 573 121 607
rect 155 573 166 607
rect 110 520 166 573
rect 110 486 121 520
rect 155 486 166 520
rect 110 437 166 486
rect 110 403 121 437
rect 155 403 166 437
rect 110 367 166 403
rect 196 599 252 619
rect 196 565 207 599
rect 241 565 252 599
rect 196 504 252 565
rect 196 470 207 504
rect 241 470 252 504
rect 196 413 252 470
rect 196 379 207 413
rect 241 379 252 413
rect 196 367 252 379
rect 282 607 338 619
rect 282 573 293 607
rect 327 573 338 607
rect 282 520 338 573
rect 282 486 293 520
rect 327 486 338 520
rect 282 437 338 486
rect 282 403 293 437
rect 327 403 338 437
rect 282 367 338 403
rect 368 599 424 619
rect 368 565 379 599
rect 413 565 424 599
rect 368 504 424 565
rect 368 470 379 504
rect 413 470 424 504
rect 368 413 424 470
rect 368 379 379 413
rect 413 379 424 413
rect 368 367 424 379
rect 454 607 510 619
rect 454 573 465 607
rect 499 573 510 607
rect 454 520 510 573
rect 454 486 465 520
rect 499 486 510 520
rect 454 437 510 486
rect 454 403 465 437
rect 499 403 510 437
rect 454 367 510 403
rect 540 599 596 619
rect 540 565 551 599
rect 585 565 596 599
rect 540 504 596 565
rect 540 470 551 504
rect 585 470 596 504
rect 540 413 596 470
rect 540 379 551 413
rect 585 379 596 413
rect 540 367 596 379
rect 626 607 682 619
rect 626 573 637 607
rect 671 573 682 607
rect 626 520 682 573
rect 626 486 637 520
rect 671 486 682 520
rect 626 437 682 486
rect 626 403 637 437
rect 671 403 682 437
rect 626 367 682 403
rect 712 599 836 619
rect 712 565 723 599
rect 757 565 791 599
rect 825 565 836 599
rect 712 518 836 565
rect 712 484 723 518
rect 757 484 791 518
rect 825 484 836 518
rect 712 434 836 484
rect 712 400 723 434
rect 757 400 791 434
rect 825 400 836 434
rect 712 367 836 400
rect 866 607 922 619
rect 866 573 877 607
rect 911 573 922 607
rect 866 495 922 573
rect 866 461 877 495
rect 911 461 922 495
rect 866 367 922 461
rect 952 599 1008 619
rect 952 565 963 599
rect 997 565 1008 599
rect 952 518 1008 565
rect 952 484 963 518
rect 997 484 1008 518
rect 952 418 1008 484
rect 952 384 963 418
rect 997 384 1008 418
rect 952 367 1008 384
rect 1038 607 1094 619
rect 1038 573 1049 607
rect 1083 573 1094 607
rect 1038 495 1094 573
rect 1038 461 1049 495
rect 1083 461 1094 495
rect 1038 367 1094 461
rect 1124 599 1180 619
rect 1124 565 1135 599
rect 1169 565 1180 599
rect 1124 518 1180 565
rect 1124 484 1135 518
rect 1169 484 1180 518
rect 1124 418 1180 484
rect 1124 384 1135 418
rect 1169 384 1180 418
rect 1124 367 1180 384
rect 1210 603 1266 619
rect 1210 569 1221 603
rect 1255 569 1266 603
rect 1210 495 1266 569
rect 1210 461 1221 495
rect 1255 461 1266 495
rect 1210 367 1266 461
rect 1296 529 1352 619
rect 1296 495 1307 529
rect 1341 495 1352 529
rect 1296 413 1352 495
rect 1296 379 1307 413
rect 1341 379 1352 413
rect 1296 367 1352 379
rect 1382 603 1438 619
rect 1382 569 1393 603
rect 1427 569 1438 603
rect 1382 529 1438 569
rect 1382 495 1393 529
rect 1427 495 1438 529
rect 1382 459 1438 495
rect 1382 425 1393 459
rect 1427 425 1438 459
rect 1382 367 1438 425
rect 1468 423 1521 619
rect 1468 389 1479 423
rect 1513 389 1521 423
rect 1468 367 1521 389
rect 1575 577 1628 619
rect 1575 543 1583 577
rect 1617 543 1628 577
rect 1575 367 1628 543
rect 1658 599 1714 619
rect 1658 565 1669 599
rect 1703 565 1714 599
rect 1658 504 1714 565
rect 1658 470 1669 504
rect 1703 470 1714 504
rect 1658 420 1714 470
rect 1658 386 1669 420
rect 1703 386 1714 420
rect 1658 367 1714 386
rect 1744 607 1800 619
rect 1744 573 1755 607
rect 1789 573 1800 607
rect 1744 494 1800 573
rect 1744 460 1755 494
rect 1789 460 1800 494
rect 1744 367 1800 460
rect 1830 599 1886 619
rect 1830 565 1841 599
rect 1875 565 1886 599
rect 1830 517 1886 565
rect 1830 483 1841 517
rect 1875 483 1886 517
rect 1830 436 1886 483
rect 1830 402 1841 436
rect 1875 402 1886 436
rect 1830 367 1886 402
rect 1916 607 1969 619
rect 1916 573 1927 607
rect 1961 573 1969 607
rect 1916 510 1969 573
rect 1916 476 1927 510
rect 1961 476 1969 510
rect 1916 420 1969 476
rect 1916 386 1927 420
rect 1961 386 1969 420
rect 1916 367 1969 386
<< ndiffc >>
rect 35 129 69 163
rect 35 59 69 93
rect 121 156 155 190
rect 207 63 241 97
rect 293 156 327 190
rect 379 165 413 199
rect 379 67 413 101
rect 465 129 499 163
rect 465 59 499 93
rect 551 147 585 181
rect 637 59 671 93
rect 723 147 757 181
rect 827 147 861 181
rect 913 135 947 169
rect 913 59 947 93
rect 999 135 1033 169
rect 1085 135 1119 169
rect 1085 59 1119 93
rect 1171 169 1205 203
rect 1171 67 1205 101
rect 1257 135 1291 169
rect 1257 59 1291 93
rect 1343 169 1377 203
rect 1343 67 1377 101
rect 1429 98 1463 132
rect 1515 173 1549 207
rect 1587 169 1621 203
rect 1515 67 1549 101
rect 1587 67 1621 101
rect 1673 133 1707 167
rect 1673 59 1707 93
rect 1759 169 1793 203
rect 1759 67 1793 101
rect 1845 133 1879 167
rect 1845 59 1879 93
rect 1931 169 1965 203
rect 1931 67 1965 101
<< pdiffc >>
rect 35 565 69 599
rect 35 470 69 504
rect 35 379 69 413
rect 121 573 155 607
rect 121 486 155 520
rect 121 403 155 437
rect 207 565 241 599
rect 207 470 241 504
rect 207 379 241 413
rect 293 573 327 607
rect 293 486 327 520
rect 293 403 327 437
rect 379 565 413 599
rect 379 470 413 504
rect 379 379 413 413
rect 465 573 499 607
rect 465 486 499 520
rect 465 403 499 437
rect 551 565 585 599
rect 551 470 585 504
rect 551 379 585 413
rect 637 573 671 607
rect 637 486 671 520
rect 637 403 671 437
rect 723 565 757 599
rect 791 565 825 599
rect 723 484 757 518
rect 791 484 825 518
rect 723 400 757 434
rect 791 400 825 434
rect 877 573 911 607
rect 877 461 911 495
rect 963 565 997 599
rect 963 484 997 518
rect 963 384 997 418
rect 1049 573 1083 607
rect 1049 461 1083 495
rect 1135 565 1169 599
rect 1135 484 1169 518
rect 1135 384 1169 418
rect 1221 569 1255 603
rect 1221 461 1255 495
rect 1307 495 1341 529
rect 1307 379 1341 413
rect 1393 569 1427 603
rect 1393 495 1427 529
rect 1393 425 1427 459
rect 1479 389 1513 423
rect 1583 543 1617 577
rect 1669 565 1703 599
rect 1669 470 1703 504
rect 1669 386 1703 420
rect 1755 573 1789 607
rect 1755 460 1789 494
rect 1841 565 1875 599
rect 1841 483 1875 517
rect 1841 402 1875 436
rect 1927 573 1961 607
rect 1927 476 1961 510
rect 1927 386 1961 420
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 252 619 282 645
rect 338 619 368 645
rect 424 619 454 645
rect 510 619 540 645
rect 596 619 626 645
rect 682 619 712 645
rect 836 619 866 645
rect 922 619 952 645
rect 1008 619 1038 645
rect 1094 619 1124 645
rect 1180 619 1210 645
rect 1266 619 1296 645
rect 1352 619 1382 645
rect 1438 619 1468 645
rect 1628 619 1658 645
rect 1714 619 1744 645
rect 1800 619 1830 645
rect 1886 619 1916 645
rect 80 317 110 367
rect 166 317 196 367
rect 252 317 282 367
rect 338 317 368 367
rect 424 317 454 367
rect 510 317 540 367
rect 596 317 626 367
rect 682 317 712 367
rect 836 346 866 367
rect 799 345 871 346
rect 922 345 952 367
rect 1008 345 1038 367
rect 1094 345 1124 367
rect 799 335 1124 345
rect 1180 345 1210 367
rect 1266 345 1296 367
rect 1352 345 1382 367
rect 1438 345 1468 367
rect 799 319 1137 335
rect 80 301 375 317
rect 80 267 121 301
rect 155 267 189 301
rect 223 267 257 301
rect 291 267 325 301
rect 359 267 375 301
rect 80 251 375 267
rect 417 301 755 317
rect 417 267 433 301
rect 467 267 501 301
rect 535 267 569 301
rect 603 267 637 301
rect 671 267 705 301
rect 739 267 755 301
rect 417 251 755 267
rect 799 285 815 319
rect 849 285 883 319
rect 917 285 951 319
rect 985 285 1019 319
rect 1053 285 1087 319
rect 1121 285 1137 319
rect 1180 321 1468 345
rect 1628 325 1658 367
rect 1714 325 1744 367
rect 1800 325 1830 367
rect 1886 325 1916 367
rect 1180 315 1504 321
rect 799 267 1137 285
rect 1202 305 1504 315
rect 1202 271 1218 305
rect 1252 271 1286 305
rect 1320 271 1354 305
rect 1388 271 1422 305
rect 1456 271 1504 305
rect 80 215 110 251
rect 166 215 196 251
rect 252 215 282 251
rect 338 215 368 251
rect 424 215 454 251
rect 510 215 540 251
rect 596 215 626 251
rect 682 215 712 251
rect 799 237 1160 267
rect 1202 255 1504 271
rect 1585 309 1991 325
rect 1585 275 1601 309
rect 1635 275 1669 309
rect 1703 275 1737 309
rect 1771 275 1805 309
rect 1839 275 1873 309
rect 1907 275 1941 309
rect 1975 275 1991 309
rect 1585 259 1991 275
rect 872 215 902 237
rect 958 215 988 237
rect 1044 215 1074 237
rect 1130 215 1160 237
rect 1216 215 1246 255
rect 1302 215 1332 255
rect 1388 215 1418 255
rect 1474 215 1504 255
rect 1632 215 1662 259
rect 1718 215 1748 259
rect 1804 215 1834 259
rect 1890 215 1920 259
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 424 21 454 47
rect 510 21 540 47
rect 596 21 626 47
rect 682 21 712 47
rect 872 21 902 47
rect 958 21 988 47
rect 1044 21 1074 47
rect 1130 21 1160 47
rect 1216 21 1246 47
rect 1302 21 1332 47
rect 1388 21 1418 47
rect 1474 21 1504 47
rect 1632 21 1662 47
rect 1718 21 1748 47
rect 1804 21 1834 47
rect 1890 21 1920 47
<< polycont >>
rect 121 267 155 301
rect 189 267 223 301
rect 257 267 291 301
rect 325 267 359 301
rect 433 267 467 301
rect 501 267 535 301
rect 569 267 603 301
rect 637 267 671 301
rect 705 267 739 301
rect 815 285 849 319
rect 883 285 917 319
rect 951 285 985 319
rect 1019 285 1053 319
rect 1087 285 1121 319
rect 1218 271 1252 305
rect 1286 271 1320 305
rect 1354 271 1388 305
rect 1422 271 1456 305
rect 1601 275 1635 309
rect 1669 275 1703 309
rect 1737 275 1771 309
rect 1805 275 1839 309
rect 1873 275 1907 309
rect 1941 275 1975 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 17 599 71 615
rect 17 565 35 599
rect 69 565 71 599
rect 17 504 71 565
rect 17 470 35 504
rect 69 470 71 504
rect 17 413 71 470
rect 17 379 35 413
rect 69 379 71 413
rect 105 607 171 649
rect 105 573 121 607
rect 155 573 171 607
rect 105 520 171 573
rect 105 486 121 520
rect 155 486 171 520
rect 105 437 171 486
rect 105 403 121 437
rect 155 403 171 437
rect 205 599 243 615
rect 205 565 207 599
rect 241 565 243 599
rect 205 504 243 565
rect 205 470 207 504
rect 241 470 243 504
rect 205 413 243 470
rect 17 369 71 379
rect 205 379 207 413
rect 241 379 243 413
rect 277 607 343 649
rect 277 573 293 607
rect 327 573 343 607
rect 277 520 343 573
rect 277 486 293 520
rect 327 486 343 520
rect 277 437 343 486
rect 277 403 293 437
rect 327 403 343 437
rect 377 599 415 615
rect 377 565 379 599
rect 413 565 415 599
rect 377 504 415 565
rect 377 470 379 504
rect 413 470 415 504
rect 377 413 415 470
rect 205 369 243 379
rect 377 379 379 413
rect 413 379 415 413
rect 449 607 515 649
rect 449 573 465 607
rect 499 573 515 607
rect 449 520 515 573
rect 449 486 465 520
rect 499 486 515 520
rect 449 437 515 486
rect 449 403 465 437
rect 499 403 515 437
rect 549 599 587 615
rect 549 565 551 599
rect 585 565 587 599
rect 549 504 587 565
rect 549 470 551 504
rect 585 470 587 504
rect 549 413 587 470
rect 377 369 415 379
rect 549 379 551 413
rect 585 379 587 413
rect 621 607 687 649
rect 621 573 637 607
rect 671 573 687 607
rect 621 520 687 573
rect 621 486 637 520
rect 671 486 687 520
rect 621 437 687 486
rect 621 403 637 437
rect 671 403 687 437
rect 721 599 826 615
rect 721 565 723 599
rect 757 565 791 599
rect 825 565 826 599
rect 721 518 826 565
rect 721 484 723 518
rect 757 484 791 518
rect 825 484 826 518
rect 721 434 826 484
rect 860 607 927 649
rect 860 573 877 607
rect 911 573 927 607
rect 860 495 927 573
rect 860 461 877 495
rect 911 461 927 495
rect 860 454 927 461
rect 961 599 999 615
rect 961 565 963 599
rect 997 565 999 599
rect 961 518 999 565
rect 961 484 963 518
rect 997 484 999 518
rect 549 369 587 379
rect 721 400 723 434
rect 757 400 791 434
rect 825 420 826 434
rect 961 420 999 484
rect 1033 607 1099 649
rect 1033 573 1049 607
rect 1083 573 1099 607
rect 1033 495 1099 573
rect 1033 461 1049 495
rect 1083 461 1099 495
rect 1033 454 1099 461
rect 1133 599 1171 615
rect 1133 565 1135 599
rect 1169 565 1171 599
rect 1133 518 1171 565
rect 1133 484 1135 518
rect 1169 484 1171 518
rect 1133 420 1171 484
rect 1205 603 1443 615
rect 1205 569 1221 603
rect 1255 579 1393 603
rect 1255 569 1271 579
rect 1205 495 1271 569
rect 1377 569 1393 579
rect 1427 569 1443 603
rect 1205 461 1221 495
rect 1255 461 1271 495
rect 1205 454 1271 461
rect 1305 529 1343 545
rect 1305 495 1307 529
rect 1341 495 1343 529
rect 1305 420 1343 495
rect 825 418 1343 420
rect 825 400 963 418
rect 721 384 963 400
rect 997 384 1135 418
rect 1169 413 1343 418
rect 1169 384 1307 413
rect 721 369 755 384
rect 17 335 755 369
rect 1302 379 1307 384
rect 1341 379 1343 413
rect 1377 529 1443 569
rect 1567 577 1633 649
rect 1567 543 1583 577
rect 1617 543 1633 577
rect 1567 533 1633 543
rect 1667 599 1705 615
rect 1667 565 1669 599
rect 1703 565 1705 599
rect 1377 495 1393 529
rect 1427 499 1443 529
rect 1667 504 1705 565
rect 1667 499 1669 504
rect 1427 495 1669 499
rect 1377 470 1669 495
rect 1703 470 1705 504
rect 1377 465 1705 470
rect 1377 459 1429 465
rect 1377 425 1393 459
rect 1427 425 1429 459
rect 1377 409 1429 425
rect 1463 423 1529 431
rect 1302 375 1343 379
rect 1463 389 1479 423
rect 1513 389 1529 423
rect 1463 375 1529 389
rect 1653 420 1705 465
rect 1739 607 1805 649
rect 1739 573 1755 607
rect 1789 573 1805 607
rect 1739 494 1805 573
rect 1739 460 1755 494
rect 1789 460 1805 494
rect 1739 454 1805 460
rect 1839 599 1877 615
rect 1839 565 1841 599
rect 1875 565 1877 599
rect 1839 517 1877 565
rect 1839 483 1841 517
rect 1875 483 1877 517
rect 1839 436 1877 483
rect 1839 420 1841 436
rect 1653 386 1669 420
rect 1703 402 1841 420
rect 1875 402 1877 436
rect 1703 386 1877 402
rect 1911 607 1977 649
rect 1911 573 1927 607
rect 1961 573 1977 607
rect 1911 510 1977 573
rect 1911 476 1927 510
rect 1961 476 1977 510
rect 1911 420 1977 476
rect 1911 386 1927 420
rect 1961 386 1977 420
rect 17 231 71 335
rect 789 319 1137 350
rect 1302 341 1529 375
rect 105 267 121 301
rect 155 267 189 301
rect 223 267 257 301
rect 291 267 325 301
rect 359 267 375 301
rect 417 267 433 301
rect 467 267 501 301
rect 535 267 569 301
rect 603 267 637 301
rect 671 267 705 301
rect 739 267 755 301
rect 789 285 815 319
rect 849 285 883 319
rect 917 285 951 319
rect 985 285 1019 319
rect 1053 285 1087 319
rect 1121 285 1137 319
rect 1585 309 1999 352
rect 789 271 1137 285
rect 1202 271 1218 305
rect 1252 271 1286 305
rect 1320 271 1354 305
rect 1388 271 1422 305
rect 1456 271 1533 305
rect 1585 275 1601 309
rect 1635 275 1669 309
rect 1703 275 1737 309
rect 1771 275 1805 309
rect 1839 275 1873 309
rect 1907 275 1941 309
rect 1975 275 1999 309
rect 189 240 337 267
rect 417 265 755 267
rect 623 231 755 265
rect 1427 241 1533 271
rect 17 206 155 231
rect 17 197 337 206
rect 119 190 337 197
rect 19 129 35 163
rect 69 129 85 163
rect 119 156 121 190
rect 155 156 293 190
rect 327 156 337 190
rect 119 140 337 156
rect 371 199 589 231
rect 371 165 379 199
rect 413 197 589 199
rect 811 207 1393 237
rect 1567 207 1981 235
rect 811 203 1515 207
rect 413 165 415 197
rect 19 106 85 129
rect 371 106 415 165
rect 549 181 761 197
rect 19 101 415 106
rect 19 97 379 101
rect 19 93 207 97
rect 19 59 35 93
rect 69 63 207 93
rect 241 67 379 97
rect 413 67 415 101
rect 241 63 415 67
rect 69 59 415 63
rect 19 51 415 59
rect 449 129 465 163
rect 499 129 515 163
rect 549 147 551 181
rect 585 147 723 181
rect 757 147 761 181
rect 549 131 761 147
rect 811 181 863 203
rect 811 147 827 181
rect 861 147 863 181
rect 997 169 1035 203
rect 1169 169 1171 203
rect 1205 169 1207 203
rect 1341 169 1343 203
rect 1377 173 1515 203
rect 1549 203 1981 207
rect 1549 173 1587 203
rect 1377 169 1379 173
rect 811 131 863 147
rect 897 135 913 169
rect 947 135 963 169
rect 449 97 515 129
rect 897 97 963 135
rect 997 135 999 169
rect 1033 135 1035 169
rect 997 119 1035 135
rect 1069 135 1085 169
rect 1119 135 1135 169
rect 449 93 963 97
rect 449 59 465 93
rect 499 59 637 93
rect 671 59 913 93
rect 947 85 963 93
rect 1069 93 1135 135
rect 1069 85 1085 93
rect 947 59 1085 85
rect 1119 59 1135 93
rect 449 51 1135 59
rect 1169 101 1207 169
rect 1169 67 1171 101
rect 1205 67 1207 101
rect 1169 51 1207 67
rect 1241 135 1257 169
rect 1291 135 1307 169
rect 1241 93 1307 135
rect 1241 59 1257 93
rect 1291 59 1307 93
rect 1241 17 1307 59
rect 1341 101 1379 169
rect 1513 169 1587 173
rect 1621 201 1759 203
rect 1621 169 1623 201
rect 1341 67 1343 101
rect 1377 67 1379 101
rect 1341 51 1379 67
rect 1413 132 1479 139
rect 1413 98 1429 132
rect 1463 98 1479 132
rect 1413 17 1479 98
rect 1513 101 1623 169
rect 1757 169 1759 201
rect 1793 201 1931 203
rect 1793 169 1795 201
rect 1513 67 1515 101
rect 1549 67 1587 101
rect 1621 67 1623 101
rect 1513 51 1623 67
rect 1657 133 1673 167
rect 1707 133 1723 167
rect 1657 93 1723 133
rect 1657 59 1673 93
rect 1707 59 1723 93
rect 1657 17 1723 59
rect 1757 101 1795 169
rect 1929 169 1931 201
rect 1965 169 1981 203
rect 1757 67 1759 101
rect 1793 67 1795 101
rect 1757 51 1795 67
rect 1829 133 1845 167
rect 1879 133 1895 167
rect 1829 93 1895 133
rect 1829 59 1845 93
rect 1879 59 1895 93
rect 1829 17 1895 59
rect 1929 101 1981 169
rect 1929 67 1931 101
rect 1965 67 1981 101
rect 1929 51 1981 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2111ai_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4727608
string GDS_START 4710040
<< end >>
