magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
<< pwell >>
rect 331 159 1241 241
rect 28 49 1241 159
rect 0 0 1248 49
<< scnmos >>
rect 107 49 137 133
rect 193 49 223 133
rect 410 47 440 215
rect 496 47 526 215
rect 584 47 614 215
rect 684 47 714 215
rect 874 47 904 215
rect 960 47 990 215
rect 1046 47 1076 215
rect 1132 47 1162 215
<< scpmoshvt >>
rect 80 373 110 457
rect 220 373 250 457
rect 426 367 456 619
rect 512 367 542 619
rect 598 367 628 619
rect 684 367 714 619
rect 770 367 800 619
rect 856 367 886 619
rect 942 367 972 619
rect 1104 367 1134 619
<< ndiff >>
rect 357 203 410 215
rect 357 169 365 203
rect 399 169 410 203
rect 54 105 107 133
rect 54 71 62 105
rect 96 71 107 105
rect 54 49 107 71
rect 137 103 193 133
rect 137 69 148 103
rect 182 69 193 103
rect 137 49 193 69
rect 223 105 276 133
rect 223 71 234 105
rect 268 71 276 105
rect 223 49 276 71
rect 357 105 410 169
rect 357 71 365 105
rect 399 71 410 105
rect 357 47 410 71
rect 440 169 496 215
rect 440 135 451 169
rect 485 135 496 169
rect 440 47 496 135
rect 526 165 584 215
rect 526 131 537 165
rect 571 131 584 165
rect 526 93 584 131
rect 526 59 537 93
rect 571 59 584 93
rect 526 47 584 59
rect 614 163 684 215
rect 614 129 639 163
rect 673 129 684 163
rect 614 47 684 129
rect 714 93 767 215
rect 714 59 725 93
rect 759 59 767 93
rect 714 47 767 59
rect 821 93 874 215
rect 821 59 829 93
rect 863 59 874 93
rect 821 47 874 59
rect 904 167 960 215
rect 904 133 915 167
rect 949 133 960 167
rect 904 47 960 133
rect 990 197 1046 215
rect 990 163 1001 197
rect 1035 163 1046 197
rect 990 101 1046 163
rect 990 67 1001 101
rect 1035 67 1046 101
rect 990 47 1046 67
rect 1076 179 1132 215
rect 1076 145 1087 179
rect 1121 145 1132 179
rect 1076 93 1132 145
rect 1076 59 1087 93
rect 1121 59 1132 93
rect 1076 47 1132 59
rect 1162 203 1215 215
rect 1162 169 1173 203
rect 1207 169 1215 203
rect 1162 101 1215 169
rect 1162 67 1173 101
rect 1207 67 1215 101
rect 1162 47 1215 67
<< pdiff >>
rect 373 581 426 619
rect 373 547 381 581
rect 415 547 426 581
rect 27 432 80 457
rect 27 398 35 432
rect 69 398 80 432
rect 27 373 80 398
rect 110 443 220 457
rect 110 409 125 443
rect 159 409 220 443
rect 110 373 220 409
rect 250 419 303 457
rect 250 385 261 419
rect 295 385 303 419
rect 250 373 303 385
rect 373 367 426 547
rect 456 599 512 619
rect 456 565 467 599
rect 501 565 512 599
rect 456 504 512 565
rect 456 470 467 504
rect 501 470 512 504
rect 456 413 512 470
rect 456 379 467 413
rect 501 379 512 413
rect 456 367 512 379
rect 542 607 598 619
rect 542 573 553 607
rect 587 573 598 607
rect 542 539 598 573
rect 542 505 553 539
rect 587 505 598 539
rect 542 471 598 505
rect 542 437 553 471
rect 587 437 598 471
rect 542 367 598 437
rect 628 599 684 619
rect 628 565 639 599
rect 673 565 684 599
rect 628 504 684 565
rect 628 470 639 504
rect 673 470 684 504
rect 628 413 684 470
rect 628 379 639 413
rect 673 379 684 413
rect 628 367 684 379
rect 714 607 770 619
rect 714 573 725 607
rect 759 573 770 607
rect 714 533 770 573
rect 714 499 725 533
rect 759 499 770 533
rect 714 452 770 499
rect 714 418 725 452
rect 759 418 770 452
rect 714 367 770 418
rect 800 599 856 619
rect 800 565 811 599
rect 845 565 856 599
rect 800 503 856 565
rect 800 469 811 503
rect 845 469 856 503
rect 800 413 856 469
rect 800 379 811 413
rect 845 379 856 413
rect 800 367 856 379
rect 886 607 942 619
rect 886 573 897 607
rect 931 573 942 607
rect 886 519 942 573
rect 886 485 897 519
rect 931 485 942 519
rect 886 423 942 485
rect 886 389 897 423
rect 931 389 942 423
rect 886 367 942 389
rect 972 599 1104 619
rect 972 565 983 599
rect 1017 565 1059 599
rect 1093 565 1104 599
rect 972 513 1104 565
rect 972 503 1059 513
rect 972 469 983 503
rect 1017 479 1059 503
rect 1093 479 1104 513
rect 1017 469 1104 479
rect 972 434 1104 469
rect 972 413 1059 434
rect 972 379 983 413
rect 1017 400 1059 413
rect 1093 400 1104 434
rect 1017 379 1104 400
rect 972 367 1104 379
rect 1134 607 1187 619
rect 1134 573 1145 607
rect 1179 573 1187 607
rect 1134 513 1187 573
rect 1134 479 1145 513
rect 1179 479 1187 513
rect 1134 418 1187 479
rect 1134 384 1145 418
rect 1179 384 1187 418
rect 1134 367 1187 384
<< ndiffc >>
rect 365 169 399 203
rect 62 71 96 105
rect 148 69 182 103
rect 234 71 268 105
rect 365 71 399 105
rect 451 135 485 169
rect 537 131 571 165
rect 537 59 571 93
rect 639 129 673 163
rect 725 59 759 93
rect 829 59 863 93
rect 915 133 949 167
rect 1001 163 1035 197
rect 1001 67 1035 101
rect 1087 145 1121 179
rect 1087 59 1121 93
rect 1173 169 1207 203
rect 1173 67 1207 101
<< pdiffc >>
rect 381 547 415 581
rect 35 398 69 432
rect 125 409 159 443
rect 261 385 295 419
rect 467 565 501 599
rect 467 470 501 504
rect 467 379 501 413
rect 553 573 587 607
rect 553 505 587 539
rect 553 437 587 471
rect 639 565 673 599
rect 639 470 673 504
rect 639 379 673 413
rect 725 573 759 607
rect 725 499 759 533
rect 725 418 759 452
rect 811 565 845 599
rect 811 469 845 503
rect 811 379 845 413
rect 897 573 931 607
rect 897 485 931 519
rect 897 389 931 423
rect 983 565 1017 599
rect 1059 565 1093 599
rect 983 469 1017 503
rect 1059 479 1093 513
rect 983 379 1017 413
rect 1059 400 1093 434
rect 1145 573 1179 607
rect 1145 479 1179 513
rect 1145 384 1179 418
<< poly >>
rect 426 619 456 645
rect 512 619 542 645
rect 598 619 628 645
rect 684 619 714 645
rect 770 619 800 645
rect 856 619 886 645
rect 942 619 972 645
rect 1104 619 1134 645
rect 80 457 110 483
rect 220 457 250 483
rect 80 289 110 373
rect 220 289 250 373
rect 426 331 456 367
rect 512 331 542 367
rect 307 315 542 331
rect 598 330 628 367
rect 684 330 714 367
rect 79 273 145 289
rect 79 239 95 273
rect 129 239 145 273
rect 79 205 145 239
rect 79 171 95 205
rect 129 171 145 205
rect 79 155 145 171
rect 193 273 259 289
rect 193 239 209 273
rect 243 239 259 273
rect 307 281 323 315
rect 357 281 542 315
rect 307 265 542 281
rect 584 314 714 330
rect 584 280 600 314
rect 634 280 714 314
rect 193 205 259 239
rect 410 215 440 265
rect 496 215 526 265
rect 584 264 714 280
rect 584 215 614 264
rect 684 215 714 264
rect 770 303 800 367
rect 856 303 886 367
rect 942 345 972 367
rect 1104 345 1134 367
rect 942 335 1134 345
rect 942 319 1170 335
rect 942 315 1120 319
rect 770 298 901 303
rect 770 295 903 298
rect 770 287 905 295
rect 770 253 787 287
rect 821 253 855 287
rect 889 267 905 287
rect 1032 285 1120 315
rect 1154 285 1170 319
rect 1032 269 1170 285
rect 889 253 990 267
rect 770 237 990 253
rect 874 215 904 237
rect 960 215 990 237
rect 1046 215 1076 269
rect 1132 215 1162 269
rect 193 171 209 205
rect 243 171 259 205
rect 193 155 259 171
rect 107 133 137 155
rect 193 133 223 155
rect 107 23 137 49
rect 193 23 223 49
rect 410 21 440 47
rect 496 21 526 47
rect 584 21 614 47
rect 684 21 714 47
rect 874 21 904 47
rect 960 21 990 47
rect 1046 21 1076 47
rect 1132 21 1162 47
<< polycont >>
rect 95 239 129 273
rect 95 171 129 205
rect 209 239 243 273
rect 323 281 357 315
rect 600 280 634 314
rect 787 253 821 287
rect 855 253 889 287
rect 1120 285 1154 319
rect 209 171 243 205
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 17 432 78 448
rect 17 398 35 432
rect 69 398 78 432
rect 17 359 78 398
rect 112 443 159 649
rect 365 581 431 649
rect 365 547 381 581
rect 415 547 431 581
rect 365 537 431 547
rect 465 599 503 615
rect 465 565 467 599
rect 501 565 503 599
rect 465 504 503 565
rect 112 409 125 443
rect 112 393 159 409
rect 193 469 431 503
rect 193 359 227 469
rect 261 419 363 435
rect 295 385 363 419
rect 261 369 363 385
rect 17 325 227 359
rect 17 121 59 325
rect 295 315 363 369
rect 93 273 169 289
rect 93 239 95 273
rect 129 239 169 273
rect 93 205 169 239
rect 93 171 95 205
rect 129 171 169 205
rect 93 155 169 171
rect 203 273 261 289
rect 203 239 209 273
rect 243 239 261 273
rect 203 205 261 239
rect 203 171 209 205
rect 243 171 261 205
rect 203 155 261 171
rect 295 281 323 315
rect 357 281 363 315
rect 295 265 363 281
rect 397 314 431 469
rect 465 470 467 504
rect 501 470 503 504
rect 465 413 503 470
rect 537 607 603 649
rect 537 573 553 607
rect 587 573 603 607
rect 537 539 603 573
rect 537 505 553 539
rect 587 505 603 539
rect 537 471 603 505
rect 537 437 553 471
rect 587 437 603 471
rect 537 421 603 437
rect 637 599 675 615
rect 637 565 639 599
rect 673 565 675 599
rect 637 504 675 565
rect 637 470 639 504
rect 673 470 675 504
rect 465 379 467 413
rect 501 384 503 413
rect 637 413 675 470
rect 709 607 775 649
rect 709 573 725 607
rect 759 573 775 607
rect 709 533 775 573
rect 709 499 725 533
rect 759 499 775 533
rect 709 452 775 499
rect 709 418 725 452
rect 759 418 775 452
rect 809 599 847 615
rect 809 565 811 599
rect 845 565 847 599
rect 809 503 847 565
rect 809 469 811 503
rect 845 469 847 503
rect 637 384 639 413
rect 501 379 639 384
rect 673 384 675 413
rect 809 413 847 469
rect 809 384 811 413
rect 673 379 811 384
rect 845 379 847 413
rect 881 607 947 649
rect 881 573 897 607
rect 931 573 947 607
rect 881 519 947 573
rect 881 485 897 519
rect 931 485 947 519
rect 881 423 947 485
rect 881 389 897 423
rect 931 389 947 423
rect 981 599 1095 615
rect 981 565 983 599
rect 1017 565 1059 599
rect 1093 565 1095 599
rect 981 513 1095 565
rect 981 503 1059 513
rect 981 469 983 503
rect 1017 479 1059 503
rect 1093 479 1095 513
rect 1017 469 1095 479
rect 981 434 1095 469
rect 981 413 1059 434
rect 465 355 847 379
rect 981 379 983 413
rect 1017 400 1059 413
rect 1093 400 1095 434
rect 1017 384 1095 400
rect 1129 607 1195 649
rect 1129 573 1145 607
rect 1179 573 1195 607
rect 1129 513 1195 573
rect 1129 479 1145 513
rect 1179 479 1195 513
rect 1129 418 1195 479
rect 1129 384 1145 418
rect 1179 384 1195 418
rect 1017 379 1053 384
rect 981 355 1053 379
rect 465 348 1053 355
rect 684 321 1053 348
rect 397 280 600 314
rect 634 280 650 314
rect 397 275 650 280
rect 295 121 329 265
rect 684 241 737 321
rect 1087 319 1217 350
rect 771 253 787 287
rect 821 253 855 287
rect 889 253 929 287
rect 1087 285 1120 319
rect 1154 285 1217 319
rect 771 242 929 253
rect 17 105 98 121
rect 17 71 62 105
rect 96 71 98 105
rect 17 55 98 71
rect 132 103 198 111
rect 132 69 148 103
rect 182 69 198 103
rect 132 17 198 69
rect 232 105 329 121
rect 232 71 234 105
rect 268 71 329 105
rect 232 55 329 71
rect 363 203 403 219
rect 363 169 365 203
rect 399 169 403 203
rect 363 105 403 169
rect 442 207 737 241
rect 999 213 1223 247
rect 442 169 487 207
rect 999 197 1037 213
rect 442 135 451 169
rect 485 135 487 169
rect 623 167 965 173
rect 442 119 487 135
rect 521 131 537 165
rect 571 131 587 165
rect 363 71 365 105
rect 399 85 403 105
rect 521 93 587 131
rect 623 163 915 167
rect 623 129 639 163
rect 673 133 915 163
rect 949 133 965 167
rect 673 129 965 133
rect 623 127 965 129
rect 999 163 1001 197
rect 1035 163 1037 197
rect 1171 203 1223 213
rect 999 101 1037 163
rect 999 93 1001 101
rect 521 85 537 93
rect 399 71 537 85
rect 363 59 537 71
rect 571 59 725 93
rect 759 59 775 93
rect 363 51 775 59
rect 813 59 829 93
rect 863 67 1001 93
rect 1035 67 1037 101
rect 863 59 1037 67
rect 813 51 1037 59
rect 1071 145 1087 179
rect 1121 145 1137 179
rect 1071 93 1137 145
rect 1071 59 1087 93
rect 1121 59 1137 93
rect 1071 17 1137 59
rect 1171 169 1173 203
rect 1207 169 1223 203
rect 1171 101 1223 169
rect 1171 67 1173 101
rect 1207 67 1223 101
rect 1171 51 1223 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4bb_2
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5651068
string GDS_START 5640360
<< end >>
