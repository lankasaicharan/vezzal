magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1288 -1260 1544 1525
use sky130_fd_pr__dfm1sd2__example_5595914180836  sky130_fd_pr__dfm1sd2__example_5595914180836_0
timestamp 1627201311
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180835  sky130_fd_pr__hvdfm1sd__example_5595914180835_0
timestamp 1627201311
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180835  sky130_fd_pr__hvdfm1sd__example_5595914180835_1
timestamp 1627201311
transform 1 0 256 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 284 265 284 265 0 FreeSans 300 0 0 0 S
flabel comment s 128 265 128 265 0 FreeSans 300 0 0 0 D
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 43661154
string GDS_START 43659714
<< end >>
