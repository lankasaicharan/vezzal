magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1490 1975
<< nwell >>
rect -38 331 230 704
<< pwell >>
rect 5 49 187 255
rect 0 0 192 49
<< psubdiff >>
rect 31 205 161 229
rect 65 171 127 205
rect 31 122 161 171
rect 65 88 127 122
rect 31 64 161 88
<< nsubdiff >>
rect 31 578 161 602
rect 65 544 127 578
rect 31 491 161 544
rect 65 457 127 491
rect 31 433 161 457
<< psubdiffcont >>
rect 31 171 65 205
rect 127 171 161 205
rect 31 88 65 122
rect 127 88 161 122
<< nsubdiffcont >>
rect 31 544 65 578
rect 127 544 161 578
rect 31 457 65 491
rect 127 457 161 491
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 18 578 174 613
rect 18 544 31 578
rect 65 544 127 578
rect 161 544 174 578
rect 18 491 174 544
rect 18 457 31 491
rect 65 457 127 491
rect 161 457 174 491
rect 18 378 174 457
rect 18 205 174 288
rect 18 171 31 205
rect 65 171 127 205
rect 161 171 174 205
rect 18 122 174 171
rect 18 88 31 122
rect 65 88 127 122
rect 161 88 174 122
rect 18 53 174 88
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 31 -17 65 17
rect 127 -17 161 17
<< metal1 >>
rect 0 683 192 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 0 617 192 649
rect 0 17 192 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
rect 0 -49 192 -17
<< labels >>
flabel pwell s 0 0 192 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew ground bidirectional
flabel nwell s 0 617 192 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew power bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 VNB
port 2 nsew ground bidirectional
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 VNB
port 2 nsew ground bidirectional
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 VNB
port 2 nsew ground bidirectional
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 VPB
port 3 nsew power bidirectional
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 VPB
port 3 nsew power bidirectional
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 VPB
port 3 nsew power bidirectional
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 VPB
port 3 nsew power bidirectional
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 VNB
port 2 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 VNB
port 2 nsew ground bidirectional
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 VPB
port 3 nsew power bidirectional
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 VPB
port 3 nsew power bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 VNB
port 2 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 tap_2
flabel metal1 s 0 617 192 666 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional
flabel metal1 s 0 0 192 49 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional
rlabel pwell s 0 0 192 49 1 VNB
port 2 nsew ground bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE WELLTAP
string FIXED_BBOX 0 0 192 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1420706
string GDS_START 1416790
<< end >>
