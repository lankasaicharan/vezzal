magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 17 49 667 250
rect 0 0 672 49
<< scnmos >>
rect 96 56 126 224
rect 264 56 294 224
rect 342 56 372 224
rect 450 56 480 224
rect 558 56 588 224
<< scpmoshvt >>
rect 80 367 110 619
rect 270 367 300 619
rect 360 367 390 619
rect 450 367 480 619
rect 558 367 588 619
<< ndiff >>
rect 43 212 96 224
rect 43 178 51 212
rect 85 178 96 212
rect 43 102 96 178
rect 43 68 51 102
rect 85 68 96 102
rect 43 56 96 68
rect 126 132 264 224
rect 126 98 137 132
rect 171 98 219 132
rect 253 98 264 132
rect 126 56 264 98
rect 294 56 342 224
rect 372 208 450 224
rect 372 174 395 208
rect 429 174 450 208
rect 372 101 450 174
rect 372 67 395 101
rect 429 67 450 101
rect 372 56 450 67
rect 480 56 558 224
rect 588 208 641 224
rect 588 174 599 208
rect 633 174 641 208
rect 588 102 641 174
rect 588 68 599 102
rect 633 68 641 102
rect 588 56 641 68
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 502 80 565
rect 27 468 35 502
rect 69 468 80 502
rect 27 420 80 468
rect 27 386 35 420
rect 69 386 80 420
rect 27 367 80 386
rect 110 607 163 619
rect 110 573 121 607
rect 155 573 163 607
rect 110 525 163 573
rect 110 491 121 525
rect 155 491 163 525
rect 110 448 163 491
rect 110 414 121 448
rect 155 414 163 448
rect 110 367 163 414
rect 217 599 270 619
rect 217 565 225 599
rect 259 565 270 599
rect 217 520 270 565
rect 217 486 225 520
rect 259 486 270 520
rect 217 448 270 486
rect 217 414 225 448
rect 259 414 270 448
rect 217 367 270 414
rect 300 547 360 619
rect 300 513 311 547
rect 345 513 360 547
rect 300 413 360 513
rect 300 379 311 413
rect 345 379 360 413
rect 300 367 360 379
rect 390 599 450 619
rect 390 565 401 599
rect 435 565 450 599
rect 390 511 450 565
rect 390 477 401 511
rect 435 477 450 511
rect 390 413 450 477
rect 390 379 401 413
rect 435 379 450 413
rect 390 367 450 379
rect 480 607 558 619
rect 480 573 503 607
rect 537 573 558 607
rect 480 529 558 573
rect 480 495 503 529
rect 537 495 558 529
rect 480 448 558 495
rect 480 414 503 448
rect 537 414 558 448
rect 480 367 558 414
rect 588 599 641 619
rect 588 565 599 599
rect 633 565 641 599
rect 588 511 641 565
rect 588 477 599 511
rect 633 477 641 511
rect 588 413 641 477
rect 588 379 599 413
rect 633 379 641 413
rect 588 367 641 379
<< ndiffc >>
rect 51 178 85 212
rect 51 68 85 102
rect 137 98 171 132
rect 219 98 253 132
rect 395 174 429 208
rect 395 67 429 101
rect 599 174 633 208
rect 599 68 633 102
<< pdiffc >>
rect 35 565 69 599
rect 35 468 69 502
rect 35 386 69 420
rect 121 573 155 607
rect 121 491 155 525
rect 121 414 155 448
rect 225 565 259 599
rect 225 486 259 520
rect 225 414 259 448
rect 311 513 345 547
rect 311 379 345 413
rect 401 565 435 599
rect 401 477 435 511
rect 401 379 435 413
rect 503 573 537 607
rect 503 495 537 529
rect 503 414 537 448
rect 599 565 633 599
rect 599 477 633 511
rect 599 379 633 413
<< poly >>
rect 80 619 110 645
rect 270 619 300 645
rect 360 619 390 645
rect 450 619 480 645
rect 558 619 588 645
rect 80 312 110 367
rect 270 312 300 367
rect 360 312 390 367
rect 450 312 480 367
rect 558 312 588 367
rect 80 296 175 312
rect 80 262 125 296
rect 159 262 175 296
rect 80 246 175 262
rect 217 296 300 312
rect 217 262 233 296
rect 267 282 300 296
rect 342 296 408 312
rect 267 262 294 282
rect 217 246 294 262
rect 96 224 126 246
rect 264 224 294 246
rect 342 262 358 296
rect 392 262 408 296
rect 342 246 408 262
rect 450 296 516 312
rect 450 262 466 296
rect 500 262 516 296
rect 450 246 516 262
rect 558 296 631 312
rect 558 262 581 296
rect 615 262 631 296
rect 558 246 631 262
rect 342 224 372 246
rect 450 224 480 246
rect 558 224 588 246
rect 96 30 126 56
rect 264 30 294 56
rect 342 30 372 56
rect 450 30 480 56
rect 558 30 588 56
<< polycont >>
rect 125 262 159 296
rect 233 262 267 296
rect 358 262 392 296
rect 466 262 500 296
rect 581 262 615 296
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 19 599 73 615
rect 19 565 35 599
rect 69 565 73 599
rect 19 502 73 565
rect 19 468 35 502
rect 69 468 73 502
rect 19 420 73 468
rect 19 386 35 420
rect 69 386 73 420
rect 117 607 171 649
rect 117 573 121 607
rect 155 573 171 607
rect 117 525 171 573
rect 117 491 121 525
rect 155 491 171 525
rect 117 448 171 491
rect 117 414 121 448
rect 155 414 171 448
rect 117 398 171 414
rect 209 599 451 615
rect 209 565 225 599
rect 259 581 401 599
rect 259 565 261 581
rect 209 520 261 565
rect 395 565 401 581
rect 435 565 451 599
rect 209 486 225 520
rect 259 486 261 520
rect 209 448 261 486
rect 209 414 225 448
rect 259 414 261 448
rect 209 398 261 414
rect 295 513 311 547
rect 345 513 361 547
rect 295 413 361 513
rect 19 228 73 386
rect 295 379 311 413
rect 345 379 361 413
rect 295 364 361 379
rect 121 330 361 364
rect 395 511 451 565
rect 395 477 401 511
rect 435 477 451 511
rect 395 413 451 477
rect 485 607 553 649
rect 485 573 503 607
rect 537 573 553 607
rect 485 529 553 573
rect 485 495 503 529
rect 537 495 553 529
rect 485 448 553 495
rect 485 414 503 448
rect 537 414 553 448
rect 587 599 649 615
rect 587 565 599 599
rect 633 565 649 599
rect 587 511 649 565
rect 587 477 599 511
rect 633 477 649 511
rect 395 379 401 413
rect 435 380 451 413
rect 587 413 649 477
rect 587 380 599 413
rect 435 379 599 380
rect 633 379 649 413
rect 395 346 649 379
rect 121 296 169 330
rect 466 296 547 312
rect 121 262 125 296
rect 159 262 169 296
rect 19 212 87 228
rect 19 178 51 212
rect 85 178 87 212
rect 19 102 87 178
rect 121 208 169 262
rect 203 262 233 296
rect 267 262 283 296
rect 203 242 283 262
rect 317 262 358 296
rect 392 262 408 296
rect 317 242 408 262
rect 500 262 547 296
rect 466 242 547 262
rect 581 296 655 312
rect 615 262 655 296
rect 581 242 655 262
rect 121 174 395 208
rect 429 174 445 208
rect 19 68 51 102
rect 85 68 87 102
rect 19 51 87 68
rect 121 132 269 140
rect 121 98 137 132
rect 171 98 219 132
rect 253 98 269 132
rect 121 17 269 98
rect 379 101 445 174
rect 379 67 395 101
rect 429 67 445 101
rect 490 79 547 242
rect 583 174 599 208
rect 633 174 649 208
rect 583 102 649 174
rect 379 51 445 67
rect 583 68 599 102
rect 633 68 649 102
rect 583 17 649 68
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a22o_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1153930
string GDS_START 1146520
<< end >>
