magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 497 241 947 261
rect 43 49 947 241
rect 0 0 960 49
<< scnmos >>
rect 122 47 152 215
rect 208 47 238 215
rect 300 47 330 215
rect 386 47 416 215
rect 580 67 610 235
rect 666 67 696 235
rect 752 67 782 235
rect 838 67 868 235
<< scpmoshvt >>
rect 156 367 186 619
rect 242 367 272 619
rect 328 367 358 619
rect 414 367 444 619
rect 516 367 546 619
rect 602 367 632 619
rect 738 367 768 619
rect 824 367 854 619
<< ndiff >>
rect 69 203 122 215
rect 69 169 77 203
rect 111 169 122 203
rect 69 101 122 169
rect 69 67 77 101
rect 111 67 122 101
rect 69 47 122 67
rect 152 157 208 215
rect 152 123 163 157
rect 197 123 208 157
rect 152 89 208 123
rect 152 55 163 89
rect 197 55 208 89
rect 152 47 208 55
rect 238 203 300 215
rect 238 169 249 203
rect 283 169 300 203
rect 238 101 300 169
rect 238 67 249 101
rect 283 67 300 101
rect 238 47 300 67
rect 330 183 386 215
rect 330 149 341 183
rect 375 149 386 183
rect 330 47 386 149
rect 416 99 469 215
rect 416 65 427 99
rect 461 65 469 99
rect 523 109 580 235
rect 523 75 535 109
rect 569 75 580 109
rect 523 67 580 75
rect 610 179 666 235
rect 610 145 621 179
rect 655 145 666 179
rect 610 67 666 145
rect 696 165 752 235
rect 696 131 707 165
rect 741 131 752 165
rect 696 67 752 131
rect 782 227 838 235
rect 782 193 793 227
rect 827 193 838 227
rect 782 153 838 193
rect 782 119 793 153
rect 827 119 838 153
rect 782 67 838 119
rect 868 223 921 235
rect 868 189 879 223
rect 913 189 921 223
rect 868 113 921 189
rect 868 79 879 113
rect 913 79 921 113
rect 868 67 921 79
rect 416 47 469 65
<< pdiff >>
rect 35 607 156 619
rect 35 573 43 607
rect 77 573 111 607
rect 145 573 156 607
rect 35 509 156 573
rect 35 475 43 509
rect 77 475 111 509
rect 145 475 156 509
rect 35 413 156 475
rect 35 379 43 413
rect 77 379 156 413
rect 35 367 156 379
rect 186 599 242 619
rect 186 565 197 599
rect 231 565 242 599
rect 186 505 242 565
rect 186 471 197 505
rect 231 471 242 505
rect 186 413 242 471
rect 186 379 197 413
rect 231 379 242 413
rect 186 367 242 379
rect 272 607 328 619
rect 272 573 283 607
rect 317 573 328 607
rect 272 530 328 573
rect 272 496 283 530
rect 317 496 328 530
rect 272 453 328 496
rect 272 419 283 453
rect 317 419 328 453
rect 272 367 328 419
rect 358 599 414 619
rect 358 565 369 599
rect 403 565 414 599
rect 358 505 414 565
rect 358 471 369 505
rect 403 471 414 505
rect 358 413 414 471
rect 358 379 369 413
rect 403 379 414 413
rect 358 367 414 379
rect 444 607 516 619
rect 444 573 464 607
rect 498 573 516 607
rect 444 493 516 573
rect 444 459 464 493
rect 498 459 516 493
rect 444 367 516 459
rect 546 599 602 619
rect 546 565 557 599
rect 591 565 602 599
rect 546 509 602 565
rect 546 475 557 509
rect 591 475 602 509
rect 546 418 602 475
rect 546 384 557 418
rect 591 384 602 418
rect 546 367 602 384
rect 632 607 738 619
rect 632 573 668 607
rect 702 573 738 607
rect 632 493 738 573
rect 632 459 668 493
rect 702 459 738 493
rect 632 367 738 459
rect 768 599 824 619
rect 768 565 779 599
rect 813 565 824 599
rect 768 509 824 565
rect 768 475 779 509
rect 813 475 824 509
rect 768 434 824 475
rect 768 400 779 434
rect 813 400 824 434
rect 768 367 824 400
rect 854 607 907 619
rect 854 573 865 607
rect 899 573 907 607
rect 854 509 907 573
rect 854 475 865 509
rect 899 475 907 509
rect 854 418 907 475
rect 854 384 865 418
rect 899 384 907 418
rect 854 367 907 384
<< ndiffc >>
rect 77 169 111 203
rect 77 67 111 101
rect 163 123 197 157
rect 163 55 197 89
rect 249 169 283 203
rect 249 67 283 101
rect 341 149 375 183
rect 427 65 461 99
rect 535 75 569 109
rect 621 145 655 179
rect 707 131 741 165
rect 793 193 827 227
rect 793 119 827 153
rect 879 189 913 223
rect 879 79 913 113
<< pdiffc >>
rect 43 573 77 607
rect 111 573 145 607
rect 43 475 77 509
rect 111 475 145 509
rect 43 379 77 413
rect 197 565 231 599
rect 197 471 231 505
rect 197 379 231 413
rect 283 573 317 607
rect 283 496 317 530
rect 283 419 317 453
rect 369 565 403 599
rect 369 471 403 505
rect 369 379 403 413
rect 464 573 498 607
rect 464 459 498 493
rect 557 565 591 599
rect 557 475 591 509
rect 557 384 591 418
rect 668 573 702 607
rect 668 459 702 493
rect 779 565 813 599
rect 779 475 813 509
rect 779 400 813 434
rect 865 573 899 607
rect 865 475 899 509
rect 865 384 899 418
<< poly >>
rect 156 619 186 645
rect 242 619 272 645
rect 328 619 358 645
rect 414 619 444 645
rect 516 619 546 645
rect 602 619 632 645
rect 738 619 768 645
rect 824 619 854 645
rect 156 345 186 367
rect 242 345 272 367
rect 111 319 272 345
rect 111 285 127 319
rect 161 315 272 319
rect 161 285 238 315
rect 111 269 238 285
rect 122 215 152 269
rect 208 215 238 269
rect 328 267 358 367
rect 414 303 444 367
rect 400 287 466 303
rect 400 267 416 287
rect 300 253 416 267
rect 450 253 466 287
rect 516 299 546 367
rect 602 335 632 367
rect 738 335 768 367
rect 824 335 854 367
rect 601 319 696 335
rect 601 299 617 319
rect 516 285 617 299
rect 651 285 696 319
rect 516 269 696 285
rect 738 319 872 335
rect 738 285 754 319
rect 788 285 822 319
rect 856 285 872 319
rect 738 269 872 285
rect 300 237 466 253
rect 300 215 330 237
rect 386 215 416 237
rect 580 235 610 269
rect 666 235 696 269
rect 752 235 782 269
rect 838 235 868 269
rect 122 21 152 47
rect 208 21 238 47
rect 300 21 330 47
rect 386 21 416 47
rect 580 41 610 67
rect 666 41 696 67
rect 752 41 782 67
rect 838 41 868 67
<< polycont >>
rect 127 285 161 319
rect 416 253 450 287
rect 617 285 651 319
rect 754 285 788 319
rect 822 285 856 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 27 607 161 649
rect 27 573 43 607
rect 77 573 111 607
rect 145 573 161 607
rect 27 509 161 573
rect 27 475 43 509
rect 77 475 111 509
rect 145 475 161 509
rect 27 459 161 475
rect 195 599 233 615
rect 195 565 197 599
rect 231 565 233 599
rect 195 505 233 565
rect 195 471 197 505
rect 231 471 233 505
rect 27 413 91 459
rect 27 379 43 413
rect 77 379 91 413
rect 27 363 91 379
rect 125 334 161 424
rect 195 413 233 471
rect 267 607 333 649
rect 267 573 283 607
rect 317 573 333 607
rect 267 530 333 573
rect 267 496 283 530
rect 317 496 333 530
rect 267 453 333 496
rect 267 419 283 453
rect 317 419 333 453
rect 367 599 403 615
rect 367 565 369 599
rect 367 505 403 565
rect 367 471 369 505
rect 195 379 197 413
rect 231 385 233 413
rect 367 418 403 471
rect 448 607 514 649
rect 448 573 464 607
rect 498 573 514 607
rect 448 493 514 573
rect 448 459 464 493
rect 498 459 514 493
rect 448 452 514 459
rect 548 599 607 615
rect 548 565 557 599
rect 591 565 607 599
rect 548 509 607 565
rect 548 475 557 509
rect 591 475 607 509
rect 548 418 607 475
rect 652 607 718 649
rect 652 573 668 607
rect 702 573 718 607
rect 652 493 718 573
rect 652 459 668 493
rect 702 459 718 493
rect 652 452 718 459
rect 763 599 815 615
rect 763 565 779 599
rect 813 565 815 599
rect 763 509 815 565
rect 763 475 779 509
rect 813 475 815 509
rect 763 434 815 475
rect 763 418 779 434
rect 367 413 557 418
rect 367 385 369 413
rect 231 379 369 385
rect 403 384 557 413
rect 591 400 779 418
rect 813 400 815 434
rect 591 384 815 400
rect 849 607 915 649
rect 849 573 865 607
rect 899 573 915 607
rect 849 509 915 573
rect 849 475 865 509
rect 899 475 915 509
rect 849 418 915 475
rect 849 384 865 418
rect 899 384 915 418
rect 403 379 567 384
rect 195 351 567 379
rect 111 328 161 334
rect 111 319 169 328
rect 403 321 567 351
rect 111 285 127 319
rect 161 285 169 319
rect 111 269 169 285
rect 317 253 416 287
rect 450 253 466 287
rect 317 233 466 253
rect 500 249 567 321
rect 601 319 667 350
rect 601 285 617 319
rect 651 285 667 319
rect 701 319 943 350
rect 701 285 754 319
rect 788 285 822 319
rect 856 285 943 319
rect 61 203 283 231
rect 500 227 843 249
rect 500 215 793 227
rect 61 169 77 203
rect 111 197 249 203
rect 111 169 113 197
rect 61 101 113 169
rect 247 169 249 197
rect 61 67 77 101
rect 111 67 113 101
rect 61 51 113 67
rect 147 157 213 161
rect 147 123 163 157
rect 197 123 213 157
rect 147 89 213 123
rect 147 55 163 89
rect 197 55 213 89
rect 147 17 213 55
rect 247 109 283 169
rect 325 183 391 199
rect 325 149 341 183
rect 375 181 391 183
rect 777 193 793 215
rect 827 193 843 227
rect 375 179 671 181
rect 375 149 621 179
rect 325 145 621 149
rect 655 145 671 179
rect 325 143 671 145
rect 705 165 743 181
rect 705 131 707 165
rect 741 131 743 165
rect 705 109 743 131
rect 777 153 843 193
rect 777 119 793 153
rect 827 119 843 153
rect 877 223 929 239
rect 877 189 879 223
rect 913 189 929 223
rect 247 101 477 109
rect 247 67 249 101
rect 283 99 477 101
rect 283 67 427 99
rect 247 65 427 67
rect 461 65 477 99
rect 247 51 477 65
rect 519 75 535 109
rect 569 85 743 109
rect 877 113 929 189
rect 877 85 879 113
rect 569 79 879 85
rect 913 79 929 113
rect 569 75 929 79
rect 519 51 929 75
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4631382
string GDS_START 4622602
<< end >>
