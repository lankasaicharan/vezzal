magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4082 1975
<< nwell >>
rect -38 331 2822 704
<< pwell >>
rect 2052 241 2366 267
rect 2052 229 2781 241
rect 773 223 1161 229
rect 1667 223 2781 229
rect 773 191 2781 223
rect 9 160 197 184
rect 376 160 2781 191
rect 9 49 2781 160
rect 0 0 2784 49
<< scnmos >>
rect 88 74 118 158
rect 278 50 308 134
rect 350 50 380 134
rect 482 81 512 165
rect 554 81 584 165
rect 643 81 673 165
rect 875 119 905 203
rect 961 119 991 203
rect 1055 119 1085 203
rect 1157 113 1187 197
rect 1290 69 1320 197
rect 1376 69 1406 197
rect 1563 113 1593 197
rect 1635 113 1665 197
rect 1779 119 1809 203
rect 1851 119 1881 203
rect 2135 73 2165 241
rect 2253 73 2283 241
rect 2484 47 2514 131
rect 2586 47 2616 215
rect 2672 47 2702 215
<< scpmoshvt >>
rect 216 468 246 596
rect 302 468 332 596
rect 374 468 404 596
rect 460 468 490 596
rect 554 468 584 596
rect 673 463 703 591
rect 778 463 808 547
rect 864 463 894 547
rect 936 463 966 547
rect 1044 463 1074 547
rect 1329 379 1359 547
rect 1415 379 1445 547
rect 1539 534 1569 618
rect 1657 534 1687 618
rect 1837 534 1867 618
rect 1923 534 1953 618
rect 2136 367 2166 619
rect 2253 367 2283 619
rect 2484 367 2514 495
rect 2586 367 2616 619
rect 2672 367 2702 619
<< ndiff >>
rect 35 133 88 158
rect 35 99 43 133
rect 77 99 88 133
rect 35 74 88 99
rect 118 130 171 158
rect 402 157 482 165
rect 402 134 414 157
rect 118 96 129 130
rect 163 96 171 130
rect 118 74 171 96
rect 225 109 278 134
rect 225 75 233 109
rect 267 75 278 109
rect 225 50 278 75
rect 308 50 350 134
rect 380 123 414 134
rect 448 123 482 157
rect 380 81 482 123
rect 512 81 554 165
rect 584 127 643 165
rect 584 93 595 127
rect 629 93 643 127
rect 584 81 643 93
rect 673 127 739 165
rect 673 93 697 127
rect 731 93 739 127
rect 673 81 739 93
rect 380 50 460 81
rect 799 178 875 203
rect 799 144 809 178
rect 843 144 875 178
rect 799 119 875 144
rect 905 178 961 203
rect 905 144 916 178
rect 950 144 961 178
rect 905 119 961 144
rect 991 119 1055 203
rect 1085 197 1135 203
rect 2078 233 2135 241
rect 1693 197 1779 203
rect 1085 119 1157 197
rect 1107 113 1157 119
rect 1187 119 1290 197
rect 1187 113 1245 119
rect 1237 85 1245 113
rect 1279 85 1290 119
rect 1237 69 1290 85
rect 1320 189 1376 197
rect 1320 155 1331 189
rect 1365 155 1376 189
rect 1320 115 1376 155
rect 1320 81 1331 115
rect 1365 81 1376 115
rect 1320 69 1376 81
rect 1406 183 1563 197
rect 1406 149 1417 183
rect 1451 169 1563 183
rect 1451 149 1518 169
rect 1406 135 1518 149
rect 1552 135 1563 169
rect 1406 115 1563 135
rect 1406 81 1417 115
rect 1451 113 1563 115
rect 1593 113 1635 197
rect 1665 175 1779 197
rect 1665 141 1710 175
rect 1744 141 1779 175
rect 1665 119 1779 141
rect 1809 119 1851 203
rect 1881 178 1934 203
rect 1881 144 1892 178
rect 1926 144 1934 178
rect 1881 119 1934 144
rect 2078 199 2090 233
rect 2124 199 2135 233
rect 1665 113 1743 119
rect 1451 81 1459 113
rect 1406 69 1459 81
rect 2078 73 2135 199
rect 2165 93 2253 241
rect 2165 73 2192 93
rect 2180 59 2192 73
rect 2226 73 2253 93
rect 2283 233 2340 241
rect 2283 199 2294 233
rect 2328 199 2340 233
rect 2283 73 2340 199
rect 2536 131 2586 215
rect 2431 93 2484 131
rect 2226 59 2238 73
rect 2180 51 2238 59
rect 2431 59 2439 93
rect 2473 59 2484 93
rect 2431 47 2484 59
rect 2514 89 2586 131
rect 2514 55 2539 89
rect 2573 55 2586 89
rect 2514 47 2586 55
rect 2616 197 2672 215
rect 2616 163 2627 197
rect 2661 163 2672 197
rect 2616 101 2672 163
rect 2616 67 2627 101
rect 2661 67 2672 101
rect 2616 47 2672 67
rect 2702 203 2755 215
rect 2702 169 2713 203
rect 2747 169 2755 203
rect 2702 93 2755 169
rect 2702 59 2713 93
rect 2747 59 2755 93
rect 2702 47 2755 59
<< pdiff >>
rect 163 584 216 596
rect 163 550 171 584
rect 205 550 216 584
rect 163 514 216 550
rect 163 480 171 514
rect 205 480 216 514
rect 163 468 216 480
rect 246 588 302 596
rect 246 554 257 588
rect 291 554 302 588
rect 246 514 302 554
rect 246 480 257 514
rect 291 480 302 514
rect 246 468 302 480
rect 332 468 374 596
rect 404 584 460 596
rect 404 550 415 584
rect 449 550 460 584
rect 404 510 460 550
rect 404 476 415 510
rect 449 476 460 510
rect 404 468 460 476
rect 490 468 554 596
rect 584 591 637 596
rect 584 570 673 591
rect 584 536 610 570
rect 644 536 673 570
rect 584 468 673 536
rect 623 463 673 468
rect 703 578 756 591
rect 703 544 714 578
rect 748 547 756 578
rect 1257 565 1307 577
rect 748 544 778 547
rect 703 510 778 544
rect 703 476 733 510
rect 767 476 778 510
rect 703 463 778 476
rect 808 523 864 547
rect 808 489 819 523
rect 853 489 864 523
rect 808 463 864 489
rect 894 463 936 547
rect 966 539 1044 547
rect 966 505 987 539
rect 1021 505 1044 539
rect 966 463 1044 505
rect 1074 523 1127 547
rect 1074 489 1085 523
rect 1119 489 1127 523
rect 1257 531 1265 565
rect 1299 547 1307 565
rect 1467 547 1539 618
rect 1299 531 1329 547
rect 1074 463 1127 489
rect 1257 379 1329 531
rect 1359 425 1415 547
rect 1359 391 1370 425
rect 1404 391 1415 425
rect 1359 379 1415 391
rect 1445 534 1539 547
rect 1569 534 1657 618
rect 1687 610 1837 618
rect 1687 576 1698 610
rect 1732 576 1778 610
rect 1812 576 1837 610
rect 1687 534 1837 576
rect 1867 609 1923 618
rect 1867 575 1878 609
rect 1912 575 1923 609
rect 1867 534 1923 575
rect 1953 591 2029 618
rect 1953 557 1985 591
rect 2019 557 2029 591
rect 1953 534 2029 557
rect 1445 455 1517 534
rect 1445 421 1464 455
rect 1498 421 1517 455
rect 1445 379 1517 421
rect 2083 413 2136 619
rect 2083 379 2091 413
rect 2125 379 2136 413
rect 2083 367 2136 379
rect 2166 583 2253 619
rect 2166 549 2186 583
rect 2220 549 2253 583
rect 2166 367 2253 549
rect 2283 570 2336 619
rect 2283 536 2294 570
rect 2328 536 2336 570
rect 2283 367 2336 536
rect 2533 607 2586 619
rect 2533 573 2541 607
rect 2575 573 2586 607
rect 2533 522 2586 573
rect 2533 495 2541 522
rect 2431 483 2484 495
rect 2431 449 2439 483
rect 2473 449 2484 483
rect 2431 413 2484 449
rect 2431 379 2439 413
rect 2473 379 2484 413
rect 2431 367 2484 379
rect 2514 488 2541 495
rect 2575 488 2586 522
rect 2514 437 2586 488
rect 2514 403 2525 437
rect 2559 403 2586 437
rect 2514 367 2586 403
rect 2616 599 2672 619
rect 2616 565 2627 599
rect 2661 565 2672 599
rect 2616 500 2672 565
rect 2616 466 2627 500
rect 2661 466 2672 500
rect 2616 409 2672 466
rect 2616 375 2627 409
rect 2661 375 2672 409
rect 2616 367 2672 375
rect 2702 607 2755 619
rect 2702 573 2713 607
rect 2747 573 2755 607
rect 2702 512 2755 573
rect 2702 478 2713 512
rect 2747 478 2755 512
rect 2702 413 2755 478
rect 2702 379 2713 413
rect 2747 379 2755 413
rect 2702 367 2755 379
<< ndiffc >>
rect 43 99 77 133
rect 129 96 163 130
rect 233 75 267 109
rect 414 123 448 157
rect 595 93 629 127
rect 697 93 731 127
rect 809 144 843 178
rect 916 144 950 178
rect 1245 85 1279 119
rect 1331 155 1365 189
rect 1331 81 1365 115
rect 1417 149 1451 183
rect 1518 135 1552 169
rect 1417 81 1451 115
rect 1710 141 1744 175
rect 1892 144 1926 178
rect 2090 199 2124 233
rect 2192 59 2226 93
rect 2294 199 2328 233
rect 2439 59 2473 93
rect 2539 55 2573 89
rect 2627 163 2661 197
rect 2627 67 2661 101
rect 2713 169 2747 203
rect 2713 59 2747 93
<< pdiffc >>
rect 171 550 205 584
rect 171 480 205 514
rect 257 554 291 588
rect 257 480 291 514
rect 415 550 449 584
rect 415 476 449 510
rect 610 536 644 570
rect 714 544 748 578
rect 733 476 767 510
rect 819 489 853 523
rect 987 505 1021 539
rect 1085 489 1119 523
rect 1265 531 1299 565
rect 1370 391 1404 425
rect 1698 576 1732 610
rect 1778 576 1812 610
rect 1878 575 1912 609
rect 1985 557 2019 591
rect 1464 421 1498 455
rect 2091 379 2125 413
rect 2186 549 2220 583
rect 2294 536 2328 570
rect 2541 573 2575 607
rect 2439 449 2473 483
rect 2439 379 2473 413
rect 2541 488 2575 522
rect 2525 403 2559 437
rect 2627 565 2661 599
rect 2627 466 2661 500
rect 2627 375 2661 409
rect 2713 573 2747 607
rect 2713 478 2747 512
rect 2713 379 2747 413
<< poly >>
rect 216 596 246 622
rect 302 596 332 622
rect 374 596 404 622
rect 460 596 490 622
rect 554 596 584 622
rect 673 591 703 617
rect 864 615 1445 645
rect 1539 618 1569 644
rect 1657 618 1687 644
rect 1837 618 1867 644
rect 1923 618 1953 644
rect 2136 619 2166 645
rect 2253 619 2283 645
rect 2586 619 2616 645
rect 2672 619 2702 645
rect 216 442 246 468
rect 302 442 332 468
rect 88 412 332 442
rect 88 276 183 412
rect 374 364 404 468
rect 460 436 490 468
rect 446 420 512 436
rect 446 386 462 420
rect 496 386 512 420
rect 446 370 512 386
rect 554 399 584 468
rect 778 547 808 573
rect 864 547 894 615
rect 936 547 966 573
rect 1044 547 1074 573
rect 1329 547 1359 573
rect 1415 547 1445 615
rect 1151 492 1225 508
rect 554 383 631 399
rect 554 369 581 383
rect 332 348 404 364
rect 332 314 348 348
rect 382 334 404 348
rect 565 349 581 369
rect 615 349 631 383
rect 382 314 398 334
rect 332 298 398 314
rect 565 315 631 349
rect 88 242 133 276
rect 167 242 183 276
rect 88 226 183 242
rect 88 158 118 226
rect 236 206 308 222
rect 236 172 252 206
rect 286 172 308 206
rect 236 156 308 172
rect 278 134 308 156
rect 350 134 380 298
rect 446 276 512 292
rect 446 242 462 276
rect 496 242 512 276
rect 565 281 581 315
rect 615 281 631 315
rect 565 267 631 281
rect 446 226 512 242
rect 482 165 512 226
rect 554 265 631 267
rect 554 237 595 265
rect 554 165 584 237
rect 673 217 703 463
rect 778 399 808 463
rect 756 383 822 399
rect 756 349 772 383
rect 806 349 822 383
rect 756 315 822 349
rect 756 281 772 315
rect 806 281 822 315
rect 756 265 822 281
rect 864 285 894 463
rect 936 399 966 463
rect 1044 441 1074 463
rect 1151 458 1175 492
rect 1209 458 1225 492
rect 1151 441 1225 458
rect 1044 424 1225 441
rect 1044 411 1175 424
rect 936 383 1002 399
rect 936 349 952 383
rect 986 369 1002 383
rect 1151 390 1175 411
rect 1209 390 1225 424
rect 1151 374 1225 390
rect 1539 485 1569 534
rect 1539 469 1615 485
rect 1539 435 1565 469
rect 1599 435 1615 469
rect 1539 419 1615 435
rect 1657 455 1687 534
rect 1837 502 1867 534
rect 1815 486 1881 502
rect 1657 439 1773 455
rect 1657 425 1723 439
rect 1707 405 1723 425
rect 1757 405 1773 439
rect 1815 452 1831 486
rect 1865 452 1881 486
rect 1815 436 1881 452
rect 1707 389 1773 405
rect 986 349 1091 369
rect 936 339 1091 349
rect 936 333 1002 339
rect 864 255 905 285
rect 643 187 784 217
rect 875 203 905 255
rect 947 275 1013 291
rect 1061 285 1091 339
rect 947 241 963 275
rect 997 241 1013 275
rect 947 225 1013 241
rect 1055 255 1091 285
rect 961 203 991 225
rect 1055 203 1085 255
rect 1151 249 1181 374
rect 1329 327 1359 379
rect 1415 357 1445 379
rect 1563 361 1665 377
rect 1563 357 1615 361
rect 1415 327 1615 357
rect 1649 327 1665 361
rect 1290 297 1359 327
rect 1563 311 1665 327
rect 1290 285 1320 297
rect 1229 269 1320 285
rect 1151 219 1187 249
rect 1229 235 1245 269
rect 1279 235 1320 269
rect 1455 269 1521 285
rect 1455 249 1471 269
rect 1229 219 1320 235
rect 643 165 673 187
rect 88 48 118 74
rect 482 55 512 81
rect 554 55 584 81
rect 643 51 673 81
rect 754 51 784 187
rect 1157 197 1187 219
rect 1290 197 1320 219
rect 1376 235 1471 249
rect 1505 235 1521 269
rect 1376 219 1521 235
rect 1376 197 1406 219
rect 1563 197 1593 311
rect 1707 249 1737 389
rect 1851 333 1881 436
rect 1635 219 1737 249
rect 1779 303 1881 333
rect 1635 197 1665 219
rect 1779 203 1809 303
rect 1923 299 1953 534
rect 2484 495 2514 521
rect 2136 335 2166 367
rect 2135 319 2211 335
rect 1923 275 1989 299
rect 1923 255 1939 275
rect 1851 241 1939 255
rect 1973 241 1989 275
rect 2135 285 2161 319
rect 2195 285 2211 319
rect 2135 269 2211 285
rect 2253 299 2283 367
rect 2328 319 2394 335
rect 2328 299 2344 319
rect 2253 285 2344 299
rect 2378 285 2394 319
rect 2484 317 2514 367
rect 2253 269 2394 285
rect 2442 301 2514 317
rect 2586 315 2616 367
rect 2672 315 2702 367
rect 2135 241 2165 269
rect 2253 241 2283 269
rect 2442 267 2458 301
rect 2492 267 2514 301
rect 1851 225 1989 241
rect 1851 203 1881 225
rect 875 93 905 119
rect 961 93 991 119
rect 1055 93 1085 119
rect 1157 51 1187 113
rect 1563 87 1593 113
rect 278 24 308 50
rect 350 24 380 50
rect 643 21 1187 51
rect 1290 43 1320 69
rect 1376 43 1406 69
rect 1635 51 1665 113
rect 1779 93 1809 119
rect 1851 93 1881 119
rect 1956 87 2022 103
rect 1956 53 1972 87
rect 2006 53 2022 87
rect 1956 51 2022 53
rect 1635 21 2022 51
rect 2135 47 2165 73
rect 2442 233 2514 267
rect 2556 299 2702 315
rect 2556 265 2572 299
rect 2606 265 2702 299
rect 2556 249 2702 265
rect 2442 199 2458 233
rect 2492 199 2514 233
rect 2586 215 2616 249
rect 2672 215 2702 249
rect 2442 171 2514 199
rect 2484 131 2514 171
rect 2253 47 2283 73
rect 2484 21 2514 47
rect 2586 21 2616 47
rect 2672 21 2702 47
<< polycont >>
rect 462 386 496 420
rect 348 314 382 348
rect 581 349 615 383
rect 133 242 167 276
rect 252 172 286 206
rect 462 242 496 276
rect 581 281 615 315
rect 772 349 806 383
rect 772 281 806 315
rect 1175 458 1209 492
rect 952 349 986 383
rect 1175 390 1209 424
rect 1565 435 1599 469
rect 1723 405 1757 439
rect 1831 452 1865 486
rect 963 241 997 275
rect 1615 327 1649 361
rect 1245 235 1279 269
rect 1471 235 1505 269
rect 1939 241 1973 275
rect 2161 285 2195 319
rect 2344 285 2378 319
rect 2458 267 2492 301
rect 1972 53 2006 87
rect 2572 265 2606 299
rect 2458 199 2492 233
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 27 584 207 600
rect 27 550 171 584
rect 205 550 207 584
rect 27 514 207 550
rect 27 480 171 514
rect 205 480 207 514
rect 27 426 207 480
rect 241 588 295 649
rect 241 554 257 588
rect 291 554 295 588
rect 241 514 295 554
rect 241 480 257 514
rect 291 480 295 514
rect 241 464 295 480
rect 399 584 465 600
rect 399 550 415 584
rect 449 550 465 584
rect 399 510 465 550
rect 594 570 660 649
rect 594 536 610 570
rect 644 536 660 570
rect 594 528 660 536
rect 702 578 777 594
rect 702 544 714 578
rect 748 544 777 578
rect 399 476 415 510
rect 449 494 465 510
rect 702 510 777 544
rect 971 539 1037 649
rect 1249 565 1315 649
rect 1682 610 1828 649
rect 1682 576 1698 610
rect 1732 576 1778 610
rect 1812 576 1828 610
rect 1682 573 1828 576
rect 1862 609 1951 615
rect 1862 575 1878 609
rect 1912 575 1951 609
rect 1862 573 1951 575
rect 702 494 733 510
rect 449 476 733 494
rect 767 476 777 510
rect 399 460 777 476
rect 811 523 877 539
rect 811 489 819 523
rect 853 489 877 523
rect 971 505 987 539
rect 1021 505 1037 539
rect 971 503 1037 505
rect 1071 523 1125 539
rect 1249 531 1265 565
rect 1299 531 1315 565
rect 1249 529 1315 531
rect 811 469 877 489
rect 1071 489 1085 523
rect 1119 489 1125 523
rect 1351 505 1881 539
rect 1351 495 1385 505
rect 1071 469 1125 489
rect 27 420 512 426
rect 27 386 462 420
rect 496 386 512 420
rect 27 206 81 386
rect 581 383 657 426
rect 115 348 547 352
rect 115 314 348 348
rect 382 314 547 348
rect 115 310 547 314
rect 615 349 657 383
rect 581 315 657 349
rect 615 281 657 315
rect 115 242 133 276
rect 167 242 462 276
rect 496 242 547 276
rect 581 242 657 281
rect 115 240 547 242
rect 27 172 252 206
rect 286 172 302 206
rect 691 201 736 460
rect 811 435 1125 469
rect 1159 492 1385 495
rect 1159 458 1175 492
rect 1209 461 1385 492
rect 1815 486 1881 505
rect 1209 458 1225 461
rect 770 383 843 399
rect 770 349 772 383
rect 806 349 843 383
rect 770 315 843 349
rect 770 281 772 315
rect 806 281 843 315
rect 770 276 843 281
rect 770 242 799 276
rect 833 242 843 276
rect 770 235 843 242
rect 398 178 843 201
rect 27 133 79 172
rect 398 167 809 178
rect 398 157 464 167
rect 27 99 43 133
rect 77 99 79 133
rect 27 83 79 99
rect 113 130 179 138
rect 113 96 129 130
rect 163 96 179 130
rect 113 17 179 96
rect 217 109 283 125
rect 398 123 414 157
rect 448 123 464 157
rect 791 144 809 167
rect 398 121 464 123
rect 579 127 645 133
rect 217 75 233 109
rect 267 87 283 109
rect 579 93 595 127
rect 629 93 645 127
rect 579 87 645 93
rect 267 75 645 87
rect 217 53 645 75
rect 681 127 747 133
rect 791 128 843 144
rect 877 199 911 435
rect 1159 424 1225 458
rect 1454 455 1511 471
rect 945 383 1002 399
rect 1159 390 1175 424
rect 1209 390 1225 424
rect 1331 425 1420 427
rect 1331 391 1370 425
rect 1404 391 1420 425
rect 945 349 952 383
rect 986 354 1002 383
rect 1331 389 1420 391
rect 1454 421 1464 455
rect 1498 421 1511 455
rect 1331 354 1367 389
rect 1454 355 1511 421
rect 986 349 1367 354
rect 945 320 1367 349
rect 947 276 1040 286
rect 947 275 991 276
rect 947 241 963 275
rect 1025 242 1040 276
rect 997 241 1040 242
rect 947 233 1040 241
rect 1229 269 1295 286
rect 1229 235 1245 269
rect 1279 235 1295 269
rect 1229 199 1295 235
rect 877 178 1295 199
rect 877 144 916 178
rect 950 157 1295 178
rect 1329 189 1367 320
rect 950 144 960 157
rect 877 128 960 144
rect 1329 155 1331 189
rect 1365 155 1367 189
rect 681 93 697 127
rect 731 93 747 127
rect 681 17 747 93
rect 1229 119 1295 123
rect 1229 85 1245 119
rect 1279 85 1295 119
rect 1229 17 1295 85
rect 1329 115 1367 155
rect 1329 81 1331 115
rect 1365 81 1367 115
rect 1329 65 1367 81
rect 1401 321 1511 355
rect 1545 469 1615 471
rect 1545 435 1565 469
rect 1599 435 1615 469
rect 1545 419 1615 435
rect 1707 439 1773 455
rect 1815 452 1831 486
rect 1865 452 1881 486
rect 1815 450 1881 452
rect 1401 185 1435 321
rect 1545 285 1579 419
rect 1707 405 1723 439
rect 1757 416 1773 439
rect 1917 416 1951 573
rect 1985 591 2035 649
rect 2019 557 2035 591
rect 1985 541 2035 557
rect 2161 583 2224 649
rect 2509 607 2589 649
rect 2161 549 2186 583
rect 2220 549 2224 583
rect 2161 533 2224 549
rect 2258 570 2344 588
rect 2258 536 2294 570
rect 2328 536 2344 570
rect 2258 532 2344 536
rect 2509 573 2541 607
rect 2575 573 2589 607
rect 2258 499 2292 532
rect 2509 522 2589 573
rect 1757 405 1951 416
rect 1707 382 1951 405
rect 1987 465 2292 499
rect 1613 361 1665 377
rect 1613 327 1615 361
rect 1649 346 1665 361
rect 1987 346 2021 465
rect 1649 327 2021 346
rect 1613 312 2021 327
rect 2075 413 2127 431
rect 2075 379 2091 413
rect 2125 379 2127 413
rect 1613 311 1649 312
rect 2075 285 2127 379
rect 1469 276 1579 285
rect 1469 235 1471 276
rect 1505 235 1579 276
rect 2042 276 2127 285
rect 1469 219 1579 235
rect 1613 241 1939 275
rect 1973 241 2000 275
rect 1613 185 1647 241
rect 1401 183 1647 185
rect 1401 149 1417 183
rect 1451 169 1647 183
rect 1451 149 1518 169
rect 1401 135 1518 149
rect 1552 135 1647 169
rect 1401 115 1647 135
rect 1401 81 1417 115
rect 1451 81 1647 115
rect 1401 65 1647 81
rect 1694 175 1760 191
rect 1694 141 1710 175
rect 1744 141 1760 175
rect 1694 17 1760 141
rect 1876 178 1932 194
rect 1876 144 1892 178
rect 1926 144 1932 178
rect 1876 95 1932 144
rect 1966 163 2000 241
rect 2042 242 2047 276
rect 2081 242 2127 276
rect 2161 319 2292 465
rect 2195 285 2292 319
rect 2161 269 2292 285
rect 2326 319 2401 498
rect 2435 483 2475 499
rect 2435 449 2439 483
rect 2473 449 2475 483
rect 2435 413 2475 449
rect 2435 379 2439 413
rect 2473 379 2475 413
rect 2509 488 2541 522
rect 2575 488 2589 522
rect 2509 437 2589 488
rect 2509 403 2525 437
rect 2559 403 2589 437
rect 2623 599 2675 615
rect 2623 565 2627 599
rect 2661 565 2675 599
rect 2623 500 2675 565
rect 2623 466 2627 500
rect 2661 466 2675 500
rect 2623 409 2675 466
rect 2435 369 2475 379
rect 2623 375 2627 409
rect 2661 375 2675 409
rect 2435 335 2578 369
rect 2623 351 2675 375
rect 2709 607 2763 649
rect 2709 573 2713 607
rect 2747 573 2763 607
rect 2709 512 2763 573
rect 2709 478 2713 512
rect 2747 478 2763 512
rect 2709 413 2763 478
rect 2709 379 2713 413
rect 2747 379 2763 413
rect 2709 363 2763 379
rect 2326 285 2344 319
rect 2378 285 2401 319
rect 2544 315 2578 335
rect 2326 283 2401 285
rect 2042 233 2127 242
rect 2258 249 2292 269
rect 2442 267 2458 301
rect 2492 267 2508 301
rect 2442 249 2508 267
rect 2258 233 2344 249
rect 2042 199 2090 233
rect 2124 199 2140 233
rect 2042 197 2140 199
rect 2258 199 2294 233
rect 2328 199 2344 233
rect 2258 197 2344 199
rect 2380 233 2508 249
rect 2380 199 2458 233
rect 2492 199 2508 233
rect 2544 299 2606 315
rect 2544 265 2572 299
rect 2544 249 2606 265
rect 2380 163 2414 199
rect 2544 163 2589 249
rect 2640 213 2675 351
rect 1966 129 2414 163
rect 2455 129 2589 163
rect 2623 197 2675 213
rect 2623 163 2627 197
rect 2661 163 2675 197
rect 1876 87 2022 95
rect 1876 53 1972 87
rect 2006 53 2022 87
rect 1876 51 2022 53
rect 2176 93 2242 95
rect 2455 93 2489 129
rect 2623 101 2675 163
rect 2176 59 2192 93
rect 2226 59 2242 93
rect 2176 17 2242 59
rect 2423 59 2439 93
rect 2473 59 2489 93
rect 2423 55 2489 59
rect 2523 89 2589 95
rect 2523 55 2539 89
rect 2573 55 2589 89
rect 2523 17 2589 55
rect 2623 67 2627 101
rect 2661 67 2675 101
rect 2623 51 2675 67
rect 2709 203 2763 219
rect 2709 169 2713 203
rect 2747 169 2763 203
rect 2709 93 2763 169
rect 2709 59 2713 93
rect 2747 59 2763 93
rect 2709 17 2763 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 799 242 833 276
rect 991 275 1025 276
rect 991 242 997 275
rect 997 242 1025 275
rect 1471 269 1505 276
rect 1471 242 1505 269
rect 2047 242 2081 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 787 276 845 282
rect 787 242 799 276
rect 833 273 845 276
rect 979 276 1037 282
rect 979 273 991 276
rect 833 245 991 273
rect 833 242 845 245
rect 787 236 845 242
rect 979 242 991 245
rect 1025 273 1037 276
rect 1459 276 1517 282
rect 1459 273 1471 276
rect 1025 245 1471 273
rect 1025 242 1037 245
rect 979 236 1037 242
rect 1459 242 1471 245
rect 1505 273 1517 276
rect 2035 276 2093 282
rect 2035 273 2047 276
rect 1505 245 2047 273
rect 1505 242 1517 245
rect 1459 236 1517 242
rect 2035 242 2047 245
rect 2081 242 2093 276
rect 2035 236 2093 242
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfrtp_2
flabel comment s 1722 326 1722 326 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 1183 390 1217 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 2335 316 2369 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2335 390 2369 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2335 464 2369 498 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2623 390 2657 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 464 2657 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 538 2657 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3289420
string GDS_START 3268418
<< end >>
