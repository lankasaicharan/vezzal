magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1260 -1253 16260 40860
<< metal3 >>
rect 100 10163 4880 10164
rect 100 10099 106 10163
rect 170 10099 188 10163
rect 252 10099 270 10163
rect 334 10099 352 10163
rect 416 10099 434 10163
rect 498 10099 516 10163
rect 580 10099 598 10163
rect 662 10099 679 10163
rect 743 10099 760 10163
rect 824 10099 841 10163
rect 905 10099 922 10163
rect 986 10099 1003 10163
rect 1067 10099 1084 10163
rect 1148 10099 1165 10163
rect 1229 10099 1246 10163
rect 1310 10099 1327 10163
rect 1391 10099 1408 10163
rect 1472 10099 1489 10163
rect 1553 10099 1570 10163
rect 1634 10099 1651 10163
rect 1715 10099 1732 10163
rect 1796 10099 1813 10163
rect 1877 10099 1894 10163
rect 1958 10099 1975 10163
rect 2039 10099 2056 10163
rect 2120 10099 2137 10163
rect 2201 10099 2218 10163
rect 2282 10099 2299 10163
rect 2363 10099 2380 10163
rect 2444 10099 2461 10163
rect 2525 10099 2542 10163
rect 2606 10099 2623 10163
rect 2687 10099 2704 10163
rect 2768 10099 2785 10163
rect 2849 10099 2866 10163
rect 2930 10099 2947 10163
rect 3011 10099 3028 10163
rect 3092 10099 3109 10163
rect 3173 10099 3190 10163
rect 3254 10099 3271 10163
rect 3335 10099 3352 10163
rect 3416 10099 3433 10163
rect 3497 10099 3514 10163
rect 3578 10099 3595 10163
rect 3659 10099 3676 10163
rect 3740 10099 3757 10163
rect 3821 10099 3838 10163
rect 3902 10099 3919 10163
rect 3983 10099 4000 10163
rect 4064 10099 4081 10163
rect 4145 10099 4162 10163
rect 4226 10099 4243 10163
rect 4307 10099 4324 10163
rect 4388 10099 4405 10163
rect 4469 10099 4486 10163
rect 4550 10099 4567 10163
rect 4631 10099 4648 10163
rect 4712 10099 4729 10163
rect 4793 10099 4810 10163
rect 4874 10099 4880 10163
rect 100 10079 4880 10099
rect 100 10015 106 10079
rect 170 10015 188 10079
rect 252 10015 270 10079
rect 334 10015 352 10079
rect 416 10015 434 10079
rect 498 10015 516 10079
rect 580 10015 598 10079
rect 662 10015 679 10079
rect 743 10015 760 10079
rect 824 10015 841 10079
rect 905 10015 922 10079
rect 986 10015 1003 10079
rect 1067 10015 1084 10079
rect 1148 10015 1165 10079
rect 1229 10015 1246 10079
rect 1310 10015 1327 10079
rect 1391 10015 1408 10079
rect 1472 10015 1489 10079
rect 1553 10015 1570 10079
rect 1634 10015 1651 10079
rect 1715 10015 1732 10079
rect 1796 10015 1813 10079
rect 1877 10015 1894 10079
rect 1958 10015 1975 10079
rect 2039 10015 2056 10079
rect 2120 10015 2137 10079
rect 2201 10015 2218 10079
rect 2282 10015 2299 10079
rect 2363 10015 2380 10079
rect 2444 10015 2461 10079
rect 2525 10015 2542 10079
rect 2606 10015 2623 10079
rect 2687 10015 2704 10079
rect 2768 10015 2785 10079
rect 2849 10015 2866 10079
rect 2930 10015 2947 10079
rect 3011 10015 3028 10079
rect 3092 10015 3109 10079
rect 3173 10015 3190 10079
rect 3254 10015 3271 10079
rect 3335 10015 3352 10079
rect 3416 10015 3433 10079
rect 3497 10015 3514 10079
rect 3578 10015 3595 10079
rect 3659 10015 3676 10079
rect 3740 10015 3757 10079
rect 3821 10015 3838 10079
rect 3902 10015 3919 10079
rect 3983 10015 4000 10079
rect 4064 10015 4081 10079
rect 4145 10015 4162 10079
rect 4226 10015 4243 10079
rect 4307 10015 4324 10079
rect 4388 10015 4405 10079
rect 4469 10015 4486 10079
rect 4550 10015 4567 10079
rect 4631 10015 4648 10079
rect 4712 10015 4729 10079
rect 4793 10015 4810 10079
rect 4874 10015 4880 10079
rect 100 9995 4880 10015
rect 100 9931 106 9995
rect 170 9931 188 9995
rect 252 9931 270 9995
rect 334 9931 352 9995
rect 416 9931 434 9995
rect 498 9931 516 9995
rect 580 9931 598 9995
rect 662 9931 679 9995
rect 743 9931 760 9995
rect 824 9931 841 9995
rect 905 9931 922 9995
rect 986 9931 1003 9995
rect 1067 9931 1084 9995
rect 1148 9931 1165 9995
rect 1229 9931 1246 9995
rect 1310 9931 1327 9995
rect 1391 9931 1408 9995
rect 1472 9931 1489 9995
rect 1553 9931 1570 9995
rect 1634 9931 1651 9995
rect 1715 9931 1732 9995
rect 1796 9931 1813 9995
rect 1877 9931 1894 9995
rect 1958 9931 1975 9995
rect 2039 9931 2056 9995
rect 2120 9931 2137 9995
rect 2201 9931 2218 9995
rect 2282 9931 2299 9995
rect 2363 9931 2380 9995
rect 2444 9931 2461 9995
rect 2525 9931 2542 9995
rect 2606 9931 2623 9995
rect 2687 9931 2704 9995
rect 2768 9931 2785 9995
rect 2849 9931 2866 9995
rect 2930 9931 2947 9995
rect 3011 9931 3028 9995
rect 3092 9931 3109 9995
rect 3173 9931 3190 9995
rect 3254 9931 3271 9995
rect 3335 9931 3352 9995
rect 3416 9931 3433 9995
rect 3497 9931 3514 9995
rect 3578 9931 3595 9995
rect 3659 9931 3676 9995
rect 3740 9931 3757 9995
rect 3821 9931 3838 9995
rect 3902 9931 3919 9995
rect 3983 9931 4000 9995
rect 4064 9931 4081 9995
rect 4145 9931 4162 9995
rect 4226 9931 4243 9995
rect 4307 9931 4324 9995
rect 4388 9931 4405 9995
rect 4469 9931 4486 9995
rect 4550 9931 4567 9995
rect 4631 9931 4648 9995
rect 4712 9931 4729 9995
rect 4793 9931 4810 9995
rect 4874 9931 4880 9995
rect 100 9930 4880 9931
rect 10151 10163 14931 10164
rect 10151 10099 10157 10163
rect 10221 10099 10239 10163
rect 10303 10099 10321 10163
rect 10385 10099 10403 10163
rect 10467 10099 10485 10163
rect 10549 10099 10567 10163
rect 10631 10099 10649 10163
rect 10713 10099 10730 10163
rect 10794 10099 10811 10163
rect 10875 10099 10892 10163
rect 10956 10099 10973 10163
rect 11037 10099 11054 10163
rect 11118 10099 11135 10163
rect 11199 10099 11216 10163
rect 11280 10099 11297 10163
rect 11361 10099 11378 10163
rect 11442 10099 11459 10163
rect 11523 10099 11540 10163
rect 11604 10099 11621 10163
rect 11685 10099 11702 10163
rect 11766 10099 11783 10163
rect 11847 10099 11864 10163
rect 11928 10099 11945 10163
rect 12009 10099 12026 10163
rect 12090 10099 12107 10163
rect 12171 10099 12188 10163
rect 12252 10099 12269 10163
rect 12333 10099 12350 10163
rect 12414 10099 12431 10163
rect 12495 10099 12512 10163
rect 12576 10099 12593 10163
rect 12657 10099 12674 10163
rect 12738 10099 12755 10163
rect 12819 10099 12836 10163
rect 12900 10099 12917 10163
rect 12981 10099 12998 10163
rect 13062 10099 13079 10163
rect 13143 10099 13160 10163
rect 13224 10099 13241 10163
rect 13305 10099 13322 10163
rect 13386 10099 13403 10163
rect 13467 10099 13484 10163
rect 13548 10099 13565 10163
rect 13629 10099 13646 10163
rect 13710 10099 13727 10163
rect 13791 10099 13808 10163
rect 13872 10099 13889 10163
rect 13953 10099 13970 10163
rect 14034 10099 14051 10163
rect 14115 10099 14132 10163
rect 14196 10099 14213 10163
rect 14277 10099 14294 10163
rect 14358 10099 14375 10163
rect 14439 10099 14456 10163
rect 14520 10099 14537 10163
rect 14601 10099 14618 10163
rect 14682 10099 14699 10163
rect 14763 10099 14780 10163
rect 14844 10099 14861 10163
rect 14925 10099 14931 10163
rect 10151 10079 14931 10099
rect 10151 10015 10157 10079
rect 10221 10015 10239 10079
rect 10303 10015 10321 10079
rect 10385 10015 10403 10079
rect 10467 10015 10485 10079
rect 10549 10015 10567 10079
rect 10631 10015 10649 10079
rect 10713 10015 10730 10079
rect 10794 10015 10811 10079
rect 10875 10015 10892 10079
rect 10956 10015 10973 10079
rect 11037 10015 11054 10079
rect 11118 10015 11135 10079
rect 11199 10015 11216 10079
rect 11280 10015 11297 10079
rect 11361 10015 11378 10079
rect 11442 10015 11459 10079
rect 11523 10015 11540 10079
rect 11604 10015 11621 10079
rect 11685 10015 11702 10079
rect 11766 10015 11783 10079
rect 11847 10015 11864 10079
rect 11928 10015 11945 10079
rect 12009 10015 12026 10079
rect 12090 10015 12107 10079
rect 12171 10015 12188 10079
rect 12252 10015 12269 10079
rect 12333 10015 12350 10079
rect 12414 10015 12431 10079
rect 12495 10015 12512 10079
rect 12576 10015 12593 10079
rect 12657 10015 12674 10079
rect 12738 10015 12755 10079
rect 12819 10015 12836 10079
rect 12900 10015 12917 10079
rect 12981 10015 12998 10079
rect 13062 10015 13079 10079
rect 13143 10015 13160 10079
rect 13224 10015 13241 10079
rect 13305 10015 13322 10079
rect 13386 10015 13403 10079
rect 13467 10015 13484 10079
rect 13548 10015 13565 10079
rect 13629 10015 13646 10079
rect 13710 10015 13727 10079
rect 13791 10015 13808 10079
rect 13872 10015 13889 10079
rect 13953 10015 13970 10079
rect 14034 10015 14051 10079
rect 14115 10015 14132 10079
rect 14196 10015 14213 10079
rect 14277 10015 14294 10079
rect 14358 10015 14375 10079
rect 14439 10015 14456 10079
rect 14520 10015 14537 10079
rect 14601 10015 14618 10079
rect 14682 10015 14699 10079
rect 14763 10015 14780 10079
rect 14844 10015 14861 10079
rect 14925 10015 14931 10079
rect 10151 9995 14931 10015
rect 10151 9931 10157 9995
rect 10221 9931 10239 9995
rect 10303 9931 10321 9995
rect 10385 9931 10403 9995
rect 10467 9931 10485 9995
rect 10549 9931 10567 9995
rect 10631 9931 10649 9995
rect 10713 9931 10730 9995
rect 10794 9931 10811 9995
rect 10875 9931 10892 9995
rect 10956 9931 10973 9995
rect 11037 9931 11054 9995
rect 11118 9931 11135 9995
rect 11199 9931 11216 9995
rect 11280 9931 11297 9995
rect 11361 9931 11378 9995
rect 11442 9931 11459 9995
rect 11523 9931 11540 9995
rect 11604 9931 11621 9995
rect 11685 9931 11702 9995
rect 11766 9931 11783 9995
rect 11847 9931 11864 9995
rect 11928 9931 11945 9995
rect 12009 9931 12026 9995
rect 12090 9931 12107 9995
rect 12171 9931 12188 9995
rect 12252 9931 12269 9995
rect 12333 9931 12350 9995
rect 12414 9931 12431 9995
rect 12495 9931 12512 9995
rect 12576 9931 12593 9995
rect 12657 9931 12674 9995
rect 12738 9931 12755 9995
rect 12819 9931 12836 9995
rect 12900 9931 12917 9995
rect 12981 9931 12998 9995
rect 13062 9931 13079 9995
rect 13143 9931 13160 9995
rect 13224 9931 13241 9995
rect 13305 9931 13322 9995
rect 13386 9931 13403 9995
rect 13467 9931 13484 9995
rect 13548 9931 13565 9995
rect 13629 9931 13646 9995
rect 13710 9931 13727 9995
rect 13791 9931 13808 9995
rect 13872 9931 13889 9995
rect 13953 9931 13970 9995
rect 14034 9931 14051 9995
rect 14115 9931 14132 9995
rect 14196 9931 14213 9995
rect 14277 9931 14294 9995
rect 14358 9931 14375 9995
rect 14439 9931 14456 9995
rect 14520 9931 14537 9995
rect 14601 9931 14618 9995
rect 14682 9931 14699 9995
rect 14763 9931 14780 9995
rect 14844 9931 14861 9995
rect 14925 9931 14931 9995
rect 10151 9930 14931 9931
rect 100 7632 4880 7636
rect 100 7568 106 7632
rect 170 7568 188 7632
rect 252 7568 270 7632
rect 334 7568 352 7632
rect 416 7568 434 7632
rect 498 7568 516 7632
rect 580 7568 598 7632
rect 662 7568 679 7632
rect 743 7568 760 7632
rect 824 7568 841 7632
rect 905 7568 922 7632
rect 986 7568 1003 7632
rect 1067 7568 1084 7632
rect 1148 7568 1165 7632
rect 1229 7568 1246 7632
rect 1310 7568 1327 7632
rect 1391 7568 1408 7632
rect 1472 7568 1489 7632
rect 1553 7568 1570 7632
rect 1634 7568 1651 7632
rect 1715 7568 1732 7632
rect 1796 7568 1813 7632
rect 1877 7568 1894 7632
rect 1958 7568 1975 7632
rect 2039 7568 2056 7632
rect 2120 7568 2137 7632
rect 2201 7568 2218 7632
rect 2282 7568 2299 7632
rect 2363 7568 2380 7632
rect 2444 7568 2461 7632
rect 2525 7568 2542 7632
rect 2606 7568 2623 7632
rect 2687 7568 2704 7632
rect 2768 7568 2785 7632
rect 2849 7568 2866 7632
rect 2930 7568 2947 7632
rect 3011 7568 3028 7632
rect 3092 7568 3109 7632
rect 3173 7568 3190 7632
rect 3254 7568 3271 7632
rect 3335 7568 3352 7632
rect 3416 7568 3433 7632
rect 3497 7568 3514 7632
rect 3578 7568 3595 7632
rect 3659 7568 3676 7632
rect 3740 7568 3757 7632
rect 3821 7568 3838 7632
rect 3902 7568 3919 7632
rect 3983 7568 4000 7632
rect 4064 7568 4081 7632
rect 4145 7568 4162 7632
rect 4226 7568 4243 7632
rect 4307 7568 4324 7632
rect 4388 7568 4405 7632
rect 4469 7568 4486 7632
rect 4550 7568 4567 7632
rect 4631 7568 4648 7632
rect 4712 7568 4729 7632
rect 4793 7568 4810 7632
rect 4874 7568 4880 7632
rect 100 7544 4880 7568
rect 100 7480 106 7544
rect 170 7480 188 7544
rect 252 7480 270 7544
rect 334 7480 352 7544
rect 416 7480 434 7544
rect 498 7480 516 7544
rect 580 7480 598 7544
rect 662 7480 679 7544
rect 743 7480 760 7544
rect 824 7480 841 7544
rect 905 7480 922 7544
rect 986 7480 1003 7544
rect 1067 7480 1084 7544
rect 1148 7480 1165 7544
rect 1229 7480 1246 7544
rect 1310 7480 1327 7544
rect 1391 7480 1408 7544
rect 1472 7480 1489 7544
rect 1553 7480 1570 7544
rect 1634 7480 1651 7544
rect 1715 7480 1732 7544
rect 1796 7480 1813 7544
rect 1877 7480 1894 7544
rect 1958 7480 1975 7544
rect 2039 7480 2056 7544
rect 2120 7480 2137 7544
rect 2201 7480 2218 7544
rect 2282 7480 2299 7544
rect 2363 7480 2380 7544
rect 2444 7480 2461 7544
rect 2525 7480 2542 7544
rect 2606 7480 2623 7544
rect 2687 7480 2704 7544
rect 2768 7480 2785 7544
rect 2849 7480 2866 7544
rect 2930 7480 2947 7544
rect 3011 7480 3028 7544
rect 3092 7480 3109 7544
rect 3173 7480 3190 7544
rect 3254 7480 3271 7544
rect 3335 7480 3352 7544
rect 3416 7480 3433 7544
rect 3497 7480 3514 7544
rect 3578 7480 3595 7544
rect 3659 7480 3676 7544
rect 3740 7480 3757 7544
rect 3821 7480 3838 7544
rect 3902 7480 3919 7544
rect 3983 7480 4000 7544
rect 4064 7480 4081 7544
rect 4145 7480 4162 7544
rect 4226 7480 4243 7544
rect 4307 7480 4324 7544
rect 4388 7480 4405 7544
rect 4469 7480 4486 7544
rect 4550 7480 4567 7544
rect 4631 7480 4648 7544
rect 4712 7480 4729 7544
rect 4793 7480 4810 7544
rect 4874 7480 4880 7544
rect 100 7456 4880 7480
rect 100 7392 106 7456
rect 170 7392 188 7456
rect 252 7392 270 7456
rect 334 7392 352 7456
rect 416 7392 434 7456
rect 498 7392 516 7456
rect 580 7392 598 7456
rect 662 7392 679 7456
rect 743 7392 760 7456
rect 824 7392 841 7456
rect 905 7392 922 7456
rect 986 7392 1003 7456
rect 1067 7392 1084 7456
rect 1148 7392 1165 7456
rect 1229 7392 1246 7456
rect 1310 7392 1327 7456
rect 1391 7392 1408 7456
rect 1472 7392 1489 7456
rect 1553 7392 1570 7456
rect 1634 7392 1651 7456
rect 1715 7392 1732 7456
rect 1796 7392 1813 7456
rect 1877 7392 1894 7456
rect 1958 7392 1975 7456
rect 2039 7392 2056 7456
rect 2120 7392 2137 7456
rect 2201 7392 2218 7456
rect 2282 7392 2299 7456
rect 2363 7392 2380 7456
rect 2444 7392 2461 7456
rect 2525 7392 2542 7456
rect 2606 7392 2623 7456
rect 2687 7392 2704 7456
rect 2768 7392 2785 7456
rect 2849 7392 2866 7456
rect 2930 7392 2947 7456
rect 3011 7392 3028 7456
rect 3092 7392 3109 7456
rect 3173 7392 3190 7456
rect 3254 7392 3271 7456
rect 3335 7392 3352 7456
rect 3416 7392 3433 7456
rect 3497 7392 3514 7456
rect 3578 7392 3595 7456
rect 3659 7392 3676 7456
rect 3740 7392 3757 7456
rect 3821 7392 3838 7456
rect 3902 7392 3919 7456
rect 3983 7392 4000 7456
rect 4064 7392 4081 7456
rect 4145 7392 4162 7456
rect 4226 7392 4243 7456
rect 4307 7392 4324 7456
rect 4388 7392 4405 7456
rect 4469 7392 4486 7456
rect 4550 7392 4567 7456
rect 4631 7392 4648 7456
rect 4712 7392 4729 7456
rect 4793 7392 4810 7456
rect 4874 7392 4880 7456
rect 100 7368 4880 7392
rect 100 7304 106 7368
rect 170 7304 188 7368
rect 252 7304 270 7368
rect 334 7304 352 7368
rect 416 7304 434 7368
rect 498 7304 516 7368
rect 580 7304 598 7368
rect 662 7304 679 7368
rect 743 7304 760 7368
rect 824 7304 841 7368
rect 905 7304 922 7368
rect 986 7304 1003 7368
rect 1067 7304 1084 7368
rect 1148 7304 1165 7368
rect 1229 7304 1246 7368
rect 1310 7304 1327 7368
rect 1391 7304 1408 7368
rect 1472 7304 1489 7368
rect 1553 7304 1570 7368
rect 1634 7304 1651 7368
rect 1715 7304 1732 7368
rect 1796 7304 1813 7368
rect 1877 7304 1894 7368
rect 1958 7304 1975 7368
rect 2039 7304 2056 7368
rect 2120 7304 2137 7368
rect 2201 7304 2218 7368
rect 2282 7304 2299 7368
rect 2363 7304 2380 7368
rect 2444 7304 2461 7368
rect 2525 7304 2542 7368
rect 2606 7304 2623 7368
rect 2687 7304 2704 7368
rect 2768 7304 2785 7368
rect 2849 7304 2866 7368
rect 2930 7304 2947 7368
rect 3011 7304 3028 7368
rect 3092 7304 3109 7368
rect 3173 7304 3190 7368
rect 3254 7304 3271 7368
rect 3335 7304 3352 7368
rect 3416 7304 3433 7368
rect 3497 7304 3514 7368
rect 3578 7304 3595 7368
rect 3659 7304 3676 7368
rect 3740 7304 3757 7368
rect 3821 7304 3838 7368
rect 3902 7304 3919 7368
rect 3983 7304 4000 7368
rect 4064 7304 4081 7368
rect 4145 7304 4162 7368
rect 4226 7304 4243 7368
rect 4307 7304 4324 7368
rect 4388 7304 4405 7368
rect 4469 7304 4486 7368
rect 4550 7304 4567 7368
rect 4631 7304 4648 7368
rect 4712 7304 4729 7368
rect 4793 7304 4810 7368
rect 4874 7304 4880 7368
rect 100 7280 4880 7304
rect 100 7216 106 7280
rect 170 7216 188 7280
rect 252 7216 270 7280
rect 334 7216 352 7280
rect 416 7216 434 7280
rect 498 7216 516 7280
rect 580 7216 598 7280
rect 662 7216 679 7280
rect 743 7216 760 7280
rect 824 7216 841 7280
rect 905 7216 922 7280
rect 986 7216 1003 7280
rect 1067 7216 1084 7280
rect 1148 7216 1165 7280
rect 1229 7216 1246 7280
rect 1310 7216 1327 7280
rect 1391 7216 1408 7280
rect 1472 7216 1489 7280
rect 1553 7216 1570 7280
rect 1634 7216 1651 7280
rect 1715 7216 1732 7280
rect 1796 7216 1813 7280
rect 1877 7216 1894 7280
rect 1958 7216 1975 7280
rect 2039 7216 2056 7280
rect 2120 7216 2137 7280
rect 2201 7216 2218 7280
rect 2282 7216 2299 7280
rect 2363 7216 2380 7280
rect 2444 7216 2461 7280
rect 2525 7216 2542 7280
rect 2606 7216 2623 7280
rect 2687 7216 2704 7280
rect 2768 7216 2785 7280
rect 2849 7216 2866 7280
rect 2930 7216 2947 7280
rect 3011 7216 3028 7280
rect 3092 7216 3109 7280
rect 3173 7216 3190 7280
rect 3254 7216 3271 7280
rect 3335 7216 3352 7280
rect 3416 7216 3433 7280
rect 3497 7216 3514 7280
rect 3578 7216 3595 7280
rect 3659 7216 3676 7280
rect 3740 7216 3757 7280
rect 3821 7216 3838 7280
rect 3902 7216 3919 7280
rect 3983 7216 4000 7280
rect 4064 7216 4081 7280
rect 4145 7216 4162 7280
rect 4226 7216 4243 7280
rect 4307 7216 4324 7280
rect 4388 7216 4405 7280
rect 4469 7216 4486 7280
rect 4550 7216 4567 7280
rect 4631 7216 4648 7280
rect 4712 7216 4729 7280
rect 4793 7216 4810 7280
rect 4874 7216 4880 7280
rect 100 7192 4880 7216
rect 100 7128 106 7192
rect 170 7128 188 7192
rect 252 7128 270 7192
rect 334 7128 352 7192
rect 416 7128 434 7192
rect 498 7128 516 7192
rect 580 7128 598 7192
rect 662 7128 679 7192
rect 743 7128 760 7192
rect 824 7128 841 7192
rect 905 7128 922 7192
rect 986 7128 1003 7192
rect 1067 7128 1084 7192
rect 1148 7128 1165 7192
rect 1229 7128 1246 7192
rect 1310 7128 1327 7192
rect 1391 7128 1408 7192
rect 1472 7128 1489 7192
rect 1553 7128 1570 7192
rect 1634 7128 1651 7192
rect 1715 7128 1732 7192
rect 1796 7128 1813 7192
rect 1877 7128 1894 7192
rect 1958 7128 1975 7192
rect 2039 7128 2056 7192
rect 2120 7128 2137 7192
rect 2201 7128 2218 7192
rect 2282 7128 2299 7192
rect 2363 7128 2380 7192
rect 2444 7128 2461 7192
rect 2525 7128 2542 7192
rect 2606 7128 2623 7192
rect 2687 7128 2704 7192
rect 2768 7128 2785 7192
rect 2849 7128 2866 7192
rect 2930 7128 2947 7192
rect 3011 7128 3028 7192
rect 3092 7128 3109 7192
rect 3173 7128 3190 7192
rect 3254 7128 3271 7192
rect 3335 7128 3352 7192
rect 3416 7128 3433 7192
rect 3497 7128 3514 7192
rect 3578 7128 3595 7192
rect 3659 7128 3676 7192
rect 3740 7128 3757 7192
rect 3821 7128 3838 7192
rect 3902 7128 3919 7192
rect 3983 7128 4000 7192
rect 4064 7128 4081 7192
rect 4145 7128 4162 7192
rect 4226 7128 4243 7192
rect 4307 7128 4324 7192
rect 4388 7128 4405 7192
rect 4469 7128 4486 7192
rect 4550 7128 4567 7192
rect 4631 7128 4648 7192
rect 4712 7128 4729 7192
rect 4793 7128 4810 7192
rect 4874 7128 4880 7192
rect 100 7104 4880 7128
rect 100 7040 106 7104
rect 170 7040 188 7104
rect 252 7040 270 7104
rect 334 7040 352 7104
rect 416 7040 434 7104
rect 498 7040 516 7104
rect 580 7040 598 7104
rect 662 7040 679 7104
rect 743 7040 760 7104
rect 824 7040 841 7104
rect 905 7040 922 7104
rect 986 7040 1003 7104
rect 1067 7040 1084 7104
rect 1148 7040 1165 7104
rect 1229 7040 1246 7104
rect 1310 7040 1327 7104
rect 1391 7040 1408 7104
rect 1472 7040 1489 7104
rect 1553 7040 1570 7104
rect 1634 7040 1651 7104
rect 1715 7040 1732 7104
rect 1796 7040 1813 7104
rect 1877 7040 1894 7104
rect 1958 7040 1975 7104
rect 2039 7040 2056 7104
rect 2120 7040 2137 7104
rect 2201 7040 2218 7104
rect 2282 7040 2299 7104
rect 2363 7040 2380 7104
rect 2444 7040 2461 7104
rect 2525 7040 2542 7104
rect 2606 7040 2623 7104
rect 2687 7040 2704 7104
rect 2768 7040 2785 7104
rect 2849 7040 2866 7104
rect 2930 7040 2947 7104
rect 3011 7040 3028 7104
rect 3092 7040 3109 7104
rect 3173 7040 3190 7104
rect 3254 7040 3271 7104
rect 3335 7040 3352 7104
rect 3416 7040 3433 7104
rect 3497 7040 3514 7104
rect 3578 7040 3595 7104
rect 3659 7040 3676 7104
rect 3740 7040 3757 7104
rect 3821 7040 3838 7104
rect 3902 7040 3919 7104
rect 3983 7040 4000 7104
rect 4064 7040 4081 7104
rect 4145 7040 4162 7104
rect 4226 7040 4243 7104
rect 4307 7040 4324 7104
rect 4388 7040 4405 7104
rect 4469 7040 4486 7104
rect 4550 7040 4567 7104
rect 4631 7040 4648 7104
rect 4712 7040 4729 7104
rect 4793 7040 4810 7104
rect 4874 7040 4880 7104
rect 100 7016 4880 7040
rect 100 6952 106 7016
rect 170 6952 188 7016
rect 252 6952 270 7016
rect 334 6952 352 7016
rect 416 6952 434 7016
rect 498 6952 516 7016
rect 580 6952 598 7016
rect 662 6952 679 7016
rect 743 6952 760 7016
rect 824 6952 841 7016
rect 905 6952 922 7016
rect 986 6952 1003 7016
rect 1067 6952 1084 7016
rect 1148 6952 1165 7016
rect 1229 6952 1246 7016
rect 1310 6952 1327 7016
rect 1391 6952 1408 7016
rect 1472 6952 1489 7016
rect 1553 6952 1570 7016
rect 1634 6952 1651 7016
rect 1715 6952 1732 7016
rect 1796 6952 1813 7016
rect 1877 6952 1894 7016
rect 1958 6952 1975 7016
rect 2039 6952 2056 7016
rect 2120 6952 2137 7016
rect 2201 6952 2218 7016
rect 2282 6952 2299 7016
rect 2363 6952 2380 7016
rect 2444 6952 2461 7016
rect 2525 6952 2542 7016
rect 2606 6952 2623 7016
rect 2687 6952 2704 7016
rect 2768 6952 2785 7016
rect 2849 6952 2866 7016
rect 2930 6952 2947 7016
rect 3011 6952 3028 7016
rect 3092 6952 3109 7016
rect 3173 6952 3190 7016
rect 3254 6952 3271 7016
rect 3335 6952 3352 7016
rect 3416 6952 3433 7016
rect 3497 6952 3514 7016
rect 3578 6952 3595 7016
rect 3659 6952 3676 7016
rect 3740 6952 3757 7016
rect 3821 6952 3838 7016
rect 3902 6952 3919 7016
rect 3983 6952 4000 7016
rect 4064 6952 4081 7016
rect 4145 6952 4162 7016
rect 4226 6952 4243 7016
rect 4307 6952 4324 7016
rect 4388 6952 4405 7016
rect 4469 6952 4486 7016
rect 4550 6952 4567 7016
rect 4631 6952 4648 7016
rect 4712 6952 4729 7016
rect 4793 6952 4810 7016
rect 4874 6952 4880 7016
rect 100 6948 4880 6952
rect 10151 7632 14931 7636
rect 10151 7568 10157 7632
rect 10221 7568 10239 7632
rect 10303 7568 10321 7632
rect 10385 7568 10403 7632
rect 10467 7568 10485 7632
rect 10549 7568 10567 7632
rect 10631 7568 10649 7632
rect 10713 7568 10730 7632
rect 10794 7568 10811 7632
rect 10875 7568 10892 7632
rect 10956 7568 10973 7632
rect 11037 7568 11054 7632
rect 11118 7568 11135 7632
rect 11199 7568 11216 7632
rect 11280 7568 11297 7632
rect 11361 7568 11378 7632
rect 11442 7568 11459 7632
rect 11523 7568 11540 7632
rect 11604 7568 11621 7632
rect 11685 7568 11702 7632
rect 11766 7568 11783 7632
rect 11847 7568 11864 7632
rect 11928 7568 11945 7632
rect 12009 7568 12026 7632
rect 12090 7568 12107 7632
rect 12171 7568 12188 7632
rect 12252 7568 12269 7632
rect 12333 7568 12350 7632
rect 12414 7568 12431 7632
rect 12495 7568 12512 7632
rect 12576 7568 12593 7632
rect 12657 7568 12674 7632
rect 12738 7568 12755 7632
rect 12819 7568 12836 7632
rect 12900 7568 12917 7632
rect 12981 7568 12998 7632
rect 13062 7568 13079 7632
rect 13143 7568 13160 7632
rect 13224 7568 13241 7632
rect 13305 7568 13322 7632
rect 13386 7568 13403 7632
rect 13467 7568 13484 7632
rect 13548 7568 13565 7632
rect 13629 7568 13646 7632
rect 13710 7568 13727 7632
rect 13791 7568 13808 7632
rect 13872 7568 13889 7632
rect 13953 7568 13970 7632
rect 14034 7568 14051 7632
rect 14115 7568 14132 7632
rect 14196 7568 14213 7632
rect 14277 7568 14294 7632
rect 14358 7568 14375 7632
rect 14439 7568 14456 7632
rect 14520 7568 14537 7632
rect 14601 7568 14618 7632
rect 14682 7568 14699 7632
rect 14763 7568 14780 7632
rect 14844 7568 14861 7632
rect 14925 7568 14931 7632
rect 10151 7544 14931 7568
rect 10151 7480 10157 7544
rect 10221 7480 10239 7544
rect 10303 7480 10321 7544
rect 10385 7480 10403 7544
rect 10467 7480 10485 7544
rect 10549 7480 10567 7544
rect 10631 7480 10649 7544
rect 10713 7480 10730 7544
rect 10794 7480 10811 7544
rect 10875 7480 10892 7544
rect 10956 7480 10973 7544
rect 11037 7480 11054 7544
rect 11118 7480 11135 7544
rect 11199 7480 11216 7544
rect 11280 7480 11297 7544
rect 11361 7480 11378 7544
rect 11442 7480 11459 7544
rect 11523 7480 11540 7544
rect 11604 7480 11621 7544
rect 11685 7480 11702 7544
rect 11766 7480 11783 7544
rect 11847 7480 11864 7544
rect 11928 7480 11945 7544
rect 12009 7480 12026 7544
rect 12090 7480 12107 7544
rect 12171 7480 12188 7544
rect 12252 7480 12269 7544
rect 12333 7480 12350 7544
rect 12414 7480 12431 7544
rect 12495 7480 12512 7544
rect 12576 7480 12593 7544
rect 12657 7480 12674 7544
rect 12738 7480 12755 7544
rect 12819 7480 12836 7544
rect 12900 7480 12917 7544
rect 12981 7480 12998 7544
rect 13062 7480 13079 7544
rect 13143 7480 13160 7544
rect 13224 7480 13241 7544
rect 13305 7480 13322 7544
rect 13386 7480 13403 7544
rect 13467 7480 13484 7544
rect 13548 7480 13565 7544
rect 13629 7480 13646 7544
rect 13710 7480 13727 7544
rect 13791 7480 13808 7544
rect 13872 7480 13889 7544
rect 13953 7480 13970 7544
rect 14034 7480 14051 7544
rect 14115 7480 14132 7544
rect 14196 7480 14213 7544
rect 14277 7480 14294 7544
rect 14358 7480 14375 7544
rect 14439 7480 14456 7544
rect 14520 7480 14537 7544
rect 14601 7480 14618 7544
rect 14682 7480 14699 7544
rect 14763 7480 14780 7544
rect 14844 7480 14861 7544
rect 14925 7480 14931 7544
rect 10151 7456 14931 7480
rect 10151 7392 10157 7456
rect 10221 7392 10239 7456
rect 10303 7392 10321 7456
rect 10385 7392 10403 7456
rect 10467 7392 10485 7456
rect 10549 7392 10567 7456
rect 10631 7392 10649 7456
rect 10713 7392 10730 7456
rect 10794 7392 10811 7456
rect 10875 7392 10892 7456
rect 10956 7392 10973 7456
rect 11037 7392 11054 7456
rect 11118 7392 11135 7456
rect 11199 7392 11216 7456
rect 11280 7392 11297 7456
rect 11361 7392 11378 7456
rect 11442 7392 11459 7456
rect 11523 7392 11540 7456
rect 11604 7392 11621 7456
rect 11685 7392 11702 7456
rect 11766 7392 11783 7456
rect 11847 7392 11864 7456
rect 11928 7392 11945 7456
rect 12009 7392 12026 7456
rect 12090 7392 12107 7456
rect 12171 7392 12188 7456
rect 12252 7392 12269 7456
rect 12333 7392 12350 7456
rect 12414 7392 12431 7456
rect 12495 7392 12512 7456
rect 12576 7392 12593 7456
rect 12657 7392 12674 7456
rect 12738 7392 12755 7456
rect 12819 7392 12836 7456
rect 12900 7392 12917 7456
rect 12981 7392 12998 7456
rect 13062 7392 13079 7456
rect 13143 7392 13160 7456
rect 13224 7392 13241 7456
rect 13305 7392 13322 7456
rect 13386 7392 13403 7456
rect 13467 7392 13484 7456
rect 13548 7392 13565 7456
rect 13629 7392 13646 7456
rect 13710 7392 13727 7456
rect 13791 7392 13808 7456
rect 13872 7392 13889 7456
rect 13953 7392 13970 7456
rect 14034 7392 14051 7456
rect 14115 7392 14132 7456
rect 14196 7392 14213 7456
rect 14277 7392 14294 7456
rect 14358 7392 14375 7456
rect 14439 7392 14456 7456
rect 14520 7392 14537 7456
rect 14601 7392 14618 7456
rect 14682 7392 14699 7456
rect 14763 7392 14780 7456
rect 14844 7392 14861 7456
rect 14925 7392 14931 7456
rect 10151 7368 14931 7392
rect 10151 7304 10157 7368
rect 10221 7304 10239 7368
rect 10303 7304 10321 7368
rect 10385 7304 10403 7368
rect 10467 7304 10485 7368
rect 10549 7304 10567 7368
rect 10631 7304 10649 7368
rect 10713 7304 10730 7368
rect 10794 7304 10811 7368
rect 10875 7304 10892 7368
rect 10956 7304 10973 7368
rect 11037 7304 11054 7368
rect 11118 7304 11135 7368
rect 11199 7304 11216 7368
rect 11280 7304 11297 7368
rect 11361 7304 11378 7368
rect 11442 7304 11459 7368
rect 11523 7304 11540 7368
rect 11604 7304 11621 7368
rect 11685 7304 11702 7368
rect 11766 7304 11783 7368
rect 11847 7304 11864 7368
rect 11928 7304 11945 7368
rect 12009 7304 12026 7368
rect 12090 7304 12107 7368
rect 12171 7304 12188 7368
rect 12252 7304 12269 7368
rect 12333 7304 12350 7368
rect 12414 7304 12431 7368
rect 12495 7304 12512 7368
rect 12576 7304 12593 7368
rect 12657 7304 12674 7368
rect 12738 7304 12755 7368
rect 12819 7304 12836 7368
rect 12900 7304 12917 7368
rect 12981 7304 12998 7368
rect 13062 7304 13079 7368
rect 13143 7304 13160 7368
rect 13224 7304 13241 7368
rect 13305 7304 13322 7368
rect 13386 7304 13403 7368
rect 13467 7304 13484 7368
rect 13548 7304 13565 7368
rect 13629 7304 13646 7368
rect 13710 7304 13727 7368
rect 13791 7304 13808 7368
rect 13872 7304 13889 7368
rect 13953 7304 13970 7368
rect 14034 7304 14051 7368
rect 14115 7304 14132 7368
rect 14196 7304 14213 7368
rect 14277 7304 14294 7368
rect 14358 7304 14375 7368
rect 14439 7304 14456 7368
rect 14520 7304 14537 7368
rect 14601 7304 14618 7368
rect 14682 7304 14699 7368
rect 14763 7304 14780 7368
rect 14844 7304 14861 7368
rect 14925 7304 14931 7368
rect 10151 7280 14931 7304
rect 10151 7216 10157 7280
rect 10221 7216 10239 7280
rect 10303 7216 10321 7280
rect 10385 7216 10403 7280
rect 10467 7216 10485 7280
rect 10549 7216 10567 7280
rect 10631 7216 10649 7280
rect 10713 7216 10730 7280
rect 10794 7216 10811 7280
rect 10875 7216 10892 7280
rect 10956 7216 10973 7280
rect 11037 7216 11054 7280
rect 11118 7216 11135 7280
rect 11199 7216 11216 7280
rect 11280 7216 11297 7280
rect 11361 7216 11378 7280
rect 11442 7216 11459 7280
rect 11523 7216 11540 7280
rect 11604 7216 11621 7280
rect 11685 7216 11702 7280
rect 11766 7216 11783 7280
rect 11847 7216 11864 7280
rect 11928 7216 11945 7280
rect 12009 7216 12026 7280
rect 12090 7216 12107 7280
rect 12171 7216 12188 7280
rect 12252 7216 12269 7280
rect 12333 7216 12350 7280
rect 12414 7216 12431 7280
rect 12495 7216 12512 7280
rect 12576 7216 12593 7280
rect 12657 7216 12674 7280
rect 12738 7216 12755 7280
rect 12819 7216 12836 7280
rect 12900 7216 12917 7280
rect 12981 7216 12998 7280
rect 13062 7216 13079 7280
rect 13143 7216 13160 7280
rect 13224 7216 13241 7280
rect 13305 7216 13322 7280
rect 13386 7216 13403 7280
rect 13467 7216 13484 7280
rect 13548 7216 13565 7280
rect 13629 7216 13646 7280
rect 13710 7216 13727 7280
rect 13791 7216 13808 7280
rect 13872 7216 13889 7280
rect 13953 7216 13970 7280
rect 14034 7216 14051 7280
rect 14115 7216 14132 7280
rect 14196 7216 14213 7280
rect 14277 7216 14294 7280
rect 14358 7216 14375 7280
rect 14439 7216 14456 7280
rect 14520 7216 14537 7280
rect 14601 7216 14618 7280
rect 14682 7216 14699 7280
rect 14763 7216 14780 7280
rect 14844 7216 14861 7280
rect 14925 7216 14931 7280
rect 10151 7192 14931 7216
rect 10151 7128 10157 7192
rect 10221 7128 10239 7192
rect 10303 7128 10321 7192
rect 10385 7128 10403 7192
rect 10467 7128 10485 7192
rect 10549 7128 10567 7192
rect 10631 7128 10649 7192
rect 10713 7128 10730 7192
rect 10794 7128 10811 7192
rect 10875 7128 10892 7192
rect 10956 7128 10973 7192
rect 11037 7128 11054 7192
rect 11118 7128 11135 7192
rect 11199 7128 11216 7192
rect 11280 7128 11297 7192
rect 11361 7128 11378 7192
rect 11442 7128 11459 7192
rect 11523 7128 11540 7192
rect 11604 7128 11621 7192
rect 11685 7128 11702 7192
rect 11766 7128 11783 7192
rect 11847 7128 11864 7192
rect 11928 7128 11945 7192
rect 12009 7128 12026 7192
rect 12090 7128 12107 7192
rect 12171 7128 12188 7192
rect 12252 7128 12269 7192
rect 12333 7128 12350 7192
rect 12414 7128 12431 7192
rect 12495 7128 12512 7192
rect 12576 7128 12593 7192
rect 12657 7128 12674 7192
rect 12738 7128 12755 7192
rect 12819 7128 12836 7192
rect 12900 7128 12917 7192
rect 12981 7128 12998 7192
rect 13062 7128 13079 7192
rect 13143 7128 13160 7192
rect 13224 7128 13241 7192
rect 13305 7128 13322 7192
rect 13386 7128 13403 7192
rect 13467 7128 13484 7192
rect 13548 7128 13565 7192
rect 13629 7128 13646 7192
rect 13710 7128 13727 7192
rect 13791 7128 13808 7192
rect 13872 7128 13889 7192
rect 13953 7128 13970 7192
rect 14034 7128 14051 7192
rect 14115 7128 14132 7192
rect 14196 7128 14213 7192
rect 14277 7128 14294 7192
rect 14358 7128 14375 7192
rect 14439 7128 14456 7192
rect 14520 7128 14537 7192
rect 14601 7128 14618 7192
rect 14682 7128 14699 7192
rect 14763 7128 14780 7192
rect 14844 7128 14861 7192
rect 14925 7128 14931 7192
rect 10151 7104 14931 7128
rect 10151 7040 10157 7104
rect 10221 7040 10239 7104
rect 10303 7040 10321 7104
rect 10385 7040 10403 7104
rect 10467 7040 10485 7104
rect 10549 7040 10567 7104
rect 10631 7040 10649 7104
rect 10713 7040 10730 7104
rect 10794 7040 10811 7104
rect 10875 7040 10892 7104
rect 10956 7040 10973 7104
rect 11037 7040 11054 7104
rect 11118 7040 11135 7104
rect 11199 7040 11216 7104
rect 11280 7040 11297 7104
rect 11361 7040 11378 7104
rect 11442 7040 11459 7104
rect 11523 7040 11540 7104
rect 11604 7040 11621 7104
rect 11685 7040 11702 7104
rect 11766 7040 11783 7104
rect 11847 7040 11864 7104
rect 11928 7040 11945 7104
rect 12009 7040 12026 7104
rect 12090 7040 12107 7104
rect 12171 7040 12188 7104
rect 12252 7040 12269 7104
rect 12333 7040 12350 7104
rect 12414 7040 12431 7104
rect 12495 7040 12512 7104
rect 12576 7040 12593 7104
rect 12657 7040 12674 7104
rect 12738 7040 12755 7104
rect 12819 7040 12836 7104
rect 12900 7040 12917 7104
rect 12981 7040 12998 7104
rect 13062 7040 13079 7104
rect 13143 7040 13160 7104
rect 13224 7040 13241 7104
rect 13305 7040 13322 7104
rect 13386 7040 13403 7104
rect 13467 7040 13484 7104
rect 13548 7040 13565 7104
rect 13629 7040 13646 7104
rect 13710 7040 13727 7104
rect 13791 7040 13808 7104
rect 13872 7040 13889 7104
rect 13953 7040 13970 7104
rect 14034 7040 14051 7104
rect 14115 7040 14132 7104
rect 14196 7040 14213 7104
rect 14277 7040 14294 7104
rect 14358 7040 14375 7104
rect 14439 7040 14456 7104
rect 14520 7040 14537 7104
rect 14601 7040 14618 7104
rect 14682 7040 14699 7104
rect 14763 7040 14780 7104
rect 14844 7040 14861 7104
rect 14925 7040 14931 7104
rect 10151 7016 14931 7040
rect 10151 6952 10157 7016
rect 10221 6952 10239 7016
rect 10303 6952 10321 7016
rect 10385 6952 10403 7016
rect 10467 6952 10485 7016
rect 10549 6952 10567 7016
rect 10631 6952 10649 7016
rect 10713 6952 10730 7016
rect 10794 6952 10811 7016
rect 10875 6952 10892 7016
rect 10956 6952 10973 7016
rect 11037 6952 11054 7016
rect 11118 6952 11135 7016
rect 11199 6952 11216 7016
rect 11280 6952 11297 7016
rect 11361 6952 11378 7016
rect 11442 6952 11459 7016
rect 11523 6952 11540 7016
rect 11604 6952 11621 7016
rect 11685 6952 11702 7016
rect 11766 6952 11783 7016
rect 11847 6952 11864 7016
rect 11928 6952 11945 7016
rect 12009 6952 12026 7016
rect 12090 6952 12107 7016
rect 12171 6952 12188 7016
rect 12252 6952 12269 7016
rect 12333 6952 12350 7016
rect 12414 6952 12431 7016
rect 12495 6952 12512 7016
rect 12576 6952 12593 7016
rect 12657 6952 12674 7016
rect 12738 6952 12755 7016
rect 12819 6952 12836 7016
rect 12900 6952 12917 7016
rect 12981 6952 12998 7016
rect 13062 6952 13079 7016
rect 13143 6952 13160 7016
rect 13224 6952 13241 7016
rect 13305 6952 13322 7016
rect 13386 6952 13403 7016
rect 13467 6952 13484 7016
rect 13548 6952 13565 7016
rect 13629 6952 13646 7016
rect 13710 6952 13727 7016
rect 13791 6952 13808 7016
rect 13872 6952 13889 7016
rect 13953 6952 13970 7016
rect 14034 6952 14051 7016
rect 14115 6952 14132 7016
rect 14196 6952 14213 7016
rect 14277 6952 14294 7016
rect 14358 6952 14375 7016
rect 14439 6952 14456 7016
rect 14520 6952 14537 7016
rect 14601 6952 14618 7016
rect 14682 6952 14699 7016
rect 14763 6952 14780 7016
rect 14844 6952 14861 7016
rect 14925 6952 14931 7016
rect 10151 6948 14931 6952
<< via3 >>
rect 106 10099 170 10163
rect 188 10099 252 10163
rect 270 10099 334 10163
rect 352 10099 416 10163
rect 434 10099 498 10163
rect 516 10099 580 10163
rect 598 10099 662 10163
rect 679 10099 743 10163
rect 760 10099 824 10163
rect 841 10099 905 10163
rect 922 10099 986 10163
rect 1003 10099 1067 10163
rect 1084 10099 1148 10163
rect 1165 10099 1229 10163
rect 1246 10099 1310 10163
rect 1327 10099 1391 10163
rect 1408 10099 1472 10163
rect 1489 10099 1553 10163
rect 1570 10099 1634 10163
rect 1651 10099 1715 10163
rect 1732 10099 1796 10163
rect 1813 10099 1877 10163
rect 1894 10099 1958 10163
rect 1975 10099 2039 10163
rect 2056 10099 2120 10163
rect 2137 10099 2201 10163
rect 2218 10099 2282 10163
rect 2299 10099 2363 10163
rect 2380 10099 2444 10163
rect 2461 10099 2525 10163
rect 2542 10099 2606 10163
rect 2623 10099 2687 10163
rect 2704 10099 2768 10163
rect 2785 10099 2849 10163
rect 2866 10099 2930 10163
rect 2947 10099 3011 10163
rect 3028 10099 3092 10163
rect 3109 10099 3173 10163
rect 3190 10099 3254 10163
rect 3271 10099 3335 10163
rect 3352 10099 3416 10163
rect 3433 10099 3497 10163
rect 3514 10099 3578 10163
rect 3595 10099 3659 10163
rect 3676 10099 3740 10163
rect 3757 10099 3821 10163
rect 3838 10099 3902 10163
rect 3919 10099 3983 10163
rect 4000 10099 4064 10163
rect 4081 10099 4145 10163
rect 4162 10099 4226 10163
rect 4243 10099 4307 10163
rect 4324 10099 4388 10163
rect 4405 10099 4469 10163
rect 4486 10099 4550 10163
rect 4567 10099 4631 10163
rect 4648 10099 4712 10163
rect 4729 10099 4793 10163
rect 4810 10099 4874 10163
rect 106 10015 170 10079
rect 188 10015 252 10079
rect 270 10015 334 10079
rect 352 10015 416 10079
rect 434 10015 498 10079
rect 516 10015 580 10079
rect 598 10015 662 10079
rect 679 10015 743 10079
rect 760 10015 824 10079
rect 841 10015 905 10079
rect 922 10015 986 10079
rect 1003 10015 1067 10079
rect 1084 10015 1148 10079
rect 1165 10015 1229 10079
rect 1246 10015 1310 10079
rect 1327 10015 1391 10079
rect 1408 10015 1472 10079
rect 1489 10015 1553 10079
rect 1570 10015 1634 10079
rect 1651 10015 1715 10079
rect 1732 10015 1796 10079
rect 1813 10015 1877 10079
rect 1894 10015 1958 10079
rect 1975 10015 2039 10079
rect 2056 10015 2120 10079
rect 2137 10015 2201 10079
rect 2218 10015 2282 10079
rect 2299 10015 2363 10079
rect 2380 10015 2444 10079
rect 2461 10015 2525 10079
rect 2542 10015 2606 10079
rect 2623 10015 2687 10079
rect 2704 10015 2768 10079
rect 2785 10015 2849 10079
rect 2866 10015 2930 10079
rect 2947 10015 3011 10079
rect 3028 10015 3092 10079
rect 3109 10015 3173 10079
rect 3190 10015 3254 10079
rect 3271 10015 3335 10079
rect 3352 10015 3416 10079
rect 3433 10015 3497 10079
rect 3514 10015 3578 10079
rect 3595 10015 3659 10079
rect 3676 10015 3740 10079
rect 3757 10015 3821 10079
rect 3838 10015 3902 10079
rect 3919 10015 3983 10079
rect 4000 10015 4064 10079
rect 4081 10015 4145 10079
rect 4162 10015 4226 10079
rect 4243 10015 4307 10079
rect 4324 10015 4388 10079
rect 4405 10015 4469 10079
rect 4486 10015 4550 10079
rect 4567 10015 4631 10079
rect 4648 10015 4712 10079
rect 4729 10015 4793 10079
rect 4810 10015 4874 10079
rect 106 9931 170 9995
rect 188 9931 252 9995
rect 270 9931 334 9995
rect 352 9931 416 9995
rect 434 9931 498 9995
rect 516 9931 580 9995
rect 598 9931 662 9995
rect 679 9931 743 9995
rect 760 9931 824 9995
rect 841 9931 905 9995
rect 922 9931 986 9995
rect 1003 9931 1067 9995
rect 1084 9931 1148 9995
rect 1165 9931 1229 9995
rect 1246 9931 1310 9995
rect 1327 9931 1391 9995
rect 1408 9931 1472 9995
rect 1489 9931 1553 9995
rect 1570 9931 1634 9995
rect 1651 9931 1715 9995
rect 1732 9931 1796 9995
rect 1813 9931 1877 9995
rect 1894 9931 1958 9995
rect 1975 9931 2039 9995
rect 2056 9931 2120 9995
rect 2137 9931 2201 9995
rect 2218 9931 2282 9995
rect 2299 9931 2363 9995
rect 2380 9931 2444 9995
rect 2461 9931 2525 9995
rect 2542 9931 2606 9995
rect 2623 9931 2687 9995
rect 2704 9931 2768 9995
rect 2785 9931 2849 9995
rect 2866 9931 2930 9995
rect 2947 9931 3011 9995
rect 3028 9931 3092 9995
rect 3109 9931 3173 9995
rect 3190 9931 3254 9995
rect 3271 9931 3335 9995
rect 3352 9931 3416 9995
rect 3433 9931 3497 9995
rect 3514 9931 3578 9995
rect 3595 9931 3659 9995
rect 3676 9931 3740 9995
rect 3757 9931 3821 9995
rect 3838 9931 3902 9995
rect 3919 9931 3983 9995
rect 4000 9931 4064 9995
rect 4081 9931 4145 9995
rect 4162 9931 4226 9995
rect 4243 9931 4307 9995
rect 4324 9931 4388 9995
rect 4405 9931 4469 9995
rect 4486 9931 4550 9995
rect 4567 9931 4631 9995
rect 4648 9931 4712 9995
rect 4729 9931 4793 9995
rect 4810 9931 4874 9995
rect 10157 10099 10221 10163
rect 10239 10099 10303 10163
rect 10321 10099 10385 10163
rect 10403 10099 10467 10163
rect 10485 10099 10549 10163
rect 10567 10099 10631 10163
rect 10649 10099 10713 10163
rect 10730 10099 10794 10163
rect 10811 10099 10875 10163
rect 10892 10099 10956 10163
rect 10973 10099 11037 10163
rect 11054 10099 11118 10163
rect 11135 10099 11199 10163
rect 11216 10099 11280 10163
rect 11297 10099 11361 10163
rect 11378 10099 11442 10163
rect 11459 10099 11523 10163
rect 11540 10099 11604 10163
rect 11621 10099 11685 10163
rect 11702 10099 11766 10163
rect 11783 10099 11847 10163
rect 11864 10099 11928 10163
rect 11945 10099 12009 10163
rect 12026 10099 12090 10163
rect 12107 10099 12171 10163
rect 12188 10099 12252 10163
rect 12269 10099 12333 10163
rect 12350 10099 12414 10163
rect 12431 10099 12495 10163
rect 12512 10099 12576 10163
rect 12593 10099 12657 10163
rect 12674 10099 12738 10163
rect 12755 10099 12819 10163
rect 12836 10099 12900 10163
rect 12917 10099 12981 10163
rect 12998 10099 13062 10163
rect 13079 10099 13143 10163
rect 13160 10099 13224 10163
rect 13241 10099 13305 10163
rect 13322 10099 13386 10163
rect 13403 10099 13467 10163
rect 13484 10099 13548 10163
rect 13565 10099 13629 10163
rect 13646 10099 13710 10163
rect 13727 10099 13791 10163
rect 13808 10099 13872 10163
rect 13889 10099 13953 10163
rect 13970 10099 14034 10163
rect 14051 10099 14115 10163
rect 14132 10099 14196 10163
rect 14213 10099 14277 10163
rect 14294 10099 14358 10163
rect 14375 10099 14439 10163
rect 14456 10099 14520 10163
rect 14537 10099 14601 10163
rect 14618 10099 14682 10163
rect 14699 10099 14763 10163
rect 14780 10099 14844 10163
rect 14861 10099 14925 10163
rect 10157 10015 10221 10079
rect 10239 10015 10303 10079
rect 10321 10015 10385 10079
rect 10403 10015 10467 10079
rect 10485 10015 10549 10079
rect 10567 10015 10631 10079
rect 10649 10015 10713 10079
rect 10730 10015 10794 10079
rect 10811 10015 10875 10079
rect 10892 10015 10956 10079
rect 10973 10015 11037 10079
rect 11054 10015 11118 10079
rect 11135 10015 11199 10079
rect 11216 10015 11280 10079
rect 11297 10015 11361 10079
rect 11378 10015 11442 10079
rect 11459 10015 11523 10079
rect 11540 10015 11604 10079
rect 11621 10015 11685 10079
rect 11702 10015 11766 10079
rect 11783 10015 11847 10079
rect 11864 10015 11928 10079
rect 11945 10015 12009 10079
rect 12026 10015 12090 10079
rect 12107 10015 12171 10079
rect 12188 10015 12252 10079
rect 12269 10015 12333 10079
rect 12350 10015 12414 10079
rect 12431 10015 12495 10079
rect 12512 10015 12576 10079
rect 12593 10015 12657 10079
rect 12674 10015 12738 10079
rect 12755 10015 12819 10079
rect 12836 10015 12900 10079
rect 12917 10015 12981 10079
rect 12998 10015 13062 10079
rect 13079 10015 13143 10079
rect 13160 10015 13224 10079
rect 13241 10015 13305 10079
rect 13322 10015 13386 10079
rect 13403 10015 13467 10079
rect 13484 10015 13548 10079
rect 13565 10015 13629 10079
rect 13646 10015 13710 10079
rect 13727 10015 13791 10079
rect 13808 10015 13872 10079
rect 13889 10015 13953 10079
rect 13970 10015 14034 10079
rect 14051 10015 14115 10079
rect 14132 10015 14196 10079
rect 14213 10015 14277 10079
rect 14294 10015 14358 10079
rect 14375 10015 14439 10079
rect 14456 10015 14520 10079
rect 14537 10015 14601 10079
rect 14618 10015 14682 10079
rect 14699 10015 14763 10079
rect 14780 10015 14844 10079
rect 14861 10015 14925 10079
rect 10157 9931 10221 9995
rect 10239 9931 10303 9995
rect 10321 9931 10385 9995
rect 10403 9931 10467 9995
rect 10485 9931 10549 9995
rect 10567 9931 10631 9995
rect 10649 9931 10713 9995
rect 10730 9931 10794 9995
rect 10811 9931 10875 9995
rect 10892 9931 10956 9995
rect 10973 9931 11037 9995
rect 11054 9931 11118 9995
rect 11135 9931 11199 9995
rect 11216 9931 11280 9995
rect 11297 9931 11361 9995
rect 11378 9931 11442 9995
rect 11459 9931 11523 9995
rect 11540 9931 11604 9995
rect 11621 9931 11685 9995
rect 11702 9931 11766 9995
rect 11783 9931 11847 9995
rect 11864 9931 11928 9995
rect 11945 9931 12009 9995
rect 12026 9931 12090 9995
rect 12107 9931 12171 9995
rect 12188 9931 12252 9995
rect 12269 9931 12333 9995
rect 12350 9931 12414 9995
rect 12431 9931 12495 9995
rect 12512 9931 12576 9995
rect 12593 9931 12657 9995
rect 12674 9931 12738 9995
rect 12755 9931 12819 9995
rect 12836 9931 12900 9995
rect 12917 9931 12981 9995
rect 12998 9931 13062 9995
rect 13079 9931 13143 9995
rect 13160 9931 13224 9995
rect 13241 9931 13305 9995
rect 13322 9931 13386 9995
rect 13403 9931 13467 9995
rect 13484 9931 13548 9995
rect 13565 9931 13629 9995
rect 13646 9931 13710 9995
rect 13727 9931 13791 9995
rect 13808 9931 13872 9995
rect 13889 9931 13953 9995
rect 13970 9931 14034 9995
rect 14051 9931 14115 9995
rect 14132 9931 14196 9995
rect 14213 9931 14277 9995
rect 14294 9931 14358 9995
rect 14375 9931 14439 9995
rect 14456 9931 14520 9995
rect 14537 9931 14601 9995
rect 14618 9931 14682 9995
rect 14699 9931 14763 9995
rect 14780 9931 14844 9995
rect 14861 9931 14925 9995
rect 106 7568 170 7632
rect 188 7568 252 7632
rect 270 7568 334 7632
rect 352 7568 416 7632
rect 434 7568 498 7632
rect 516 7568 580 7632
rect 598 7568 662 7632
rect 679 7568 743 7632
rect 760 7568 824 7632
rect 841 7568 905 7632
rect 922 7568 986 7632
rect 1003 7568 1067 7632
rect 1084 7568 1148 7632
rect 1165 7568 1229 7632
rect 1246 7568 1310 7632
rect 1327 7568 1391 7632
rect 1408 7568 1472 7632
rect 1489 7568 1553 7632
rect 1570 7568 1634 7632
rect 1651 7568 1715 7632
rect 1732 7568 1796 7632
rect 1813 7568 1877 7632
rect 1894 7568 1958 7632
rect 1975 7568 2039 7632
rect 2056 7568 2120 7632
rect 2137 7568 2201 7632
rect 2218 7568 2282 7632
rect 2299 7568 2363 7632
rect 2380 7568 2444 7632
rect 2461 7568 2525 7632
rect 2542 7568 2606 7632
rect 2623 7568 2687 7632
rect 2704 7568 2768 7632
rect 2785 7568 2849 7632
rect 2866 7568 2930 7632
rect 2947 7568 3011 7632
rect 3028 7568 3092 7632
rect 3109 7568 3173 7632
rect 3190 7568 3254 7632
rect 3271 7568 3335 7632
rect 3352 7568 3416 7632
rect 3433 7568 3497 7632
rect 3514 7568 3578 7632
rect 3595 7568 3659 7632
rect 3676 7568 3740 7632
rect 3757 7568 3821 7632
rect 3838 7568 3902 7632
rect 3919 7568 3983 7632
rect 4000 7568 4064 7632
rect 4081 7568 4145 7632
rect 4162 7568 4226 7632
rect 4243 7568 4307 7632
rect 4324 7568 4388 7632
rect 4405 7568 4469 7632
rect 4486 7568 4550 7632
rect 4567 7568 4631 7632
rect 4648 7568 4712 7632
rect 4729 7568 4793 7632
rect 4810 7568 4874 7632
rect 106 7480 170 7544
rect 188 7480 252 7544
rect 270 7480 334 7544
rect 352 7480 416 7544
rect 434 7480 498 7544
rect 516 7480 580 7544
rect 598 7480 662 7544
rect 679 7480 743 7544
rect 760 7480 824 7544
rect 841 7480 905 7544
rect 922 7480 986 7544
rect 1003 7480 1067 7544
rect 1084 7480 1148 7544
rect 1165 7480 1229 7544
rect 1246 7480 1310 7544
rect 1327 7480 1391 7544
rect 1408 7480 1472 7544
rect 1489 7480 1553 7544
rect 1570 7480 1634 7544
rect 1651 7480 1715 7544
rect 1732 7480 1796 7544
rect 1813 7480 1877 7544
rect 1894 7480 1958 7544
rect 1975 7480 2039 7544
rect 2056 7480 2120 7544
rect 2137 7480 2201 7544
rect 2218 7480 2282 7544
rect 2299 7480 2363 7544
rect 2380 7480 2444 7544
rect 2461 7480 2525 7544
rect 2542 7480 2606 7544
rect 2623 7480 2687 7544
rect 2704 7480 2768 7544
rect 2785 7480 2849 7544
rect 2866 7480 2930 7544
rect 2947 7480 3011 7544
rect 3028 7480 3092 7544
rect 3109 7480 3173 7544
rect 3190 7480 3254 7544
rect 3271 7480 3335 7544
rect 3352 7480 3416 7544
rect 3433 7480 3497 7544
rect 3514 7480 3578 7544
rect 3595 7480 3659 7544
rect 3676 7480 3740 7544
rect 3757 7480 3821 7544
rect 3838 7480 3902 7544
rect 3919 7480 3983 7544
rect 4000 7480 4064 7544
rect 4081 7480 4145 7544
rect 4162 7480 4226 7544
rect 4243 7480 4307 7544
rect 4324 7480 4388 7544
rect 4405 7480 4469 7544
rect 4486 7480 4550 7544
rect 4567 7480 4631 7544
rect 4648 7480 4712 7544
rect 4729 7480 4793 7544
rect 4810 7480 4874 7544
rect 106 7392 170 7456
rect 188 7392 252 7456
rect 270 7392 334 7456
rect 352 7392 416 7456
rect 434 7392 498 7456
rect 516 7392 580 7456
rect 598 7392 662 7456
rect 679 7392 743 7456
rect 760 7392 824 7456
rect 841 7392 905 7456
rect 922 7392 986 7456
rect 1003 7392 1067 7456
rect 1084 7392 1148 7456
rect 1165 7392 1229 7456
rect 1246 7392 1310 7456
rect 1327 7392 1391 7456
rect 1408 7392 1472 7456
rect 1489 7392 1553 7456
rect 1570 7392 1634 7456
rect 1651 7392 1715 7456
rect 1732 7392 1796 7456
rect 1813 7392 1877 7456
rect 1894 7392 1958 7456
rect 1975 7392 2039 7456
rect 2056 7392 2120 7456
rect 2137 7392 2201 7456
rect 2218 7392 2282 7456
rect 2299 7392 2363 7456
rect 2380 7392 2444 7456
rect 2461 7392 2525 7456
rect 2542 7392 2606 7456
rect 2623 7392 2687 7456
rect 2704 7392 2768 7456
rect 2785 7392 2849 7456
rect 2866 7392 2930 7456
rect 2947 7392 3011 7456
rect 3028 7392 3092 7456
rect 3109 7392 3173 7456
rect 3190 7392 3254 7456
rect 3271 7392 3335 7456
rect 3352 7392 3416 7456
rect 3433 7392 3497 7456
rect 3514 7392 3578 7456
rect 3595 7392 3659 7456
rect 3676 7392 3740 7456
rect 3757 7392 3821 7456
rect 3838 7392 3902 7456
rect 3919 7392 3983 7456
rect 4000 7392 4064 7456
rect 4081 7392 4145 7456
rect 4162 7392 4226 7456
rect 4243 7392 4307 7456
rect 4324 7392 4388 7456
rect 4405 7392 4469 7456
rect 4486 7392 4550 7456
rect 4567 7392 4631 7456
rect 4648 7392 4712 7456
rect 4729 7392 4793 7456
rect 4810 7392 4874 7456
rect 106 7304 170 7368
rect 188 7304 252 7368
rect 270 7304 334 7368
rect 352 7304 416 7368
rect 434 7304 498 7368
rect 516 7304 580 7368
rect 598 7304 662 7368
rect 679 7304 743 7368
rect 760 7304 824 7368
rect 841 7304 905 7368
rect 922 7304 986 7368
rect 1003 7304 1067 7368
rect 1084 7304 1148 7368
rect 1165 7304 1229 7368
rect 1246 7304 1310 7368
rect 1327 7304 1391 7368
rect 1408 7304 1472 7368
rect 1489 7304 1553 7368
rect 1570 7304 1634 7368
rect 1651 7304 1715 7368
rect 1732 7304 1796 7368
rect 1813 7304 1877 7368
rect 1894 7304 1958 7368
rect 1975 7304 2039 7368
rect 2056 7304 2120 7368
rect 2137 7304 2201 7368
rect 2218 7304 2282 7368
rect 2299 7304 2363 7368
rect 2380 7304 2444 7368
rect 2461 7304 2525 7368
rect 2542 7304 2606 7368
rect 2623 7304 2687 7368
rect 2704 7304 2768 7368
rect 2785 7304 2849 7368
rect 2866 7304 2930 7368
rect 2947 7304 3011 7368
rect 3028 7304 3092 7368
rect 3109 7304 3173 7368
rect 3190 7304 3254 7368
rect 3271 7304 3335 7368
rect 3352 7304 3416 7368
rect 3433 7304 3497 7368
rect 3514 7304 3578 7368
rect 3595 7304 3659 7368
rect 3676 7304 3740 7368
rect 3757 7304 3821 7368
rect 3838 7304 3902 7368
rect 3919 7304 3983 7368
rect 4000 7304 4064 7368
rect 4081 7304 4145 7368
rect 4162 7304 4226 7368
rect 4243 7304 4307 7368
rect 4324 7304 4388 7368
rect 4405 7304 4469 7368
rect 4486 7304 4550 7368
rect 4567 7304 4631 7368
rect 4648 7304 4712 7368
rect 4729 7304 4793 7368
rect 4810 7304 4874 7368
rect 106 7216 170 7280
rect 188 7216 252 7280
rect 270 7216 334 7280
rect 352 7216 416 7280
rect 434 7216 498 7280
rect 516 7216 580 7280
rect 598 7216 662 7280
rect 679 7216 743 7280
rect 760 7216 824 7280
rect 841 7216 905 7280
rect 922 7216 986 7280
rect 1003 7216 1067 7280
rect 1084 7216 1148 7280
rect 1165 7216 1229 7280
rect 1246 7216 1310 7280
rect 1327 7216 1391 7280
rect 1408 7216 1472 7280
rect 1489 7216 1553 7280
rect 1570 7216 1634 7280
rect 1651 7216 1715 7280
rect 1732 7216 1796 7280
rect 1813 7216 1877 7280
rect 1894 7216 1958 7280
rect 1975 7216 2039 7280
rect 2056 7216 2120 7280
rect 2137 7216 2201 7280
rect 2218 7216 2282 7280
rect 2299 7216 2363 7280
rect 2380 7216 2444 7280
rect 2461 7216 2525 7280
rect 2542 7216 2606 7280
rect 2623 7216 2687 7280
rect 2704 7216 2768 7280
rect 2785 7216 2849 7280
rect 2866 7216 2930 7280
rect 2947 7216 3011 7280
rect 3028 7216 3092 7280
rect 3109 7216 3173 7280
rect 3190 7216 3254 7280
rect 3271 7216 3335 7280
rect 3352 7216 3416 7280
rect 3433 7216 3497 7280
rect 3514 7216 3578 7280
rect 3595 7216 3659 7280
rect 3676 7216 3740 7280
rect 3757 7216 3821 7280
rect 3838 7216 3902 7280
rect 3919 7216 3983 7280
rect 4000 7216 4064 7280
rect 4081 7216 4145 7280
rect 4162 7216 4226 7280
rect 4243 7216 4307 7280
rect 4324 7216 4388 7280
rect 4405 7216 4469 7280
rect 4486 7216 4550 7280
rect 4567 7216 4631 7280
rect 4648 7216 4712 7280
rect 4729 7216 4793 7280
rect 4810 7216 4874 7280
rect 106 7128 170 7192
rect 188 7128 252 7192
rect 270 7128 334 7192
rect 352 7128 416 7192
rect 434 7128 498 7192
rect 516 7128 580 7192
rect 598 7128 662 7192
rect 679 7128 743 7192
rect 760 7128 824 7192
rect 841 7128 905 7192
rect 922 7128 986 7192
rect 1003 7128 1067 7192
rect 1084 7128 1148 7192
rect 1165 7128 1229 7192
rect 1246 7128 1310 7192
rect 1327 7128 1391 7192
rect 1408 7128 1472 7192
rect 1489 7128 1553 7192
rect 1570 7128 1634 7192
rect 1651 7128 1715 7192
rect 1732 7128 1796 7192
rect 1813 7128 1877 7192
rect 1894 7128 1958 7192
rect 1975 7128 2039 7192
rect 2056 7128 2120 7192
rect 2137 7128 2201 7192
rect 2218 7128 2282 7192
rect 2299 7128 2363 7192
rect 2380 7128 2444 7192
rect 2461 7128 2525 7192
rect 2542 7128 2606 7192
rect 2623 7128 2687 7192
rect 2704 7128 2768 7192
rect 2785 7128 2849 7192
rect 2866 7128 2930 7192
rect 2947 7128 3011 7192
rect 3028 7128 3092 7192
rect 3109 7128 3173 7192
rect 3190 7128 3254 7192
rect 3271 7128 3335 7192
rect 3352 7128 3416 7192
rect 3433 7128 3497 7192
rect 3514 7128 3578 7192
rect 3595 7128 3659 7192
rect 3676 7128 3740 7192
rect 3757 7128 3821 7192
rect 3838 7128 3902 7192
rect 3919 7128 3983 7192
rect 4000 7128 4064 7192
rect 4081 7128 4145 7192
rect 4162 7128 4226 7192
rect 4243 7128 4307 7192
rect 4324 7128 4388 7192
rect 4405 7128 4469 7192
rect 4486 7128 4550 7192
rect 4567 7128 4631 7192
rect 4648 7128 4712 7192
rect 4729 7128 4793 7192
rect 4810 7128 4874 7192
rect 106 7040 170 7104
rect 188 7040 252 7104
rect 270 7040 334 7104
rect 352 7040 416 7104
rect 434 7040 498 7104
rect 516 7040 580 7104
rect 598 7040 662 7104
rect 679 7040 743 7104
rect 760 7040 824 7104
rect 841 7040 905 7104
rect 922 7040 986 7104
rect 1003 7040 1067 7104
rect 1084 7040 1148 7104
rect 1165 7040 1229 7104
rect 1246 7040 1310 7104
rect 1327 7040 1391 7104
rect 1408 7040 1472 7104
rect 1489 7040 1553 7104
rect 1570 7040 1634 7104
rect 1651 7040 1715 7104
rect 1732 7040 1796 7104
rect 1813 7040 1877 7104
rect 1894 7040 1958 7104
rect 1975 7040 2039 7104
rect 2056 7040 2120 7104
rect 2137 7040 2201 7104
rect 2218 7040 2282 7104
rect 2299 7040 2363 7104
rect 2380 7040 2444 7104
rect 2461 7040 2525 7104
rect 2542 7040 2606 7104
rect 2623 7040 2687 7104
rect 2704 7040 2768 7104
rect 2785 7040 2849 7104
rect 2866 7040 2930 7104
rect 2947 7040 3011 7104
rect 3028 7040 3092 7104
rect 3109 7040 3173 7104
rect 3190 7040 3254 7104
rect 3271 7040 3335 7104
rect 3352 7040 3416 7104
rect 3433 7040 3497 7104
rect 3514 7040 3578 7104
rect 3595 7040 3659 7104
rect 3676 7040 3740 7104
rect 3757 7040 3821 7104
rect 3838 7040 3902 7104
rect 3919 7040 3983 7104
rect 4000 7040 4064 7104
rect 4081 7040 4145 7104
rect 4162 7040 4226 7104
rect 4243 7040 4307 7104
rect 4324 7040 4388 7104
rect 4405 7040 4469 7104
rect 4486 7040 4550 7104
rect 4567 7040 4631 7104
rect 4648 7040 4712 7104
rect 4729 7040 4793 7104
rect 4810 7040 4874 7104
rect 106 6952 170 7016
rect 188 6952 252 7016
rect 270 6952 334 7016
rect 352 6952 416 7016
rect 434 6952 498 7016
rect 516 6952 580 7016
rect 598 6952 662 7016
rect 679 6952 743 7016
rect 760 6952 824 7016
rect 841 6952 905 7016
rect 922 6952 986 7016
rect 1003 6952 1067 7016
rect 1084 6952 1148 7016
rect 1165 6952 1229 7016
rect 1246 6952 1310 7016
rect 1327 6952 1391 7016
rect 1408 6952 1472 7016
rect 1489 6952 1553 7016
rect 1570 6952 1634 7016
rect 1651 6952 1715 7016
rect 1732 6952 1796 7016
rect 1813 6952 1877 7016
rect 1894 6952 1958 7016
rect 1975 6952 2039 7016
rect 2056 6952 2120 7016
rect 2137 6952 2201 7016
rect 2218 6952 2282 7016
rect 2299 6952 2363 7016
rect 2380 6952 2444 7016
rect 2461 6952 2525 7016
rect 2542 6952 2606 7016
rect 2623 6952 2687 7016
rect 2704 6952 2768 7016
rect 2785 6952 2849 7016
rect 2866 6952 2930 7016
rect 2947 6952 3011 7016
rect 3028 6952 3092 7016
rect 3109 6952 3173 7016
rect 3190 6952 3254 7016
rect 3271 6952 3335 7016
rect 3352 6952 3416 7016
rect 3433 6952 3497 7016
rect 3514 6952 3578 7016
rect 3595 6952 3659 7016
rect 3676 6952 3740 7016
rect 3757 6952 3821 7016
rect 3838 6952 3902 7016
rect 3919 6952 3983 7016
rect 4000 6952 4064 7016
rect 4081 6952 4145 7016
rect 4162 6952 4226 7016
rect 4243 6952 4307 7016
rect 4324 6952 4388 7016
rect 4405 6952 4469 7016
rect 4486 6952 4550 7016
rect 4567 6952 4631 7016
rect 4648 6952 4712 7016
rect 4729 6952 4793 7016
rect 4810 6952 4874 7016
rect 10157 7568 10221 7632
rect 10239 7568 10303 7632
rect 10321 7568 10385 7632
rect 10403 7568 10467 7632
rect 10485 7568 10549 7632
rect 10567 7568 10631 7632
rect 10649 7568 10713 7632
rect 10730 7568 10794 7632
rect 10811 7568 10875 7632
rect 10892 7568 10956 7632
rect 10973 7568 11037 7632
rect 11054 7568 11118 7632
rect 11135 7568 11199 7632
rect 11216 7568 11280 7632
rect 11297 7568 11361 7632
rect 11378 7568 11442 7632
rect 11459 7568 11523 7632
rect 11540 7568 11604 7632
rect 11621 7568 11685 7632
rect 11702 7568 11766 7632
rect 11783 7568 11847 7632
rect 11864 7568 11928 7632
rect 11945 7568 12009 7632
rect 12026 7568 12090 7632
rect 12107 7568 12171 7632
rect 12188 7568 12252 7632
rect 12269 7568 12333 7632
rect 12350 7568 12414 7632
rect 12431 7568 12495 7632
rect 12512 7568 12576 7632
rect 12593 7568 12657 7632
rect 12674 7568 12738 7632
rect 12755 7568 12819 7632
rect 12836 7568 12900 7632
rect 12917 7568 12981 7632
rect 12998 7568 13062 7632
rect 13079 7568 13143 7632
rect 13160 7568 13224 7632
rect 13241 7568 13305 7632
rect 13322 7568 13386 7632
rect 13403 7568 13467 7632
rect 13484 7568 13548 7632
rect 13565 7568 13629 7632
rect 13646 7568 13710 7632
rect 13727 7568 13791 7632
rect 13808 7568 13872 7632
rect 13889 7568 13953 7632
rect 13970 7568 14034 7632
rect 14051 7568 14115 7632
rect 14132 7568 14196 7632
rect 14213 7568 14277 7632
rect 14294 7568 14358 7632
rect 14375 7568 14439 7632
rect 14456 7568 14520 7632
rect 14537 7568 14601 7632
rect 14618 7568 14682 7632
rect 14699 7568 14763 7632
rect 14780 7568 14844 7632
rect 14861 7568 14925 7632
rect 10157 7480 10221 7544
rect 10239 7480 10303 7544
rect 10321 7480 10385 7544
rect 10403 7480 10467 7544
rect 10485 7480 10549 7544
rect 10567 7480 10631 7544
rect 10649 7480 10713 7544
rect 10730 7480 10794 7544
rect 10811 7480 10875 7544
rect 10892 7480 10956 7544
rect 10973 7480 11037 7544
rect 11054 7480 11118 7544
rect 11135 7480 11199 7544
rect 11216 7480 11280 7544
rect 11297 7480 11361 7544
rect 11378 7480 11442 7544
rect 11459 7480 11523 7544
rect 11540 7480 11604 7544
rect 11621 7480 11685 7544
rect 11702 7480 11766 7544
rect 11783 7480 11847 7544
rect 11864 7480 11928 7544
rect 11945 7480 12009 7544
rect 12026 7480 12090 7544
rect 12107 7480 12171 7544
rect 12188 7480 12252 7544
rect 12269 7480 12333 7544
rect 12350 7480 12414 7544
rect 12431 7480 12495 7544
rect 12512 7480 12576 7544
rect 12593 7480 12657 7544
rect 12674 7480 12738 7544
rect 12755 7480 12819 7544
rect 12836 7480 12900 7544
rect 12917 7480 12981 7544
rect 12998 7480 13062 7544
rect 13079 7480 13143 7544
rect 13160 7480 13224 7544
rect 13241 7480 13305 7544
rect 13322 7480 13386 7544
rect 13403 7480 13467 7544
rect 13484 7480 13548 7544
rect 13565 7480 13629 7544
rect 13646 7480 13710 7544
rect 13727 7480 13791 7544
rect 13808 7480 13872 7544
rect 13889 7480 13953 7544
rect 13970 7480 14034 7544
rect 14051 7480 14115 7544
rect 14132 7480 14196 7544
rect 14213 7480 14277 7544
rect 14294 7480 14358 7544
rect 14375 7480 14439 7544
rect 14456 7480 14520 7544
rect 14537 7480 14601 7544
rect 14618 7480 14682 7544
rect 14699 7480 14763 7544
rect 14780 7480 14844 7544
rect 14861 7480 14925 7544
rect 10157 7392 10221 7456
rect 10239 7392 10303 7456
rect 10321 7392 10385 7456
rect 10403 7392 10467 7456
rect 10485 7392 10549 7456
rect 10567 7392 10631 7456
rect 10649 7392 10713 7456
rect 10730 7392 10794 7456
rect 10811 7392 10875 7456
rect 10892 7392 10956 7456
rect 10973 7392 11037 7456
rect 11054 7392 11118 7456
rect 11135 7392 11199 7456
rect 11216 7392 11280 7456
rect 11297 7392 11361 7456
rect 11378 7392 11442 7456
rect 11459 7392 11523 7456
rect 11540 7392 11604 7456
rect 11621 7392 11685 7456
rect 11702 7392 11766 7456
rect 11783 7392 11847 7456
rect 11864 7392 11928 7456
rect 11945 7392 12009 7456
rect 12026 7392 12090 7456
rect 12107 7392 12171 7456
rect 12188 7392 12252 7456
rect 12269 7392 12333 7456
rect 12350 7392 12414 7456
rect 12431 7392 12495 7456
rect 12512 7392 12576 7456
rect 12593 7392 12657 7456
rect 12674 7392 12738 7456
rect 12755 7392 12819 7456
rect 12836 7392 12900 7456
rect 12917 7392 12981 7456
rect 12998 7392 13062 7456
rect 13079 7392 13143 7456
rect 13160 7392 13224 7456
rect 13241 7392 13305 7456
rect 13322 7392 13386 7456
rect 13403 7392 13467 7456
rect 13484 7392 13548 7456
rect 13565 7392 13629 7456
rect 13646 7392 13710 7456
rect 13727 7392 13791 7456
rect 13808 7392 13872 7456
rect 13889 7392 13953 7456
rect 13970 7392 14034 7456
rect 14051 7392 14115 7456
rect 14132 7392 14196 7456
rect 14213 7392 14277 7456
rect 14294 7392 14358 7456
rect 14375 7392 14439 7456
rect 14456 7392 14520 7456
rect 14537 7392 14601 7456
rect 14618 7392 14682 7456
rect 14699 7392 14763 7456
rect 14780 7392 14844 7456
rect 14861 7392 14925 7456
rect 10157 7304 10221 7368
rect 10239 7304 10303 7368
rect 10321 7304 10385 7368
rect 10403 7304 10467 7368
rect 10485 7304 10549 7368
rect 10567 7304 10631 7368
rect 10649 7304 10713 7368
rect 10730 7304 10794 7368
rect 10811 7304 10875 7368
rect 10892 7304 10956 7368
rect 10973 7304 11037 7368
rect 11054 7304 11118 7368
rect 11135 7304 11199 7368
rect 11216 7304 11280 7368
rect 11297 7304 11361 7368
rect 11378 7304 11442 7368
rect 11459 7304 11523 7368
rect 11540 7304 11604 7368
rect 11621 7304 11685 7368
rect 11702 7304 11766 7368
rect 11783 7304 11847 7368
rect 11864 7304 11928 7368
rect 11945 7304 12009 7368
rect 12026 7304 12090 7368
rect 12107 7304 12171 7368
rect 12188 7304 12252 7368
rect 12269 7304 12333 7368
rect 12350 7304 12414 7368
rect 12431 7304 12495 7368
rect 12512 7304 12576 7368
rect 12593 7304 12657 7368
rect 12674 7304 12738 7368
rect 12755 7304 12819 7368
rect 12836 7304 12900 7368
rect 12917 7304 12981 7368
rect 12998 7304 13062 7368
rect 13079 7304 13143 7368
rect 13160 7304 13224 7368
rect 13241 7304 13305 7368
rect 13322 7304 13386 7368
rect 13403 7304 13467 7368
rect 13484 7304 13548 7368
rect 13565 7304 13629 7368
rect 13646 7304 13710 7368
rect 13727 7304 13791 7368
rect 13808 7304 13872 7368
rect 13889 7304 13953 7368
rect 13970 7304 14034 7368
rect 14051 7304 14115 7368
rect 14132 7304 14196 7368
rect 14213 7304 14277 7368
rect 14294 7304 14358 7368
rect 14375 7304 14439 7368
rect 14456 7304 14520 7368
rect 14537 7304 14601 7368
rect 14618 7304 14682 7368
rect 14699 7304 14763 7368
rect 14780 7304 14844 7368
rect 14861 7304 14925 7368
rect 10157 7216 10221 7280
rect 10239 7216 10303 7280
rect 10321 7216 10385 7280
rect 10403 7216 10467 7280
rect 10485 7216 10549 7280
rect 10567 7216 10631 7280
rect 10649 7216 10713 7280
rect 10730 7216 10794 7280
rect 10811 7216 10875 7280
rect 10892 7216 10956 7280
rect 10973 7216 11037 7280
rect 11054 7216 11118 7280
rect 11135 7216 11199 7280
rect 11216 7216 11280 7280
rect 11297 7216 11361 7280
rect 11378 7216 11442 7280
rect 11459 7216 11523 7280
rect 11540 7216 11604 7280
rect 11621 7216 11685 7280
rect 11702 7216 11766 7280
rect 11783 7216 11847 7280
rect 11864 7216 11928 7280
rect 11945 7216 12009 7280
rect 12026 7216 12090 7280
rect 12107 7216 12171 7280
rect 12188 7216 12252 7280
rect 12269 7216 12333 7280
rect 12350 7216 12414 7280
rect 12431 7216 12495 7280
rect 12512 7216 12576 7280
rect 12593 7216 12657 7280
rect 12674 7216 12738 7280
rect 12755 7216 12819 7280
rect 12836 7216 12900 7280
rect 12917 7216 12981 7280
rect 12998 7216 13062 7280
rect 13079 7216 13143 7280
rect 13160 7216 13224 7280
rect 13241 7216 13305 7280
rect 13322 7216 13386 7280
rect 13403 7216 13467 7280
rect 13484 7216 13548 7280
rect 13565 7216 13629 7280
rect 13646 7216 13710 7280
rect 13727 7216 13791 7280
rect 13808 7216 13872 7280
rect 13889 7216 13953 7280
rect 13970 7216 14034 7280
rect 14051 7216 14115 7280
rect 14132 7216 14196 7280
rect 14213 7216 14277 7280
rect 14294 7216 14358 7280
rect 14375 7216 14439 7280
rect 14456 7216 14520 7280
rect 14537 7216 14601 7280
rect 14618 7216 14682 7280
rect 14699 7216 14763 7280
rect 14780 7216 14844 7280
rect 14861 7216 14925 7280
rect 10157 7128 10221 7192
rect 10239 7128 10303 7192
rect 10321 7128 10385 7192
rect 10403 7128 10467 7192
rect 10485 7128 10549 7192
rect 10567 7128 10631 7192
rect 10649 7128 10713 7192
rect 10730 7128 10794 7192
rect 10811 7128 10875 7192
rect 10892 7128 10956 7192
rect 10973 7128 11037 7192
rect 11054 7128 11118 7192
rect 11135 7128 11199 7192
rect 11216 7128 11280 7192
rect 11297 7128 11361 7192
rect 11378 7128 11442 7192
rect 11459 7128 11523 7192
rect 11540 7128 11604 7192
rect 11621 7128 11685 7192
rect 11702 7128 11766 7192
rect 11783 7128 11847 7192
rect 11864 7128 11928 7192
rect 11945 7128 12009 7192
rect 12026 7128 12090 7192
rect 12107 7128 12171 7192
rect 12188 7128 12252 7192
rect 12269 7128 12333 7192
rect 12350 7128 12414 7192
rect 12431 7128 12495 7192
rect 12512 7128 12576 7192
rect 12593 7128 12657 7192
rect 12674 7128 12738 7192
rect 12755 7128 12819 7192
rect 12836 7128 12900 7192
rect 12917 7128 12981 7192
rect 12998 7128 13062 7192
rect 13079 7128 13143 7192
rect 13160 7128 13224 7192
rect 13241 7128 13305 7192
rect 13322 7128 13386 7192
rect 13403 7128 13467 7192
rect 13484 7128 13548 7192
rect 13565 7128 13629 7192
rect 13646 7128 13710 7192
rect 13727 7128 13791 7192
rect 13808 7128 13872 7192
rect 13889 7128 13953 7192
rect 13970 7128 14034 7192
rect 14051 7128 14115 7192
rect 14132 7128 14196 7192
rect 14213 7128 14277 7192
rect 14294 7128 14358 7192
rect 14375 7128 14439 7192
rect 14456 7128 14520 7192
rect 14537 7128 14601 7192
rect 14618 7128 14682 7192
rect 14699 7128 14763 7192
rect 14780 7128 14844 7192
rect 14861 7128 14925 7192
rect 10157 7040 10221 7104
rect 10239 7040 10303 7104
rect 10321 7040 10385 7104
rect 10403 7040 10467 7104
rect 10485 7040 10549 7104
rect 10567 7040 10631 7104
rect 10649 7040 10713 7104
rect 10730 7040 10794 7104
rect 10811 7040 10875 7104
rect 10892 7040 10956 7104
rect 10973 7040 11037 7104
rect 11054 7040 11118 7104
rect 11135 7040 11199 7104
rect 11216 7040 11280 7104
rect 11297 7040 11361 7104
rect 11378 7040 11442 7104
rect 11459 7040 11523 7104
rect 11540 7040 11604 7104
rect 11621 7040 11685 7104
rect 11702 7040 11766 7104
rect 11783 7040 11847 7104
rect 11864 7040 11928 7104
rect 11945 7040 12009 7104
rect 12026 7040 12090 7104
rect 12107 7040 12171 7104
rect 12188 7040 12252 7104
rect 12269 7040 12333 7104
rect 12350 7040 12414 7104
rect 12431 7040 12495 7104
rect 12512 7040 12576 7104
rect 12593 7040 12657 7104
rect 12674 7040 12738 7104
rect 12755 7040 12819 7104
rect 12836 7040 12900 7104
rect 12917 7040 12981 7104
rect 12998 7040 13062 7104
rect 13079 7040 13143 7104
rect 13160 7040 13224 7104
rect 13241 7040 13305 7104
rect 13322 7040 13386 7104
rect 13403 7040 13467 7104
rect 13484 7040 13548 7104
rect 13565 7040 13629 7104
rect 13646 7040 13710 7104
rect 13727 7040 13791 7104
rect 13808 7040 13872 7104
rect 13889 7040 13953 7104
rect 13970 7040 14034 7104
rect 14051 7040 14115 7104
rect 14132 7040 14196 7104
rect 14213 7040 14277 7104
rect 14294 7040 14358 7104
rect 14375 7040 14439 7104
rect 14456 7040 14520 7104
rect 14537 7040 14601 7104
rect 14618 7040 14682 7104
rect 14699 7040 14763 7104
rect 14780 7040 14844 7104
rect 14861 7040 14925 7104
rect 10157 6952 10221 7016
rect 10239 6952 10303 7016
rect 10321 6952 10385 7016
rect 10403 6952 10467 7016
rect 10485 6952 10549 7016
rect 10567 6952 10631 7016
rect 10649 6952 10713 7016
rect 10730 6952 10794 7016
rect 10811 6952 10875 7016
rect 10892 6952 10956 7016
rect 10973 6952 11037 7016
rect 11054 6952 11118 7016
rect 11135 6952 11199 7016
rect 11216 6952 11280 7016
rect 11297 6952 11361 7016
rect 11378 6952 11442 7016
rect 11459 6952 11523 7016
rect 11540 6952 11604 7016
rect 11621 6952 11685 7016
rect 11702 6952 11766 7016
rect 11783 6952 11847 7016
rect 11864 6952 11928 7016
rect 11945 6952 12009 7016
rect 12026 6952 12090 7016
rect 12107 6952 12171 7016
rect 12188 6952 12252 7016
rect 12269 6952 12333 7016
rect 12350 6952 12414 7016
rect 12431 6952 12495 7016
rect 12512 6952 12576 7016
rect 12593 6952 12657 7016
rect 12674 6952 12738 7016
rect 12755 6952 12819 7016
rect 12836 6952 12900 7016
rect 12917 6952 12981 7016
rect 12998 6952 13062 7016
rect 13079 6952 13143 7016
rect 13160 6952 13224 7016
rect 13241 6952 13305 7016
rect 13322 6952 13386 7016
rect 13403 6952 13467 7016
rect 13484 6952 13548 7016
rect 13565 6952 13629 7016
rect 13646 6952 13710 7016
rect 13727 6952 13791 7016
rect 13808 6952 13872 7016
rect 13889 6952 13953 7016
rect 13970 6952 14034 7016
rect 14051 6952 14115 7016
rect 14132 6952 14196 7016
rect 14213 6952 14277 7016
rect 14294 6952 14358 7016
rect 14375 6952 14439 7016
rect 14456 6952 14520 7016
rect 14537 6952 14601 7016
rect 14618 6952 14682 7016
rect 14699 6952 14763 7016
rect 14780 6952 14844 7016
rect 14861 6952 14925 7016
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 254 10947
rect 14746 10881 15000 10947
rect 0 10225 254 10821
rect 14746 10225 15000 10821
rect 0 10163 4875 10165
rect 0 10099 106 10163
rect 170 10099 188 10163
rect 252 10099 270 10163
rect 334 10099 352 10163
rect 416 10099 434 10163
rect 498 10099 516 10163
rect 580 10099 598 10163
rect 662 10099 679 10163
rect 743 10099 760 10163
rect 824 10099 841 10163
rect 905 10099 922 10163
rect 986 10099 1003 10163
rect 1067 10099 1084 10163
rect 1148 10099 1165 10163
rect 1229 10099 1246 10163
rect 1310 10099 1327 10163
rect 1391 10099 1408 10163
rect 1472 10099 1489 10163
rect 1553 10099 1570 10163
rect 1634 10099 1651 10163
rect 1715 10099 1732 10163
rect 1796 10099 1813 10163
rect 1877 10099 1894 10163
rect 1958 10099 1975 10163
rect 2039 10099 2056 10163
rect 2120 10099 2137 10163
rect 2201 10099 2218 10163
rect 2282 10099 2299 10163
rect 2363 10099 2380 10163
rect 2444 10099 2461 10163
rect 2525 10099 2542 10163
rect 2606 10099 2623 10163
rect 2687 10099 2704 10163
rect 2768 10099 2785 10163
rect 2849 10099 2866 10163
rect 2930 10099 2947 10163
rect 3011 10099 3028 10163
rect 3092 10099 3109 10163
rect 3173 10099 3190 10163
rect 3254 10099 3271 10163
rect 3335 10099 3352 10163
rect 3416 10099 3433 10163
rect 3497 10099 3514 10163
rect 3578 10099 3595 10163
rect 3659 10099 3676 10163
rect 3740 10099 3757 10163
rect 3821 10099 3838 10163
rect 3902 10099 3919 10163
rect 3983 10099 4000 10163
rect 4064 10099 4081 10163
rect 4145 10099 4162 10163
rect 4226 10099 4243 10163
rect 4307 10099 4324 10163
rect 4388 10099 4405 10163
rect 4469 10099 4486 10163
rect 4550 10099 4567 10163
rect 4631 10099 4648 10163
rect 4712 10099 4729 10163
rect 4793 10099 4810 10163
rect 4874 10099 4875 10163
rect 0 10079 4875 10099
rect 0 10015 106 10079
rect 170 10015 188 10079
rect 252 10015 270 10079
rect 334 10015 352 10079
rect 416 10015 434 10079
rect 498 10015 516 10079
rect 580 10015 598 10079
rect 662 10015 679 10079
rect 743 10015 760 10079
rect 824 10015 841 10079
rect 905 10015 922 10079
rect 986 10015 1003 10079
rect 1067 10015 1084 10079
rect 1148 10015 1165 10079
rect 1229 10015 1246 10079
rect 1310 10015 1327 10079
rect 1391 10015 1408 10079
rect 1472 10015 1489 10079
rect 1553 10015 1570 10079
rect 1634 10015 1651 10079
rect 1715 10015 1732 10079
rect 1796 10015 1813 10079
rect 1877 10015 1894 10079
rect 1958 10015 1975 10079
rect 2039 10015 2056 10079
rect 2120 10015 2137 10079
rect 2201 10015 2218 10079
rect 2282 10015 2299 10079
rect 2363 10015 2380 10079
rect 2444 10015 2461 10079
rect 2525 10015 2542 10079
rect 2606 10015 2623 10079
rect 2687 10015 2704 10079
rect 2768 10015 2785 10079
rect 2849 10015 2866 10079
rect 2930 10015 2947 10079
rect 3011 10015 3028 10079
rect 3092 10015 3109 10079
rect 3173 10015 3190 10079
rect 3254 10015 3271 10079
rect 3335 10015 3352 10079
rect 3416 10015 3433 10079
rect 3497 10015 3514 10079
rect 3578 10015 3595 10079
rect 3659 10015 3676 10079
rect 3740 10015 3757 10079
rect 3821 10015 3838 10079
rect 3902 10015 3919 10079
rect 3983 10015 4000 10079
rect 4064 10015 4081 10079
rect 4145 10015 4162 10079
rect 4226 10015 4243 10079
rect 4307 10015 4324 10079
rect 4388 10015 4405 10079
rect 4469 10015 4486 10079
rect 4550 10015 4567 10079
rect 4631 10015 4648 10079
rect 4712 10015 4729 10079
rect 4793 10015 4810 10079
rect 4874 10015 4875 10079
rect 0 9995 4875 10015
rect 0 9931 106 9995
rect 170 9931 188 9995
rect 252 9931 270 9995
rect 334 9931 352 9995
rect 416 9931 434 9995
rect 498 9931 516 9995
rect 580 9931 598 9995
rect 662 9931 679 9995
rect 743 9931 760 9995
rect 824 9931 841 9995
rect 905 9931 922 9995
rect 986 9931 1003 9995
rect 1067 9931 1084 9995
rect 1148 9931 1165 9995
rect 1229 9931 1246 9995
rect 1310 9931 1327 9995
rect 1391 9931 1408 9995
rect 1472 9931 1489 9995
rect 1553 9931 1570 9995
rect 1634 9931 1651 9995
rect 1715 9931 1732 9995
rect 1796 9931 1813 9995
rect 1877 9931 1894 9995
rect 1958 9931 1975 9995
rect 2039 9931 2056 9995
rect 2120 9931 2137 9995
rect 2201 9931 2218 9995
rect 2282 9931 2299 9995
rect 2363 9931 2380 9995
rect 2444 9931 2461 9995
rect 2525 9931 2542 9995
rect 2606 9931 2623 9995
rect 2687 9931 2704 9995
rect 2768 9931 2785 9995
rect 2849 9931 2866 9995
rect 2930 9931 2947 9995
rect 3011 9931 3028 9995
rect 3092 9931 3109 9995
rect 3173 9931 3190 9995
rect 3254 9931 3271 9995
rect 3335 9931 3352 9995
rect 3416 9931 3433 9995
rect 3497 9931 3514 9995
rect 3578 9931 3595 9995
rect 3659 9931 3676 9995
rect 3740 9931 3757 9995
rect 3821 9931 3838 9995
rect 3902 9931 3919 9995
rect 3983 9931 4000 9995
rect 4064 9931 4081 9995
rect 4145 9931 4162 9995
rect 4226 9931 4243 9995
rect 4307 9931 4324 9995
rect 4388 9931 4405 9995
rect 4469 9931 4486 9995
rect 4550 9931 4567 9995
rect 4631 9931 4648 9995
rect 4712 9931 4729 9995
rect 4793 9931 4810 9995
rect 4874 9931 4875 9995
rect 0 9929 4875 9931
rect 10156 10163 15000 10165
rect 10156 10099 10157 10163
rect 10221 10099 10239 10163
rect 10303 10099 10321 10163
rect 10385 10099 10403 10163
rect 10467 10099 10485 10163
rect 10549 10099 10567 10163
rect 10631 10099 10649 10163
rect 10713 10099 10730 10163
rect 10794 10099 10811 10163
rect 10875 10099 10892 10163
rect 10956 10099 10973 10163
rect 11037 10099 11054 10163
rect 11118 10099 11135 10163
rect 11199 10099 11216 10163
rect 11280 10099 11297 10163
rect 11361 10099 11378 10163
rect 11442 10099 11459 10163
rect 11523 10099 11540 10163
rect 11604 10099 11621 10163
rect 11685 10099 11702 10163
rect 11766 10099 11783 10163
rect 11847 10099 11864 10163
rect 11928 10099 11945 10163
rect 12009 10099 12026 10163
rect 12090 10099 12107 10163
rect 12171 10099 12188 10163
rect 12252 10099 12269 10163
rect 12333 10099 12350 10163
rect 12414 10099 12431 10163
rect 12495 10099 12512 10163
rect 12576 10099 12593 10163
rect 12657 10099 12674 10163
rect 12738 10099 12755 10163
rect 12819 10099 12836 10163
rect 12900 10099 12917 10163
rect 12981 10099 12998 10163
rect 13062 10099 13079 10163
rect 13143 10099 13160 10163
rect 13224 10099 13241 10163
rect 13305 10099 13322 10163
rect 13386 10099 13403 10163
rect 13467 10099 13484 10163
rect 13548 10099 13565 10163
rect 13629 10099 13646 10163
rect 13710 10099 13727 10163
rect 13791 10099 13808 10163
rect 13872 10099 13889 10163
rect 13953 10099 13970 10163
rect 14034 10099 14051 10163
rect 14115 10099 14132 10163
rect 14196 10099 14213 10163
rect 14277 10099 14294 10163
rect 14358 10099 14375 10163
rect 14439 10099 14456 10163
rect 14520 10099 14537 10163
rect 14601 10099 14618 10163
rect 14682 10099 14699 10163
rect 14763 10099 14780 10163
rect 14844 10099 14861 10163
rect 14925 10099 15000 10163
rect 10156 10079 15000 10099
rect 10156 10015 10157 10079
rect 10221 10015 10239 10079
rect 10303 10015 10321 10079
rect 10385 10015 10403 10079
rect 10467 10015 10485 10079
rect 10549 10015 10567 10079
rect 10631 10015 10649 10079
rect 10713 10015 10730 10079
rect 10794 10015 10811 10079
rect 10875 10015 10892 10079
rect 10956 10015 10973 10079
rect 11037 10015 11054 10079
rect 11118 10015 11135 10079
rect 11199 10015 11216 10079
rect 11280 10015 11297 10079
rect 11361 10015 11378 10079
rect 11442 10015 11459 10079
rect 11523 10015 11540 10079
rect 11604 10015 11621 10079
rect 11685 10015 11702 10079
rect 11766 10015 11783 10079
rect 11847 10015 11864 10079
rect 11928 10015 11945 10079
rect 12009 10015 12026 10079
rect 12090 10015 12107 10079
rect 12171 10015 12188 10079
rect 12252 10015 12269 10079
rect 12333 10015 12350 10079
rect 12414 10015 12431 10079
rect 12495 10015 12512 10079
rect 12576 10015 12593 10079
rect 12657 10015 12674 10079
rect 12738 10015 12755 10079
rect 12819 10015 12836 10079
rect 12900 10015 12917 10079
rect 12981 10015 12998 10079
rect 13062 10015 13079 10079
rect 13143 10015 13160 10079
rect 13224 10015 13241 10079
rect 13305 10015 13322 10079
rect 13386 10015 13403 10079
rect 13467 10015 13484 10079
rect 13548 10015 13565 10079
rect 13629 10015 13646 10079
rect 13710 10015 13727 10079
rect 13791 10015 13808 10079
rect 13872 10015 13889 10079
rect 13953 10015 13970 10079
rect 14034 10015 14051 10079
rect 14115 10015 14132 10079
rect 14196 10015 14213 10079
rect 14277 10015 14294 10079
rect 14358 10015 14375 10079
rect 14439 10015 14456 10079
rect 14520 10015 14537 10079
rect 14601 10015 14618 10079
rect 14682 10015 14699 10079
rect 14763 10015 14780 10079
rect 14844 10015 14861 10079
rect 14925 10015 15000 10079
rect 10156 9995 15000 10015
rect 10156 9931 10157 9995
rect 10221 9931 10239 9995
rect 10303 9931 10321 9995
rect 10385 9931 10403 9995
rect 10467 9931 10485 9995
rect 10549 9931 10567 9995
rect 10631 9931 10649 9995
rect 10713 9931 10730 9995
rect 10794 9931 10811 9995
rect 10875 9931 10892 9995
rect 10956 9931 10973 9995
rect 11037 9931 11054 9995
rect 11118 9931 11135 9995
rect 11199 9931 11216 9995
rect 11280 9931 11297 9995
rect 11361 9931 11378 9995
rect 11442 9931 11459 9995
rect 11523 9931 11540 9995
rect 11604 9931 11621 9995
rect 11685 9931 11702 9995
rect 11766 9931 11783 9995
rect 11847 9931 11864 9995
rect 11928 9931 11945 9995
rect 12009 9931 12026 9995
rect 12090 9931 12107 9995
rect 12171 9931 12188 9995
rect 12252 9931 12269 9995
rect 12333 9931 12350 9995
rect 12414 9931 12431 9995
rect 12495 9931 12512 9995
rect 12576 9931 12593 9995
rect 12657 9931 12674 9995
rect 12738 9931 12755 9995
rect 12819 9931 12836 9995
rect 12900 9931 12917 9995
rect 12981 9931 12998 9995
rect 13062 9931 13079 9995
rect 13143 9931 13160 9995
rect 13224 9931 13241 9995
rect 13305 9931 13322 9995
rect 13386 9931 13403 9995
rect 13467 9931 13484 9995
rect 13548 9931 13565 9995
rect 13629 9931 13646 9995
rect 13710 9931 13727 9995
rect 13791 9931 13808 9995
rect 13872 9931 13889 9995
rect 13953 9931 13970 9995
rect 14034 9931 14051 9995
rect 14115 9931 14132 9995
rect 14196 9931 14213 9995
rect 14277 9931 14294 9995
rect 14358 9931 14375 9995
rect 14439 9931 14456 9995
rect 14520 9931 14537 9995
rect 14601 9931 14618 9995
rect 14682 9931 14699 9995
rect 14763 9931 14780 9995
rect 14844 9931 14861 9995
rect 14925 9931 15000 9995
rect 10156 9929 15000 9931
rect 0 9273 254 9869
rect 14746 9273 15000 9869
rect 0 9147 254 9213
rect 14746 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 7632 4875 7637
rect 0 7568 106 7632
rect 170 7568 188 7632
rect 252 7568 270 7632
rect 334 7568 352 7632
rect 416 7568 434 7632
rect 498 7568 516 7632
rect 580 7568 598 7632
rect 662 7568 679 7632
rect 743 7568 760 7632
rect 824 7568 841 7632
rect 905 7568 922 7632
rect 986 7568 1003 7632
rect 1067 7568 1084 7632
rect 1148 7568 1165 7632
rect 1229 7568 1246 7632
rect 1310 7568 1327 7632
rect 1391 7568 1408 7632
rect 1472 7568 1489 7632
rect 1553 7568 1570 7632
rect 1634 7568 1651 7632
rect 1715 7568 1732 7632
rect 1796 7568 1813 7632
rect 1877 7568 1894 7632
rect 1958 7568 1975 7632
rect 2039 7568 2056 7632
rect 2120 7568 2137 7632
rect 2201 7568 2218 7632
rect 2282 7568 2299 7632
rect 2363 7568 2380 7632
rect 2444 7568 2461 7632
rect 2525 7568 2542 7632
rect 2606 7568 2623 7632
rect 2687 7568 2704 7632
rect 2768 7568 2785 7632
rect 2849 7568 2866 7632
rect 2930 7568 2947 7632
rect 3011 7568 3028 7632
rect 3092 7568 3109 7632
rect 3173 7568 3190 7632
rect 3254 7568 3271 7632
rect 3335 7568 3352 7632
rect 3416 7568 3433 7632
rect 3497 7568 3514 7632
rect 3578 7568 3595 7632
rect 3659 7568 3676 7632
rect 3740 7568 3757 7632
rect 3821 7568 3838 7632
rect 3902 7568 3919 7632
rect 3983 7568 4000 7632
rect 4064 7568 4081 7632
rect 4145 7568 4162 7632
rect 4226 7568 4243 7632
rect 4307 7568 4324 7632
rect 4388 7568 4405 7632
rect 4469 7568 4486 7632
rect 4550 7568 4567 7632
rect 4631 7568 4648 7632
rect 4712 7568 4729 7632
rect 4793 7568 4810 7632
rect 4874 7568 4875 7632
rect 0 7544 4875 7568
rect 0 7480 106 7544
rect 170 7480 188 7544
rect 252 7480 270 7544
rect 334 7480 352 7544
rect 416 7480 434 7544
rect 498 7480 516 7544
rect 580 7480 598 7544
rect 662 7480 679 7544
rect 743 7480 760 7544
rect 824 7480 841 7544
rect 905 7480 922 7544
rect 986 7480 1003 7544
rect 1067 7480 1084 7544
rect 1148 7480 1165 7544
rect 1229 7480 1246 7544
rect 1310 7480 1327 7544
rect 1391 7480 1408 7544
rect 1472 7480 1489 7544
rect 1553 7480 1570 7544
rect 1634 7480 1651 7544
rect 1715 7480 1732 7544
rect 1796 7480 1813 7544
rect 1877 7480 1894 7544
rect 1958 7480 1975 7544
rect 2039 7480 2056 7544
rect 2120 7480 2137 7544
rect 2201 7480 2218 7544
rect 2282 7480 2299 7544
rect 2363 7480 2380 7544
rect 2444 7480 2461 7544
rect 2525 7480 2542 7544
rect 2606 7480 2623 7544
rect 2687 7480 2704 7544
rect 2768 7480 2785 7544
rect 2849 7480 2866 7544
rect 2930 7480 2947 7544
rect 3011 7480 3028 7544
rect 3092 7480 3109 7544
rect 3173 7480 3190 7544
rect 3254 7480 3271 7544
rect 3335 7480 3352 7544
rect 3416 7480 3433 7544
rect 3497 7480 3514 7544
rect 3578 7480 3595 7544
rect 3659 7480 3676 7544
rect 3740 7480 3757 7544
rect 3821 7480 3838 7544
rect 3902 7480 3919 7544
rect 3983 7480 4000 7544
rect 4064 7480 4081 7544
rect 4145 7480 4162 7544
rect 4226 7480 4243 7544
rect 4307 7480 4324 7544
rect 4388 7480 4405 7544
rect 4469 7480 4486 7544
rect 4550 7480 4567 7544
rect 4631 7480 4648 7544
rect 4712 7480 4729 7544
rect 4793 7480 4810 7544
rect 4874 7480 4875 7544
rect 0 7456 4875 7480
rect 0 7392 106 7456
rect 170 7392 188 7456
rect 252 7392 270 7456
rect 334 7392 352 7456
rect 416 7392 434 7456
rect 498 7392 516 7456
rect 580 7392 598 7456
rect 662 7392 679 7456
rect 743 7392 760 7456
rect 824 7392 841 7456
rect 905 7392 922 7456
rect 986 7392 1003 7456
rect 1067 7392 1084 7456
rect 1148 7392 1165 7456
rect 1229 7392 1246 7456
rect 1310 7392 1327 7456
rect 1391 7392 1408 7456
rect 1472 7392 1489 7456
rect 1553 7392 1570 7456
rect 1634 7392 1651 7456
rect 1715 7392 1732 7456
rect 1796 7392 1813 7456
rect 1877 7392 1894 7456
rect 1958 7392 1975 7456
rect 2039 7392 2056 7456
rect 2120 7392 2137 7456
rect 2201 7392 2218 7456
rect 2282 7392 2299 7456
rect 2363 7392 2380 7456
rect 2444 7392 2461 7456
rect 2525 7392 2542 7456
rect 2606 7392 2623 7456
rect 2687 7392 2704 7456
rect 2768 7392 2785 7456
rect 2849 7392 2866 7456
rect 2930 7392 2947 7456
rect 3011 7392 3028 7456
rect 3092 7392 3109 7456
rect 3173 7392 3190 7456
rect 3254 7392 3271 7456
rect 3335 7392 3352 7456
rect 3416 7392 3433 7456
rect 3497 7392 3514 7456
rect 3578 7392 3595 7456
rect 3659 7392 3676 7456
rect 3740 7392 3757 7456
rect 3821 7392 3838 7456
rect 3902 7392 3919 7456
rect 3983 7392 4000 7456
rect 4064 7392 4081 7456
rect 4145 7392 4162 7456
rect 4226 7392 4243 7456
rect 4307 7392 4324 7456
rect 4388 7392 4405 7456
rect 4469 7392 4486 7456
rect 4550 7392 4567 7456
rect 4631 7392 4648 7456
rect 4712 7392 4729 7456
rect 4793 7392 4810 7456
rect 4874 7392 4875 7456
rect 0 7368 4875 7392
rect 0 7304 106 7368
rect 170 7304 188 7368
rect 252 7304 270 7368
rect 334 7304 352 7368
rect 416 7304 434 7368
rect 498 7304 516 7368
rect 580 7304 598 7368
rect 662 7304 679 7368
rect 743 7304 760 7368
rect 824 7304 841 7368
rect 905 7304 922 7368
rect 986 7304 1003 7368
rect 1067 7304 1084 7368
rect 1148 7304 1165 7368
rect 1229 7304 1246 7368
rect 1310 7304 1327 7368
rect 1391 7304 1408 7368
rect 1472 7304 1489 7368
rect 1553 7304 1570 7368
rect 1634 7304 1651 7368
rect 1715 7304 1732 7368
rect 1796 7304 1813 7368
rect 1877 7304 1894 7368
rect 1958 7304 1975 7368
rect 2039 7304 2056 7368
rect 2120 7304 2137 7368
rect 2201 7304 2218 7368
rect 2282 7304 2299 7368
rect 2363 7304 2380 7368
rect 2444 7304 2461 7368
rect 2525 7304 2542 7368
rect 2606 7304 2623 7368
rect 2687 7304 2704 7368
rect 2768 7304 2785 7368
rect 2849 7304 2866 7368
rect 2930 7304 2947 7368
rect 3011 7304 3028 7368
rect 3092 7304 3109 7368
rect 3173 7304 3190 7368
rect 3254 7304 3271 7368
rect 3335 7304 3352 7368
rect 3416 7304 3433 7368
rect 3497 7304 3514 7368
rect 3578 7304 3595 7368
rect 3659 7304 3676 7368
rect 3740 7304 3757 7368
rect 3821 7304 3838 7368
rect 3902 7304 3919 7368
rect 3983 7304 4000 7368
rect 4064 7304 4081 7368
rect 4145 7304 4162 7368
rect 4226 7304 4243 7368
rect 4307 7304 4324 7368
rect 4388 7304 4405 7368
rect 4469 7304 4486 7368
rect 4550 7304 4567 7368
rect 4631 7304 4648 7368
rect 4712 7304 4729 7368
rect 4793 7304 4810 7368
rect 4874 7304 4875 7368
rect 0 7280 4875 7304
rect 0 7216 106 7280
rect 170 7216 188 7280
rect 252 7216 270 7280
rect 334 7216 352 7280
rect 416 7216 434 7280
rect 498 7216 516 7280
rect 580 7216 598 7280
rect 662 7216 679 7280
rect 743 7216 760 7280
rect 824 7216 841 7280
rect 905 7216 922 7280
rect 986 7216 1003 7280
rect 1067 7216 1084 7280
rect 1148 7216 1165 7280
rect 1229 7216 1246 7280
rect 1310 7216 1327 7280
rect 1391 7216 1408 7280
rect 1472 7216 1489 7280
rect 1553 7216 1570 7280
rect 1634 7216 1651 7280
rect 1715 7216 1732 7280
rect 1796 7216 1813 7280
rect 1877 7216 1894 7280
rect 1958 7216 1975 7280
rect 2039 7216 2056 7280
rect 2120 7216 2137 7280
rect 2201 7216 2218 7280
rect 2282 7216 2299 7280
rect 2363 7216 2380 7280
rect 2444 7216 2461 7280
rect 2525 7216 2542 7280
rect 2606 7216 2623 7280
rect 2687 7216 2704 7280
rect 2768 7216 2785 7280
rect 2849 7216 2866 7280
rect 2930 7216 2947 7280
rect 3011 7216 3028 7280
rect 3092 7216 3109 7280
rect 3173 7216 3190 7280
rect 3254 7216 3271 7280
rect 3335 7216 3352 7280
rect 3416 7216 3433 7280
rect 3497 7216 3514 7280
rect 3578 7216 3595 7280
rect 3659 7216 3676 7280
rect 3740 7216 3757 7280
rect 3821 7216 3838 7280
rect 3902 7216 3919 7280
rect 3983 7216 4000 7280
rect 4064 7216 4081 7280
rect 4145 7216 4162 7280
rect 4226 7216 4243 7280
rect 4307 7216 4324 7280
rect 4388 7216 4405 7280
rect 4469 7216 4486 7280
rect 4550 7216 4567 7280
rect 4631 7216 4648 7280
rect 4712 7216 4729 7280
rect 4793 7216 4810 7280
rect 4874 7216 4875 7280
rect 0 7192 4875 7216
rect 0 7128 106 7192
rect 170 7128 188 7192
rect 252 7128 270 7192
rect 334 7128 352 7192
rect 416 7128 434 7192
rect 498 7128 516 7192
rect 580 7128 598 7192
rect 662 7128 679 7192
rect 743 7128 760 7192
rect 824 7128 841 7192
rect 905 7128 922 7192
rect 986 7128 1003 7192
rect 1067 7128 1084 7192
rect 1148 7128 1165 7192
rect 1229 7128 1246 7192
rect 1310 7128 1327 7192
rect 1391 7128 1408 7192
rect 1472 7128 1489 7192
rect 1553 7128 1570 7192
rect 1634 7128 1651 7192
rect 1715 7128 1732 7192
rect 1796 7128 1813 7192
rect 1877 7128 1894 7192
rect 1958 7128 1975 7192
rect 2039 7128 2056 7192
rect 2120 7128 2137 7192
rect 2201 7128 2218 7192
rect 2282 7128 2299 7192
rect 2363 7128 2380 7192
rect 2444 7128 2461 7192
rect 2525 7128 2542 7192
rect 2606 7128 2623 7192
rect 2687 7128 2704 7192
rect 2768 7128 2785 7192
rect 2849 7128 2866 7192
rect 2930 7128 2947 7192
rect 3011 7128 3028 7192
rect 3092 7128 3109 7192
rect 3173 7128 3190 7192
rect 3254 7128 3271 7192
rect 3335 7128 3352 7192
rect 3416 7128 3433 7192
rect 3497 7128 3514 7192
rect 3578 7128 3595 7192
rect 3659 7128 3676 7192
rect 3740 7128 3757 7192
rect 3821 7128 3838 7192
rect 3902 7128 3919 7192
rect 3983 7128 4000 7192
rect 4064 7128 4081 7192
rect 4145 7128 4162 7192
rect 4226 7128 4243 7192
rect 4307 7128 4324 7192
rect 4388 7128 4405 7192
rect 4469 7128 4486 7192
rect 4550 7128 4567 7192
rect 4631 7128 4648 7192
rect 4712 7128 4729 7192
rect 4793 7128 4810 7192
rect 4874 7128 4875 7192
rect 0 7104 4875 7128
rect 0 7040 106 7104
rect 170 7040 188 7104
rect 252 7040 270 7104
rect 334 7040 352 7104
rect 416 7040 434 7104
rect 498 7040 516 7104
rect 580 7040 598 7104
rect 662 7040 679 7104
rect 743 7040 760 7104
rect 824 7040 841 7104
rect 905 7040 922 7104
rect 986 7040 1003 7104
rect 1067 7040 1084 7104
rect 1148 7040 1165 7104
rect 1229 7040 1246 7104
rect 1310 7040 1327 7104
rect 1391 7040 1408 7104
rect 1472 7040 1489 7104
rect 1553 7040 1570 7104
rect 1634 7040 1651 7104
rect 1715 7040 1732 7104
rect 1796 7040 1813 7104
rect 1877 7040 1894 7104
rect 1958 7040 1975 7104
rect 2039 7040 2056 7104
rect 2120 7040 2137 7104
rect 2201 7040 2218 7104
rect 2282 7040 2299 7104
rect 2363 7040 2380 7104
rect 2444 7040 2461 7104
rect 2525 7040 2542 7104
rect 2606 7040 2623 7104
rect 2687 7040 2704 7104
rect 2768 7040 2785 7104
rect 2849 7040 2866 7104
rect 2930 7040 2947 7104
rect 3011 7040 3028 7104
rect 3092 7040 3109 7104
rect 3173 7040 3190 7104
rect 3254 7040 3271 7104
rect 3335 7040 3352 7104
rect 3416 7040 3433 7104
rect 3497 7040 3514 7104
rect 3578 7040 3595 7104
rect 3659 7040 3676 7104
rect 3740 7040 3757 7104
rect 3821 7040 3838 7104
rect 3902 7040 3919 7104
rect 3983 7040 4000 7104
rect 4064 7040 4081 7104
rect 4145 7040 4162 7104
rect 4226 7040 4243 7104
rect 4307 7040 4324 7104
rect 4388 7040 4405 7104
rect 4469 7040 4486 7104
rect 4550 7040 4567 7104
rect 4631 7040 4648 7104
rect 4712 7040 4729 7104
rect 4793 7040 4810 7104
rect 4874 7040 4875 7104
rect 0 7016 4875 7040
rect 0 6952 106 7016
rect 170 6952 188 7016
rect 252 6952 270 7016
rect 334 6952 352 7016
rect 416 6952 434 7016
rect 498 6952 516 7016
rect 580 6952 598 7016
rect 662 6952 679 7016
rect 743 6952 760 7016
rect 824 6952 841 7016
rect 905 6952 922 7016
rect 986 6952 1003 7016
rect 1067 6952 1084 7016
rect 1148 6952 1165 7016
rect 1229 6952 1246 7016
rect 1310 6952 1327 7016
rect 1391 6952 1408 7016
rect 1472 6952 1489 7016
rect 1553 6952 1570 7016
rect 1634 6952 1651 7016
rect 1715 6952 1732 7016
rect 1796 6952 1813 7016
rect 1877 6952 1894 7016
rect 1958 6952 1975 7016
rect 2039 6952 2056 7016
rect 2120 6952 2137 7016
rect 2201 6952 2218 7016
rect 2282 6952 2299 7016
rect 2363 6952 2380 7016
rect 2444 6952 2461 7016
rect 2525 6952 2542 7016
rect 2606 6952 2623 7016
rect 2687 6952 2704 7016
rect 2768 6952 2785 7016
rect 2849 6952 2866 7016
rect 2930 6952 2947 7016
rect 3011 6952 3028 7016
rect 3092 6952 3109 7016
rect 3173 6952 3190 7016
rect 3254 6952 3271 7016
rect 3335 6952 3352 7016
rect 3416 6952 3433 7016
rect 3497 6952 3514 7016
rect 3578 6952 3595 7016
rect 3659 6952 3676 7016
rect 3740 6952 3757 7016
rect 3821 6952 3838 7016
rect 3902 6952 3919 7016
rect 3983 6952 4000 7016
rect 4064 6952 4081 7016
rect 4145 6952 4162 7016
rect 4226 6952 4243 7016
rect 4307 6952 4324 7016
rect 4388 6952 4405 7016
rect 4469 6952 4486 7016
rect 4550 6952 4567 7016
rect 4631 6952 4648 7016
rect 4712 6952 4729 7016
rect 4793 6952 4810 7016
rect 4874 6952 4875 7016
rect 0 6947 4875 6952
rect 10156 7632 15000 7637
rect 10156 7568 10157 7632
rect 10221 7568 10239 7632
rect 10303 7568 10321 7632
rect 10385 7568 10403 7632
rect 10467 7568 10485 7632
rect 10549 7568 10567 7632
rect 10631 7568 10649 7632
rect 10713 7568 10730 7632
rect 10794 7568 10811 7632
rect 10875 7568 10892 7632
rect 10956 7568 10973 7632
rect 11037 7568 11054 7632
rect 11118 7568 11135 7632
rect 11199 7568 11216 7632
rect 11280 7568 11297 7632
rect 11361 7568 11378 7632
rect 11442 7568 11459 7632
rect 11523 7568 11540 7632
rect 11604 7568 11621 7632
rect 11685 7568 11702 7632
rect 11766 7568 11783 7632
rect 11847 7568 11864 7632
rect 11928 7568 11945 7632
rect 12009 7568 12026 7632
rect 12090 7568 12107 7632
rect 12171 7568 12188 7632
rect 12252 7568 12269 7632
rect 12333 7568 12350 7632
rect 12414 7568 12431 7632
rect 12495 7568 12512 7632
rect 12576 7568 12593 7632
rect 12657 7568 12674 7632
rect 12738 7568 12755 7632
rect 12819 7568 12836 7632
rect 12900 7568 12917 7632
rect 12981 7568 12998 7632
rect 13062 7568 13079 7632
rect 13143 7568 13160 7632
rect 13224 7568 13241 7632
rect 13305 7568 13322 7632
rect 13386 7568 13403 7632
rect 13467 7568 13484 7632
rect 13548 7568 13565 7632
rect 13629 7568 13646 7632
rect 13710 7568 13727 7632
rect 13791 7568 13808 7632
rect 13872 7568 13889 7632
rect 13953 7568 13970 7632
rect 14034 7568 14051 7632
rect 14115 7568 14132 7632
rect 14196 7568 14213 7632
rect 14277 7568 14294 7632
rect 14358 7568 14375 7632
rect 14439 7568 14456 7632
rect 14520 7568 14537 7632
rect 14601 7568 14618 7632
rect 14682 7568 14699 7632
rect 14763 7568 14780 7632
rect 14844 7568 14861 7632
rect 14925 7568 15000 7632
rect 10156 7544 15000 7568
rect 10156 7480 10157 7544
rect 10221 7480 10239 7544
rect 10303 7480 10321 7544
rect 10385 7480 10403 7544
rect 10467 7480 10485 7544
rect 10549 7480 10567 7544
rect 10631 7480 10649 7544
rect 10713 7480 10730 7544
rect 10794 7480 10811 7544
rect 10875 7480 10892 7544
rect 10956 7480 10973 7544
rect 11037 7480 11054 7544
rect 11118 7480 11135 7544
rect 11199 7480 11216 7544
rect 11280 7480 11297 7544
rect 11361 7480 11378 7544
rect 11442 7480 11459 7544
rect 11523 7480 11540 7544
rect 11604 7480 11621 7544
rect 11685 7480 11702 7544
rect 11766 7480 11783 7544
rect 11847 7480 11864 7544
rect 11928 7480 11945 7544
rect 12009 7480 12026 7544
rect 12090 7480 12107 7544
rect 12171 7480 12188 7544
rect 12252 7480 12269 7544
rect 12333 7480 12350 7544
rect 12414 7480 12431 7544
rect 12495 7480 12512 7544
rect 12576 7480 12593 7544
rect 12657 7480 12674 7544
rect 12738 7480 12755 7544
rect 12819 7480 12836 7544
rect 12900 7480 12917 7544
rect 12981 7480 12998 7544
rect 13062 7480 13079 7544
rect 13143 7480 13160 7544
rect 13224 7480 13241 7544
rect 13305 7480 13322 7544
rect 13386 7480 13403 7544
rect 13467 7480 13484 7544
rect 13548 7480 13565 7544
rect 13629 7480 13646 7544
rect 13710 7480 13727 7544
rect 13791 7480 13808 7544
rect 13872 7480 13889 7544
rect 13953 7480 13970 7544
rect 14034 7480 14051 7544
rect 14115 7480 14132 7544
rect 14196 7480 14213 7544
rect 14277 7480 14294 7544
rect 14358 7480 14375 7544
rect 14439 7480 14456 7544
rect 14520 7480 14537 7544
rect 14601 7480 14618 7544
rect 14682 7480 14699 7544
rect 14763 7480 14780 7544
rect 14844 7480 14861 7544
rect 14925 7480 15000 7544
rect 10156 7456 15000 7480
rect 10156 7392 10157 7456
rect 10221 7392 10239 7456
rect 10303 7392 10321 7456
rect 10385 7392 10403 7456
rect 10467 7392 10485 7456
rect 10549 7392 10567 7456
rect 10631 7392 10649 7456
rect 10713 7392 10730 7456
rect 10794 7392 10811 7456
rect 10875 7392 10892 7456
rect 10956 7392 10973 7456
rect 11037 7392 11054 7456
rect 11118 7392 11135 7456
rect 11199 7392 11216 7456
rect 11280 7392 11297 7456
rect 11361 7392 11378 7456
rect 11442 7392 11459 7456
rect 11523 7392 11540 7456
rect 11604 7392 11621 7456
rect 11685 7392 11702 7456
rect 11766 7392 11783 7456
rect 11847 7392 11864 7456
rect 11928 7392 11945 7456
rect 12009 7392 12026 7456
rect 12090 7392 12107 7456
rect 12171 7392 12188 7456
rect 12252 7392 12269 7456
rect 12333 7392 12350 7456
rect 12414 7392 12431 7456
rect 12495 7392 12512 7456
rect 12576 7392 12593 7456
rect 12657 7392 12674 7456
rect 12738 7392 12755 7456
rect 12819 7392 12836 7456
rect 12900 7392 12917 7456
rect 12981 7392 12998 7456
rect 13062 7392 13079 7456
rect 13143 7392 13160 7456
rect 13224 7392 13241 7456
rect 13305 7392 13322 7456
rect 13386 7392 13403 7456
rect 13467 7392 13484 7456
rect 13548 7392 13565 7456
rect 13629 7392 13646 7456
rect 13710 7392 13727 7456
rect 13791 7392 13808 7456
rect 13872 7392 13889 7456
rect 13953 7392 13970 7456
rect 14034 7392 14051 7456
rect 14115 7392 14132 7456
rect 14196 7392 14213 7456
rect 14277 7392 14294 7456
rect 14358 7392 14375 7456
rect 14439 7392 14456 7456
rect 14520 7392 14537 7456
rect 14601 7392 14618 7456
rect 14682 7392 14699 7456
rect 14763 7392 14780 7456
rect 14844 7392 14861 7456
rect 14925 7392 15000 7456
rect 10156 7368 15000 7392
rect 10156 7304 10157 7368
rect 10221 7304 10239 7368
rect 10303 7304 10321 7368
rect 10385 7304 10403 7368
rect 10467 7304 10485 7368
rect 10549 7304 10567 7368
rect 10631 7304 10649 7368
rect 10713 7304 10730 7368
rect 10794 7304 10811 7368
rect 10875 7304 10892 7368
rect 10956 7304 10973 7368
rect 11037 7304 11054 7368
rect 11118 7304 11135 7368
rect 11199 7304 11216 7368
rect 11280 7304 11297 7368
rect 11361 7304 11378 7368
rect 11442 7304 11459 7368
rect 11523 7304 11540 7368
rect 11604 7304 11621 7368
rect 11685 7304 11702 7368
rect 11766 7304 11783 7368
rect 11847 7304 11864 7368
rect 11928 7304 11945 7368
rect 12009 7304 12026 7368
rect 12090 7304 12107 7368
rect 12171 7304 12188 7368
rect 12252 7304 12269 7368
rect 12333 7304 12350 7368
rect 12414 7304 12431 7368
rect 12495 7304 12512 7368
rect 12576 7304 12593 7368
rect 12657 7304 12674 7368
rect 12738 7304 12755 7368
rect 12819 7304 12836 7368
rect 12900 7304 12917 7368
rect 12981 7304 12998 7368
rect 13062 7304 13079 7368
rect 13143 7304 13160 7368
rect 13224 7304 13241 7368
rect 13305 7304 13322 7368
rect 13386 7304 13403 7368
rect 13467 7304 13484 7368
rect 13548 7304 13565 7368
rect 13629 7304 13646 7368
rect 13710 7304 13727 7368
rect 13791 7304 13808 7368
rect 13872 7304 13889 7368
rect 13953 7304 13970 7368
rect 14034 7304 14051 7368
rect 14115 7304 14132 7368
rect 14196 7304 14213 7368
rect 14277 7304 14294 7368
rect 14358 7304 14375 7368
rect 14439 7304 14456 7368
rect 14520 7304 14537 7368
rect 14601 7304 14618 7368
rect 14682 7304 14699 7368
rect 14763 7304 14780 7368
rect 14844 7304 14861 7368
rect 14925 7304 15000 7368
rect 10156 7280 15000 7304
rect 10156 7216 10157 7280
rect 10221 7216 10239 7280
rect 10303 7216 10321 7280
rect 10385 7216 10403 7280
rect 10467 7216 10485 7280
rect 10549 7216 10567 7280
rect 10631 7216 10649 7280
rect 10713 7216 10730 7280
rect 10794 7216 10811 7280
rect 10875 7216 10892 7280
rect 10956 7216 10973 7280
rect 11037 7216 11054 7280
rect 11118 7216 11135 7280
rect 11199 7216 11216 7280
rect 11280 7216 11297 7280
rect 11361 7216 11378 7280
rect 11442 7216 11459 7280
rect 11523 7216 11540 7280
rect 11604 7216 11621 7280
rect 11685 7216 11702 7280
rect 11766 7216 11783 7280
rect 11847 7216 11864 7280
rect 11928 7216 11945 7280
rect 12009 7216 12026 7280
rect 12090 7216 12107 7280
rect 12171 7216 12188 7280
rect 12252 7216 12269 7280
rect 12333 7216 12350 7280
rect 12414 7216 12431 7280
rect 12495 7216 12512 7280
rect 12576 7216 12593 7280
rect 12657 7216 12674 7280
rect 12738 7216 12755 7280
rect 12819 7216 12836 7280
rect 12900 7216 12917 7280
rect 12981 7216 12998 7280
rect 13062 7216 13079 7280
rect 13143 7216 13160 7280
rect 13224 7216 13241 7280
rect 13305 7216 13322 7280
rect 13386 7216 13403 7280
rect 13467 7216 13484 7280
rect 13548 7216 13565 7280
rect 13629 7216 13646 7280
rect 13710 7216 13727 7280
rect 13791 7216 13808 7280
rect 13872 7216 13889 7280
rect 13953 7216 13970 7280
rect 14034 7216 14051 7280
rect 14115 7216 14132 7280
rect 14196 7216 14213 7280
rect 14277 7216 14294 7280
rect 14358 7216 14375 7280
rect 14439 7216 14456 7280
rect 14520 7216 14537 7280
rect 14601 7216 14618 7280
rect 14682 7216 14699 7280
rect 14763 7216 14780 7280
rect 14844 7216 14861 7280
rect 14925 7216 15000 7280
rect 10156 7192 15000 7216
rect 10156 7128 10157 7192
rect 10221 7128 10239 7192
rect 10303 7128 10321 7192
rect 10385 7128 10403 7192
rect 10467 7128 10485 7192
rect 10549 7128 10567 7192
rect 10631 7128 10649 7192
rect 10713 7128 10730 7192
rect 10794 7128 10811 7192
rect 10875 7128 10892 7192
rect 10956 7128 10973 7192
rect 11037 7128 11054 7192
rect 11118 7128 11135 7192
rect 11199 7128 11216 7192
rect 11280 7128 11297 7192
rect 11361 7128 11378 7192
rect 11442 7128 11459 7192
rect 11523 7128 11540 7192
rect 11604 7128 11621 7192
rect 11685 7128 11702 7192
rect 11766 7128 11783 7192
rect 11847 7128 11864 7192
rect 11928 7128 11945 7192
rect 12009 7128 12026 7192
rect 12090 7128 12107 7192
rect 12171 7128 12188 7192
rect 12252 7128 12269 7192
rect 12333 7128 12350 7192
rect 12414 7128 12431 7192
rect 12495 7128 12512 7192
rect 12576 7128 12593 7192
rect 12657 7128 12674 7192
rect 12738 7128 12755 7192
rect 12819 7128 12836 7192
rect 12900 7128 12917 7192
rect 12981 7128 12998 7192
rect 13062 7128 13079 7192
rect 13143 7128 13160 7192
rect 13224 7128 13241 7192
rect 13305 7128 13322 7192
rect 13386 7128 13403 7192
rect 13467 7128 13484 7192
rect 13548 7128 13565 7192
rect 13629 7128 13646 7192
rect 13710 7128 13727 7192
rect 13791 7128 13808 7192
rect 13872 7128 13889 7192
rect 13953 7128 13970 7192
rect 14034 7128 14051 7192
rect 14115 7128 14132 7192
rect 14196 7128 14213 7192
rect 14277 7128 14294 7192
rect 14358 7128 14375 7192
rect 14439 7128 14456 7192
rect 14520 7128 14537 7192
rect 14601 7128 14618 7192
rect 14682 7128 14699 7192
rect 14763 7128 14780 7192
rect 14844 7128 14861 7192
rect 14925 7128 15000 7192
rect 10156 7104 15000 7128
rect 10156 7040 10157 7104
rect 10221 7040 10239 7104
rect 10303 7040 10321 7104
rect 10385 7040 10403 7104
rect 10467 7040 10485 7104
rect 10549 7040 10567 7104
rect 10631 7040 10649 7104
rect 10713 7040 10730 7104
rect 10794 7040 10811 7104
rect 10875 7040 10892 7104
rect 10956 7040 10973 7104
rect 11037 7040 11054 7104
rect 11118 7040 11135 7104
rect 11199 7040 11216 7104
rect 11280 7040 11297 7104
rect 11361 7040 11378 7104
rect 11442 7040 11459 7104
rect 11523 7040 11540 7104
rect 11604 7040 11621 7104
rect 11685 7040 11702 7104
rect 11766 7040 11783 7104
rect 11847 7040 11864 7104
rect 11928 7040 11945 7104
rect 12009 7040 12026 7104
rect 12090 7040 12107 7104
rect 12171 7040 12188 7104
rect 12252 7040 12269 7104
rect 12333 7040 12350 7104
rect 12414 7040 12431 7104
rect 12495 7040 12512 7104
rect 12576 7040 12593 7104
rect 12657 7040 12674 7104
rect 12738 7040 12755 7104
rect 12819 7040 12836 7104
rect 12900 7040 12917 7104
rect 12981 7040 12998 7104
rect 13062 7040 13079 7104
rect 13143 7040 13160 7104
rect 13224 7040 13241 7104
rect 13305 7040 13322 7104
rect 13386 7040 13403 7104
rect 13467 7040 13484 7104
rect 13548 7040 13565 7104
rect 13629 7040 13646 7104
rect 13710 7040 13727 7104
rect 13791 7040 13808 7104
rect 13872 7040 13889 7104
rect 13953 7040 13970 7104
rect 14034 7040 14051 7104
rect 14115 7040 14132 7104
rect 14196 7040 14213 7104
rect 14277 7040 14294 7104
rect 14358 7040 14375 7104
rect 14439 7040 14456 7104
rect 14520 7040 14537 7104
rect 14601 7040 14618 7104
rect 14682 7040 14699 7104
rect 14763 7040 14780 7104
rect 14844 7040 14861 7104
rect 14925 7040 15000 7104
rect 10156 7016 15000 7040
rect 10156 6952 10157 7016
rect 10221 6952 10239 7016
rect 10303 6952 10321 7016
rect 10385 6952 10403 7016
rect 10467 6952 10485 7016
rect 10549 6952 10567 7016
rect 10631 6952 10649 7016
rect 10713 6952 10730 7016
rect 10794 6952 10811 7016
rect 10875 6952 10892 7016
rect 10956 6952 10973 7016
rect 11037 6952 11054 7016
rect 11118 6952 11135 7016
rect 11199 6952 11216 7016
rect 11280 6952 11297 7016
rect 11361 6952 11378 7016
rect 11442 6952 11459 7016
rect 11523 6952 11540 7016
rect 11604 6952 11621 7016
rect 11685 6952 11702 7016
rect 11766 6952 11783 7016
rect 11847 6952 11864 7016
rect 11928 6952 11945 7016
rect 12009 6952 12026 7016
rect 12090 6952 12107 7016
rect 12171 6952 12188 7016
rect 12252 6952 12269 7016
rect 12333 6952 12350 7016
rect 12414 6952 12431 7016
rect 12495 6952 12512 7016
rect 12576 6952 12593 7016
rect 12657 6952 12674 7016
rect 12738 6952 12755 7016
rect 12819 6952 12836 7016
rect 12900 6952 12917 7016
rect 12981 6952 12998 7016
rect 13062 6952 13079 7016
rect 13143 6952 13160 7016
rect 13224 6952 13241 7016
rect 13305 6952 13322 7016
rect 13386 6952 13403 7016
rect 13467 6952 13484 7016
rect 13548 6952 13565 7016
rect 13629 6952 13646 7016
rect 13710 6952 13727 7016
rect 13791 6952 13808 7016
rect 13872 6952 13889 7016
rect 13953 6952 13970 7016
rect 14034 6952 14051 7016
rect 14115 6952 14132 7016
rect 14196 6952 14213 7016
rect 14277 6952 14294 7016
rect 14358 6952 14375 7016
rect 14439 6952 14456 7016
rect 14520 6952 14537 7016
rect 14601 6952 14618 7016
rect 14682 6952 14699 7016
rect 14763 6952 14780 7016
rect 14844 6952 14861 7016
rect 14925 6952 15000 7016
rect 10156 6947 15000 6952
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 14746 13607 15000 18597
rect 0 12437 254 13287
rect 14746 12437 15000 13287
rect 0 11267 254 12117
rect 14746 11267 15000 12117
rect 0 9147 254 10947
rect 14746 9147 15000 10947
rect 0 7937 254 8827
rect 14746 7937 15000 8827
rect 0 6968 254 7617
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 14746 5997 15000 6647
rect 0 4787 254 5677
rect 14746 4787 15000 5677
rect 0 3577 254 4467
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 14746 1397 15000 2287
rect 0 27 254 1077
rect 14746 27 15000 1077
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1627201311
transform 1 0 0 0 1 149
box 0 -142 15000 39451
<< labels >>
flabel metal5 s 0 12437 254 13287 3 FreeSans 520 0 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal5 s 14746 9147 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal5 s 14746 6968 15000 7617 3 FreeSans 520 180 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal5 s 0 27 254 1077 3 FreeSans 520 0 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal5 s 0 9147 254 10947 3 FreeSans 520 0 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal5 s 0 6968 254 7617 3 FreeSans 520 0 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal5 s 14746 7937 15000 8827 3 FreeSans 520 180 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal5 s 0 7937 254 8827 3 FreeSans 520 0 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal5 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 14746 4787 15000 5677 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 0 4787 254 5677 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal5 s 14746 11267 15000 12117 3 FreeSans 520 180 0 0 VSSIO_Q
port 6 nsew ground bidirectional
flabel metal5 s 0 11267 254 12117 3 FreeSans 520 0 0 0 VSSIO_Q
port 6 nsew ground bidirectional
flabel metal5 s 14746 1397 15000 2287 3 FreeSans 520 180 0 0 VCCD
port 7 nsew power bidirectional
flabel metal5 s 0 1397 254 2287 3 FreeSans 520 0 0 0 VCCD
port 7 nsew power bidirectional
flabel metal5 s 14746 27 15000 1077 3 FreeSans 520 180 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal5 s 14807 2607 15000 3257 3 FreeSans 520 180 0 0 VDDA
port 8 nsew power bidirectional
flabel metal5 s 0 2607 193 3257 3 FreeSans 520 0 0 0 VDDA
port 8 nsew power bidirectional
flabel metal5 s 14746 13607 15000 18597 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal5 s 14746 3577 15000 4467 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal5 s 0 13607 254 18597 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal5 s 0 3577 254 4467 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal5 s 14746 5997 15000 6647 3 FreeSans 520 180 0 0 VSWITCH
port 10 nsew power bidirectional
flabel metal5 s 14746 12437 15000 13287 3 FreeSans 520 180 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal5 s 0 5997 254 6647 3 FreeSans 520 0 0 0 VSWITCH
port 10 nsew power bidirectional
flabel metal4 s 14746 10225 15000 10821 3 FreeSans 520 180 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 0 1377 254 2307 3 FreeSans 520 0 0 0 VCCD
port 7 nsew power bidirectional
flabel metal4 s 14746 6947 15000 7637 3 FreeSans 520 180 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal4 s 14746 9147 15000 9213 3 FreeSans 520 180 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal4 s 14746 10881 15000 10947 3 FreeSans 520 180 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal4 s 14746 9929 15000 10165 3 FreeSans 520 180 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal4 s 0 9147 254 9213 3 FreeSans 520 0 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal4 s 14807 2587 15000 3277 3 FreeSans 520 180 0 0 VDDA
port 8 nsew power bidirectional
flabel metal4 s 0 10881 254 10947 3 FreeSans 520 0 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal4 s 0 9929 254 10165 3 FreeSans 520 0 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal4 s 0 6947 254 7637 3 FreeSans 520 0 0 0 VSSA
port 2 nsew ground bidirectional
flabel metal4 s 14746 7917 15000 8847 3 FreeSans 520 180 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal4 s 0 7917 254 8847 3 FreeSans 520 0 0 0 VSSD
port 4 nsew ground bidirectional
flabel metal4 s 14746 34757 15000 39600 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 14746 4767 15000 5697 3 FreeSans 520 180 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 0 34757 254 39600 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 0 4767 254 5697 3 FreeSans 520 0 0 0 VSSIO
port 5 nsew ground bidirectional
flabel metal4 s 14746 11247 15000 12137 3 FreeSans 520 180 0 0 VSSIO_Q
port 6 nsew ground bidirectional
flabel metal4 s 0 11247 254 12137 3 FreeSans 520 0 0 0 VSSIO_Q
port 6 nsew ground bidirectional
flabel metal4 s 0 10225 254 10821 3 FreeSans 520 0 0 0 AMUXBUS_A
port 11 nsew signal bidirectional
flabel metal4 s 14746 9273 15000 9869 3 FreeSans 520 180 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
flabel metal4 s 0 9273 254 9869 3 FreeSans 520 0 0 0 AMUXBUS_B
port 12 nsew signal bidirectional
flabel metal4 s 14746 1377 15000 2307 3 FreeSans 520 180 0 0 VCCD
port 7 nsew power bidirectional
flabel metal4 s 14746 7 15000 1097 3 FreeSans 520 180 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal4 s 0 7 254 1097 3 FreeSans 520 0 0 0 VCCHIB
port 3 nsew power bidirectional
flabel metal4 s 0 2587 193 3277 3 FreeSans 520 0 0 0 VDDA
port 8 nsew power bidirectional
flabel metal4 s 14746 3557 15000 4487 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal4 s 14746 13607 15000 18600 3 FreeSans 520 180 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal4 s 0 3557 254 4487 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal4 s 0 13607 254 18600 3 FreeSans 520 0 0 0 VDDIO
port 9 nsew power bidirectional
flabel metal4 s 14746 12417 15000 13307 3 FreeSans 520 180 0 0 VDDIO_Q
port 1 nsew power bidirectional
flabel metal4 s 14746 5977 15000 6667 3 FreeSans 520 180 0 0 VSWITCH
port 10 nsew power bidirectional
flabel metal4 s 0 5977 254 6667 3 FreeSans 520 0 0 0 VSWITCH
port 10 nsew power bidirectional
flabel metal4 s 0 12417 254 13307 3 FreeSans 520 0 0 0 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14746 10225 15000 10821 1 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 14746 9273 15000 9869 1 AMUXBUS_B
port 12 nsew signal bidirectional
rlabel metal4 s 14746 1377 15000 2307 1 VCCD
port 7 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 1 VCCD
port 7 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 1 VCCD
port 7 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 1 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 1 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 1 VCCHIB
port 3 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 1 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 1 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 1 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 1 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 1 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 1 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 1 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 1 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 1 VDDIO
port 9 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 1 VDDIO
port 9 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 1 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 100 9930 4880 10164 1 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10151 6948 14931 7636 1 VSSA
port 2 nsew ground bidirectional
rlabel metal3 s 10151 9930 14931 10164 1 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 0 6947 4875 7637 1 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 0 9147 254 9213 1 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 0 9929 4875 10165 1 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 0 10881 254 10947 1 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 10156 6947 15000 7637 1 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 10156 9929 15000 10165 1 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 14746 9147 15000 9213 1 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 14746 10881 15000 10947 1 VSSA
port 2 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 1 VSSA
port 2 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 1 VSSA
port 2 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 1 VSSA
port 2 nsew ground bidirectional
rlabel metal5 s 14746 9147 15000 10947 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14873 10111 14913 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14873 10027 14913 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14873 9943 14913 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14873 7580 14913 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14873 7492 14913 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14873 7404 14913 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14873 7316 14913 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14873 7228 14913 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14873 7140 14913 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14873 7052 14913 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14873 6964 14913 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14792 10111 14832 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14792 10027 14832 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14792 9943 14832 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14792 7580 14832 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14792 7492 14832 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14792 7404 14832 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14792 7316 14832 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14792 7228 14832 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14792 7140 14832 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14792 7052 14832 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14792 6964 14832 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14711 10111 14751 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14711 10027 14751 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14711 9943 14751 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14711 7580 14751 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14711 7492 14751 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14711 7404 14751 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14711 7316 14751 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14711 7228 14751 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14711 7140 14751 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14711 7052 14751 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14711 6964 14751 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14630 10111 14670 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14630 10027 14670 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14630 9943 14670 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14630 7580 14670 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14630 7492 14670 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14630 7404 14670 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14630 7316 14670 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14630 7228 14670 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14630 7140 14670 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14630 7052 14670 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14630 6964 14670 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14549 10111 14589 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14549 10027 14589 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14549 9943 14589 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14549 7580 14589 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14549 7492 14589 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14549 7404 14589 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14549 7316 14589 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14549 7228 14589 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14549 7140 14589 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14549 7052 14589 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14549 6964 14589 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14468 10111 14508 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14468 10027 14508 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14468 9943 14508 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14468 7580 14508 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14468 7492 14508 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14468 7404 14508 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14468 7316 14508 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14468 7228 14508 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14468 7140 14508 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14468 7052 14508 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14468 6964 14508 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14387 10111 14427 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14387 10027 14427 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14387 9943 14427 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14387 7580 14427 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14387 7492 14427 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14387 7404 14427 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14387 7316 14427 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14387 7228 14427 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14387 7140 14427 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14387 7052 14427 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14387 6964 14427 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14306 10111 14346 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14306 10027 14346 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14306 9943 14346 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14306 7580 14346 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14306 7492 14346 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14306 7404 14346 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14306 7316 14346 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14306 7228 14346 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14306 7140 14346 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14306 7052 14346 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14306 6964 14346 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14225 10111 14265 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14225 10027 14265 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14225 9943 14265 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14225 7580 14265 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14225 7492 14265 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14225 7404 14265 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14225 7316 14265 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14225 7228 14265 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14225 7140 14265 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14225 7052 14265 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14225 6964 14265 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14144 10111 14184 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14144 10027 14184 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14144 9943 14184 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14144 7580 14184 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14144 7492 14184 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14144 7404 14184 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14144 7316 14184 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14144 7228 14184 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14144 7140 14184 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14144 7052 14184 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14144 6964 14184 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14063 10111 14103 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14063 10027 14103 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14063 9943 14103 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14063 7580 14103 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14063 7492 14103 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14063 7404 14103 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14063 7316 14103 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14063 7228 14103 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14063 7140 14103 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14063 7052 14103 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 14063 6964 14103 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13982 10111 14022 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13982 10027 14022 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13982 9943 14022 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13982 7580 14022 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13982 7492 14022 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13982 7404 14022 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13982 7316 14022 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13982 7228 14022 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13982 7140 14022 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13982 7052 14022 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13982 6964 14022 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13901 10111 13941 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13901 10027 13941 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13901 9943 13941 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13901 7580 13941 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13901 7492 13941 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13901 7404 13941 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13901 7316 13941 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13901 7228 13941 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13901 7140 13941 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13901 7052 13941 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13901 6964 13941 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13820 10111 13860 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13820 10027 13860 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13820 9943 13860 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13820 7580 13860 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13820 7492 13860 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13820 7404 13860 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13820 7316 13860 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13820 7228 13860 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13820 7140 13860 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13820 7052 13860 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13820 6964 13860 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13739 10111 13779 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13739 10027 13779 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13739 9943 13779 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13739 7580 13779 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13739 7492 13779 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13739 7404 13779 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13739 7316 13779 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13739 7228 13779 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13739 7140 13779 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13739 7052 13779 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13739 6964 13779 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13658 10111 13698 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13658 10027 13698 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13658 9943 13698 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13658 7580 13698 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13658 7492 13698 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13658 7404 13698 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13658 7316 13698 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13658 7228 13698 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13658 7140 13698 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13658 7052 13698 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13658 6964 13698 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13577 10111 13617 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13577 10027 13617 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13577 9943 13617 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13577 7580 13617 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13577 7492 13617 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13577 7404 13617 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13577 7316 13617 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13577 7228 13617 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13577 7140 13617 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13577 7052 13617 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13577 6964 13617 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13496 10111 13536 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13496 10027 13536 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13496 9943 13536 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13496 7580 13536 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13496 7492 13536 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13496 7404 13536 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13496 7316 13536 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13496 7228 13536 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13496 7140 13536 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13496 7052 13536 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13496 6964 13536 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13415 10111 13455 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13415 10027 13455 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13415 9943 13455 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13415 7580 13455 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13415 7492 13455 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13415 7404 13455 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13415 7316 13455 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13415 7228 13455 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13415 7140 13455 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13415 7052 13455 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13415 6964 13455 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13334 10111 13374 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13334 10027 13374 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13334 9943 13374 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13334 7580 13374 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13334 7492 13374 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13334 7404 13374 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13334 7316 13374 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13334 7228 13374 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13334 7140 13374 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13334 7052 13374 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13334 6964 13374 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13253 10111 13293 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13253 10027 13293 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13253 9943 13293 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13253 7580 13293 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13253 7492 13293 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13253 7404 13293 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13253 7316 13293 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13253 7228 13293 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13253 7140 13293 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13253 7052 13293 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13253 6964 13293 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13172 10111 13212 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13172 10027 13212 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13172 9943 13212 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13172 7580 13212 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13172 7492 13212 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13172 7404 13212 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13172 7316 13212 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13172 7228 13212 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13172 7140 13212 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13172 7052 13212 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13172 6964 13212 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13091 10111 13131 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13091 10027 13131 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13091 9943 13131 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13091 7580 13131 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13091 7492 13131 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13091 7404 13131 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13091 7316 13131 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13091 7228 13131 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13091 7140 13131 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13091 7052 13131 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13091 6964 13131 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13010 10111 13050 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13010 10027 13050 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13010 9943 13050 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13010 7580 13050 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13010 7492 13050 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13010 7404 13050 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13010 7316 13050 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13010 7228 13050 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13010 7140 13050 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13010 7052 13050 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 13010 6964 13050 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12929 10111 12969 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12929 10027 12969 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12929 9943 12969 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12929 7580 12969 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12929 7492 12969 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12929 7404 12969 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12929 7316 12969 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12929 7228 12969 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12929 7140 12969 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12929 7052 12969 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12929 6964 12969 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12848 10111 12888 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12848 10027 12888 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12848 9943 12888 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12848 7580 12888 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12848 7492 12888 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12848 7404 12888 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12848 7316 12888 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12848 7228 12888 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12848 7140 12888 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12848 7052 12888 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12848 6964 12888 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12767 10111 12807 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12767 10027 12807 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12767 9943 12807 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12767 7580 12807 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12767 7492 12807 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12767 7404 12807 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12767 7316 12807 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12767 7228 12807 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12767 7140 12807 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12767 7052 12807 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12767 6964 12807 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12686 10111 12726 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12686 10027 12726 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12686 9943 12726 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12686 7580 12726 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12686 7492 12726 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12686 7404 12726 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12686 7316 12726 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12686 7228 12726 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12686 7140 12726 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12686 7052 12726 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12686 6964 12726 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12605 10111 12645 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12605 10027 12645 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12605 9943 12645 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12605 7580 12645 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12605 7492 12645 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12605 7404 12645 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12605 7316 12645 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12605 7228 12645 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12605 7140 12645 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12605 7052 12645 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12605 6964 12645 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12524 10111 12564 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12524 10027 12564 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12524 9943 12564 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12524 7580 12564 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12524 7492 12564 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12524 7404 12564 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12524 7316 12564 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12524 7228 12564 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12524 7140 12564 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12524 7052 12564 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12524 6964 12564 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12443 10111 12483 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12443 10027 12483 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12443 9943 12483 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12443 7580 12483 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12443 7492 12483 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12443 7404 12483 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12443 7316 12483 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12443 7228 12483 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12443 7140 12483 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12443 7052 12483 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12443 6964 12483 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12362 10111 12402 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12362 10027 12402 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12362 9943 12402 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12362 7580 12402 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12362 7492 12402 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12362 7404 12402 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12362 7316 12402 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12362 7228 12402 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12362 7140 12402 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12362 7052 12402 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12362 6964 12402 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12281 10111 12321 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12281 10027 12321 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12281 9943 12321 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12281 7580 12321 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12281 7492 12321 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12281 7404 12321 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12281 7316 12321 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12281 7228 12321 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12281 7140 12321 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12281 7052 12321 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12281 6964 12321 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12200 10111 12240 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12200 10027 12240 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12200 9943 12240 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12200 7580 12240 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12200 7492 12240 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12200 7404 12240 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12200 7316 12240 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12200 7228 12240 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12200 7140 12240 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12200 7052 12240 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12200 6964 12240 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12119 10111 12159 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12119 10027 12159 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12119 9943 12159 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12119 7580 12159 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12119 7492 12159 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12119 7404 12159 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12119 7316 12159 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12119 7228 12159 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12119 7140 12159 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12119 7052 12159 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12119 6964 12159 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12038 10111 12078 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12038 10027 12078 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12038 9943 12078 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12038 7580 12078 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12038 7492 12078 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12038 7404 12078 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12038 7316 12078 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12038 7228 12078 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12038 7140 12078 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12038 7052 12078 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 12038 6964 12078 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11957 10111 11997 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11957 10027 11997 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11957 9943 11997 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11957 7580 11997 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11957 7492 11997 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11957 7404 11997 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11957 7316 11997 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11957 7228 11997 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11957 7140 11997 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11957 7052 11997 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11957 6964 11997 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11876 10111 11916 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11876 10027 11916 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11876 9943 11916 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11876 7580 11916 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11876 7492 11916 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11876 7404 11916 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11876 7316 11916 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11876 7228 11916 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11876 7140 11916 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11876 7052 11916 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11876 6964 11916 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11795 10111 11835 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11795 10027 11835 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11795 9943 11835 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11795 7580 11835 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11795 7492 11835 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11795 7404 11835 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11795 7316 11835 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11795 7228 11835 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11795 7140 11835 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11795 7052 11835 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11795 6964 11835 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11714 10111 11754 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11714 10027 11754 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11714 9943 11754 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11714 7580 11754 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11714 7492 11754 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11714 7404 11754 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11714 7316 11754 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11714 7228 11754 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11714 7140 11754 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11714 7052 11754 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11714 6964 11754 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11633 10111 11673 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11633 10027 11673 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11633 9943 11673 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11633 7580 11673 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11633 7492 11673 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11633 7404 11673 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11633 7316 11673 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11633 7228 11673 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11633 7140 11673 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11633 7052 11673 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11633 6964 11673 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11552 10111 11592 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11552 10027 11592 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11552 9943 11592 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11552 7580 11592 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11552 7492 11592 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11552 7404 11592 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11552 7316 11592 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11552 7228 11592 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11552 7140 11592 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11552 7052 11592 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11552 6964 11592 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11471 10111 11511 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11471 10027 11511 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11471 9943 11511 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11471 7580 11511 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11471 7492 11511 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11471 7404 11511 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11471 7316 11511 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11471 7228 11511 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11471 7140 11511 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11471 7052 11511 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11471 6964 11511 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11390 10111 11430 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11390 10027 11430 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11390 9943 11430 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11390 7580 11430 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11390 7492 11430 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11390 7404 11430 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11390 7316 11430 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11390 7228 11430 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11390 7140 11430 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11390 7052 11430 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11390 6964 11430 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11309 10111 11349 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11309 10027 11349 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11309 9943 11349 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11309 7580 11349 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11309 7492 11349 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11309 7404 11349 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11309 7316 11349 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11309 7228 11349 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11309 7140 11349 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11309 7052 11349 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11309 6964 11349 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11228 10111 11268 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11228 10027 11268 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11228 9943 11268 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11228 7580 11268 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11228 7492 11268 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11228 7404 11268 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11228 7316 11268 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11228 7228 11268 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11228 7140 11268 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11228 7052 11268 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11228 6964 11268 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11147 10111 11187 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11147 10027 11187 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11147 9943 11187 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11147 7580 11187 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11147 7492 11187 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11147 7404 11187 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11147 7316 11187 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11147 7228 11187 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11147 7140 11187 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11147 7052 11187 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11147 6964 11187 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11066 10111 11106 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11066 10027 11106 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11066 9943 11106 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11066 7580 11106 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11066 7492 11106 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11066 7404 11106 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11066 7316 11106 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11066 7228 11106 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11066 7140 11106 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11066 7052 11106 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 11066 6964 11106 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10985 10111 11025 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10985 10027 11025 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10985 9943 11025 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10985 7580 11025 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10985 7492 11025 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10985 7404 11025 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10985 7316 11025 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10985 7228 11025 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10985 7140 11025 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10985 7052 11025 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10985 6964 11025 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10904 10111 10944 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10904 10027 10944 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10904 9943 10944 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10904 7580 10944 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10904 7492 10944 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10904 7404 10944 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10904 7316 10944 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10904 7228 10944 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10904 7140 10944 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10904 7052 10944 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10904 6964 10944 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10823 10111 10863 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10823 10027 10863 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10823 9943 10863 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10823 7580 10863 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10823 7492 10863 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10823 7404 10863 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10823 7316 10863 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10823 7228 10863 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10823 7140 10863 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10823 7052 10863 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10823 6964 10863 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10742 10111 10782 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10742 10027 10782 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10742 9943 10782 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10742 7580 10782 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10742 7492 10782 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10742 7404 10782 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10742 7316 10782 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10742 7228 10782 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10742 7140 10782 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10742 7052 10782 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10742 6964 10782 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10661 10111 10701 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10661 10027 10701 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10661 9943 10701 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10661 7580 10701 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10661 7492 10701 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10661 7404 10701 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10661 7316 10701 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10661 7228 10701 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10661 7140 10701 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10661 7052 10701 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10661 6964 10701 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10579 10111 10619 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10579 10027 10619 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10579 9943 10619 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10579 7580 10619 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10579 7492 10619 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10579 7404 10619 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10579 7316 10619 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10579 7228 10619 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10579 7140 10619 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10579 7052 10619 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10579 6964 10619 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10497 10111 10537 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10497 10027 10537 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10497 9943 10537 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10497 7580 10537 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10497 7492 10537 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10497 7404 10537 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10497 7316 10537 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10497 7228 10537 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10497 7140 10537 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10497 7052 10537 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10497 6964 10537 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10415 10111 10455 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10415 10027 10455 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10415 9943 10455 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10415 7580 10455 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10415 7492 10455 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10415 7404 10455 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10415 7316 10455 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10415 7228 10455 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10415 7140 10455 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10415 7052 10455 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10415 6964 10455 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10333 10111 10373 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10333 10027 10373 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10333 9943 10373 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10333 7580 10373 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10333 7492 10373 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10333 7404 10373 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10333 7316 10373 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10333 7228 10373 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10333 7140 10373 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10333 7052 10373 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10333 6964 10373 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10251 10111 10291 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10251 10027 10291 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10251 9943 10291 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10251 7580 10291 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10251 7492 10291 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10251 7404 10291 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10251 7316 10291 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10251 7228 10291 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10251 7140 10291 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10251 7052 10291 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10251 6964 10291 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10169 10111 10209 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10169 10027 10209 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10169 9943 10209 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10169 7580 10209 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10169 7492 10209 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10169 7404 10209 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10169 7316 10209 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10169 7228 10209 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10169 7140 10209 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10169 7052 10209 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 10169 6964 10209 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4822 10111 4862 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4822 10027 4862 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4822 9943 4862 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4822 7580 4862 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4822 7492 4862 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4822 7404 4862 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4822 7316 4862 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4822 7228 4862 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4822 7140 4862 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4822 7052 4862 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4822 6964 4862 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4741 10111 4781 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4741 10027 4781 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4741 9943 4781 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4741 7580 4781 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4741 7492 4781 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4741 7404 4781 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4741 7316 4781 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4741 7228 4781 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4741 7140 4781 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4741 7052 4781 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4741 6964 4781 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4660 10111 4700 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4660 10027 4700 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4660 9943 4700 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4660 7580 4700 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4660 7492 4700 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4660 7404 4700 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4660 7316 4700 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4660 7228 4700 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4660 7140 4700 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4660 7052 4700 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4660 6964 4700 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4579 10111 4619 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4579 10027 4619 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4579 9943 4619 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4579 7580 4619 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4579 7492 4619 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4579 7404 4619 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4579 7316 4619 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4579 7228 4619 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4579 7140 4619 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4579 7052 4619 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4579 6964 4619 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4498 10111 4538 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4498 10027 4538 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4498 9943 4538 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4498 7580 4538 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4498 7492 4538 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4498 7404 4538 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4498 7316 4538 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4498 7228 4538 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4498 7140 4538 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4498 7052 4538 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4498 6964 4538 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4417 10111 4457 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4417 10027 4457 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4417 9943 4457 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4417 7580 4457 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4417 7492 4457 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4417 7404 4457 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4417 7316 4457 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4417 7228 4457 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4417 7140 4457 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4417 7052 4457 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4417 6964 4457 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4336 10111 4376 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4336 10027 4376 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4336 9943 4376 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4336 7580 4376 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4336 7492 4376 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4336 7404 4376 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4336 7316 4376 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4336 7228 4376 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4336 7140 4376 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4336 7052 4376 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4336 6964 4376 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4255 10111 4295 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4255 10027 4295 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4255 9943 4295 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4255 7580 4295 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4255 7492 4295 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4255 7404 4295 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4255 7316 4295 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4255 7228 4295 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4255 7140 4295 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4255 7052 4295 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4255 6964 4295 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4174 10111 4214 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4174 10027 4214 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4174 9943 4214 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4174 7580 4214 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4174 7492 4214 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4174 7404 4214 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4174 7316 4214 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4174 7228 4214 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4174 7140 4214 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4174 7052 4214 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4174 6964 4214 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4093 10111 4133 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4093 10027 4133 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4093 9943 4133 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4093 7580 4133 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4093 7492 4133 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4093 7404 4133 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4093 7316 4133 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4093 7228 4133 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4093 7140 4133 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4093 7052 4133 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4093 6964 4133 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4012 10111 4052 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4012 10027 4052 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4012 9943 4052 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4012 7580 4052 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4012 7492 4052 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4012 7404 4052 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4012 7316 4052 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4012 7228 4052 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4012 7140 4052 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4012 7052 4052 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 4012 6964 4052 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3931 10111 3971 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3931 10027 3971 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3931 9943 3971 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3931 7580 3971 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3931 7492 3971 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3931 7404 3971 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3931 7316 3971 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3931 7228 3971 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3931 7140 3971 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3931 7052 3971 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3931 6964 3971 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3850 10111 3890 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3850 10027 3890 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3850 9943 3890 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3850 7580 3890 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3850 7492 3890 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3850 7404 3890 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3850 7316 3890 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3850 7228 3890 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3850 7140 3890 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3850 7052 3890 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3850 6964 3890 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3769 10111 3809 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3769 10027 3809 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3769 9943 3809 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3769 7580 3809 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3769 7492 3809 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3769 7404 3809 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3769 7316 3809 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3769 7228 3809 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3769 7140 3809 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3769 7052 3809 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3769 6964 3809 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3688 10111 3728 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3688 10027 3728 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3688 9943 3728 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3688 7580 3728 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3688 7492 3728 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3688 7404 3728 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3688 7316 3728 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3688 7228 3728 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3688 7140 3728 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3688 7052 3728 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3688 6964 3728 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3607 10111 3647 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3607 10027 3647 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3607 9943 3647 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3607 7580 3647 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3607 7492 3647 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3607 7404 3647 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3607 7316 3647 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3607 7228 3647 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3607 7140 3647 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3607 7052 3647 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3607 6964 3647 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3526 10111 3566 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3526 10027 3566 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3526 9943 3566 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3526 7580 3566 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3526 7492 3566 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3526 7404 3566 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3526 7316 3566 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3526 7228 3566 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3526 7140 3566 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3526 7052 3566 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3526 6964 3566 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3445 10111 3485 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3445 10027 3485 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3445 9943 3485 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3445 7580 3485 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3445 7492 3485 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3445 7404 3485 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3445 7316 3485 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3445 7228 3485 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3445 7140 3485 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3445 7052 3485 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3445 6964 3485 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3364 10111 3404 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3364 10027 3404 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3364 9943 3404 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3364 7580 3404 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3364 7492 3404 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3364 7404 3404 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3364 7316 3404 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3364 7228 3404 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3364 7140 3404 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3364 7052 3404 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3364 6964 3404 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3283 10111 3323 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3283 10027 3323 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3283 9943 3323 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3283 7580 3323 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3283 7492 3323 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3283 7404 3323 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3283 7316 3323 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3283 7228 3323 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3283 7140 3323 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3283 7052 3323 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3283 6964 3323 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3202 10111 3242 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3202 10027 3242 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3202 9943 3242 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3202 7580 3242 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3202 7492 3242 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3202 7404 3242 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3202 7316 3242 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3202 7228 3242 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3202 7140 3242 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3202 7052 3242 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3202 6964 3242 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3121 10111 3161 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3121 10027 3161 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3121 9943 3161 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3121 7580 3161 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3121 7492 3161 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3121 7404 3161 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3121 7316 3161 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3121 7228 3161 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3121 7140 3161 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3121 7052 3161 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3121 6964 3161 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3040 10111 3080 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3040 10027 3080 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3040 9943 3080 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3040 7580 3080 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3040 7492 3080 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3040 7404 3080 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3040 7316 3080 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3040 7228 3080 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3040 7140 3080 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3040 7052 3080 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 3040 6964 3080 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2959 10111 2999 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2959 10027 2999 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2959 9943 2999 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2959 7580 2999 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2959 7492 2999 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2959 7404 2999 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2959 7316 2999 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2959 7228 2999 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2959 7140 2999 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2959 7052 2999 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2959 6964 2999 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2878 10111 2918 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2878 10027 2918 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2878 9943 2918 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2878 7580 2918 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2878 7492 2918 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2878 7404 2918 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2878 7316 2918 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2878 7228 2918 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2878 7140 2918 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2878 7052 2918 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2878 6964 2918 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2797 10111 2837 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2797 10027 2837 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2797 9943 2837 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2797 7580 2837 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2797 7492 2837 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2797 7404 2837 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2797 7316 2837 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2797 7228 2837 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2797 7140 2837 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2797 7052 2837 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2797 6964 2837 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2716 10111 2756 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2716 10027 2756 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2716 9943 2756 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2716 7580 2756 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2716 7492 2756 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2716 7404 2756 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2716 7316 2756 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2716 7228 2756 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2716 7140 2756 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2716 7052 2756 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2716 6964 2756 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2635 10111 2675 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2635 10027 2675 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2635 9943 2675 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2635 7580 2675 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2635 7492 2675 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2635 7404 2675 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2635 7316 2675 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2635 7228 2675 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2635 7140 2675 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2635 7052 2675 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2635 6964 2675 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2554 10111 2594 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2554 10027 2594 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2554 9943 2594 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2554 7580 2594 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2554 7492 2594 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2554 7404 2594 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2554 7316 2594 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2554 7228 2594 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2554 7140 2594 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2554 7052 2594 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2554 6964 2594 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2473 10111 2513 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2473 10027 2513 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2473 9943 2513 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2473 7580 2513 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2473 7492 2513 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2473 7404 2513 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2473 7316 2513 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2473 7228 2513 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2473 7140 2513 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2473 7052 2513 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2473 6964 2513 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2392 10111 2432 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2392 10027 2432 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2392 9943 2432 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2392 7580 2432 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2392 7492 2432 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2392 7404 2432 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2392 7316 2432 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2392 7228 2432 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2392 7140 2432 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2392 7052 2432 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2392 6964 2432 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2311 10111 2351 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2311 10027 2351 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2311 9943 2351 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2311 7580 2351 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2311 7492 2351 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2311 7404 2351 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2311 7316 2351 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2311 7228 2351 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2311 7140 2351 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2311 7052 2351 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2311 6964 2351 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2230 10111 2270 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2230 10027 2270 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2230 9943 2270 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2230 7580 2270 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2230 7492 2270 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2230 7404 2270 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2230 7316 2270 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2230 7228 2270 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2230 7140 2270 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2230 7052 2270 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2230 6964 2270 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2149 10111 2189 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2149 10027 2189 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2149 9943 2189 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2149 7580 2189 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2149 7492 2189 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2149 7404 2189 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2149 7316 2189 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2149 7228 2189 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2149 7140 2189 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2149 7052 2189 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2149 6964 2189 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2068 10111 2108 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2068 10027 2108 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2068 9943 2108 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2068 7580 2108 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2068 7492 2108 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2068 7404 2108 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2068 7316 2108 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2068 7228 2108 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2068 7140 2108 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2068 7052 2108 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 2068 6964 2108 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1987 10111 2027 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1987 10027 2027 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1987 9943 2027 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1987 7580 2027 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1987 7492 2027 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1987 7404 2027 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1987 7316 2027 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1987 7228 2027 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1987 7140 2027 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1987 7052 2027 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1987 6964 2027 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1906 10111 1946 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1906 10027 1946 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1906 9943 1946 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1906 7580 1946 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1906 7492 1946 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1906 7404 1946 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1906 7316 1946 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1906 7228 1946 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1906 7140 1946 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1906 7052 1946 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1906 6964 1946 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1825 10111 1865 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1825 10027 1865 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1825 9943 1865 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1825 7580 1865 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1825 7492 1865 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1825 7404 1865 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1825 7316 1865 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1825 7228 1865 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1825 7140 1865 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1825 7052 1865 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1825 6964 1865 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1744 10111 1784 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1744 10027 1784 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1744 9943 1784 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1744 7580 1784 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1744 7492 1784 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1744 7404 1784 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1744 7316 1784 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1744 7228 1784 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1744 7140 1784 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1744 7052 1784 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1744 6964 1784 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1663 10111 1703 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1663 10027 1703 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1663 9943 1703 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1663 7580 1703 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1663 7492 1703 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1663 7404 1703 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1663 7316 1703 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1663 7228 1703 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1663 7140 1703 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1663 7052 1703 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1663 6964 1703 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1582 10111 1622 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1582 10027 1622 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1582 9943 1622 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1582 7580 1622 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1582 7492 1622 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1582 7404 1622 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1582 7316 1622 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1582 7228 1622 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1582 7140 1622 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1582 7052 1622 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1582 6964 1622 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1501 10111 1541 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1501 10027 1541 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1501 9943 1541 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1501 7580 1541 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1501 7492 1541 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1501 7404 1541 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1501 7316 1541 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1501 7228 1541 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1501 7140 1541 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1501 7052 1541 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1501 6964 1541 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1420 10111 1460 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1420 10027 1460 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1420 9943 1460 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1420 7580 1460 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1420 7492 1460 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1420 7404 1460 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1420 7316 1460 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1420 7228 1460 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1420 7140 1460 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1420 7052 1460 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1420 6964 1460 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1339 10111 1379 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1339 10027 1379 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1339 9943 1379 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1339 7580 1379 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1339 7492 1379 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1339 7404 1379 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1339 7316 1379 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1339 7228 1379 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1339 7140 1379 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1339 7052 1379 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1339 6964 1379 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1258 10111 1298 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1258 10027 1298 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1258 9943 1298 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1258 7580 1298 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1258 7492 1298 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1258 7404 1298 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1258 7316 1298 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1258 7228 1298 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1258 7140 1298 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1258 7052 1298 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1258 6964 1298 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1177 10111 1217 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1177 10027 1217 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1177 9943 1217 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1177 7580 1217 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1177 7492 1217 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1177 7404 1217 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1177 7316 1217 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1177 7228 1217 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1177 7140 1217 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1177 7052 1217 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1177 6964 1217 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1096 10111 1136 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1096 10027 1136 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1096 9943 1136 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1096 7580 1136 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1096 7492 1136 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1096 7404 1136 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1096 7316 1136 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1096 7228 1136 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1096 7140 1136 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1096 7052 1136 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1096 6964 1136 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1015 10111 1055 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1015 10027 1055 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1015 9943 1055 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1015 7580 1055 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1015 7492 1055 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1015 7404 1055 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1015 7316 1055 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1015 7228 1055 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1015 7140 1055 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1015 7052 1055 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 1015 6964 1055 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 934 10111 974 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 934 10027 974 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 934 9943 974 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 934 7580 974 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 934 7492 974 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 934 7404 974 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 934 7316 974 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 934 7228 974 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 934 7140 974 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 934 7052 974 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 934 6964 974 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 853 10111 893 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 853 10027 893 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 853 9943 893 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 853 7580 893 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 853 7492 893 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 853 7404 893 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 853 7316 893 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 853 7228 893 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 853 7140 893 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 853 7052 893 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 853 6964 893 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 772 10111 812 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 772 10027 812 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 772 9943 812 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 772 7580 812 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 772 7492 812 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 772 7404 812 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 772 7316 812 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 772 7228 812 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 772 7140 812 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 772 7052 812 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 772 6964 812 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 691 10111 731 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 691 10027 731 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 691 9943 731 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 691 7580 731 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 691 7492 731 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 691 7404 731 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 691 7316 731 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 691 7228 731 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 691 7140 731 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 691 7052 731 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 691 6964 731 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 610 10111 650 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 610 10027 650 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 610 9943 650 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 610 7580 650 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 610 7492 650 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 610 7404 650 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 610 7316 650 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 610 7228 650 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 610 7140 650 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 610 7052 650 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 610 6964 650 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 528 10111 568 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 528 10027 568 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 528 9943 568 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 528 7580 568 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 528 7492 568 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 528 7404 568 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 528 7316 568 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 528 7228 568 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 528 7140 568 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 528 7052 568 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 528 6964 568 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 446 10111 486 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 446 10027 486 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 446 9943 486 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 446 7580 486 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 446 7492 486 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 446 7404 486 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 446 7316 486 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 446 7228 486 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 446 7140 486 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 446 7052 486 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 446 6964 486 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 364 10111 404 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 364 10027 404 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 364 9943 404 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 364 7580 404 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 364 7492 404 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 364 7404 404 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 364 7316 404 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 364 7228 404 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 364 7140 404 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 364 7052 404 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 364 6964 404 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 282 10111 322 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 282 10027 322 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 282 9943 322 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 282 7580 322 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 282 7492 322 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 282 7404 322 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 282 7316 322 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 282 7228 322 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 282 7140 322 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 282 7052 322 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 282 6964 322 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 200 10111 240 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 200 10027 240 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 200 9943 240 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 200 7580 240 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 200 7492 240 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 200 7404 240 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 200 7316 240 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 200 7228 240 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 200 7140 240 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 200 7052 240 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 200 6964 240 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 118 10111 158 10151 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 118 10027 158 10067 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 118 9943 158 9983 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 118 7580 158 7620 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 118 7492 158 7532 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 118 7404 158 7444 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 118 7316 158 7356 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 118 7228 158 7268 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 118 7140 158 7180 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 118 7052 158 7092 1 VSSA
port 2 nsew ground bidirectional
rlabel via3 s 118 6964 158 7004 1 VSSA
port 2 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 1 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 1 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 1 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 1 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 1 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 1 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 1 VSSIO_Q
port 6 nsew ground bidirectional
rlabel metal4 s 14746 5977 15000 6667 1 VSWITCH
port 10 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 1 VSWITCH
port 10 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 1 VSWITCH
port 10 nsew power bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 39600
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string LEFsymmetry X Y R90
string GDS_END 446478
string GDS_START 354686
<< end >>
