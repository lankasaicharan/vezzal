magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
rect 889 315 1097 331
<< pwell >>
rect 17 157 295 242
rect 862 157 1529 241
rect 17 49 1529 157
rect 0 0 1536 49
<< scnmos >>
rect 96 132 126 216
rect 186 132 216 216
rect 458 47 488 131
rect 544 47 574 131
rect 616 47 646 131
rect 724 47 754 131
rect 832 47 862 131
rect 941 47 971 215
rect 1162 47 1192 215
rect 1248 47 1278 215
rect 1334 47 1364 215
rect 1420 47 1450 215
<< scpmoshvt >>
rect 84 481 114 609
rect 170 481 200 609
rect 367 485 397 613
rect 507 485 537 613
rect 579 485 609 613
rect 687 485 717 569
rect 795 485 825 569
rect 978 351 1008 603
rect 1168 367 1198 619
rect 1254 367 1284 619
rect 1340 367 1370 619
rect 1426 367 1456 619
<< ndiff >>
rect 43 186 96 216
rect 43 152 51 186
rect 85 152 96 186
rect 43 132 96 152
rect 126 188 186 216
rect 126 154 137 188
rect 171 154 186 188
rect 126 132 186 154
rect 216 198 269 216
rect 216 164 227 198
rect 261 164 269 198
rect 216 132 269 164
rect 888 161 941 215
rect 888 131 896 161
rect 405 104 458 131
rect 405 70 413 104
rect 447 70 458 104
rect 405 47 458 70
rect 488 89 544 131
rect 488 55 499 89
rect 533 55 544 89
rect 488 47 544 55
rect 574 47 616 131
rect 646 89 724 131
rect 646 55 666 89
rect 700 55 724 89
rect 646 47 724 55
rect 754 47 832 131
rect 862 127 896 131
rect 930 127 941 161
rect 862 93 941 127
rect 862 59 896 93
rect 930 59 941 93
rect 862 47 941 59
rect 971 199 1024 215
rect 971 165 982 199
rect 1016 165 1024 199
rect 971 101 1024 165
rect 971 67 982 101
rect 1016 67 1024 101
rect 971 47 1024 67
rect 1109 203 1162 215
rect 1109 169 1117 203
rect 1151 169 1162 203
rect 1109 93 1162 169
rect 1109 59 1117 93
rect 1151 59 1162 93
rect 1109 47 1162 59
rect 1192 203 1248 215
rect 1192 169 1203 203
rect 1237 169 1248 203
rect 1192 101 1248 169
rect 1192 67 1203 101
rect 1237 67 1248 101
rect 1192 47 1248 67
rect 1278 167 1334 215
rect 1278 133 1289 167
rect 1323 133 1334 167
rect 1278 93 1334 133
rect 1278 59 1289 93
rect 1323 59 1334 93
rect 1278 47 1334 59
rect 1364 203 1420 215
rect 1364 169 1375 203
rect 1409 169 1420 203
rect 1364 101 1420 169
rect 1364 67 1375 101
rect 1409 67 1420 101
rect 1364 47 1420 67
rect 1450 203 1503 215
rect 1450 169 1461 203
rect 1495 169 1503 203
rect 1450 93 1503 169
rect 1450 59 1461 93
rect 1495 59 1503 93
rect 1450 47 1503 59
<< pdiff >>
rect 27 595 84 609
rect 27 561 35 595
rect 69 561 84 595
rect 27 527 84 561
rect 27 493 35 527
rect 69 493 84 527
rect 27 481 84 493
rect 114 597 170 609
rect 114 563 125 597
rect 159 563 170 597
rect 114 529 170 563
rect 114 495 125 529
rect 159 495 170 529
rect 114 481 170 495
rect 200 597 253 609
rect 200 563 211 597
rect 245 563 253 597
rect 200 529 253 563
rect 200 495 211 529
rect 245 495 253 529
rect 200 481 253 495
rect 310 531 367 613
rect 310 497 322 531
rect 356 497 367 531
rect 310 485 367 497
rect 397 598 507 613
rect 397 564 462 598
rect 496 564 507 598
rect 397 485 507 564
rect 537 485 579 613
rect 609 588 662 613
rect 1115 607 1168 619
rect 609 554 620 588
rect 654 569 662 588
rect 925 591 978 603
rect 925 569 933 591
rect 654 554 687 569
rect 609 485 687 554
rect 717 485 795 569
rect 825 557 933 569
rect 967 557 978 591
rect 825 544 978 557
rect 825 510 841 544
rect 875 513 978 544
rect 875 510 933 513
rect 825 485 933 510
rect 925 479 933 485
rect 967 479 978 513
rect 925 437 978 479
rect 925 403 933 437
rect 967 403 978 437
rect 925 351 978 403
rect 1008 591 1061 603
rect 1008 557 1019 591
rect 1053 557 1061 591
rect 1008 494 1061 557
rect 1008 460 1019 494
rect 1053 460 1061 494
rect 1008 397 1061 460
rect 1008 363 1019 397
rect 1053 363 1061 397
rect 1115 573 1123 607
rect 1157 573 1168 607
rect 1115 507 1168 573
rect 1115 473 1123 507
rect 1157 473 1168 507
rect 1115 413 1168 473
rect 1115 379 1123 413
rect 1157 379 1168 413
rect 1115 367 1168 379
rect 1198 599 1254 619
rect 1198 565 1209 599
rect 1243 565 1254 599
rect 1198 503 1254 565
rect 1198 469 1209 503
rect 1243 469 1254 503
rect 1198 413 1254 469
rect 1198 379 1209 413
rect 1243 379 1254 413
rect 1198 367 1254 379
rect 1284 607 1340 619
rect 1284 573 1295 607
rect 1329 573 1340 607
rect 1284 531 1340 573
rect 1284 497 1295 531
rect 1329 497 1340 531
rect 1284 455 1340 497
rect 1284 421 1295 455
rect 1329 421 1340 455
rect 1284 367 1340 421
rect 1370 599 1426 619
rect 1370 565 1381 599
rect 1415 565 1426 599
rect 1370 503 1426 565
rect 1370 469 1381 503
rect 1415 469 1426 503
rect 1370 413 1426 469
rect 1370 379 1381 413
rect 1415 379 1426 413
rect 1370 367 1426 379
rect 1456 607 1509 619
rect 1456 573 1467 607
rect 1501 573 1509 607
rect 1456 513 1509 573
rect 1456 479 1467 513
rect 1501 479 1509 513
rect 1456 413 1509 479
rect 1456 379 1467 413
rect 1501 379 1509 413
rect 1456 367 1509 379
rect 1008 351 1061 363
<< ndiffc >>
rect 51 152 85 186
rect 137 154 171 188
rect 227 164 261 198
rect 413 70 447 104
rect 499 55 533 89
rect 666 55 700 89
rect 896 127 930 161
rect 896 59 930 93
rect 982 165 1016 199
rect 982 67 1016 101
rect 1117 169 1151 203
rect 1117 59 1151 93
rect 1203 169 1237 203
rect 1203 67 1237 101
rect 1289 133 1323 167
rect 1289 59 1323 93
rect 1375 169 1409 203
rect 1375 67 1409 101
rect 1461 169 1495 203
rect 1461 59 1495 93
<< pdiffc >>
rect 35 561 69 595
rect 35 493 69 527
rect 125 563 159 597
rect 125 495 159 529
rect 211 563 245 597
rect 211 495 245 529
rect 322 497 356 531
rect 462 564 496 598
rect 620 554 654 588
rect 933 557 967 591
rect 841 510 875 544
rect 933 479 967 513
rect 933 403 967 437
rect 1019 557 1053 591
rect 1019 460 1053 494
rect 1019 363 1053 397
rect 1123 573 1157 607
rect 1123 473 1157 507
rect 1123 379 1157 413
rect 1209 565 1243 599
rect 1209 469 1243 503
rect 1209 379 1243 413
rect 1295 573 1329 607
rect 1295 497 1329 531
rect 1295 421 1329 455
rect 1381 565 1415 599
rect 1381 469 1415 503
rect 1381 379 1415 413
rect 1467 573 1501 607
rect 1467 479 1501 513
rect 1467 379 1501 413
<< poly >>
rect 84 609 114 635
rect 170 609 200 635
rect 367 613 397 639
rect 507 613 537 639
rect 579 613 609 639
rect 978 603 1008 629
rect 1168 619 1198 645
rect 1254 619 1284 645
rect 1340 619 1370 645
rect 1426 619 1456 645
rect 687 569 717 595
rect 795 569 825 595
rect 84 304 114 481
rect 170 382 200 481
rect 170 352 216 382
rect 72 288 138 304
rect 72 254 88 288
rect 122 254 138 288
rect 72 238 138 254
rect 186 268 216 352
rect 367 313 397 485
rect 507 390 537 485
rect 471 374 537 390
rect 471 340 487 374
rect 521 340 537 374
rect 362 297 428 313
rect 186 238 314 268
rect 96 216 126 238
rect 186 216 216 238
rect 96 106 126 132
rect 186 106 216 132
rect 284 106 314 238
rect 362 263 378 297
rect 412 263 428 297
rect 362 229 428 263
rect 471 306 537 340
rect 579 453 609 485
rect 579 437 645 453
rect 579 403 595 437
rect 629 403 645 437
rect 579 369 645 403
rect 687 442 717 485
rect 795 453 825 485
rect 687 426 753 442
rect 687 392 703 426
rect 737 392 753 426
rect 795 437 893 453
rect 795 423 843 437
rect 687 376 753 392
rect 827 403 843 423
rect 877 403 893 437
rect 579 335 595 369
rect 629 335 645 369
rect 579 328 645 335
rect 827 369 893 403
rect 827 335 843 369
rect 877 335 893 369
rect 579 319 754 328
rect 827 319 893 335
rect 471 272 487 306
rect 521 272 537 306
rect 615 298 754 319
rect 471 256 537 272
rect 724 268 754 298
rect 832 268 868 319
rect 978 303 1008 351
rect 1168 319 1198 367
rect 1254 319 1284 367
rect 1340 319 1370 367
rect 1426 319 1456 367
rect 941 287 1008 303
rect 362 195 378 229
rect 412 195 428 229
rect 507 250 566 256
rect 507 226 574 250
rect 536 220 574 226
rect 362 184 428 195
rect 362 154 488 184
rect 458 131 488 154
rect 544 131 574 220
rect 616 229 682 245
rect 616 195 632 229
rect 666 195 682 229
rect 616 179 682 195
rect 724 213 790 268
rect 724 179 740 213
rect 774 179 790 213
rect 616 131 646 179
rect 724 163 790 179
rect 724 131 754 163
rect 832 131 862 268
rect 941 253 957 287
rect 991 253 1008 287
rect 1069 303 1456 319
rect 1069 269 1085 303
rect 1119 269 1153 303
rect 1187 269 1221 303
rect 1255 269 1289 303
rect 1323 289 1456 303
rect 1323 269 1450 289
rect 1069 253 1450 269
rect 941 237 1008 253
rect 941 215 971 237
rect 1162 215 1192 253
rect 1248 215 1278 253
rect 1334 215 1364 253
rect 1420 215 1450 253
rect 284 90 350 106
rect 284 56 300 90
rect 334 56 350 90
rect 284 40 350 56
rect 458 21 488 47
rect 544 21 574 47
rect 616 21 646 47
rect 724 21 754 47
rect 832 21 862 47
rect 941 21 971 47
rect 1162 21 1192 47
rect 1248 21 1278 47
rect 1334 21 1364 47
rect 1420 21 1450 47
<< polycont >>
rect 88 254 122 288
rect 487 340 521 374
rect 378 263 412 297
rect 595 403 629 437
rect 703 392 737 426
rect 843 403 877 437
rect 595 335 629 369
rect 843 335 877 369
rect 487 272 521 306
rect 378 195 412 229
rect 632 195 666 229
rect 740 179 774 213
rect 957 253 991 287
rect 1085 269 1119 303
rect 1153 269 1187 303
rect 1221 269 1255 303
rect 1289 269 1323 303
rect 300 56 334 90
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 18 595 82 611
rect 18 561 35 595
rect 69 561 82 595
rect 18 527 82 561
rect 18 493 35 527
rect 69 493 82 527
rect 18 376 82 493
rect 116 597 167 649
rect 116 563 125 597
rect 159 563 167 597
rect 116 529 167 563
rect 116 495 125 529
rect 159 495 167 529
rect 116 479 167 495
rect 201 597 426 615
rect 201 563 211 597
rect 245 581 426 597
rect 245 563 261 581
rect 201 529 261 563
rect 201 495 211 529
rect 245 495 261 529
rect 201 479 261 495
rect 306 531 356 547
rect 306 497 322 531
rect 306 444 356 497
rect 392 514 426 581
rect 460 598 512 649
rect 460 564 462 598
rect 496 564 512 598
rect 460 548 512 564
rect 604 588 807 604
rect 604 554 620 588
rect 654 554 807 588
rect 604 548 807 554
rect 392 480 739 514
rect 306 437 645 444
rect 306 410 595 437
rect 579 403 595 410
rect 629 403 645 437
rect 18 374 537 376
rect 18 340 487 374
rect 521 340 537 374
rect 18 202 52 340
rect 471 306 537 340
rect 579 369 645 403
rect 579 335 595 369
rect 629 335 645 369
rect 687 426 739 480
rect 687 392 703 426
rect 737 392 739 426
rect 86 288 257 304
rect 86 254 88 288
rect 122 254 257 288
rect 86 238 257 254
rect 339 297 428 306
rect 339 263 378 297
rect 412 263 428 297
rect 471 272 487 306
rect 521 272 537 306
rect 687 299 739 392
rect 471 263 537 272
rect 616 265 739 299
rect 773 283 807 548
rect 841 591 983 649
rect 1109 607 1166 649
rect 841 557 933 591
rect 967 557 983 591
rect 841 544 983 557
rect 875 513 983 544
rect 875 510 933 513
rect 841 487 933 510
rect 917 479 933 487
rect 967 479 983 513
rect 841 437 883 453
rect 841 403 843 437
rect 877 403 883 437
rect 917 437 983 479
rect 917 403 933 437
rect 967 403 983 437
rect 1017 591 1075 607
rect 1017 557 1019 591
rect 1053 557 1075 591
rect 1017 494 1075 557
rect 1017 460 1019 494
rect 1053 460 1075 494
rect 841 369 883 403
rect 1017 397 1075 460
rect 1017 369 1019 397
rect 841 335 843 369
rect 877 363 1019 369
rect 1053 363 1075 397
rect 1109 573 1123 607
rect 1157 573 1166 607
rect 1109 507 1166 573
rect 1109 473 1123 507
rect 1157 473 1166 507
rect 1109 413 1166 473
rect 1109 379 1123 413
rect 1157 379 1166 413
rect 1109 363 1166 379
rect 1200 599 1245 615
rect 1200 565 1209 599
rect 1243 565 1245 599
rect 1200 503 1245 565
rect 1200 469 1209 503
rect 1243 469 1245 503
rect 1200 413 1245 469
rect 1200 379 1209 413
rect 1243 379 1245 413
rect 1279 607 1338 649
rect 1279 573 1295 607
rect 1329 573 1338 607
rect 1279 531 1338 573
rect 1279 497 1295 531
rect 1329 497 1338 531
rect 1279 455 1338 497
rect 1279 421 1295 455
rect 1329 421 1338 455
rect 1279 405 1338 421
rect 1372 599 1419 615
rect 1372 565 1381 599
rect 1415 565 1419 599
rect 1372 503 1419 565
rect 1372 469 1381 503
rect 1415 469 1419 503
rect 1372 413 1419 469
rect 1200 371 1245 379
rect 1372 379 1381 413
rect 1415 379 1419 413
rect 1372 371 1419 379
rect 877 335 1075 363
rect 1200 337 1419 371
rect 1453 607 1517 649
rect 1453 573 1467 607
rect 1501 573 1517 607
rect 1453 513 1517 573
rect 1453 479 1467 513
rect 1501 479 1517 513
rect 1453 413 1517 479
rect 1453 379 1467 413
rect 1501 379 1517 413
rect 1453 363 1517 379
rect 841 319 877 335
rect 1041 303 1075 335
rect 941 287 1007 301
rect 941 283 957 287
rect 339 229 428 263
rect 616 229 682 265
rect 773 253 957 283
rect 991 253 1007 287
rect 773 249 1007 253
rect 1041 269 1085 303
rect 1119 269 1153 303
rect 1187 269 1221 303
rect 1255 269 1289 303
rect 1323 269 1339 303
rect 18 186 94 202
rect 18 152 51 186
rect 85 152 94 186
rect 18 136 94 152
rect 128 188 177 204
rect 339 202 378 229
rect 128 154 137 188
rect 171 154 177 188
rect 211 198 378 202
rect 211 164 227 198
rect 261 195 378 198
rect 412 195 632 229
rect 666 195 682 229
rect 261 193 682 195
rect 261 164 373 193
rect 724 179 740 213
rect 774 179 790 213
rect 724 159 790 179
rect 128 17 177 154
rect 211 90 369 130
rect 211 56 300 90
rect 334 56 369 90
rect 407 125 790 159
rect 407 104 447 125
rect 407 70 413 104
rect 826 91 860 249
rect 1041 215 1077 269
rect 1373 235 1419 337
rect 978 199 1077 215
rect 407 51 447 70
rect 483 89 549 91
rect 483 55 499 89
rect 533 55 549 89
rect 483 17 549 55
rect 650 89 860 91
rect 650 55 666 89
rect 700 55 860 89
rect 650 51 860 55
rect 894 161 944 177
rect 894 127 896 161
rect 930 127 944 161
rect 894 93 944 127
rect 894 59 896 93
rect 930 59 944 93
rect 894 17 944 59
rect 978 165 982 199
rect 1016 165 1077 199
rect 978 101 1077 165
rect 978 67 982 101
rect 1016 67 1077 101
rect 978 51 1077 67
rect 1111 203 1160 219
rect 1111 169 1117 203
rect 1151 169 1160 203
rect 1111 93 1160 169
rect 1111 59 1117 93
rect 1151 59 1160 93
rect 1111 17 1160 59
rect 1194 203 1419 235
rect 1194 169 1203 203
rect 1237 201 1375 203
rect 1237 169 1239 201
rect 1194 101 1239 169
rect 1409 169 1419 203
rect 1194 67 1203 101
rect 1237 67 1239 101
rect 1194 51 1239 67
rect 1273 133 1289 167
rect 1323 133 1339 167
rect 1273 93 1339 133
rect 1273 59 1289 93
rect 1323 59 1339 93
rect 1273 17 1339 59
rect 1375 101 1419 169
rect 1409 67 1419 101
rect 1375 51 1419 67
rect 1453 203 1499 219
rect 1453 169 1461 203
rect 1495 169 1499 203
rect 1453 93 1499 169
rect 1453 59 1461 93
rect 1495 59 1499 93
rect 1453 17 1499 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlxtn_4
flabel comment s 695 317 695 317 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1375 168 1409 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1375 390 1409 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 614594
string GDS_START 601744
<< end >>
