magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1288 -1260 2080 1731
use sky130_fd_pr__dfl1sd2__example_55959141808191  sky130_fd_pr__dfl1sd2__example_55959141808191_0
timestamp 1627201311
transform 1 0 50 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808191  sky130_fd_pr__dfl1sd2__example_55959141808191_1
timestamp 1627201311
transform 1 0 156 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808191  sky130_fd_pr__dfl1sd2__example_55959141808191_2
timestamp 1627201311
transform 1 0 262 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808191  sky130_fd_pr__dfl1sd2__example_55959141808191_3
timestamp 1627201311
transform 1 0 368 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808191  sky130_fd_pr__dfl1sd2__example_55959141808191_4
timestamp 1627201311
transform 1 0 474 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808191  sky130_fd_pr__dfl1sd2__example_55959141808191_5
timestamp 1627201311
transform 1 0 580 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808191  sky130_fd_pr__dfl1sd2__example_55959141808191_6
timestamp 1627201311
transform 1 0 686 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808190  sky130_fd_pr__dfl1sd__example_55959141808190_0
timestamp 1627201311
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808190  sky130_fd_pr__dfl1sd__example_55959141808190_1
timestamp 1627201311
transform 1 0 792 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 820 471 820 471 0 FreeSans 300 0 0 0 S
flabel comment s 714 471 714 471 0 FreeSans 300 0 0 0 D
flabel comment s 608 471 608 471 0 FreeSans 300 0 0 0 S
flabel comment s 502 471 502 471 0 FreeSans 300 0 0 0 D
flabel comment s 396 471 396 471 0 FreeSans 300 0 0 0 S
flabel comment s 290 471 290 471 0 FreeSans 300 0 0 0 D
flabel comment s 184 471 184 471 0 FreeSans 300 0 0 0 S
flabel comment s 78 471 78 471 0 FreeSans 300 0 0 0 D
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 35975314
string GDS_START 35970780
<< end >>
