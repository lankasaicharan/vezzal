magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 332 2054 704
<< pwell >>
rect 8 49 1812 248
rect 0 0 2016 49
<< scpmos >>
rect 81 368 117 592
rect 171 368 207 592
rect 261 368 297 592
rect 351 368 387 592
rect 441 368 477 592
rect 531 368 567 592
rect 621 368 657 592
rect 711 368 747 592
rect 801 368 837 592
rect 891 368 927 592
rect 981 368 1017 592
rect 1071 368 1107 592
rect 1265 368 1301 592
rect 1355 368 1391 592
rect 1445 368 1481 592
rect 1535 368 1571 592
rect 1625 368 1661 592
rect 1715 368 1751 592
rect 1805 368 1841 592
rect 1895 368 1931 592
<< nmoslvt >>
rect 91 74 121 222
rect 177 74 207 222
rect 263 74 293 222
rect 349 74 379 222
rect 435 74 465 222
rect 521 74 551 222
rect 607 74 637 222
rect 693 74 723 222
rect 927 74 957 222
rect 1013 74 1043 222
rect 1099 74 1129 222
rect 1185 74 1215 222
rect 1271 74 1301 222
rect 1527 74 1557 222
rect 1613 74 1643 222
rect 1699 74 1729 222
<< ndiff >>
rect 34 210 91 222
rect 34 176 46 210
rect 80 176 91 210
rect 34 120 91 176
rect 34 86 46 120
rect 80 86 91 120
rect 34 74 91 86
rect 121 152 177 222
rect 121 118 132 152
rect 166 118 177 152
rect 121 74 177 118
rect 207 210 263 222
rect 207 176 218 210
rect 252 176 263 210
rect 207 120 263 176
rect 207 86 218 120
rect 252 86 263 120
rect 207 74 263 86
rect 293 152 349 222
rect 293 118 304 152
rect 338 118 349 152
rect 293 74 349 118
rect 379 210 435 222
rect 379 176 390 210
rect 424 176 435 210
rect 379 120 435 176
rect 379 86 390 120
rect 424 86 435 120
rect 379 74 435 86
rect 465 120 521 222
rect 465 86 476 120
rect 510 86 521 120
rect 465 74 521 86
rect 551 207 607 222
rect 551 173 562 207
rect 596 173 607 207
rect 551 74 607 173
rect 637 120 693 222
rect 637 86 648 120
rect 682 86 693 120
rect 637 74 693 86
rect 723 207 776 222
rect 723 173 734 207
rect 768 173 776 207
rect 723 74 776 173
rect 874 207 927 222
rect 874 173 882 207
rect 916 173 927 207
rect 874 74 927 173
rect 957 120 1013 222
rect 957 86 968 120
rect 1002 86 1013 120
rect 957 74 1013 86
rect 1043 207 1099 222
rect 1043 173 1054 207
rect 1088 173 1099 207
rect 1043 74 1099 173
rect 1129 120 1185 222
rect 1129 86 1140 120
rect 1174 86 1185 120
rect 1129 74 1185 86
rect 1215 210 1271 222
rect 1215 176 1226 210
rect 1260 176 1271 210
rect 1215 120 1271 176
rect 1215 86 1226 120
rect 1260 86 1271 120
rect 1215 74 1271 86
rect 1301 127 1527 222
rect 1301 93 1326 127
rect 1360 93 1397 127
rect 1431 93 1468 127
rect 1502 93 1527 127
rect 1301 74 1527 93
rect 1557 194 1613 222
rect 1557 160 1568 194
rect 1602 160 1613 194
rect 1557 120 1613 160
rect 1557 86 1568 120
rect 1602 86 1613 120
rect 1557 74 1613 86
rect 1643 127 1699 222
rect 1643 93 1654 127
rect 1688 93 1699 127
rect 1643 74 1699 93
rect 1729 202 1786 222
rect 1729 168 1740 202
rect 1774 168 1786 202
rect 1729 120 1786 168
rect 1729 86 1740 120
rect 1774 86 1786 120
rect 1729 74 1786 86
<< pdiff >>
rect 29 580 81 592
rect 29 546 37 580
rect 71 546 81 580
rect 29 497 81 546
rect 29 463 37 497
rect 71 463 81 497
rect 29 414 81 463
rect 29 380 37 414
rect 71 380 81 414
rect 29 368 81 380
rect 117 580 171 592
rect 117 546 127 580
rect 161 546 171 580
rect 117 510 171 546
rect 117 476 127 510
rect 161 476 171 510
rect 117 440 171 476
rect 117 406 127 440
rect 161 406 171 440
rect 117 368 171 406
rect 207 580 261 592
rect 207 546 217 580
rect 251 546 261 580
rect 207 508 261 546
rect 207 474 217 508
rect 251 474 261 508
rect 207 368 261 474
rect 297 580 351 592
rect 297 546 307 580
rect 341 546 351 580
rect 297 510 351 546
rect 297 476 307 510
rect 341 476 351 510
rect 297 440 351 476
rect 297 406 307 440
rect 341 406 351 440
rect 297 368 351 406
rect 387 580 441 592
rect 387 546 397 580
rect 431 546 441 580
rect 387 508 441 546
rect 387 474 397 508
rect 431 474 441 508
rect 387 368 441 474
rect 477 580 531 592
rect 477 546 487 580
rect 521 546 531 580
rect 477 510 531 546
rect 477 476 487 510
rect 521 476 531 510
rect 477 440 531 476
rect 477 406 487 440
rect 521 406 531 440
rect 477 368 531 406
rect 567 580 621 592
rect 567 546 577 580
rect 611 546 621 580
rect 567 508 621 546
rect 567 474 577 508
rect 611 474 621 508
rect 567 368 621 474
rect 657 580 711 592
rect 657 546 667 580
rect 701 546 711 580
rect 657 510 711 546
rect 657 476 667 510
rect 701 476 711 510
rect 657 440 711 476
rect 657 406 667 440
rect 701 406 711 440
rect 657 368 711 406
rect 747 580 801 592
rect 747 546 757 580
rect 791 546 801 580
rect 747 508 801 546
rect 747 474 757 508
rect 791 474 801 508
rect 747 368 801 474
rect 837 580 891 592
rect 837 546 847 580
rect 881 546 891 580
rect 837 497 891 546
rect 837 463 847 497
rect 881 463 891 497
rect 837 414 891 463
rect 837 380 847 414
rect 881 380 891 414
rect 837 368 891 380
rect 927 580 981 592
rect 927 546 937 580
rect 971 546 981 580
rect 927 508 981 546
rect 927 474 937 508
rect 971 474 981 508
rect 927 368 981 474
rect 1017 580 1071 592
rect 1017 546 1027 580
rect 1061 546 1071 580
rect 1017 510 1071 546
rect 1017 476 1027 510
rect 1061 476 1071 510
rect 1017 440 1071 476
rect 1017 406 1027 440
rect 1061 406 1071 440
rect 1017 368 1071 406
rect 1107 580 1159 592
rect 1107 546 1117 580
rect 1151 546 1159 580
rect 1107 508 1159 546
rect 1107 474 1117 508
rect 1151 474 1159 508
rect 1107 368 1159 474
rect 1213 580 1265 592
rect 1213 546 1221 580
rect 1255 546 1265 580
rect 1213 498 1265 546
rect 1213 464 1221 498
rect 1255 464 1265 498
rect 1213 368 1265 464
rect 1301 531 1355 592
rect 1301 497 1311 531
rect 1345 497 1355 531
rect 1301 414 1355 497
rect 1301 380 1311 414
rect 1345 380 1355 414
rect 1301 368 1355 380
rect 1391 580 1445 592
rect 1391 546 1401 580
rect 1435 546 1445 580
rect 1391 498 1445 546
rect 1391 464 1401 498
rect 1435 464 1445 498
rect 1391 368 1445 464
rect 1481 531 1535 592
rect 1481 497 1491 531
rect 1525 497 1535 531
rect 1481 414 1535 497
rect 1481 380 1491 414
rect 1525 380 1535 414
rect 1481 368 1535 380
rect 1571 580 1625 592
rect 1571 546 1581 580
rect 1615 546 1625 580
rect 1571 497 1625 546
rect 1571 463 1581 497
rect 1615 463 1625 497
rect 1571 414 1625 463
rect 1571 380 1581 414
rect 1615 380 1625 414
rect 1571 368 1625 380
rect 1661 531 1715 592
rect 1661 497 1671 531
rect 1705 497 1715 531
rect 1661 414 1715 497
rect 1661 380 1671 414
rect 1705 380 1715 414
rect 1661 368 1715 380
rect 1751 580 1805 592
rect 1751 546 1761 580
rect 1795 546 1805 580
rect 1751 462 1805 546
rect 1751 428 1761 462
rect 1795 428 1805 462
rect 1751 368 1805 428
rect 1841 531 1895 592
rect 1841 497 1851 531
rect 1885 497 1895 531
rect 1841 414 1895 497
rect 1841 380 1851 414
rect 1885 380 1895 414
rect 1841 368 1895 380
rect 1931 580 1987 592
rect 1931 546 1941 580
rect 1975 546 1987 580
rect 1931 497 1987 546
rect 1931 463 1941 497
rect 1975 463 1987 497
rect 1931 414 1987 463
rect 1931 380 1941 414
rect 1975 380 1987 414
rect 1931 368 1987 380
<< ndiffc >>
rect 46 176 80 210
rect 46 86 80 120
rect 132 118 166 152
rect 218 176 252 210
rect 218 86 252 120
rect 304 118 338 152
rect 390 176 424 210
rect 390 86 424 120
rect 476 86 510 120
rect 562 173 596 207
rect 648 86 682 120
rect 734 173 768 207
rect 882 173 916 207
rect 968 86 1002 120
rect 1054 173 1088 207
rect 1140 86 1174 120
rect 1226 176 1260 210
rect 1226 86 1260 120
rect 1326 93 1360 127
rect 1397 93 1431 127
rect 1468 93 1502 127
rect 1568 160 1602 194
rect 1568 86 1602 120
rect 1654 93 1688 127
rect 1740 168 1774 202
rect 1740 86 1774 120
<< pdiffc >>
rect 37 546 71 580
rect 37 463 71 497
rect 37 380 71 414
rect 127 546 161 580
rect 127 476 161 510
rect 127 406 161 440
rect 217 546 251 580
rect 217 474 251 508
rect 307 546 341 580
rect 307 476 341 510
rect 307 406 341 440
rect 397 546 431 580
rect 397 474 431 508
rect 487 546 521 580
rect 487 476 521 510
rect 487 406 521 440
rect 577 546 611 580
rect 577 474 611 508
rect 667 546 701 580
rect 667 476 701 510
rect 667 406 701 440
rect 757 546 791 580
rect 757 474 791 508
rect 847 546 881 580
rect 847 463 881 497
rect 847 380 881 414
rect 937 546 971 580
rect 937 474 971 508
rect 1027 546 1061 580
rect 1027 476 1061 510
rect 1027 406 1061 440
rect 1117 546 1151 580
rect 1117 474 1151 508
rect 1221 546 1255 580
rect 1221 464 1255 498
rect 1311 497 1345 531
rect 1311 380 1345 414
rect 1401 546 1435 580
rect 1401 464 1435 498
rect 1491 497 1525 531
rect 1491 380 1525 414
rect 1581 546 1615 580
rect 1581 463 1615 497
rect 1581 380 1615 414
rect 1671 497 1705 531
rect 1671 380 1705 414
rect 1761 546 1795 580
rect 1761 428 1795 462
rect 1851 497 1885 531
rect 1851 380 1885 414
rect 1941 546 1975 580
rect 1941 463 1975 497
rect 1941 380 1975 414
<< poly >>
rect 81 592 117 618
rect 171 592 207 618
rect 261 592 297 618
rect 351 592 387 618
rect 441 592 477 618
rect 531 592 567 618
rect 621 592 657 618
rect 711 592 747 618
rect 801 592 837 618
rect 891 592 927 618
rect 981 592 1017 618
rect 1071 592 1107 618
rect 1265 592 1301 618
rect 1355 592 1391 618
rect 1445 592 1481 618
rect 1535 592 1571 618
rect 1625 592 1661 618
rect 1715 592 1751 618
rect 1805 592 1841 618
rect 1895 592 1931 618
rect 81 336 117 368
rect 171 336 207 368
rect 261 336 297 368
rect 351 336 387 368
rect 81 320 387 336
rect 81 286 121 320
rect 155 286 189 320
rect 223 286 257 320
rect 291 286 325 320
rect 359 286 387 320
rect 441 336 477 368
rect 531 336 567 368
rect 621 336 657 368
rect 711 336 747 368
rect 441 320 747 336
rect 441 300 457 320
rect 81 270 387 286
rect 435 286 457 300
rect 491 286 525 320
rect 559 286 593 320
rect 627 286 661 320
rect 695 286 747 320
rect 801 336 837 368
rect 891 336 927 368
rect 981 336 1017 368
rect 1071 336 1107 368
rect 801 320 1215 336
rect 801 306 943 320
rect 435 270 747 286
rect 927 286 943 306
rect 977 286 1023 320
rect 1057 286 1097 320
rect 1131 286 1165 320
rect 1199 286 1215 320
rect 927 270 1215 286
rect 91 222 121 270
rect 177 222 207 270
rect 263 222 293 270
rect 349 222 379 270
rect 435 222 465 270
rect 521 222 551 270
rect 607 222 637 270
rect 693 222 723 270
rect 927 222 957 270
rect 1013 222 1043 270
rect 1099 222 1129 270
rect 1185 222 1215 270
rect 1265 330 1301 368
rect 1355 330 1391 368
rect 1445 330 1481 368
rect 1535 330 1571 368
rect 1265 314 1571 330
rect 1265 280 1371 314
rect 1405 280 1439 314
rect 1473 280 1507 314
rect 1541 300 1571 314
rect 1625 310 1661 368
rect 1715 310 1751 368
rect 1805 310 1841 368
rect 1541 280 1557 300
rect 1265 264 1557 280
rect 1271 222 1301 264
rect 1527 222 1557 264
rect 1613 294 1841 310
rect 1895 294 1931 368
rect 1613 260 1629 294
rect 1663 260 1697 294
rect 1731 260 1765 294
rect 1799 260 1931 294
rect 1613 244 1931 260
rect 1613 222 1643 244
rect 1699 222 1729 244
rect 91 48 121 74
rect 177 48 207 74
rect 263 48 293 74
rect 349 48 379 74
rect 435 48 465 74
rect 521 48 551 74
rect 607 48 637 74
rect 693 48 723 74
rect 927 48 957 74
rect 1013 48 1043 74
rect 1099 48 1129 74
rect 1185 48 1215 74
rect 1271 48 1301 74
rect 1527 48 1557 74
rect 1613 48 1643 74
rect 1699 48 1729 74
<< polycont >>
rect 121 286 155 320
rect 189 286 223 320
rect 257 286 291 320
rect 325 286 359 320
rect 457 286 491 320
rect 525 286 559 320
rect 593 286 627 320
rect 661 286 695 320
rect 943 286 977 320
rect 1023 286 1057 320
rect 1097 286 1131 320
rect 1165 286 1199 320
rect 1371 280 1405 314
rect 1439 280 1473 314
rect 1507 280 1541 314
rect 1629 260 1663 294
rect 1697 260 1731 294
rect 1765 260 1799 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 21 580 71 649
rect 21 546 37 580
rect 21 497 71 546
rect 21 463 37 497
rect 21 414 71 463
rect 21 380 37 414
rect 111 580 161 596
rect 111 546 127 580
rect 111 510 161 546
rect 111 476 127 510
rect 111 440 161 476
rect 201 580 267 649
rect 201 546 217 580
rect 251 546 267 580
rect 201 508 267 546
rect 201 474 217 508
rect 251 474 267 508
rect 201 458 267 474
rect 307 580 341 596
rect 307 510 341 546
rect 111 406 127 440
rect 307 440 341 476
rect 381 580 447 649
rect 381 546 397 580
rect 431 546 447 580
rect 381 508 447 546
rect 381 474 397 508
rect 431 474 447 508
rect 381 458 447 474
rect 487 580 521 596
rect 487 510 521 546
rect 161 406 307 424
rect 487 440 521 476
rect 561 580 627 649
rect 561 546 577 580
rect 611 546 627 580
rect 561 508 627 546
rect 561 474 577 508
rect 611 474 627 508
rect 561 458 627 474
rect 667 580 701 596
rect 667 510 701 546
rect 341 406 487 424
rect 667 440 701 476
rect 741 580 807 649
rect 741 546 757 580
rect 791 546 807 580
rect 741 508 807 546
rect 741 474 757 508
rect 791 474 807 508
rect 741 458 807 474
rect 847 580 881 596
rect 847 497 881 546
rect 521 406 667 424
rect 847 424 881 463
rect 921 580 971 649
rect 921 546 937 580
rect 921 508 971 546
rect 921 474 937 508
rect 921 458 971 474
rect 1011 580 1061 596
rect 1011 546 1027 580
rect 1011 510 1061 546
rect 1011 476 1027 510
rect 1011 440 1061 476
rect 1101 580 1167 649
rect 1101 546 1117 580
rect 1151 546 1167 580
rect 1101 508 1167 546
rect 1101 474 1117 508
rect 1151 474 1167 508
rect 1101 458 1167 474
rect 1205 581 1991 615
rect 1205 580 1271 581
rect 1205 546 1221 580
rect 1255 546 1271 580
rect 1385 580 1451 581
rect 1205 498 1271 546
rect 1205 464 1221 498
rect 1255 464 1271 498
rect 1305 531 1351 547
rect 1305 497 1311 531
rect 1345 497 1351 531
rect 1011 424 1027 440
rect 701 414 1027 424
rect 701 406 847 414
rect 111 390 847 406
rect 21 364 71 380
rect 881 406 1027 414
rect 1305 430 1351 497
rect 1385 546 1401 580
rect 1435 546 1451 580
rect 1565 580 1631 581
rect 1385 498 1451 546
rect 1385 464 1401 498
rect 1435 464 1451 498
rect 1485 531 1531 547
rect 1485 497 1491 531
rect 1525 497 1531 531
rect 1485 430 1531 497
rect 1295 424 1531 430
rect 1061 414 1531 424
rect 1061 406 1311 414
rect 881 390 1311 406
rect 847 364 881 380
rect 1295 380 1311 390
rect 1345 380 1491 414
rect 1525 380 1531 414
rect 1295 364 1531 380
rect 1565 546 1581 580
rect 1615 546 1631 580
rect 1745 580 1811 581
rect 1565 497 1631 546
rect 1565 463 1581 497
rect 1615 463 1631 497
rect 1565 414 1631 463
rect 1565 380 1581 414
rect 1615 380 1631 414
rect 1565 364 1631 380
rect 1671 531 1705 547
rect 1671 414 1705 497
rect 1745 546 1761 580
rect 1795 546 1811 580
rect 1925 580 1991 581
rect 1745 462 1811 546
rect 1745 428 1761 462
rect 1795 428 1811 462
rect 1745 412 1811 428
rect 1851 531 1885 547
rect 1851 414 1885 497
rect 1671 378 1705 380
rect 1851 378 1885 380
rect 105 320 375 356
rect 105 286 121 320
rect 155 286 189 320
rect 223 286 257 320
rect 291 286 325 320
rect 359 286 375 320
rect 105 270 375 286
rect 409 320 743 356
rect 409 286 457 320
rect 491 286 525 320
rect 559 286 593 320
rect 627 286 661 320
rect 695 286 743 320
rect 409 270 743 286
rect 927 320 1223 356
rect 1671 344 1885 378
rect 1925 546 1941 580
rect 1975 546 1991 580
rect 1925 497 1991 546
rect 1925 463 1941 497
rect 1975 463 1991 497
rect 1925 414 1991 463
rect 1925 380 1941 414
rect 1975 380 1991 414
rect 1925 364 1991 380
rect 927 286 943 320
rect 977 286 1023 320
rect 1057 286 1097 320
rect 1131 286 1165 320
rect 1199 286 1223 320
rect 927 270 1223 286
rect 1355 314 1557 330
rect 1355 280 1371 314
rect 1405 280 1439 314
rect 1473 280 1507 314
rect 1541 280 1557 314
rect 1355 264 1557 280
rect 1613 294 1815 310
rect 1355 236 1511 264
rect 1613 260 1629 294
rect 1663 260 1697 294
rect 1731 260 1765 294
rect 1799 260 1815 294
rect 1613 244 1815 260
rect 1657 236 1815 244
rect 30 210 784 236
rect 30 176 46 210
rect 80 202 218 210
rect 30 120 80 176
rect 202 176 218 202
rect 252 202 390 210
rect 30 86 46 120
rect 30 70 80 86
rect 116 152 166 168
rect 116 118 132 152
rect 116 17 166 118
rect 202 120 252 176
rect 424 207 784 210
rect 424 195 562 207
rect 202 86 218 120
rect 202 70 252 86
rect 288 152 354 168
rect 288 118 304 152
rect 338 118 354 152
rect 288 17 354 118
rect 390 120 424 176
rect 546 173 562 195
rect 596 195 734 207
rect 596 173 612 195
rect 546 154 612 173
rect 718 173 734 195
rect 768 173 784 207
rect 718 154 784 173
rect 866 210 1276 226
rect 866 207 1226 210
rect 866 173 882 207
rect 916 173 1054 207
rect 1088 176 1226 207
rect 1260 202 1276 210
rect 1552 202 1602 210
rect 1851 202 1885 344
rect 1260 194 1740 202
rect 1260 176 1568 194
rect 1088 173 1568 176
rect 866 170 1568 173
rect 866 154 932 170
rect 1226 168 1568 170
rect 390 70 424 86
rect 460 120 512 136
rect 646 120 684 136
rect 1124 120 1190 136
rect 460 86 476 120
rect 510 86 648 120
rect 682 86 968 120
rect 1002 86 1140 120
rect 1174 86 1190 120
rect 460 70 1190 86
rect 1226 120 1276 168
rect 1552 160 1568 168
rect 1602 168 1740 194
rect 1774 168 1885 202
rect 1260 86 1276 120
rect 1226 70 1276 86
rect 1310 127 1518 134
rect 1310 93 1326 127
rect 1360 93 1397 127
rect 1431 93 1468 127
rect 1502 93 1518 127
rect 1310 17 1518 93
rect 1552 120 1602 160
rect 1740 134 1885 168
rect 1552 86 1568 120
rect 1552 70 1602 86
rect 1638 127 1704 134
rect 1638 93 1654 127
rect 1688 93 1704 127
rect 1638 17 1704 93
rect 1740 120 1991 134
rect 1774 86 1991 120
rect 1740 70 1991 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a311oi_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1759 94 1793 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1855 94 1889 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1951 94 1985 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 2124910
string GDS_START 2109152
<< end >>
