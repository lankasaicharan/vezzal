magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4946 1975
<< nwell >>
rect -38 383 3686 704
rect -38 331 534 383
rect 1396 331 3686 383
rect 1396 286 2020 331
rect 2316 311 2965 331
rect 2703 307 2965 311
<< pwell >>
rect 640 233 746 341
rect 983 233 1354 325
rect 640 207 1354 233
rect 194 187 1354 207
rect 2062 207 2172 275
rect 3451 209 3647 251
rect 2643 207 3647 209
rect 194 165 1534 187
rect 1 157 1534 165
rect 2062 157 3647 207
rect 1 49 3647 157
rect 0 0 3648 49
<< scnmos >>
rect 82 55 112 139
rect 275 97 305 181
rect 361 97 391 181
rect 439 97 469 181
rect 525 97 555 181
rect 742 89 772 173
rect 849 123 879 207
rect 1085 215 1115 299
rect 1171 215 1201 299
rect 1243 215 1273 299
rect 1343 77 1373 161
rect 1423 77 1453 161
rect 1638 47 1668 131
rect 1724 47 1754 131
rect 1810 47 1840 131
rect 1882 47 1912 131
rect 2168 97 2198 181
rect 2246 97 2276 181
rect 2318 97 2348 181
rect 2450 97 2480 181
rect 2528 97 2558 181
rect 2733 55 2763 183
rect 2849 99 2879 183
rect 2921 99 2951 183
rect 2999 99 3029 183
rect 3085 99 3115 183
rect 3163 99 3193 183
rect 3425 57 3455 141
rect 3534 57 3564 225
<< scpmoshvt >>
rect 117 491 147 619
rect 217 491 247 619
rect 295 491 325 619
rect 381 491 411 619
rect 509 491 539 619
rect 742 419 772 547
rect 902 419 932 547
rect 1011 419 1041 503
rect 1083 419 1113 503
rect 1192 419 1242 619
rect 1345 419 1395 619
rect 1632 341 1682 541
rect 1724 341 1774 541
rect 1862 341 1912 541
rect 2214 419 2244 547
rect 2300 419 2330 547
rect 2405 347 2455 547
rect 2615 427 2645 511
rect 2687 427 2717 511
rect 2792 343 2822 511
rect 3064 463 3094 547
rect 3150 463 3180 547
rect 3236 463 3266 547
rect 3429 491 3459 619
rect 3536 367 3566 619
<< ndiff >>
rect 666 303 720 315
rect 666 269 676 303
rect 710 269 720 303
rect 220 156 275 181
rect 27 114 82 139
rect 27 80 37 114
rect 71 80 82 114
rect 27 55 82 80
rect 112 114 166 139
rect 112 80 123 114
rect 157 80 166 114
rect 220 122 230 156
rect 264 122 275 156
rect 220 97 275 122
rect 305 169 361 181
rect 305 135 316 169
rect 350 135 361 169
rect 305 97 361 135
rect 391 97 439 181
rect 469 169 525 181
rect 469 135 480 169
rect 514 135 525 169
rect 469 97 525 135
rect 555 147 612 181
rect 555 113 566 147
rect 600 113 612 147
rect 555 97 612 113
rect 666 173 720 269
rect 799 173 849 207
rect 112 55 166 80
rect 666 89 742 173
rect 772 135 849 173
rect 772 101 783 135
rect 817 123 849 135
rect 879 182 936 207
rect 879 148 890 182
rect 924 148 936 182
rect 879 123 936 148
rect 817 101 827 123
rect 772 89 827 101
rect 1009 215 1085 299
rect 1115 289 1171 299
rect 1115 255 1126 289
rect 1160 255 1171 289
rect 1115 215 1171 255
rect 1201 215 1243 299
rect 1273 266 1328 299
rect 1273 232 1284 266
rect 1318 232 1328 266
rect 1273 215 1328 232
rect 1009 153 1063 215
rect 1009 119 1019 153
rect 1053 119 1063 153
rect 1009 107 1063 119
rect 1284 153 1343 161
rect 1284 119 1296 153
rect 1330 119 1343 153
rect 1284 77 1343 119
rect 1373 77 1423 161
rect 1453 124 1508 161
rect 2088 237 2146 249
rect 2088 203 2100 237
rect 2134 203 2146 237
rect 2088 181 2146 203
rect 3477 213 3534 225
rect 1453 90 1464 124
rect 1498 90 1508 124
rect 1453 77 1508 90
rect 1562 73 1638 131
rect 1562 39 1572 73
rect 1606 47 1638 73
rect 1668 110 1724 131
rect 1668 76 1679 110
rect 1713 76 1724 110
rect 1668 47 1724 76
rect 1754 106 1810 131
rect 1754 72 1765 106
rect 1799 72 1810 106
rect 1754 47 1810 72
rect 1840 47 1882 131
rect 1912 110 1969 131
rect 1912 76 1923 110
rect 1957 76 1969 110
rect 2088 97 2168 181
rect 2198 97 2246 181
rect 2276 97 2318 181
rect 2348 97 2450 181
rect 2480 97 2528 181
rect 2558 169 2615 181
rect 2558 135 2569 169
rect 2603 135 2615 169
rect 2558 97 2615 135
rect 2669 104 2733 183
rect 1912 47 1969 76
rect 2370 73 2428 97
rect 1606 39 1616 47
rect 1562 27 1616 39
rect 2370 39 2382 73
rect 2416 39 2428 73
rect 2669 70 2681 104
rect 2715 70 2733 104
rect 2669 55 2733 70
rect 2763 170 2849 183
rect 2763 136 2781 170
rect 2815 136 2849 170
rect 2763 99 2849 136
rect 2879 99 2921 183
rect 2951 99 2999 183
rect 3029 158 3085 183
rect 3029 124 3040 158
rect 3074 124 3085 158
rect 3029 99 3085 124
rect 3115 99 3163 183
rect 3193 170 3273 183
rect 3193 136 3227 170
rect 3261 136 3273 170
rect 3477 179 3489 213
rect 3523 179 3534 213
rect 3477 141 3534 179
rect 3193 99 3273 136
rect 3368 116 3425 141
rect 2763 55 2827 99
rect 3368 82 3380 116
rect 3414 82 3425 116
rect 3368 57 3425 82
rect 3455 103 3534 141
rect 3455 69 3489 103
rect 3523 69 3534 103
rect 3455 57 3534 69
rect 3564 213 3621 225
rect 3564 179 3575 213
rect 3609 179 3621 213
rect 3564 103 3621 179
rect 3564 69 3575 103
rect 3609 69 3621 103
rect 3564 57 3621 69
rect 2370 27 2428 39
<< pdiff >>
rect 60 568 117 619
rect 60 534 72 568
rect 106 534 117 568
rect 60 491 117 534
rect 147 607 217 619
rect 147 573 172 607
rect 206 573 217 607
rect 147 537 217 573
rect 147 503 172 537
rect 206 503 217 537
rect 147 491 217 503
rect 247 491 295 619
rect 325 569 381 619
rect 325 535 336 569
rect 370 535 381 569
rect 325 491 381 535
rect 411 491 509 619
rect 539 607 596 619
rect 539 573 550 607
rect 584 573 596 607
rect 539 491 596 573
rect 685 498 742 547
rect 685 464 697 498
rect 731 464 742 498
rect 685 419 742 464
rect 772 535 902 547
rect 772 501 857 535
rect 891 501 902 535
rect 772 465 902 501
rect 772 431 857 465
rect 891 431 902 465
rect 772 419 902 431
rect 932 503 989 547
rect 1135 503 1192 619
rect 932 469 943 503
rect 977 469 1011 503
rect 932 419 1011 469
rect 1041 419 1083 503
rect 1113 498 1192 503
rect 1113 464 1147 498
rect 1181 464 1192 498
rect 1113 419 1192 464
rect 1242 419 1345 619
rect 1395 593 1525 619
rect 1395 559 1483 593
rect 1517 559 1525 593
rect 1395 419 1525 559
rect 1789 588 1840 600
rect 1789 554 1798 588
rect 1832 554 1840 588
rect 1789 541 1840 554
rect 3374 568 3429 619
rect 1579 430 1632 541
rect 1579 396 1587 430
rect 1621 396 1632 430
rect 1579 341 1632 396
rect 1682 341 1724 541
rect 1774 341 1862 541
rect 1912 368 1984 541
rect 2157 527 2214 547
rect 1912 341 1942 368
rect 1934 334 1942 341
rect 1976 334 1984 368
rect 1934 322 1984 334
rect 2157 493 2169 527
rect 2203 493 2214 527
rect 2157 419 2214 493
rect 2244 498 2300 547
rect 2244 464 2255 498
rect 2289 464 2300 498
rect 2244 419 2300 464
rect 2330 521 2405 547
rect 2330 487 2360 521
rect 2394 487 2405 521
rect 2330 419 2405 487
rect 2352 347 2405 419
rect 2455 535 2508 547
rect 2455 501 2466 535
rect 2500 501 2508 535
rect 3007 523 3064 547
rect 2455 464 2508 501
rect 2455 430 2466 464
rect 2500 430 2508 464
rect 2455 393 2508 430
rect 2562 499 2615 511
rect 2562 465 2570 499
rect 2604 465 2615 499
rect 2562 427 2615 465
rect 2645 427 2687 511
rect 2717 499 2792 511
rect 2717 465 2747 499
rect 2781 465 2792 499
rect 2717 427 2792 465
rect 2455 359 2466 393
rect 2500 359 2508 393
rect 2455 347 2508 359
rect 2739 389 2792 427
rect 2739 355 2747 389
rect 2781 355 2792 389
rect 2739 343 2792 355
rect 2822 463 2929 511
rect 3007 489 3019 523
rect 3053 489 3064 523
rect 3007 463 3064 489
rect 3094 523 3150 547
rect 3094 489 3105 523
rect 3139 489 3150 523
rect 3094 463 3150 489
rect 3180 522 3236 547
rect 3180 488 3191 522
rect 3225 488 3236 522
rect 3180 463 3236 488
rect 3266 522 3320 547
rect 3266 488 3277 522
rect 3311 488 3320 522
rect 3374 534 3384 568
rect 3418 534 3429 568
rect 3374 491 3429 534
rect 3459 607 3536 619
rect 3459 573 3491 607
rect 3525 573 3536 607
rect 3459 510 3536 573
rect 3459 491 3491 510
rect 3266 463 3320 488
rect 2822 429 2883 463
rect 2917 429 2929 463
rect 2822 389 2929 429
rect 2822 355 2883 389
rect 2917 355 2929 389
rect 2822 343 2929 355
rect 3481 476 3491 491
rect 3525 476 3536 510
rect 3481 413 3536 476
rect 3481 379 3491 413
rect 3525 379 3536 413
rect 3481 367 3536 379
rect 3566 599 3621 619
rect 3566 565 3577 599
rect 3611 565 3621 599
rect 3566 506 3621 565
rect 3566 472 3577 506
rect 3611 472 3621 506
rect 3566 413 3621 472
rect 3566 379 3577 413
rect 3611 379 3621 413
rect 3566 367 3621 379
<< ndiffc >>
rect 676 269 710 303
rect 37 80 71 114
rect 123 80 157 114
rect 230 122 264 156
rect 316 135 350 169
rect 480 135 514 169
rect 566 113 600 147
rect 783 101 817 135
rect 890 148 924 182
rect 1126 255 1160 289
rect 1284 232 1318 266
rect 1019 119 1053 153
rect 1296 119 1330 153
rect 2100 203 2134 237
rect 1464 90 1498 124
rect 1572 39 1606 73
rect 1679 76 1713 110
rect 1765 72 1799 106
rect 1923 76 1957 110
rect 2569 135 2603 169
rect 2382 39 2416 73
rect 2681 70 2715 104
rect 2781 136 2815 170
rect 3040 124 3074 158
rect 3227 136 3261 170
rect 3489 179 3523 213
rect 3380 82 3414 116
rect 3489 69 3523 103
rect 3575 179 3609 213
rect 3575 69 3609 103
<< pdiffc >>
rect 72 534 106 568
rect 172 573 206 607
rect 172 503 206 537
rect 336 535 370 569
rect 550 573 584 607
rect 697 464 731 498
rect 857 501 891 535
rect 857 431 891 465
rect 943 469 977 503
rect 1147 464 1181 498
rect 1483 559 1517 593
rect 1798 554 1832 588
rect 1587 396 1621 430
rect 1942 334 1976 368
rect 2169 493 2203 527
rect 2255 464 2289 498
rect 2360 487 2394 521
rect 2466 501 2500 535
rect 2466 430 2500 464
rect 2570 465 2604 499
rect 2747 465 2781 499
rect 2466 359 2500 393
rect 2747 355 2781 389
rect 3019 489 3053 523
rect 3105 489 3139 523
rect 3191 488 3225 522
rect 3277 488 3311 522
rect 3384 534 3418 568
rect 3491 573 3525 607
rect 2883 429 2917 463
rect 2883 355 2917 389
rect 3491 476 3525 510
rect 3491 379 3525 413
rect 3577 565 3611 599
rect 3577 472 3611 506
rect 3577 379 3611 413
<< poly >>
rect 117 619 147 645
rect 217 619 247 645
rect 295 619 325 645
rect 381 619 411 645
rect 509 619 539 645
rect 742 615 1113 645
rect 1192 619 1242 645
rect 1345 619 1395 645
rect 742 547 772 615
rect 902 547 932 573
rect 117 353 147 491
rect 217 353 247 491
rect 117 337 247 353
rect 117 303 133 337
rect 167 323 247 337
rect 295 341 325 491
rect 381 455 411 491
rect 509 461 539 491
rect 381 439 461 455
rect 381 405 411 439
rect 445 405 461 439
rect 509 439 577 461
rect 509 431 527 439
rect 381 389 461 405
rect 431 383 461 389
rect 511 405 527 431
rect 561 405 577 439
rect 1011 503 1041 615
rect 1083 503 1113 615
rect 1632 615 3180 645
rect 3429 619 3459 645
rect 3536 619 3566 645
rect 1632 541 1682 615
rect 1724 541 1774 567
rect 1862 541 1912 567
rect 2214 547 2244 573
rect 2300 547 2330 573
rect 2405 547 2455 573
rect 3064 547 3094 573
rect 3150 547 3180 615
rect 3236 547 3266 573
rect 431 353 463 383
rect 295 325 383 341
rect 167 303 183 323
rect 117 269 183 303
rect 295 291 311 325
rect 345 305 383 325
rect 345 291 391 305
rect 295 275 391 291
rect 117 235 133 269
rect 167 235 183 269
rect 117 233 183 235
rect 82 203 305 233
rect 82 139 112 203
rect 275 181 305 203
rect 361 181 391 275
rect 433 273 463 353
rect 511 371 577 405
rect 511 337 527 371
rect 561 337 577 371
rect 511 321 577 337
rect 433 243 469 273
rect 439 181 469 243
rect 525 181 555 321
rect 742 173 772 419
rect 902 259 932 419
rect 1011 387 1041 419
rect 1083 387 1113 419
rect 1192 387 1242 419
rect 1010 371 1115 387
rect 1010 337 1026 371
rect 1060 337 1115 371
rect 1192 371 1297 387
rect 1192 351 1247 371
rect 1010 321 1115 337
rect 1085 299 1115 321
rect 1171 337 1247 351
rect 1281 337 1297 371
rect 1171 321 1297 337
rect 1171 299 1201 321
rect 1243 299 1273 321
rect 849 229 987 259
rect 849 207 879 229
rect 275 71 305 97
rect 361 71 391 97
rect 439 71 469 97
rect 525 71 555 97
rect 849 97 879 123
rect 957 101 987 229
rect 1345 291 1395 419
rect 1632 309 1682 341
rect 1562 293 1682 309
rect 1345 272 1514 291
rect 1345 261 1464 272
rect 1085 189 1115 215
rect 1171 189 1201 215
rect 1243 189 1273 215
rect 1345 213 1375 261
rect 1343 183 1375 213
rect 1423 238 1464 261
rect 1498 238 1514 272
rect 1562 259 1578 293
rect 1612 279 1682 293
rect 1724 304 1774 341
rect 1724 288 1805 304
rect 1612 259 1668 279
rect 1562 243 1668 259
rect 1423 222 1514 238
rect 1343 161 1373 183
rect 1423 161 1453 222
rect 742 63 772 89
rect 921 85 987 101
rect 82 29 112 55
rect 921 51 937 85
rect 971 51 987 85
rect 1638 131 1668 243
rect 1724 254 1755 288
rect 1789 254 1805 288
rect 1724 238 1805 254
rect 1724 131 1754 238
rect 1862 213 1912 341
rect 1999 495 2082 511
rect 1999 461 2032 495
rect 2066 461 2082 495
rect 1999 445 2082 461
rect 1999 213 2029 445
rect 2214 397 2244 419
rect 2071 367 2244 397
rect 2071 356 2198 367
rect 2071 322 2087 356
rect 2121 322 2198 356
rect 2300 325 2330 419
rect 2615 511 2645 537
rect 2687 511 2717 537
rect 2792 511 2822 537
rect 2615 347 2645 427
rect 2405 325 2455 347
rect 2071 306 2198 322
rect 1862 183 2029 213
rect 1810 153 1912 183
rect 1810 131 1840 153
rect 1882 131 1912 153
rect 2168 181 2198 306
rect 2246 309 2455 325
rect 2246 275 2262 309
rect 2296 275 2455 309
rect 2563 331 2645 347
rect 2563 297 2579 331
rect 2613 311 2645 331
rect 2687 311 2717 427
rect 3064 427 3094 463
rect 2999 411 3108 427
rect 2999 377 3058 411
rect 3092 377 3108 411
rect 2999 361 3108 377
rect 2613 297 2717 311
rect 2563 281 2717 297
rect 2792 313 2822 343
rect 2792 283 2879 313
rect 2246 233 2455 275
rect 2687 235 2717 281
rect 2811 275 2879 283
rect 2811 241 2827 275
rect 2861 255 2879 275
rect 2861 241 2951 255
rect 2246 203 2558 233
rect 2687 205 2763 235
rect 2811 225 2951 241
rect 2246 181 2276 203
rect 2318 181 2348 203
rect 2450 181 2480 203
rect 2528 181 2558 203
rect 2733 183 2763 205
rect 2849 183 2879 225
rect 2921 183 2951 225
rect 2999 183 3029 361
rect 3150 313 3180 463
rect 3085 283 3180 313
rect 3236 313 3266 463
rect 3429 407 3459 491
rect 3335 377 3459 407
rect 3335 313 3365 377
rect 3536 329 3566 367
rect 3236 297 3365 313
rect 3085 183 3115 283
rect 3236 263 3312 297
rect 3346 263 3365 297
rect 3459 313 3566 329
rect 3459 279 3475 313
rect 3509 279 3566 313
rect 3459 263 3566 279
rect 3236 235 3365 263
rect 3163 229 3365 235
rect 3163 205 3312 229
rect 3163 183 3193 205
rect 3296 195 3312 205
rect 3346 209 3365 229
rect 3534 225 3564 263
rect 3346 195 3455 209
rect 1343 51 1373 77
rect 1423 51 1453 77
rect 921 35 987 51
rect 2168 71 2198 97
rect 2246 71 2276 97
rect 2318 71 2348 97
rect 1638 21 1668 47
rect 1724 21 1754 47
rect 1810 21 1840 47
rect 1882 21 1912 47
rect 2450 71 2480 97
rect 2528 71 2558 97
rect 3296 179 3455 195
rect 3425 141 3455 179
rect 2849 73 2879 99
rect 2921 73 2951 99
rect 2999 73 3029 99
rect 3085 73 3115 99
rect 3163 73 3193 99
rect 2733 29 2763 55
rect 3425 31 3455 57
rect 3534 31 3564 57
<< polycont >>
rect 133 303 167 337
rect 411 405 445 439
rect 527 405 561 439
rect 311 291 345 325
rect 133 235 167 269
rect 527 337 561 371
rect 1026 337 1060 371
rect 1247 337 1281 371
rect 1464 238 1498 272
rect 1578 259 1612 293
rect 937 51 971 85
rect 1755 254 1789 288
rect 2032 461 2066 495
rect 2087 322 2121 356
rect 2262 275 2296 309
rect 2579 297 2613 331
rect 3058 377 3092 411
rect 2827 241 2861 275
rect 3312 263 3346 297
rect 3475 279 3509 313
rect 3312 195 3346 229
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3648 683
rect 21 568 122 615
rect 21 534 72 568
rect 106 534 122 568
rect 21 424 122 534
rect 156 607 222 649
rect 156 573 172 607
rect 206 573 222 607
rect 156 537 222 573
rect 156 503 172 537
rect 206 503 222 537
rect 156 487 222 503
rect 320 569 386 615
rect 320 535 336 569
rect 370 535 386 569
rect 534 607 584 649
rect 534 573 550 607
rect 534 557 584 573
rect 618 581 823 615
rect 320 523 386 535
rect 618 523 652 581
rect 320 489 652 523
rect 697 498 747 547
rect 395 439 461 455
rect 395 424 411 439
rect 21 405 411 424
rect 445 405 461 439
rect 21 390 461 405
rect 21 114 71 390
rect 395 389 461 390
rect 505 439 574 455
rect 505 405 527 439
rect 561 405 574 439
rect 505 371 574 405
rect 117 337 183 356
rect 117 303 133 337
rect 167 303 183 337
rect 117 269 183 303
rect 117 235 133 269
rect 167 235 183 269
rect 217 325 361 356
rect 217 291 311 325
rect 345 291 361 325
rect 505 337 527 371
rect 561 337 574 371
rect 505 321 574 337
rect 217 236 361 291
rect 608 287 642 489
rect 731 464 747 498
rect 697 424 747 464
rect 697 390 703 424
rect 737 390 747 424
rect 697 319 747 390
rect 789 381 823 581
rect 857 535 891 649
rect 1042 581 1449 615
rect 857 465 891 501
rect 857 415 891 431
rect 927 503 993 551
rect 927 469 943 503
rect 977 469 993 503
rect 927 421 993 469
rect 927 381 961 421
rect 1042 387 1076 581
rect 789 347 961 381
rect 395 253 642 287
rect 676 303 747 319
rect 710 269 747 303
rect 676 253 747 269
rect 927 287 961 347
rect 1010 371 1076 387
rect 1010 337 1026 371
rect 1060 337 1076 371
rect 1010 321 1076 337
rect 1110 498 1197 547
rect 1415 504 1449 581
rect 1483 593 1607 615
rect 1517 572 1607 593
rect 1517 559 1567 572
rect 1483 538 1567 559
rect 1601 538 1607 572
rect 1657 588 1848 604
rect 1657 572 1798 588
rect 1657 538 1663 572
rect 1697 554 1798 572
rect 1832 554 1848 588
rect 2169 581 2410 615
rect 1697 538 1848 554
rect 1882 545 2135 579
rect 1882 504 1916 545
rect 1110 464 1147 498
rect 1181 464 1381 498
rect 1415 470 1916 504
rect 2016 495 2067 511
rect 1110 289 1197 464
rect 1347 436 1381 464
rect 2016 461 2032 495
rect 2066 461 2067 495
rect 2016 436 2067 461
rect 1347 430 2067 436
rect 1231 424 1313 430
rect 1231 390 1279 424
rect 1347 396 1587 430
rect 1621 402 2067 430
rect 2101 436 2135 545
rect 2169 527 2203 581
rect 2329 572 2410 581
rect 2169 470 2203 493
rect 2239 498 2289 547
rect 2239 464 2255 498
rect 2239 436 2289 464
rect 2329 538 2335 572
rect 2369 538 2410 572
rect 2554 581 3053 615
rect 2329 521 2410 538
rect 2329 487 2360 521
rect 2394 487 2410 521
rect 2329 458 2410 487
rect 2450 535 2516 551
rect 2450 501 2466 535
rect 2500 501 2516 535
rect 2450 464 2516 501
rect 2101 424 2289 436
rect 2450 430 2466 464
rect 2500 430 2516 464
rect 2554 499 2620 581
rect 2554 465 2570 499
rect 2604 465 2620 499
rect 2554 449 2620 465
rect 2731 513 2985 547
rect 2731 499 2781 513
rect 2731 465 2747 499
rect 2101 402 2416 424
rect 1621 396 1637 402
rect 1347 390 1637 396
rect 1231 371 1313 390
rect 1231 337 1247 371
rect 1281 337 1313 371
rect 1231 321 1313 337
rect 1380 322 1628 356
rect 927 253 1076 287
rect 1110 255 1126 289
rect 1160 255 1197 289
rect 1268 266 1334 287
rect 117 219 183 235
rect 395 185 429 253
rect 1042 221 1076 253
rect 1268 232 1284 266
rect 1318 232 1334 266
rect 1268 221 1334 232
rect 214 156 264 185
rect 21 80 37 114
rect 21 51 71 80
rect 107 114 173 143
rect 107 80 123 114
rect 157 80 173 114
rect 107 17 173 80
rect 214 122 230 156
rect 214 85 264 122
rect 300 169 429 185
rect 300 135 316 169
rect 350 135 429 169
rect 300 119 429 135
rect 480 185 940 219
rect 1042 187 1334 221
rect 480 169 514 185
rect 874 182 940 185
rect 480 119 514 135
rect 550 147 616 151
rect 550 113 566 147
rect 600 113 616 147
rect 550 85 616 113
rect 214 51 616 85
rect 767 135 833 151
rect 767 101 783 135
rect 817 101 833 135
rect 874 148 890 182
rect 924 148 940 182
rect 874 119 940 148
rect 1003 119 1019 153
rect 1053 119 1296 153
rect 1330 119 1346 153
rect 767 17 833 101
rect 1380 85 1414 322
rect 1561 293 1628 322
rect 1448 272 1514 288
rect 1448 238 1464 272
rect 1498 238 1514 272
rect 1561 259 1578 293
rect 1612 259 1628 293
rect 1561 243 1628 259
rect 1671 334 1942 368
rect 1976 334 1992 368
rect 1448 209 1514 238
rect 1671 209 1705 334
rect 1926 318 1992 334
rect 2041 356 2137 368
rect 2041 322 2087 356
rect 2121 322 2137 356
rect 2041 311 2137 322
rect 1739 288 1805 300
rect 1739 254 1755 288
rect 1789 277 1805 288
rect 1789 254 2041 277
rect 1739 243 2041 254
rect 2171 253 2205 402
rect 2239 390 2416 402
rect 2239 309 2312 356
rect 2239 275 2262 309
rect 2296 275 2312 309
rect 2382 309 2416 390
rect 2450 415 2516 430
rect 2450 393 2697 415
rect 2450 359 2466 393
rect 2500 381 2697 393
rect 2500 359 2516 381
rect 2450 343 2516 359
rect 2550 331 2629 347
rect 2550 309 2579 331
rect 2382 297 2579 309
rect 2613 297 2629 331
rect 2382 275 2629 297
rect 2239 259 2312 275
rect 1448 175 1973 209
rect 921 51 937 85
rect 971 51 1414 85
rect 1448 124 1729 141
rect 1448 90 1464 124
rect 1498 110 1729 124
rect 1498 107 1679 110
rect 1498 90 1514 107
rect 1448 73 1514 90
rect 1663 76 1679 107
rect 1713 76 1729 110
rect 1556 39 1572 73
rect 1606 39 1622 73
rect 1663 51 1729 76
rect 1765 106 1815 135
rect 1799 72 1815 106
rect 1556 17 1622 39
rect 1765 17 1815 72
rect 1907 110 1973 175
rect 2007 153 2041 243
rect 2084 237 2205 253
rect 2084 203 2100 237
rect 2134 203 2205 237
rect 2663 225 2697 381
rect 2084 187 2205 203
rect 2239 191 2697 225
rect 2731 389 2781 465
rect 2883 463 2917 479
rect 2731 355 2747 389
rect 2731 191 2781 355
rect 2815 424 2849 430
rect 2815 291 2849 390
rect 2883 389 2917 429
rect 2951 427 2985 513
rect 3019 523 3053 581
rect 3019 461 3053 489
rect 3089 523 3139 649
rect 3089 489 3105 523
rect 3089 461 3139 489
rect 3175 522 3241 551
rect 3175 488 3191 522
rect 3225 488 3241 522
rect 3175 427 3241 488
rect 3277 522 3327 649
rect 3311 488 3327 522
rect 3277 459 3327 488
rect 3368 568 3434 615
rect 3368 534 3384 568
rect 3418 534 3434 568
rect 3368 487 3434 534
rect 2951 393 3008 427
rect 2917 355 2940 359
rect 2883 325 2940 355
rect 2815 275 2872 291
rect 2815 241 2827 275
rect 2861 241 2872 275
rect 2815 225 2872 241
rect 2239 153 2273 191
rect 2553 169 2619 191
rect 2007 119 2273 153
rect 2307 123 2519 157
rect 1907 76 1923 110
rect 1957 85 1973 110
rect 2307 85 2341 123
rect 1957 76 2341 85
rect 1907 51 2341 76
rect 2382 73 2432 89
rect 2416 39 2432 73
rect 2485 85 2519 123
rect 2553 135 2569 169
rect 2603 135 2619 169
rect 2731 170 2831 191
rect 2731 157 2781 170
rect 2553 119 2619 135
rect 2765 136 2781 157
rect 2815 136 2831 170
rect 2665 104 2731 123
rect 2765 119 2831 136
rect 2665 85 2681 104
rect 2485 70 2681 85
rect 2715 85 2731 104
rect 2906 85 2940 325
rect 2974 255 3008 393
rect 3042 411 3241 427
rect 3042 377 3058 411
rect 3092 377 3241 411
rect 3042 361 3241 377
rect 2974 221 3158 255
rect 2715 70 2940 85
rect 2485 51 2940 70
rect 3024 158 3090 187
rect 3024 124 3040 158
rect 3074 124 3090 158
rect 2382 17 2432 39
rect 3024 17 3090 124
rect 3124 85 3158 221
rect 3207 187 3241 361
rect 3396 329 3434 487
rect 3475 607 3525 649
rect 3475 573 3491 607
rect 3475 510 3525 573
rect 3475 476 3491 510
rect 3475 413 3525 476
rect 3475 379 3491 413
rect 3475 363 3525 379
rect 3559 599 3627 615
rect 3559 565 3577 599
rect 3611 565 3627 599
rect 3559 506 3627 565
rect 3559 472 3577 506
rect 3611 472 3627 506
rect 3559 413 3627 472
rect 3559 379 3577 413
rect 3611 379 3627 413
rect 3396 313 3525 329
rect 3296 297 3362 313
rect 3296 263 3312 297
rect 3346 263 3362 297
rect 3296 229 3362 263
rect 3296 195 3312 229
rect 3346 195 3362 229
rect 3207 170 3261 187
rect 3207 136 3227 170
rect 3207 119 3261 136
rect 3296 179 3362 195
rect 3396 279 3475 313
rect 3509 279 3525 313
rect 3396 263 3525 279
rect 3296 85 3330 179
rect 3396 145 3430 263
rect 3124 51 3330 85
rect 3364 116 3430 145
rect 3364 82 3380 116
rect 3414 82 3430 116
rect 3364 53 3430 82
rect 3473 213 3523 229
rect 3473 179 3489 213
rect 3473 103 3523 179
rect 3473 69 3489 103
rect 3473 17 3523 69
rect 3559 213 3627 379
rect 3559 179 3575 213
rect 3609 179 3627 213
rect 3559 103 3627 179
rect 3559 69 3575 103
rect 3609 69 3627 103
rect 3559 53 3627 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3648 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 3583 649 3617 683
rect 703 390 737 424
rect 1567 538 1601 572
rect 1663 538 1697 572
rect 1279 390 1313 424
rect 2335 538 2369 572
rect 2815 390 2849 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
<< metal1 >>
rect 0 683 3648 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3648 683
rect 0 617 3648 649
rect 14 572 3634 589
rect 14 538 1567 572
rect 1601 538 1663 572
rect 1697 538 2335 572
rect 2369 538 3634 572
rect 14 535 3634 538
rect 1555 532 1613 535
rect 1651 532 1709 535
rect 2323 532 2381 535
rect 691 424 749 430
rect 691 390 703 424
rect 737 421 749 424
rect 1267 424 1325 430
rect 1267 421 1279 424
rect 737 393 1279 421
rect 737 390 749 393
rect 691 384 749 390
rect 1267 390 1279 393
rect 1313 421 1325 424
rect 2803 424 2861 430
rect 2803 421 2815 424
rect 1313 393 2815 421
rect 1313 390 1325 393
rect 1267 384 1325 390
rect 2803 390 2815 393
rect 2849 390 2861 424
rect 2803 384 2861 390
rect 0 17 3648 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3648 17
rect 0 -49 3648 -17
<< labels >>
flabel pwell s 0 0 3648 49 0 FreeSans 200 0 0 0 VNB
port 9 nsew ground bidirectional
flabel nwell s 0 617 3648 666 0 FreeSans 200 0 0 0 VPB
port 10 nsew power bidirectional
rlabel comment s 0 0 0 0 4 srsdfrtn_1
flabel metal1 s 14 535 3634 589 0 FreeSans 200 0 0 0 KAPWR
port 7 nsew power bidirectional
flabel metal1 s 0 617 3648 666 0 FreeSans 340 0 0 0 VPWR
port 11 nsew power bidirectional
flabel metal1 s 0 0 3648 49 0 FreeSans 340 0 0 0 VGND
port 8 nsew ground bidirectional
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 3583 94 3617 128 0 FreeSans 340 0 0 0 Q
port 12 nsew signal output
flabel locali s 3583 168 3617 202 0 FreeSans 340 0 0 0 Q
port 12 nsew signal output
flabel locali s 3583 242 3617 276 0 FreeSans 340 0 0 0 Q
port 12 nsew signal output
flabel locali s 3583 316 3617 350 0 FreeSans 340 0 0 0 Q
port 12 nsew signal output
flabel locali s 3583 390 3617 424 0 FreeSans 340 0 0 0 Q
port 12 nsew signal output
flabel locali s 2239 316 2273 350 0 FreeSans 340 0 0 0 SLEEP_B
port 6 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3648 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2632006
string GDS_START 2607980
<< end >>
