magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 463 243 957 259
rect 15 49 957 243
rect 0 0 960 49
<< scnmos >>
rect 94 49 124 217
rect 180 49 210 217
rect 266 49 296 217
rect 352 49 382 217
rect 542 65 572 233
rect 660 65 690 233
rect 746 65 776 233
rect 848 65 878 233
<< scpmoshvt >>
rect 94 367 124 619
rect 180 367 210 619
rect 266 367 296 619
rect 352 367 382 619
rect 574 367 604 619
rect 660 367 690 619
rect 746 367 776 619
rect 832 367 862 619
<< ndiff >>
rect 41 192 94 217
rect 41 158 49 192
rect 83 158 94 192
rect 41 95 94 158
rect 41 61 49 95
rect 83 61 94 95
rect 41 49 94 61
rect 124 199 180 217
rect 124 165 135 199
rect 169 165 180 199
rect 124 101 180 165
rect 124 67 135 101
rect 169 67 180 101
rect 124 49 180 67
rect 210 181 266 217
rect 210 147 221 181
rect 255 147 266 181
rect 210 95 266 147
rect 210 61 221 95
rect 255 61 266 95
rect 210 49 266 61
rect 296 205 352 217
rect 296 171 307 205
rect 341 171 352 205
rect 296 101 352 171
rect 296 67 307 101
rect 341 67 352 101
rect 296 49 352 67
rect 382 165 435 217
rect 382 131 393 165
rect 427 131 435 165
rect 382 95 435 131
rect 382 61 393 95
rect 427 61 435 95
rect 489 181 542 233
rect 489 147 497 181
rect 531 147 542 181
rect 489 111 542 147
rect 489 77 497 111
rect 531 77 542 111
rect 489 65 542 77
rect 572 107 660 233
rect 572 73 599 107
rect 633 73 660 107
rect 572 65 660 73
rect 690 181 746 233
rect 690 147 701 181
rect 735 147 746 181
rect 690 107 746 147
rect 690 73 701 107
rect 735 73 746 107
rect 690 65 746 73
rect 776 225 848 233
rect 776 191 803 225
rect 837 191 848 225
rect 776 153 848 191
rect 776 119 803 153
rect 837 119 848 153
rect 776 65 848 119
rect 878 192 931 233
rect 878 158 889 192
rect 923 158 931 192
rect 878 111 931 158
rect 878 77 889 111
rect 923 77 931 111
rect 878 65 931 77
rect 382 49 435 61
<< pdiff >>
rect 41 599 94 619
rect 41 565 49 599
rect 83 565 94 599
rect 41 515 94 565
rect 41 481 49 515
rect 83 481 94 515
rect 41 434 94 481
rect 41 400 49 434
rect 83 400 94 434
rect 41 367 94 400
rect 124 547 180 619
rect 124 513 135 547
rect 169 513 180 547
rect 124 479 180 513
rect 124 445 135 479
rect 169 445 180 479
rect 124 411 180 445
rect 124 377 135 411
rect 169 377 180 411
rect 124 367 180 377
rect 210 599 266 619
rect 210 565 221 599
rect 255 565 266 599
rect 210 514 266 565
rect 210 480 221 514
rect 255 480 266 514
rect 210 434 266 480
rect 210 400 221 434
rect 255 400 266 434
rect 210 367 266 400
rect 296 540 352 619
rect 296 506 307 540
rect 341 506 352 540
rect 296 436 352 506
rect 296 402 307 436
rect 341 402 352 436
rect 296 367 352 402
rect 382 599 435 619
rect 382 565 393 599
rect 427 565 435 599
rect 382 502 435 565
rect 382 468 393 502
rect 427 468 435 502
rect 382 367 435 468
rect 521 607 574 619
rect 521 573 529 607
rect 563 573 574 607
rect 521 493 574 573
rect 521 459 529 493
rect 563 459 574 493
rect 521 367 574 459
rect 604 599 660 619
rect 604 565 615 599
rect 649 565 660 599
rect 604 508 660 565
rect 604 474 615 508
rect 649 474 660 508
rect 604 413 660 474
rect 604 379 615 413
rect 649 379 660 413
rect 604 367 660 379
rect 690 607 746 619
rect 690 573 701 607
rect 735 573 746 607
rect 690 530 746 573
rect 690 496 701 530
rect 735 496 746 530
rect 690 455 746 496
rect 690 421 701 455
rect 735 421 746 455
rect 690 367 746 421
rect 776 599 832 619
rect 776 565 787 599
rect 821 565 832 599
rect 776 508 832 565
rect 776 474 787 508
rect 821 474 832 508
rect 776 413 832 474
rect 776 379 787 413
rect 821 379 832 413
rect 776 367 832 379
rect 862 607 915 619
rect 862 573 873 607
rect 907 573 915 607
rect 862 511 915 573
rect 862 477 873 511
rect 907 477 915 511
rect 862 418 915 477
rect 862 384 873 418
rect 907 384 915 418
rect 862 367 915 384
<< ndiffc >>
rect 49 158 83 192
rect 49 61 83 95
rect 135 165 169 199
rect 135 67 169 101
rect 221 147 255 181
rect 221 61 255 95
rect 307 171 341 205
rect 307 67 341 101
rect 393 131 427 165
rect 393 61 427 95
rect 497 147 531 181
rect 497 77 531 111
rect 599 73 633 107
rect 701 147 735 181
rect 701 73 735 107
rect 803 191 837 225
rect 803 119 837 153
rect 889 158 923 192
rect 889 77 923 111
<< pdiffc >>
rect 49 565 83 599
rect 49 481 83 515
rect 49 400 83 434
rect 135 513 169 547
rect 135 445 169 479
rect 135 377 169 411
rect 221 565 255 599
rect 221 480 255 514
rect 221 400 255 434
rect 307 506 341 540
rect 307 402 341 436
rect 393 565 427 599
rect 393 468 427 502
rect 529 573 563 607
rect 529 459 563 493
rect 615 565 649 599
rect 615 474 649 508
rect 615 379 649 413
rect 701 573 735 607
rect 701 496 735 530
rect 701 421 735 455
rect 787 565 821 599
rect 787 474 821 508
rect 787 379 821 413
rect 873 573 907 607
rect 873 477 907 511
rect 873 384 907 418
<< poly >>
rect 94 619 124 645
rect 180 619 210 645
rect 266 619 296 645
rect 352 619 382 645
rect 574 619 604 645
rect 660 619 690 645
rect 746 619 776 645
rect 832 619 862 645
rect 94 308 124 367
rect 180 308 210 367
rect 35 292 210 308
rect 35 258 51 292
rect 85 258 210 292
rect 35 242 210 258
rect 94 217 124 242
rect 180 217 210 242
rect 266 335 296 367
rect 352 335 382 367
rect 574 335 604 367
rect 660 335 690 367
rect 266 319 382 335
rect 266 285 307 319
rect 341 285 382 319
rect 266 269 382 285
rect 488 319 690 335
rect 488 285 504 319
rect 538 285 572 319
rect 606 285 640 319
rect 674 285 690 319
rect 488 269 690 285
rect 266 217 296 269
rect 352 217 382 269
rect 542 233 572 269
rect 660 233 690 269
rect 746 335 776 367
rect 832 335 862 367
rect 746 321 862 335
rect 746 319 939 321
rect 746 285 762 319
rect 796 305 939 319
rect 796 285 889 305
rect 746 271 889 285
rect 923 271 939 305
rect 746 255 939 271
rect 746 233 776 255
rect 848 233 878 255
rect 94 23 124 49
rect 180 23 210 49
rect 266 23 296 49
rect 352 23 382 49
rect 542 39 572 65
rect 660 39 690 65
rect 746 39 776 65
rect 848 39 878 65
<< polycont >>
rect 51 258 85 292
rect 307 285 341 319
rect 504 285 538 319
rect 572 285 606 319
rect 640 285 674 319
rect 762 285 796 319
rect 889 271 923 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 33 599 443 615
rect 33 565 49 599
rect 83 581 221 599
rect 83 565 85 581
rect 33 515 85 565
rect 219 565 221 581
rect 255 581 393 599
rect 255 565 257 581
rect 33 481 49 515
rect 83 481 85 515
rect 33 434 85 481
rect 33 400 49 434
rect 83 400 85 434
rect 33 384 85 400
rect 119 513 135 547
rect 169 513 185 547
rect 119 479 185 513
rect 119 445 135 479
rect 169 445 185 479
rect 119 411 185 445
rect 119 377 135 411
rect 169 377 185 411
rect 219 514 257 565
rect 391 565 393 581
rect 427 565 443 599
rect 219 480 221 514
rect 255 480 257 514
rect 219 434 257 480
rect 219 400 221 434
rect 255 400 257 434
rect 219 384 257 400
rect 291 540 357 547
rect 291 506 307 540
rect 341 506 357 540
rect 291 436 357 506
rect 391 502 443 565
rect 391 468 393 502
rect 427 468 443 502
rect 391 452 443 468
rect 513 607 579 649
rect 513 573 529 607
rect 563 573 579 607
rect 513 493 579 573
rect 513 459 529 493
rect 563 459 579 493
rect 513 452 579 459
rect 613 599 651 615
rect 613 565 615 599
rect 649 565 651 599
rect 613 508 651 565
rect 613 474 615 508
rect 649 474 651 508
rect 291 402 307 436
rect 341 418 357 436
rect 613 418 651 474
rect 685 607 751 649
rect 685 573 701 607
rect 735 573 751 607
rect 685 530 751 573
rect 685 496 701 530
rect 735 496 751 530
rect 685 455 751 496
rect 685 421 701 455
rect 735 421 751 455
rect 785 599 823 615
rect 785 565 787 599
rect 821 565 823 599
rect 785 508 823 565
rect 785 474 787 508
rect 821 474 823 508
rect 341 413 651 418
rect 341 402 615 413
rect 291 384 615 402
rect 17 292 85 350
rect 17 258 51 292
rect 17 242 85 258
rect 119 249 185 377
rect 613 379 615 384
rect 649 387 651 413
rect 785 413 823 474
rect 785 387 787 413
rect 649 379 787 387
rect 821 379 823 413
rect 857 607 923 649
rect 857 573 873 607
rect 907 573 923 607
rect 857 511 923 573
rect 857 477 873 511
rect 907 477 923 511
rect 857 418 923 477
rect 857 384 873 418
rect 907 384 923 418
rect 613 353 823 379
rect 223 319 367 350
rect 223 285 307 319
rect 341 285 367 319
rect 401 319 579 350
rect 889 319 943 350
rect 401 285 504 319
rect 538 285 572 319
rect 606 285 640 319
rect 674 285 690 319
rect 401 283 690 285
rect 746 285 762 319
rect 796 305 943 319
rect 796 285 889 305
rect 746 283 889 285
rect 923 271 943 305
rect 119 225 853 249
rect 889 242 943 271
rect 119 215 803 225
rect 33 192 85 208
rect 33 158 49 192
rect 83 158 85 192
rect 33 95 85 158
rect 33 61 49 95
rect 83 61 85 95
rect 33 17 85 61
rect 119 199 171 215
rect 119 165 135 199
rect 169 165 171 199
rect 305 205 353 215
rect 119 101 171 165
rect 119 67 135 101
rect 169 67 171 101
rect 119 51 171 67
rect 205 147 221 181
rect 255 147 271 181
rect 205 95 271 147
rect 205 61 221 95
rect 255 61 271 95
rect 205 17 271 61
rect 305 171 307 205
rect 341 171 353 205
rect 787 191 803 215
rect 837 191 853 225
rect 305 101 353 171
rect 305 67 307 101
rect 341 67 353 101
rect 305 51 353 67
rect 387 165 443 181
rect 387 131 393 165
rect 427 131 443 165
rect 387 95 443 131
rect 387 61 393 95
rect 427 61 443 95
rect 481 147 497 181
rect 531 147 701 181
rect 735 147 751 181
rect 481 111 547 147
rect 481 77 497 111
rect 531 77 547 111
rect 481 61 547 77
rect 583 107 649 113
rect 583 73 599 107
rect 633 73 649 107
rect 387 17 443 61
rect 583 17 649 73
rect 685 107 751 147
rect 787 153 853 191
rect 787 119 803 153
rect 837 119 853 153
rect 887 192 939 208
rect 887 158 889 192
rect 923 158 939 192
rect 685 73 701 107
rect 735 85 751 107
rect 887 111 939 158
rect 887 85 889 111
rect 735 77 889 85
rect 923 77 939 111
rect 735 73 939 77
rect 685 51 939 73
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a211oi_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 222962
string GDS_START 213704
<< end >>
