magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 9 49 2015 259
rect 0 0 2016 49
<< scnmos >>
rect 88 65 118 233
rect 174 65 204 233
rect 260 65 290 233
rect 346 65 376 233
rect 432 65 462 233
rect 518 65 548 233
rect 604 65 634 233
rect 706 65 736 233
rect 804 65 834 233
rect 894 65 924 233
rect 996 65 1026 233
rect 1098 65 1128 233
rect 1288 65 1318 233
rect 1374 65 1404 233
rect 1460 65 1490 233
rect 1546 65 1576 233
rect 1632 65 1662 233
rect 1718 65 1748 233
rect 1804 65 1834 233
rect 1890 65 1920 233
<< scpmoshvt >>
rect 102 367 132 619
rect 188 367 218 619
rect 274 367 304 619
rect 366 367 396 619
rect 452 367 482 619
rect 538 367 568 619
rect 624 367 654 619
rect 710 367 740 619
rect 804 367 834 619
rect 890 367 920 619
rect 976 367 1006 619
rect 1062 367 1092 619
rect 1217 367 1247 619
rect 1303 367 1333 619
rect 1389 367 1419 619
rect 1475 367 1505 619
rect 1629 367 1659 619
rect 1715 367 1745 619
rect 1801 367 1831 619
rect 1887 367 1917 619
<< ndiff >>
rect 35 221 88 233
rect 35 187 43 221
rect 77 187 88 221
rect 35 111 88 187
rect 35 77 43 111
rect 77 77 88 111
rect 35 65 88 77
rect 118 177 174 233
rect 118 143 129 177
rect 163 143 174 177
rect 118 107 174 143
rect 118 73 129 107
rect 163 73 174 107
rect 118 65 174 73
rect 204 225 260 233
rect 204 191 215 225
rect 249 191 260 225
rect 204 111 260 191
rect 204 77 215 111
rect 249 77 260 111
rect 204 65 260 77
rect 290 177 346 233
rect 290 143 301 177
rect 335 143 346 177
rect 290 107 346 143
rect 290 73 301 107
rect 335 73 346 107
rect 290 65 346 73
rect 376 221 432 233
rect 376 187 387 221
rect 421 187 432 221
rect 376 111 432 187
rect 376 77 387 111
rect 421 77 432 111
rect 376 65 432 77
rect 462 177 518 233
rect 462 143 473 177
rect 507 143 518 177
rect 462 107 518 143
rect 462 73 473 107
rect 507 73 518 107
rect 462 65 518 73
rect 548 221 604 233
rect 548 187 559 221
rect 593 187 604 221
rect 548 111 604 187
rect 548 77 559 111
rect 593 77 604 111
rect 548 65 604 77
rect 634 180 706 233
rect 634 146 645 180
rect 679 146 706 180
rect 634 107 706 146
rect 634 73 645 107
rect 679 73 706 107
rect 634 65 706 73
rect 736 175 804 233
rect 736 141 747 175
rect 781 141 804 175
rect 736 107 804 141
rect 736 73 747 107
rect 781 73 804 107
rect 736 65 804 73
rect 834 225 894 233
rect 834 191 849 225
rect 883 191 894 225
rect 834 157 894 191
rect 834 123 849 157
rect 883 123 894 157
rect 834 65 894 123
rect 924 175 996 233
rect 924 141 951 175
rect 985 141 996 175
rect 924 107 996 141
rect 924 73 951 107
rect 985 73 996 107
rect 924 65 996 73
rect 1026 225 1098 233
rect 1026 191 1053 225
rect 1087 191 1098 225
rect 1026 157 1098 191
rect 1026 123 1053 157
rect 1087 123 1098 157
rect 1026 65 1098 123
rect 1128 192 1181 233
rect 1128 158 1139 192
rect 1173 158 1181 192
rect 1128 111 1181 158
rect 1128 77 1139 111
rect 1173 77 1181 111
rect 1128 65 1181 77
rect 1235 208 1288 233
rect 1235 174 1243 208
rect 1277 174 1288 208
rect 1235 111 1288 174
rect 1235 77 1243 111
rect 1277 77 1288 111
rect 1235 65 1288 77
rect 1318 133 1374 233
rect 1318 99 1329 133
rect 1363 99 1374 133
rect 1318 65 1374 99
rect 1404 221 1460 233
rect 1404 187 1415 221
rect 1449 187 1460 221
rect 1404 111 1460 187
rect 1404 77 1415 111
rect 1449 77 1460 111
rect 1404 65 1460 77
rect 1490 179 1546 233
rect 1490 145 1501 179
rect 1535 145 1546 179
rect 1490 107 1546 145
rect 1490 73 1501 107
rect 1535 73 1546 107
rect 1490 65 1546 73
rect 1576 225 1632 233
rect 1576 191 1587 225
rect 1621 191 1632 225
rect 1576 111 1632 191
rect 1576 77 1587 111
rect 1621 77 1632 111
rect 1576 65 1632 77
rect 1662 171 1718 233
rect 1662 137 1673 171
rect 1707 137 1718 171
rect 1662 65 1718 137
rect 1748 111 1804 233
rect 1748 77 1759 111
rect 1793 77 1804 111
rect 1748 65 1804 77
rect 1834 225 1890 233
rect 1834 191 1845 225
rect 1879 191 1890 225
rect 1834 157 1890 191
rect 1834 123 1845 157
rect 1879 123 1890 157
rect 1834 65 1890 123
rect 1920 179 1989 233
rect 1920 145 1947 179
rect 1981 145 1989 179
rect 1920 111 1989 145
rect 1920 77 1947 111
rect 1981 77 1989 111
rect 1920 65 1989 77
<< pdiff >>
rect 49 607 102 619
rect 49 573 57 607
rect 91 573 102 607
rect 49 504 102 573
rect 49 470 57 504
rect 91 470 102 504
rect 49 413 102 470
rect 49 379 57 413
rect 91 379 102 413
rect 49 367 102 379
rect 132 599 188 619
rect 132 565 143 599
rect 177 565 188 599
rect 132 504 188 565
rect 132 470 143 504
rect 177 470 188 504
rect 132 413 188 470
rect 132 379 143 413
rect 177 379 188 413
rect 132 367 188 379
rect 218 580 274 619
rect 218 546 229 580
rect 263 546 274 580
rect 218 367 274 546
rect 304 599 366 619
rect 304 565 319 599
rect 353 565 366 599
rect 304 520 366 565
rect 304 486 319 520
rect 353 486 366 520
rect 304 367 366 486
rect 396 510 452 619
rect 396 476 407 510
rect 441 476 452 510
rect 396 367 452 476
rect 482 600 538 619
rect 482 566 493 600
rect 527 566 538 600
rect 482 367 538 566
rect 568 510 624 619
rect 568 476 579 510
rect 613 476 624 510
rect 568 367 624 476
rect 654 600 710 619
rect 654 566 665 600
rect 699 566 710 600
rect 654 367 710 566
rect 740 610 804 619
rect 740 576 759 610
rect 793 576 804 610
rect 740 367 804 576
rect 834 599 890 619
rect 834 565 845 599
rect 879 565 890 599
rect 834 505 890 565
rect 834 471 845 505
rect 879 471 890 505
rect 834 413 890 471
rect 834 379 845 413
rect 879 379 890 413
rect 834 367 890 379
rect 920 611 976 619
rect 920 577 931 611
rect 965 577 976 611
rect 920 534 976 577
rect 920 500 931 534
rect 965 500 976 534
rect 920 459 976 500
rect 920 425 931 459
rect 965 425 976 459
rect 920 367 976 425
rect 1006 599 1062 619
rect 1006 565 1017 599
rect 1051 565 1062 599
rect 1006 505 1062 565
rect 1006 471 1017 505
rect 1051 471 1062 505
rect 1006 413 1062 471
rect 1006 379 1017 413
rect 1051 379 1062 413
rect 1006 367 1062 379
rect 1092 611 1217 619
rect 1092 577 1103 611
rect 1137 577 1172 611
rect 1206 577 1217 611
rect 1092 534 1217 577
rect 1092 500 1103 534
rect 1137 500 1172 534
rect 1206 500 1217 534
rect 1092 459 1217 500
rect 1092 425 1103 459
rect 1137 425 1172 459
rect 1206 425 1217 459
rect 1092 367 1217 425
rect 1247 599 1303 619
rect 1247 565 1258 599
rect 1292 565 1303 599
rect 1247 505 1303 565
rect 1247 471 1258 505
rect 1292 471 1303 505
rect 1247 413 1303 471
rect 1247 379 1258 413
rect 1292 379 1303 413
rect 1247 367 1303 379
rect 1333 611 1389 619
rect 1333 577 1344 611
rect 1378 577 1389 611
rect 1333 534 1389 577
rect 1333 500 1344 534
rect 1378 500 1389 534
rect 1333 459 1389 500
rect 1333 425 1344 459
rect 1378 425 1389 459
rect 1333 367 1389 425
rect 1419 599 1475 619
rect 1419 565 1430 599
rect 1464 565 1475 599
rect 1419 505 1475 565
rect 1419 471 1430 505
rect 1464 471 1475 505
rect 1419 413 1475 471
rect 1419 379 1430 413
rect 1464 379 1475 413
rect 1419 367 1475 379
rect 1505 611 1629 619
rect 1505 577 1516 611
rect 1550 577 1584 611
rect 1618 577 1629 611
rect 1505 534 1629 577
rect 1505 500 1516 534
rect 1550 500 1584 534
rect 1618 500 1629 534
rect 1505 459 1629 500
rect 1505 425 1516 459
rect 1550 425 1584 459
rect 1618 425 1629 459
rect 1505 367 1629 425
rect 1659 599 1715 619
rect 1659 565 1670 599
rect 1704 565 1715 599
rect 1659 505 1715 565
rect 1659 471 1670 505
rect 1704 471 1715 505
rect 1659 413 1715 471
rect 1659 379 1670 413
rect 1704 379 1715 413
rect 1659 367 1715 379
rect 1745 611 1801 619
rect 1745 577 1756 611
rect 1790 577 1801 611
rect 1745 534 1801 577
rect 1745 500 1756 534
rect 1790 500 1801 534
rect 1745 459 1801 500
rect 1745 425 1756 459
rect 1790 425 1801 459
rect 1745 367 1801 425
rect 1831 599 1887 619
rect 1831 565 1842 599
rect 1876 565 1887 599
rect 1831 505 1887 565
rect 1831 471 1842 505
rect 1876 471 1887 505
rect 1831 413 1887 471
rect 1831 379 1842 413
rect 1876 379 1887 413
rect 1831 367 1887 379
rect 1917 607 1970 619
rect 1917 573 1928 607
rect 1962 573 1970 607
rect 1917 534 1970 573
rect 1917 500 1928 534
rect 1962 500 1970 534
rect 1917 457 1970 500
rect 1917 423 1928 457
rect 1962 423 1970 457
rect 1917 367 1970 423
<< ndiffc >>
rect 43 187 77 221
rect 43 77 77 111
rect 129 143 163 177
rect 129 73 163 107
rect 215 191 249 225
rect 215 77 249 111
rect 301 143 335 177
rect 301 73 335 107
rect 387 187 421 221
rect 387 77 421 111
rect 473 143 507 177
rect 473 73 507 107
rect 559 187 593 221
rect 559 77 593 111
rect 645 146 679 180
rect 645 73 679 107
rect 747 141 781 175
rect 747 73 781 107
rect 849 191 883 225
rect 849 123 883 157
rect 951 141 985 175
rect 951 73 985 107
rect 1053 191 1087 225
rect 1053 123 1087 157
rect 1139 158 1173 192
rect 1139 77 1173 111
rect 1243 174 1277 208
rect 1243 77 1277 111
rect 1329 99 1363 133
rect 1415 187 1449 221
rect 1415 77 1449 111
rect 1501 145 1535 179
rect 1501 73 1535 107
rect 1587 191 1621 225
rect 1587 77 1621 111
rect 1673 137 1707 171
rect 1759 77 1793 111
rect 1845 191 1879 225
rect 1845 123 1879 157
rect 1947 145 1981 179
rect 1947 77 1981 111
<< pdiffc >>
rect 57 573 91 607
rect 57 470 91 504
rect 57 379 91 413
rect 143 565 177 599
rect 143 470 177 504
rect 143 379 177 413
rect 229 546 263 580
rect 319 565 353 599
rect 319 486 353 520
rect 407 476 441 510
rect 493 566 527 600
rect 579 476 613 510
rect 665 566 699 600
rect 759 576 793 610
rect 845 565 879 599
rect 845 471 879 505
rect 845 379 879 413
rect 931 577 965 611
rect 931 500 965 534
rect 931 425 965 459
rect 1017 565 1051 599
rect 1017 471 1051 505
rect 1017 379 1051 413
rect 1103 577 1137 611
rect 1172 577 1206 611
rect 1103 500 1137 534
rect 1172 500 1206 534
rect 1103 425 1137 459
rect 1172 425 1206 459
rect 1258 565 1292 599
rect 1258 471 1292 505
rect 1258 379 1292 413
rect 1344 577 1378 611
rect 1344 500 1378 534
rect 1344 425 1378 459
rect 1430 565 1464 599
rect 1430 471 1464 505
rect 1430 379 1464 413
rect 1516 577 1550 611
rect 1584 577 1618 611
rect 1516 500 1550 534
rect 1584 500 1618 534
rect 1516 425 1550 459
rect 1584 425 1618 459
rect 1670 565 1704 599
rect 1670 471 1704 505
rect 1670 379 1704 413
rect 1756 577 1790 611
rect 1756 500 1790 534
rect 1756 425 1790 459
rect 1842 565 1876 599
rect 1842 471 1876 505
rect 1842 379 1876 413
rect 1928 573 1962 607
rect 1928 500 1962 534
rect 1928 423 1962 457
<< poly >>
rect 102 619 132 645
rect 188 619 218 645
rect 274 619 304 645
rect 366 619 396 645
rect 452 619 482 645
rect 538 619 568 645
rect 624 619 654 645
rect 710 619 740 645
rect 804 619 834 645
rect 890 619 920 645
rect 976 619 1006 645
rect 1062 619 1092 645
rect 1217 619 1247 645
rect 1303 619 1333 645
rect 1389 619 1419 645
rect 1475 619 1505 645
rect 1629 619 1659 645
rect 1715 619 1745 645
rect 1801 619 1831 645
rect 1887 619 1917 645
rect 102 335 132 367
rect 188 335 218 367
rect 274 335 304 367
rect 366 335 396 367
rect 452 335 482 367
rect 538 335 568 367
rect 624 335 654 367
rect 710 335 740 367
rect 804 335 834 367
rect 890 335 920 367
rect 976 335 1006 367
rect 1062 335 1092 367
rect 1217 335 1247 367
rect 1303 335 1333 367
rect 1389 335 1419 367
rect 1475 335 1505 367
rect 1629 345 1659 367
rect 1715 345 1745 367
rect 1801 345 1831 367
rect 1887 345 1917 367
rect 1629 335 1917 345
rect 81 319 304 335
rect 81 285 97 319
rect 131 285 165 319
rect 199 285 233 319
rect 267 285 304 319
rect 81 269 304 285
rect 346 319 654 335
rect 346 285 362 319
rect 396 285 430 319
rect 464 285 498 319
rect 532 285 566 319
rect 600 285 654 319
rect 346 269 654 285
rect 696 319 762 335
rect 696 285 712 319
rect 746 285 762 319
rect 88 233 118 269
rect 174 233 204 269
rect 260 233 290 269
rect 346 233 376 269
rect 432 233 462 269
rect 518 233 548 269
rect 604 233 634 269
rect 696 259 762 285
rect 804 319 1139 335
rect 804 285 885 319
rect 919 285 953 319
rect 987 285 1021 319
rect 1055 285 1089 319
rect 1123 285 1139 319
rect 804 269 1139 285
rect 1217 319 1587 335
rect 1217 285 1265 319
rect 1299 285 1333 319
rect 1367 285 1401 319
rect 1435 285 1469 319
rect 1503 285 1537 319
rect 1571 285 1587 319
rect 1629 319 1927 335
rect 1629 315 1673 319
rect 1217 269 1587 285
rect 1632 285 1673 315
rect 1707 285 1741 319
rect 1775 285 1809 319
rect 1843 285 1877 319
rect 1911 285 1927 319
rect 1632 269 1927 285
rect 706 233 736 259
rect 804 233 834 269
rect 894 233 924 269
rect 996 233 1026 269
rect 1098 233 1128 269
rect 1288 233 1318 269
rect 1374 233 1404 269
rect 1460 233 1490 269
rect 1546 233 1576 269
rect 1632 233 1662 269
rect 1718 233 1748 269
rect 1804 233 1834 269
rect 1890 233 1920 269
rect 88 39 118 65
rect 174 39 204 65
rect 260 39 290 65
rect 346 39 376 65
rect 432 39 462 65
rect 518 39 548 65
rect 604 39 634 65
rect 706 39 736 65
rect 804 39 834 65
rect 894 39 924 65
rect 996 39 1026 65
rect 1098 39 1128 65
rect 1288 39 1318 65
rect 1374 39 1404 65
rect 1460 39 1490 65
rect 1546 39 1576 65
rect 1632 39 1662 65
rect 1718 39 1748 65
rect 1804 39 1834 65
rect 1890 39 1920 65
<< polycont >>
rect 97 285 131 319
rect 165 285 199 319
rect 233 285 267 319
rect 362 285 396 319
rect 430 285 464 319
rect 498 285 532 319
rect 566 285 600 319
rect 712 285 746 319
rect 885 285 919 319
rect 953 285 987 319
rect 1021 285 1055 319
rect 1089 285 1123 319
rect 1265 285 1299 319
rect 1333 285 1367 319
rect 1401 285 1435 319
rect 1469 285 1503 319
rect 1537 285 1571 319
rect 1673 285 1707 319
rect 1741 285 1775 319
rect 1809 285 1843 319
rect 1877 285 1911 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 53 607 95 649
rect 53 573 57 607
rect 91 573 95 607
rect 53 504 95 573
rect 53 470 57 504
rect 91 470 95 504
rect 53 413 95 470
rect 53 379 57 413
rect 91 379 95 413
rect 53 363 95 379
rect 139 599 179 615
rect 139 565 143 599
rect 177 565 179 599
rect 139 504 179 565
rect 213 580 279 649
rect 213 546 229 580
rect 263 546 279 580
rect 213 538 279 546
rect 315 600 715 615
rect 315 599 493 600
rect 315 565 319 599
rect 353 566 493 599
rect 527 566 665 600
rect 699 566 715 600
rect 353 565 715 566
rect 315 560 715 565
rect 749 610 809 649
rect 749 576 759 610
rect 793 576 809 610
rect 749 560 809 576
rect 843 599 881 615
rect 843 565 845 599
rect 879 565 881 599
rect 315 520 357 560
rect 843 526 881 565
rect 315 504 319 520
rect 139 470 143 504
rect 177 486 319 504
rect 353 486 357 520
rect 177 470 357 486
rect 403 510 881 526
rect 403 476 407 510
rect 441 476 579 510
rect 613 505 881 510
rect 613 476 845 505
rect 403 471 845 476
rect 879 471 881 505
rect 139 413 177 470
rect 403 460 881 471
rect 139 379 143 413
rect 139 363 177 379
rect 211 390 762 426
rect 211 329 283 390
rect 81 319 283 329
rect 81 285 97 319
rect 131 285 165 319
rect 199 285 233 319
rect 267 285 283 319
rect 319 319 641 356
rect 319 285 362 319
rect 396 285 430 319
rect 464 285 498 319
rect 532 285 566 319
rect 600 285 641 319
rect 696 319 762 390
rect 696 285 712 319
rect 746 285 762 319
rect 799 413 881 460
rect 915 611 981 649
rect 915 577 931 611
rect 965 577 981 611
rect 915 534 981 577
rect 915 500 931 534
rect 965 500 981 534
rect 915 459 981 500
rect 915 425 931 459
rect 965 425 981 459
rect 915 423 981 425
rect 1015 599 1053 615
rect 1015 565 1017 599
rect 1051 565 1053 599
rect 1015 505 1053 565
rect 1015 471 1017 505
rect 1051 471 1053 505
rect 799 379 845 413
rect 879 389 881 413
rect 1015 413 1053 471
rect 1087 611 1222 649
rect 1087 577 1103 611
rect 1137 577 1172 611
rect 1206 577 1222 611
rect 1087 534 1222 577
rect 1087 500 1103 534
rect 1137 500 1172 534
rect 1206 500 1222 534
rect 1087 459 1222 500
rect 1087 425 1103 459
rect 1137 425 1172 459
rect 1206 425 1222 459
rect 1256 599 1294 615
rect 1256 565 1258 599
rect 1292 565 1294 599
rect 1256 505 1294 565
rect 1256 471 1258 505
rect 1292 471 1294 505
rect 1015 389 1017 413
rect 879 379 1017 389
rect 1051 379 1053 413
rect 1256 413 1294 471
rect 1328 611 1394 649
rect 1328 577 1344 611
rect 1378 577 1394 611
rect 1328 534 1394 577
rect 1328 500 1344 534
rect 1378 500 1394 534
rect 1328 459 1394 500
rect 1328 425 1344 459
rect 1378 425 1394 459
rect 1428 599 1466 615
rect 1428 565 1430 599
rect 1464 565 1466 599
rect 1428 505 1466 565
rect 1428 471 1430 505
rect 1464 471 1466 505
rect 1256 389 1258 413
rect 799 355 1053 379
rect 1111 379 1258 389
rect 1292 389 1294 413
rect 1428 413 1466 471
rect 1500 611 1634 649
rect 1500 577 1516 611
rect 1550 577 1584 611
rect 1618 577 1634 611
rect 1500 534 1634 577
rect 1500 500 1516 534
rect 1550 500 1584 534
rect 1618 500 1634 534
rect 1500 459 1634 500
rect 1500 425 1516 459
rect 1550 425 1584 459
rect 1618 425 1634 459
rect 1668 599 1706 615
rect 1668 565 1670 599
rect 1704 565 1706 599
rect 1668 505 1706 565
rect 1668 471 1670 505
rect 1704 471 1706 505
rect 1428 389 1430 413
rect 1292 379 1430 389
rect 1464 389 1466 413
rect 1668 413 1706 471
rect 1740 611 1806 649
rect 1740 577 1756 611
rect 1790 577 1806 611
rect 1740 534 1806 577
rect 1740 500 1756 534
rect 1790 500 1806 534
rect 1740 459 1806 500
rect 1740 425 1756 459
rect 1790 425 1806 459
rect 1842 599 1878 615
rect 1876 565 1878 599
rect 1842 505 1878 565
rect 1876 471 1878 505
rect 1668 389 1670 413
rect 1464 379 1670 389
rect 1704 389 1706 413
rect 1842 413 1878 471
rect 1912 607 1978 649
rect 1912 573 1928 607
rect 1962 573 1978 607
rect 1912 534 1978 573
rect 1912 500 1928 534
rect 1962 500 1978 534
rect 1912 457 1978 500
rect 1912 423 1928 457
rect 1962 423 1978 457
rect 1704 379 1842 389
rect 1876 389 1878 413
rect 1876 379 1999 389
rect 27 225 765 251
rect 27 221 215 225
rect 27 187 43 221
rect 77 215 215 221
rect 27 111 77 187
rect 213 191 215 215
rect 249 221 765 225
rect 249 215 387 221
rect 249 191 251 215
rect 27 77 43 111
rect 27 61 77 77
rect 113 177 179 181
rect 113 143 129 177
rect 163 143 179 177
rect 113 107 179 143
rect 113 73 129 107
rect 163 73 179 107
rect 113 17 179 73
rect 213 111 251 191
rect 385 187 387 215
rect 421 215 559 221
rect 421 187 423 215
rect 213 77 215 111
rect 249 77 251 111
rect 213 61 251 77
rect 285 177 351 181
rect 285 143 301 177
rect 335 143 351 177
rect 285 107 351 143
rect 285 73 301 107
rect 335 73 351 107
rect 285 17 351 73
rect 385 111 423 187
rect 557 187 559 215
rect 593 217 765 221
rect 593 187 595 217
rect 385 77 387 111
rect 421 77 423 111
rect 385 61 423 77
rect 457 177 523 181
rect 457 143 473 177
rect 507 143 523 177
rect 457 107 523 143
rect 457 73 473 107
rect 507 73 523 107
rect 457 17 523 73
rect 557 111 595 187
rect 557 77 559 111
rect 593 77 595 111
rect 557 61 595 77
rect 629 180 697 183
rect 629 146 645 180
rect 679 146 697 180
rect 629 107 697 146
rect 629 73 645 107
rect 679 73 697 107
rect 629 17 697 73
rect 731 181 765 217
rect 799 249 833 355
rect 1111 353 1999 379
rect 1111 319 1145 353
rect 869 285 885 319
rect 919 285 953 319
rect 987 285 1021 319
rect 1055 285 1089 319
rect 1123 285 1145 319
rect 1181 285 1265 319
rect 1299 285 1333 319
rect 1367 285 1401 319
rect 1435 285 1469 319
rect 1503 285 1537 319
rect 1571 285 1587 319
rect 1657 285 1673 319
rect 1707 285 1741 319
rect 1775 285 1809 319
rect 1843 285 1877 319
rect 1911 285 1927 319
rect 799 225 1103 249
rect 1181 242 1313 285
rect 799 215 849 225
rect 833 191 849 215
rect 883 215 1053 225
rect 883 191 899 215
rect 731 175 797 181
rect 731 141 747 175
rect 781 141 797 175
rect 731 107 797 141
rect 833 157 899 191
rect 1037 191 1053 215
rect 1087 191 1103 225
rect 1411 225 1623 249
rect 1657 234 1795 285
rect 1963 251 1999 353
rect 1411 221 1587 225
rect 1411 208 1415 221
rect 833 123 849 157
rect 883 123 899 157
rect 833 121 899 123
rect 935 175 1001 179
rect 935 141 951 175
rect 985 141 1001 175
rect 731 73 747 107
rect 781 87 797 107
rect 935 107 1001 141
rect 1037 157 1103 191
rect 1037 123 1053 157
rect 1087 123 1103 157
rect 1137 192 1189 208
rect 1137 158 1139 192
rect 1173 158 1189 192
rect 935 87 951 107
rect 781 73 951 87
rect 985 87 1001 107
rect 1137 111 1189 158
rect 1137 87 1139 111
rect 985 77 1139 87
rect 1173 77 1189 111
rect 985 73 1189 77
rect 731 53 1189 73
rect 1227 174 1243 208
rect 1277 187 1415 208
rect 1449 215 1587 221
rect 1449 187 1451 215
rect 1277 174 1451 187
rect 1585 191 1587 215
rect 1621 191 1623 225
rect 1829 225 1999 251
rect 1829 200 1845 225
rect 1227 111 1279 174
rect 1227 77 1243 111
rect 1277 77 1279 111
rect 1227 61 1279 77
rect 1313 133 1379 140
rect 1313 99 1329 133
rect 1363 99 1379 133
rect 1313 17 1379 99
rect 1413 111 1451 174
rect 1413 77 1415 111
rect 1449 77 1451 111
rect 1413 61 1451 77
rect 1485 179 1551 181
rect 1485 145 1501 179
rect 1535 145 1551 179
rect 1485 107 1551 145
rect 1485 73 1501 107
rect 1535 73 1551 107
rect 1485 17 1551 73
rect 1585 111 1623 191
rect 1657 191 1845 200
rect 1879 215 1999 225
rect 1879 191 1895 215
rect 1657 171 1895 191
rect 1657 137 1673 171
rect 1707 163 1895 171
rect 1707 137 1717 163
rect 1657 121 1717 137
rect 1829 157 1895 163
rect 1585 77 1587 111
rect 1621 87 1623 111
rect 1751 111 1795 127
rect 1829 123 1845 157
rect 1879 123 1895 157
rect 1829 121 1895 123
rect 1931 179 1997 181
rect 1931 145 1947 179
rect 1981 145 1997 179
rect 1751 87 1759 111
rect 1621 77 1759 87
rect 1793 87 1795 111
rect 1931 111 1997 145
rect 1931 87 1947 111
rect 1793 77 1947 87
rect 1981 77 1997 111
rect 1585 53 1997 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2bb2ai_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4108062
string GDS_START 4090412
<< end >>
