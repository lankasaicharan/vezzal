magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 41 49 653 241
rect 0 0 672 49
<< scnmos >>
rect 120 47 150 215
rect 206 47 236 215
rect 304 47 334 215
rect 434 47 464 215
rect 542 47 572 215
<< scpmoshvt >>
rect 86 367 116 619
rect 172 367 202 619
rect 362 367 392 619
rect 448 367 478 619
rect 542 367 572 619
<< ndiff >>
rect 67 163 120 215
rect 67 129 75 163
rect 109 129 120 163
rect 67 93 120 129
rect 67 59 75 93
rect 109 59 120 93
rect 67 47 120 59
rect 150 203 206 215
rect 150 169 161 203
rect 195 169 206 203
rect 150 101 206 169
rect 150 67 161 101
rect 195 67 206 101
rect 150 47 206 67
rect 236 163 304 215
rect 236 129 247 163
rect 281 129 304 163
rect 236 89 304 129
rect 236 55 247 89
rect 281 55 304 89
rect 236 47 304 55
rect 334 203 434 215
rect 334 169 345 203
rect 379 169 434 203
rect 334 101 434 169
rect 334 67 345 101
rect 379 67 434 101
rect 334 47 434 67
rect 464 47 542 215
rect 572 187 627 215
rect 572 153 585 187
rect 619 153 627 187
rect 572 93 627 153
rect 572 59 585 93
rect 619 59 627 93
rect 572 47 627 59
<< pdiff >>
rect 33 607 86 619
rect 33 573 41 607
rect 75 573 86 607
rect 33 508 86 573
rect 33 474 41 508
rect 75 474 86 508
rect 33 413 86 474
rect 33 379 41 413
rect 75 379 86 413
rect 33 367 86 379
rect 116 599 172 619
rect 116 565 127 599
rect 161 565 172 599
rect 116 504 172 565
rect 116 470 127 504
rect 161 470 172 504
rect 116 413 172 470
rect 116 379 127 413
rect 161 379 172 413
rect 116 367 172 379
rect 202 607 255 619
rect 202 573 213 607
rect 247 573 255 607
rect 202 494 255 573
rect 202 460 213 494
rect 247 460 255 494
rect 202 367 255 460
rect 309 599 362 619
rect 309 565 317 599
rect 351 565 362 599
rect 309 515 362 565
rect 309 481 317 515
rect 351 481 362 515
rect 309 436 362 481
rect 309 402 317 436
rect 351 402 362 436
rect 309 367 362 402
rect 392 599 448 619
rect 392 565 403 599
rect 437 565 448 599
rect 392 509 448 565
rect 392 475 403 509
rect 437 475 448 509
rect 392 413 448 475
rect 392 379 403 413
rect 437 379 448 413
rect 392 367 448 379
rect 478 607 542 619
rect 478 573 493 607
rect 527 573 542 607
rect 478 526 542 573
rect 478 492 493 526
rect 527 492 542 526
rect 478 439 542 492
rect 478 405 493 439
rect 527 405 542 439
rect 478 367 542 405
rect 572 599 625 619
rect 572 565 583 599
rect 617 565 625 599
rect 572 509 625 565
rect 572 475 583 509
rect 617 475 625 509
rect 572 413 625 475
rect 572 379 583 413
rect 617 379 625 413
rect 572 367 625 379
<< ndiffc >>
rect 75 129 109 163
rect 75 59 109 93
rect 161 169 195 203
rect 161 67 195 101
rect 247 129 281 163
rect 247 55 281 89
rect 345 169 379 203
rect 345 67 379 101
rect 585 153 619 187
rect 585 59 619 93
<< pdiffc >>
rect 41 573 75 607
rect 41 474 75 508
rect 41 379 75 413
rect 127 565 161 599
rect 127 470 161 504
rect 127 379 161 413
rect 213 573 247 607
rect 213 460 247 494
rect 317 565 351 599
rect 317 481 351 515
rect 317 402 351 436
rect 403 565 437 599
rect 403 475 437 509
rect 403 379 437 413
rect 493 573 527 607
rect 493 492 527 526
rect 493 405 527 439
rect 583 565 617 599
rect 583 475 617 509
rect 583 379 617 413
<< poly >>
rect 86 619 116 645
rect 172 619 202 645
rect 362 619 392 645
rect 448 619 478 645
rect 542 619 572 645
rect 86 299 116 367
rect 172 335 202 367
rect 362 335 392 367
rect 172 319 256 335
rect 172 299 206 319
rect 86 285 206 299
rect 240 285 256 319
rect 86 269 256 285
rect 304 319 392 335
rect 304 285 320 319
rect 354 305 392 319
rect 354 285 370 305
rect 448 303 478 367
rect 542 303 572 367
rect 304 269 370 285
rect 434 287 500 303
rect 120 215 150 269
rect 206 215 236 269
rect 304 215 334 269
rect 434 253 450 287
rect 484 253 500 287
rect 434 237 500 253
rect 542 287 631 303
rect 542 253 581 287
rect 615 253 631 287
rect 542 237 631 253
rect 434 215 464 237
rect 542 215 572 237
rect 120 21 150 47
rect 206 21 236 47
rect 304 21 334 47
rect 434 21 464 47
rect 542 21 572 47
<< polycont >>
rect 206 285 240 319
rect 320 285 354 319
rect 450 253 484 287
rect 581 253 615 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 25 607 83 649
rect 25 573 41 607
rect 75 573 83 607
rect 25 508 83 573
rect 25 474 41 508
rect 75 474 83 508
rect 25 413 83 474
rect 25 379 41 413
rect 75 379 83 413
rect 25 363 83 379
rect 117 599 163 615
rect 117 565 127 599
rect 161 565 163 599
rect 117 504 163 565
rect 117 470 127 504
rect 161 470 163 504
rect 117 413 163 470
rect 197 607 263 649
rect 197 573 213 607
rect 247 573 263 607
rect 197 494 263 573
rect 197 460 213 494
rect 247 460 263 494
rect 197 454 263 460
rect 301 599 364 615
rect 301 565 317 599
rect 351 565 364 599
rect 301 515 364 565
rect 301 481 317 515
rect 351 481 364 515
rect 301 436 364 481
rect 301 420 317 436
rect 117 379 127 413
rect 161 379 163 413
rect 117 231 163 379
rect 197 402 317 420
rect 351 402 364 436
rect 197 386 364 402
rect 398 599 443 615
rect 398 565 403 599
rect 437 565 443 599
rect 398 509 443 565
rect 398 475 403 509
rect 437 475 443 509
rect 398 413 443 475
rect 197 319 265 386
rect 398 379 403 413
rect 437 379 443 413
rect 477 607 543 649
rect 477 573 493 607
rect 527 573 543 607
rect 477 526 543 573
rect 477 492 493 526
rect 527 492 543 526
rect 477 439 543 492
rect 477 405 493 439
rect 527 405 543 439
rect 577 599 621 615
rect 577 565 583 599
rect 617 565 621 599
rect 577 509 621 565
rect 577 475 583 509
rect 617 475 621 509
rect 577 413 621 475
rect 398 371 443 379
rect 577 379 583 413
rect 617 379 621 413
rect 577 371 621 379
rect 197 285 206 319
rect 240 285 265 319
rect 197 269 265 285
rect 299 319 364 352
rect 398 337 621 371
rect 299 285 320 319
rect 354 285 364 319
rect 299 269 364 285
rect 413 287 547 303
rect 231 231 265 269
rect 413 253 450 287
rect 484 253 547 287
rect 117 203 197 231
rect 117 197 161 203
rect 159 169 161 197
rect 195 169 197 203
rect 231 203 379 231
rect 231 197 345 203
rect 59 129 75 163
rect 109 129 125 163
rect 59 93 125 129
rect 59 59 75 93
rect 109 59 125 93
rect 59 17 125 59
rect 159 101 197 169
rect 341 169 345 197
rect 159 67 161 101
rect 195 67 197 101
rect 159 51 197 67
rect 231 129 247 163
rect 281 129 297 163
rect 231 89 297 129
rect 231 55 247 89
rect 281 55 297 89
rect 231 17 297 55
rect 341 101 379 169
rect 341 67 345 101
rect 341 51 379 67
rect 413 63 547 253
rect 581 287 654 303
rect 615 253 654 287
rect 581 237 654 253
rect 581 187 635 203
rect 581 153 585 187
rect 619 153 635 187
rect 581 93 635 153
rect 581 59 585 93
rect 619 59 635 93
rect 581 17 635 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21o_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2583068
string GDS_START 2575610
<< end >>
