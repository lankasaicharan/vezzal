magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1260 -1260 3530 1664
<< poly >>
rect 10 351 128 402
rect 10 45 26 351
rect 10 2 128 45
rect 2142 351 2260 402
rect 2244 45 2260 351
rect 2142 2 2260 45
<< polycont >>
rect 26 45 128 351
rect 2142 45 2244 351
<< npolyres >>
rect 128 2 2142 402
<< locali >>
rect 2 351 152 404
rect 2 339 26 351
rect 128 339 152 351
rect 2 305 12 339
rect 142 305 152 339
rect 2 215 26 305
rect 128 215 152 305
rect 2 181 12 215
rect 142 181 152 215
rect 2 91 26 181
rect 128 91 152 181
rect 2 57 12 91
rect 142 57 152 91
rect 2 45 26 57
rect 128 45 152 57
rect 2 0 152 45
rect 2118 351 2268 404
rect 2118 339 2142 351
rect 2244 339 2268 351
rect 2118 305 2128 339
rect 2258 305 2268 339
rect 2118 215 2142 305
rect 2244 215 2268 305
rect 2118 181 2128 215
rect 2258 181 2268 215
rect 2118 91 2142 181
rect 2244 91 2268 181
rect 2118 57 2128 91
rect 2258 57 2268 91
rect 2118 45 2142 57
rect 2244 45 2268 57
rect 2118 0 2268 45
<< viali >>
rect 12 305 26 339
rect 26 305 46 339
rect 108 305 128 339
rect 128 305 142 339
rect 12 181 26 215
rect 26 181 46 215
rect 108 181 128 215
rect 128 181 142 215
rect 12 57 26 91
rect 26 57 46 91
rect 108 57 128 91
rect 128 57 142 91
rect 2128 305 2142 339
rect 2142 305 2162 339
rect 2224 305 2244 339
rect 2244 305 2258 339
rect 2128 181 2142 215
rect 2142 181 2162 215
rect 2224 181 2244 215
rect 2244 181 2258 215
rect 2128 57 2142 91
rect 2142 57 2162 91
rect 2224 57 2244 91
rect 2244 57 2258 91
<< metal1 >>
rect 0 339 154 403
rect 0 305 12 339
rect 46 305 108 339
rect 142 305 154 339
rect 0 215 154 305
rect 0 181 12 215
rect 46 181 108 215
rect 142 181 154 215
rect 0 91 154 181
rect 0 57 12 91
rect 46 57 108 91
rect 142 57 154 91
rect 0 1 154 57
rect 2116 339 2270 403
rect 2116 305 2128 339
rect 2162 305 2224 339
rect 2258 305 2270 339
rect 2116 215 2270 305
rect 2116 181 2128 215
rect 2162 181 2224 215
rect 2258 181 2270 215
rect 2116 91 2270 181
rect 2116 57 2128 91
rect 2162 57 2224 91
rect 2258 57 2270 91
rect 2116 1 2270 57
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 1907698
string GDS_START 1904750
<< end >>
