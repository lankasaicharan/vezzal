magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 1 49 764 248
rect 0 0 768 49
<< scnmos >>
rect 82 74 112 222
rect 291 74 321 222
rect 363 74 393 222
rect 441 74 471 222
rect 543 74 573 222
rect 651 74 681 222
<< scpmoshvt >>
rect 86 368 116 592
rect 212 413 242 581
rect 312 413 342 581
rect 463 413 493 581
rect 570 381 600 581
rect 654 381 684 581
<< ndiff >>
rect 27 192 82 222
rect 27 158 37 192
rect 71 158 82 192
rect 27 120 82 158
rect 27 86 37 120
rect 71 86 82 120
rect 27 74 82 86
rect 112 192 167 222
rect 112 158 123 192
rect 157 158 167 192
rect 112 120 167 158
rect 112 86 123 120
rect 157 86 167 120
rect 112 74 167 86
rect 221 210 291 222
rect 221 176 232 210
rect 266 176 291 210
rect 221 120 291 176
rect 221 86 232 120
rect 266 86 291 120
rect 221 74 291 86
rect 321 74 363 222
rect 393 74 441 222
rect 471 210 543 222
rect 471 176 492 210
rect 526 176 543 210
rect 471 120 543 176
rect 471 86 492 120
rect 526 86 543 120
rect 471 74 543 86
rect 573 131 651 222
rect 573 97 592 131
rect 626 97 651 131
rect 573 74 651 97
rect 681 210 738 222
rect 681 176 692 210
rect 726 176 738 210
rect 681 120 738 176
rect 681 86 692 120
rect 726 86 738 120
rect 681 74 738 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 584 190 592
rect 116 550 139 584
rect 173 581 190 584
rect 173 550 212 581
rect 116 516 212 550
rect 116 482 139 516
rect 173 482 212 516
rect 116 413 212 482
rect 242 569 312 581
rect 242 535 255 569
rect 289 535 312 569
rect 242 465 312 535
rect 242 431 255 465
rect 289 431 312 465
rect 242 413 312 431
rect 342 541 463 581
rect 342 507 386 541
rect 420 507 463 541
rect 342 413 463 507
rect 493 569 570 581
rect 493 535 523 569
rect 557 535 570 569
rect 493 459 570 535
rect 493 425 523 459
rect 557 425 570 459
rect 493 413 570 425
rect 116 368 169 413
rect 511 381 570 413
rect 600 381 654 581
rect 684 569 741 581
rect 684 535 697 569
rect 731 535 741 569
rect 684 501 741 535
rect 684 467 697 501
rect 731 467 741 501
rect 684 433 741 467
rect 684 399 697 433
rect 731 399 741 433
rect 684 381 741 399
<< ndiffc >>
rect 37 158 71 192
rect 37 86 71 120
rect 123 158 157 192
rect 123 86 157 120
rect 232 176 266 210
rect 232 86 266 120
rect 492 176 526 210
rect 492 86 526 120
rect 592 97 626 131
rect 692 176 726 210
rect 692 86 726 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 550 173 584
rect 139 482 173 516
rect 255 535 289 569
rect 255 431 289 465
rect 386 507 420 541
rect 523 535 557 569
rect 523 425 557 459
rect 697 535 731 569
rect 697 467 731 501
rect 697 399 731 433
<< poly >>
rect 86 592 116 618
rect 212 581 242 607
rect 312 581 342 607
rect 463 581 493 607
rect 570 581 600 607
rect 654 581 684 607
rect 212 398 242 413
rect 312 398 342 413
rect 463 398 493 413
rect 209 376 245 398
rect 309 380 345 398
rect 86 353 116 368
rect 201 360 267 376
rect 83 310 119 353
rect 201 326 217 360
rect 251 326 267 360
rect 201 310 267 326
rect 309 364 393 380
rect 309 330 325 364
rect 359 330 393 364
rect 460 349 496 398
rect 570 366 600 381
rect 654 366 684 381
rect 567 349 603 366
rect 309 314 393 330
rect 82 294 153 310
rect 82 260 103 294
rect 137 260 153 294
rect 82 244 153 260
rect 237 267 267 310
rect 82 222 112 244
rect 237 237 321 267
rect 291 222 321 237
rect 363 222 393 314
rect 435 333 501 349
rect 435 299 451 333
rect 485 299 501 333
rect 435 283 501 299
rect 543 333 609 349
rect 543 299 559 333
rect 593 299 609 333
rect 543 283 609 299
rect 651 326 687 366
rect 651 310 747 326
rect 441 222 471 283
rect 543 222 573 283
rect 651 276 697 310
rect 731 276 747 310
rect 651 260 747 276
rect 651 222 681 260
rect 82 48 112 74
rect 291 48 321 74
rect 363 48 393 74
rect 441 48 471 74
rect 543 48 573 74
rect 651 48 681 74
<< polycont >>
rect 217 326 251 360
rect 325 330 359 364
rect 103 260 137 294
rect 451 299 485 333
rect 559 299 593 333
rect 697 276 731 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 19 580 89 596
rect 19 546 39 580
rect 73 546 89 580
rect 19 497 89 546
rect 19 463 39 497
rect 73 463 89 497
rect 123 584 189 649
rect 123 550 139 584
rect 173 550 189 584
rect 123 516 189 550
rect 123 482 139 516
rect 173 482 189 516
rect 239 569 305 585
rect 239 535 255 569
rect 289 535 305 569
rect 19 414 89 463
rect 239 465 305 535
rect 348 541 458 649
rect 348 507 386 541
rect 420 507 458 541
rect 348 491 458 507
rect 507 569 573 585
rect 507 535 523 569
rect 557 535 573 569
rect 239 448 255 465
rect 19 380 39 414
rect 73 380 89 414
rect 19 364 89 380
rect 123 431 255 448
rect 289 449 305 465
rect 507 459 573 535
rect 507 449 523 459
rect 289 431 523 449
rect 123 425 523 431
rect 557 425 573 459
rect 123 414 573 425
rect 19 208 53 364
rect 123 310 157 414
rect 507 409 573 414
rect 681 569 747 649
rect 681 535 697 569
rect 731 535 747 569
rect 681 501 747 535
rect 681 467 697 501
rect 731 467 747 501
rect 681 433 747 467
rect 681 399 697 433
rect 731 399 747 433
rect 681 390 747 399
rect 201 360 267 376
rect 201 326 217 360
rect 251 326 267 360
rect 201 310 267 326
rect 309 364 375 380
rect 309 330 325 364
rect 359 330 375 364
rect 87 294 157 310
rect 87 260 103 294
rect 137 276 157 294
rect 137 260 266 276
rect 87 242 266 260
rect 216 210 266 242
rect 19 192 71 208
rect 19 158 37 192
rect 19 120 71 158
rect 19 86 37 120
rect 19 70 71 86
rect 107 192 173 208
rect 107 158 123 192
rect 157 158 173 192
rect 107 120 173 158
rect 107 86 123 120
rect 157 86 173 120
rect 107 17 173 86
rect 216 176 232 210
rect 216 120 266 176
rect 216 86 232 120
rect 309 88 375 330
rect 409 333 501 356
rect 409 299 451 333
rect 485 299 501 333
rect 409 283 501 299
rect 543 333 647 356
rect 543 299 559 333
rect 593 299 647 333
rect 543 283 647 299
rect 681 310 747 356
rect 681 276 697 310
rect 731 276 747 310
rect 681 260 747 276
rect 476 210 742 226
rect 476 176 492 210
rect 526 192 692 210
rect 526 176 542 192
rect 476 120 542 176
rect 676 176 692 192
rect 726 176 742 210
rect 216 70 266 86
rect 476 86 492 120
rect 526 86 542 120
rect 476 70 542 86
rect 576 131 642 158
rect 576 97 592 131
rect 626 97 642 131
rect 576 17 642 97
rect 676 120 742 176
rect 676 86 692 120
rect 726 86 742 120
rect 676 70 742 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o2111a_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 2896670
string GDS_START 2888870
<< end >>
