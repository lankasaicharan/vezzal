magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3602 1975
<< nwell >>
rect -38 331 2342 704
<< pwell >>
rect 37 49 2298 243
rect 0 0 2304 49
<< scnmos >>
rect 116 49 146 217
rect 202 49 232 217
rect 288 49 318 217
rect 383 49 413 217
rect 469 49 499 217
rect 555 49 585 217
rect 641 49 671 217
rect 727 49 757 217
rect 813 49 843 217
rect 899 49 929 217
rect 985 49 1015 217
rect 1071 49 1101 217
rect 1157 49 1187 217
rect 1243 49 1273 217
rect 1329 49 1359 217
rect 1415 49 1445 217
rect 1501 49 1531 217
rect 1587 49 1617 217
rect 1673 49 1703 217
rect 1759 49 1789 217
rect 1845 49 1875 217
rect 1931 49 1961 217
rect 2017 49 2047 217
rect 2103 49 2133 217
rect 2189 49 2219 217
<< scpmoshvt >>
rect 116 367 146 619
rect 202 367 232 619
rect 288 367 318 619
rect 383 367 413 619
rect 469 367 499 619
rect 555 367 585 619
rect 641 367 671 619
rect 727 367 757 619
rect 813 367 843 619
rect 899 367 929 619
rect 985 367 1015 619
rect 1071 367 1101 619
rect 1157 367 1187 619
rect 1243 367 1273 619
rect 1329 367 1359 619
rect 1415 367 1445 619
rect 1501 367 1531 619
rect 1587 367 1617 619
rect 1673 367 1703 619
rect 1759 367 1789 619
rect 1845 367 1875 619
rect 1931 367 1961 619
rect 2017 367 2047 619
rect 2103 367 2133 619
rect 2189 367 2219 619
<< ndiff >>
rect 63 187 116 217
rect 63 153 71 187
rect 105 153 116 187
rect 63 113 116 153
rect 63 79 71 113
rect 105 79 116 113
rect 63 49 116 79
rect 146 165 202 217
rect 146 131 157 165
rect 191 131 202 165
rect 146 97 202 131
rect 146 63 157 97
rect 191 63 202 97
rect 146 49 202 63
rect 232 187 288 217
rect 232 153 243 187
rect 277 153 288 187
rect 232 113 288 153
rect 232 79 243 113
rect 277 79 288 113
rect 232 49 288 79
rect 318 165 383 217
rect 318 131 329 165
rect 363 131 383 165
rect 318 97 383 131
rect 318 63 329 97
rect 363 63 383 97
rect 318 49 383 63
rect 413 187 469 217
rect 413 153 424 187
rect 458 153 469 187
rect 413 113 469 153
rect 413 79 424 113
rect 458 79 469 113
rect 413 49 469 79
rect 499 161 555 217
rect 499 127 510 161
rect 544 127 555 161
rect 499 93 555 127
rect 499 59 510 93
rect 544 59 555 93
rect 499 49 555 59
rect 585 187 641 217
rect 585 153 596 187
rect 630 153 641 187
rect 585 113 641 153
rect 585 79 596 113
rect 630 79 641 113
rect 585 49 641 79
rect 671 161 727 217
rect 671 127 682 161
rect 716 127 727 161
rect 671 93 727 127
rect 671 59 682 93
rect 716 59 727 93
rect 671 49 727 59
rect 757 187 813 217
rect 757 153 768 187
rect 802 153 813 187
rect 757 113 813 153
rect 757 79 768 113
rect 802 79 813 113
rect 757 49 813 79
rect 843 161 899 217
rect 843 127 854 161
rect 888 127 899 161
rect 843 93 899 127
rect 843 59 854 93
rect 888 59 899 93
rect 843 49 899 59
rect 929 187 985 217
rect 929 153 940 187
rect 974 153 985 187
rect 929 113 985 153
rect 929 79 940 113
rect 974 79 985 113
rect 929 49 985 79
rect 1015 187 1071 217
rect 1015 153 1026 187
rect 1060 153 1071 187
rect 1015 113 1071 153
rect 1015 79 1026 113
rect 1060 79 1071 113
rect 1015 49 1071 79
rect 1101 187 1157 217
rect 1101 153 1112 187
rect 1146 153 1157 187
rect 1101 113 1157 153
rect 1101 79 1112 113
rect 1146 79 1157 113
rect 1101 49 1157 79
rect 1187 187 1243 217
rect 1187 153 1198 187
rect 1232 153 1243 187
rect 1187 113 1243 153
rect 1187 79 1198 113
rect 1232 79 1243 113
rect 1187 49 1243 79
rect 1273 187 1329 217
rect 1273 153 1284 187
rect 1318 153 1329 187
rect 1273 113 1329 153
rect 1273 79 1284 113
rect 1318 79 1329 113
rect 1273 49 1329 79
rect 1359 187 1415 217
rect 1359 153 1370 187
rect 1404 153 1415 187
rect 1359 113 1415 153
rect 1359 79 1370 113
rect 1404 79 1415 113
rect 1359 49 1415 79
rect 1445 187 1501 217
rect 1445 153 1456 187
rect 1490 153 1501 187
rect 1445 113 1501 153
rect 1445 79 1456 113
rect 1490 79 1501 113
rect 1445 49 1501 79
rect 1531 187 1587 217
rect 1531 153 1542 187
rect 1576 153 1587 187
rect 1531 113 1587 153
rect 1531 79 1542 113
rect 1576 79 1587 113
rect 1531 49 1587 79
rect 1617 187 1673 217
rect 1617 153 1628 187
rect 1662 153 1673 187
rect 1617 113 1673 153
rect 1617 79 1628 113
rect 1662 79 1673 113
rect 1617 49 1673 79
rect 1703 187 1759 217
rect 1703 153 1714 187
rect 1748 153 1759 187
rect 1703 113 1759 153
rect 1703 79 1714 113
rect 1748 79 1759 113
rect 1703 49 1759 79
rect 1789 187 1845 217
rect 1789 153 1800 187
rect 1834 153 1845 187
rect 1789 113 1845 153
rect 1789 79 1800 113
rect 1834 79 1845 113
rect 1789 49 1845 79
rect 1875 187 1931 217
rect 1875 153 1886 187
rect 1920 153 1931 187
rect 1875 113 1931 153
rect 1875 79 1886 113
rect 1920 79 1931 113
rect 1875 49 1931 79
rect 1961 187 2017 217
rect 1961 153 1972 187
rect 2006 153 2017 187
rect 1961 113 2017 153
rect 1961 79 1972 113
rect 2006 79 2017 113
rect 1961 49 2017 79
rect 2047 187 2103 217
rect 2047 153 2058 187
rect 2092 153 2103 187
rect 2047 113 2103 153
rect 2047 79 2058 113
rect 2092 79 2103 113
rect 2047 49 2103 79
rect 2133 187 2189 217
rect 2133 153 2144 187
rect 2178 153 2189 187
rect 2133 113 2189 153
rect 2133 79 2144 113
rect 2178 79 2189 113
rect 2133 49 2189 79
rect 2219 187 2272 217
rect 2219 153 2230 187
rect 2264 153 2272 187
rect 2219 113 2272 153
rect 2219 79 2230 113
rect 2264 79 2272 113
rect 2219 49 2272 79
<< pdiff >>
rect 63 589 116 619
rect 63 555 71 589
rect 105 555 116 589
rect 63 510 116 555
rect 63 476 71 510
rect 105 476 116 510
rect 63 436 116 476
rect 63 402 71 436
rect 105 402 116 436
rect 63 367 116 402
rect 146 572 202 619
rect 146 538 157 572
rect 191 538 202 572
rect 146 504 202 538
rect 146 470 157 504
rect 191 470 202 504
rect 146 367 202 470
rect 232 589 288 619
rect 232 555 243 589
rect 277 555 288 589
rect 232 510 288 555
rect 232 476 243 510
rect 277 476 288 510
rect 232 436 288 476
rect 232 402 243 436
rect 277 402 288 436
rect 232 367 288 402
rect 318 572 383 619
rect 318 538 333 572
rect 367 538 383 572
rect 318 504 383 538
rect 318 470 333 504
rect 367 470 383 504
rect 318 367 383 470
rect 413 589 469 619
rect 413 555 424 589
rect 458 555 469 589
rect 413 510 469 555
rect 413 476 424 510
rect 458 476 469 510
rect 413 436 469 476
rect 413 402 424 436
rect 458 402 469 436
rect 413 367 469 402
rect 499 607 555 619
rect 499 573 510 607
rect 544 573 555 607
rect 499 539 555 573
rect 499 505 510 539
rect 544 505 555 539
rect 499 471 555 505
rect 499 437 510 471
rect 544 437 555 471
rect 499 367 555 437
rect 585 589 641 619
rect 585 555 596 589
rect 630 555 641 589
rect 585 510 641 555
rect 585 476 596 510
rect 630 476 641 510
rect 585 436 641 476
rect 585 402 596 436
rect 630 402 641 436
rect 585 367 641 402
rect 671 607 727 619
rect 671 573 682 607
rect 716 573 727 607
rect 671 539 727 573
rect 671 505 682 539
rect 716 505 727 539
rect 671 471 727 505
rect 671 437 682 471
rect 716 437 727 471
rect 671 367 727 437
rect 757 589 813 619
rect 757 555 768 589
rect 802 555 813 589
rect 757 510 813 555
rect 757 476 768 510
rect 802 476 813 510
rect 757 436 813 476
rect 757 402 768 436
rect 802 402 813 436
rect 757 367 813 402
rect 843 607 899 619
rect 843 573 854 607
rect 888 573 899 607
rect 843 539 899 573
rect 843 505 854 539
rect 888 505 899 539
rect 843 471 899 505
rect 843 437 854 471
rect 888 437 899 471
rect 843 367 899 437
rect 929 589 985 619
rect 929 555 940 589
rect 974 555 985 589
rect 929 510 985 555
rect 929 476 940 510
rect 974 476 985 510
rect 929 431 985 476
rect 929 397 940 431
rect 974 397 985 431
rect 929 367 985 397
rect 1015 599 1071 619
rect 1015 565 1026 599
rect 1060 565 1071 599
rect 1015 520 1071 565
rect 1015 486 1026 520
rect 1060 486 1071 520
rect 1015 441 1071 486
rect 1015 407 1026 441
rect 1060 407 1071 441
rect 1015 367 1071 407
rect 1101 589 1157 619
rect 1101 555 1112 589
rect 1146 555 1157 589
rect 1101 510 1157 555
rect 1101 476 1112 510
rect 1146 476 1157 510
rect 1101 431 1157 476
rect 1101 397 1112 431
rect 1146 397 1157 431
rect 1101 367 1157 397
rect 1187 599 1243 619
rect 1187 565 1198 599
rect 1232 565 1243 599
rect 1187 520 1243 565
rect 1187 486 1198 520
rect 1232 486 1243 520
rect 1187 441 1243 486
rect 1187 407 1198 441
rect 1232 407 1243 441
rect 1187 367 1243 407
rect 1273 589 1329 619
rect 1273 555 1284 589
rect 1318 555 1329 589
rect 1273 510 1329 555
rect 1273 476 1284 510
rect 1318 476 1329 510
rect 1273 431 1329 476
rect 1273 397 1284 431
rect 1318 397 1329 431
rect 1273 367 1329 397
rect 1359 599 1415 619
rect 1359 565 1370 599
rect 1404 565 1415 599
rect 1359 520 1415 565
rect 1359 486 1370 520
rect 1404 486 1415 520
rect 1359 441 1415 486
rect 1359 407 1370 441
rect 1404 407 1415 441
rect 1359 367 1415 407
rect 1445 589 1501 619
rect 1445 555 1456 589
rect 1490 555 1501 589
rect 1445 510 1501 555
rect 1445 476 1456 510
rect 1490 476 1501 510
rect 1445 431 1501 476
rect 1445 397 1456 431
rect 1490 397 1501 431
rect 1445 367 1501 397
rect 1531 599 1587 619
rect 1531 565 1542 599
rect 1576 565 1587 599
rect 1531 520 1587 565
rect 1531 486 1542 520
rect 1576 486 1587 520
rect 1531 441 1587 486
rect 1531 407 1542 441
rect 1576 407 1587 441
rect 1531 367 1587 407
rect 1617 589 1673 619
rect 1617 555 1628 589
rect 1662 555 1673 589
rect 1617 510 1673 555
rect 1617 476 1628 510
rect 1662 476 1673 510
rect 1617 431 1673 476
rect 1617 397 1628 431
rect 1662 397 1673 431
rect 1617 367 1673 397
rect 1703 599 1759 619
rect 1703 565 1714 599
rect 1748 565 1759 599
rect 1703 520 1759 565
rect 1703 486 1714 520
rect 1748 486 1759 520
rect 1703 441 1759 486
rect 1703 407 1714 441
rect 1748 407 1759 441
rect 1703 367 1759 407
rect 1789 589 1845 619
rect 1789 555 1800 589
rect 1834 555 1845 589
rect 1789 510 1845 555
rect 1789 476 1800 510
rect 1834 476 1845 510
rect 1789 431 1845 476
rect 1789 397 1800 431
rect 1834 397 1845 431
rect 1789 367 1845 397
rect 1875 599 1931 619
rect 1875 565 1886 599
rect 1920 565 1931 599
rect 1875 520 1931 565
rect 1875 486 1886 520
rect 1920 486 1931 520
rect 1875 441 1931 486
rect 1875 407 1886 441
rect 1920 407 1931 441
rect 1875 367 1931 407
rect 1961 589 2017 619
rect 1961 555 1972 589
rect 2006 555 2017 589
rect 1961 510 2017 555
rect 1961 476 1972 510
rect 2006 476 2017 510
rect 1961 431 2017 476
rect 1961 397 1972 431
rect 2006 397 2017 431
rect 1961 367 2017 397
rect 2047 599 2103 619
rect 2047 565 2058 599
rect 2092 565 2103 599
rect 2047 520 2103 565
rect 2047 486 2058 520
rect 2092 486 2103 520
rect 2047 441 2103 486
rect 2047 407 2058 441
rect 2092 407 2103 441
rect 2047 367 2103 407
rect 2133 589 2189 619
rect 2133 555 2144 589
rect 2178 555 2189 589
rect 2133 510 2189 555
rect 2133 476 2144 510
rect 2178 476 2189 510
rect 2133 431 2189 476
rect 2133 397 2144 431
rect 2178 397 2189 431
rect 2133 367 2189 397
rect 2219 599 2272 619
rect 2219 565 2230 599
rect 2264 565 2272 599
rect 2219 520 2272 565
rect 2219 486 2230 520
rect 2264 486 2272 520
rect 2219 441 2272 486
rect 2219 407 2230 441
rect 2264 407 2272 441
rect 2219 367 2272 407
<< ndiffc >>
rect 71 153 105 187
rect 71 79 105 113
rect 157 131 191 165
rect 157 63 191 97
rect 243 153 277 187
rect 243 79 277 113
rect 329 131 363 165
rect 329 63 363 97
rect 424 153 458 187
rect 424 79 458 113
rect 510 127 544 161
rect 510 59 544 93
rect 596 153 630 187
rect 596 79 630 113
rect 682 127 716 161
rect 682 59 716 93
rect 768 153 802 187
rect 768 79 802 113
rect 854 127 888 161
rect 854 59 888 93
rect 940 153 974 187
rect 940 79 974 113
rect 1026 153 1060 187
rect 1026 79 1060 113
rect 1112 153 1146 187
rect 1112 79 1146 113
rect 1198 153 1232 187
rect 1198 79 1232 113
rect 1284 153 1318 187
rect 1284 79 1318 113
rect 1370 153 1404 187
rect 1370 79 1404 113
rect 1456 153 1490 187
rect 1456 79 1490 113
rect 1542 153 1576 187
rect 1542 79 1576 113
rect 1628 153 1662 187
rect 1628 79 1662 113
rect 1714 153 1748 187
rect 1714 79 1748 113
rect 1800 153 1834 187
rect 1800 79 1834 113
rect 1886 153 1920 187
rect 1886 79 1920 113
rect 1972 153 2006 187
rect 1972 79 2006 113
rect 2058 153 2092 187
rect 2058 79 2092 113
rect 2144 153 2178 187
rect 2144 79 2178 113
rect 2230 153 2264 187
rect 2230 79 2264 113
<< pdiffc >>
rect 71 555 105 589
rect 71 476 105 510
rect 71 402 105 436
rect 157 538 191 572
rect 157 470 191 504
rect 243 555 277 589
rect 243 476 277 510
rect 243 402 277 436
rect 333 538 367 572
rect 333 470 367 504
rect 424 555 458 589
rect 424 476 458 510
rect 424 402 458 436
rect 510 573 544 607
rect 510 505 544 539
rect 510 437 544 471
rect 596 555 630 589
rect 596 476 630 510
rect 596 402 630 436
rect 682 573 716 607
rect 682 505 716 539
rect 682 437 716 471
rect 768 555 802 589
rect 768 476 802 510
rect 768 402 802 436
rect 854 573 888 607
rect 854 505 888 539
rect 854 437 888 471
rect 940 555 974 589
rect 940 476 974 510
rect 940 397 974 431
rect 1026 565 1060 599
rect 1026 486 1060 520
rect 1026 407 1060 441
rect 1112 555 1146 589
rect 1112 476 1146 510
rect 1112 397 1146 431
rect 1198 565 1232 599
rect 1198 486 1232 520
rect 1198 407 1232 441
rect 1284 555 1318 589
rect 1284 476 1318 510
rect 1284 397 1318 431
rect 1370 565 1404 599
rect 1370 486 1404 520
rect 1370 407 1404 441
rect 1456 555 1490 589
rect 1456 476 1490 510
rect 1456 397 1490 431
rect 1542 565 1576 599
rect 1542 486 1576 520
rect 1542 407 1576 441
rect 1628 555 1662 589
rect 1628 476 1662 510
rect 1628 397 1662 431
rect 1714 565 1748 599
rect 1714 486 1748 520
rect 1714 407 1748 441
rect 1800 555 1834 589
rect 1800 476 1834 510
rect 1800 397 1834 431
rect 1886 565 1920 599
rect 1886 486 1920 520
rect 1886 407 1920 441
rect 1972 555 2006 589
rect 1972 476 2006 510
rect 1972 397 2006 431
rect 2058 565 2092 599
rect 2058 486 2092 520
rect 2058 407 2092 441
rect 2144 555 2178 589
rect 2144 476 2178 510
rect 2144 397 2178 431
rect 2230 565 2264 599
rect 2230 486 2264 520
rect 2230 407 2264 441
<< poly >>
rect 116 619 146 645
rect 202 619 232 645
rect 288 619 318 645
rect 383 619 413 645
rect 469 619 499 645
rect 555 619 585 645
rect 641 619 671 645
rect 727 619 757 645
rect 813 619 843 645
rect 899 619 929 645
rect 985 619 1015 645
rect 1071 619 1101 645
rect 1157 619 1187 645
rect 1243 619 1273 645
rect 1329 619 1359 645
rect 1415 619 1445 645
rect 1501 619 1531 645
rect 1587 619 1617 645
rect 1673 619 1703 645
rect 1759 619 1789 645
rect 1845 619 1875 645
rect 1931 619 1961 645
rect 2017 619 2047 645
rect 2103 619 2133 645
rect 2189 619 2219 645
rect 116 335 146 367
rect 202 335 232 367
rect 288 335 318 367
rect 44 319 318 335
rect 383 331 413 367
rect 469 331 499 367
rect 555 331 585 367
rect 641 331 671 367
rect 727 331 757 367
rect 813 331 843 367
rect 44 285 60 319
rect 94 285 128 319
rect 162 285 196 319
rect 230 285 264 319
rect 298 285 318 319
rect 44 269 318 285
rect 116 217 146 269
rect 202 217 232 269
rect 288 217 318 269
rect 360 315 843 331
rect 360 281 376 315
rect 410 281 444 315
rect 478 281 512 315
rect 546 281 580 315
rect 614 281 648 315
rect 682 281 716 315
rect 750 281 784 315
rect 818 281 843 315
rect 360 265 843 281
rect 383 217 413 265
rect 469 217 499 265
rect 555 217 585 265
rect 641 217 671 265
rect 727 217 757 265
rect 813 217 843 265
rect 899 335 929 367
rect 985 335 1015 367
rect 1071 335 1101 367
rect 1157 335 1187 367
rect 1243 335 1273 367
rect 1329 335 1359 367
rect 1415 335 1445 367
rect 1501 335 1531 367
rect 1587 335 1617 367
rect 1673 335 1703 367
rect 1759 335 1789 367
rect 1845 335 1875 367
rect 1931 335 1961 367
rect 2017 335 2047 367
rect 2103 335 2133 367
rect 2189 335 2219 367
rect 899 319 2219 335
rect 899 285 1026 319
rect 1060 285 1198 319
rect 1232 285 1370 319
rect 1404 285 1542 319
rect 1576 285 1714 319
rect 1748 285 1886 319
rect 1920 285 2058 319
rect 2092 285 2219 319
rect 899 269 2219 285
rect 899 217 929 269
rect 985 217 1015 269
rect 1071 217 1101 269
rect 1157 217 1187 269
rect 1243 217 1273 269
rect 1329 217 1359 269
rect 1415 217 1445 269
rect 1501 217 1531 269
rect 1587 217 1617 269
rect 1673 217 1703 269
rect 1759 217 1789 269
rect 1845 217 1875 269
rect 1931 217 1961 269
rect 2017 217 2047 269
rect 2103 217 2133 269
rect 2189 217 2219 269
rect 116 23 146 49
rect 202 23 232 49
rect 288 23 318 49
rect 383 23 413 49
rect 469 23 499 49
rect 555 23 585 49
rect 641 23 671 49
rect 727 23 757 49
rect 813 23 843 49
rect 899 23 929 49
rect 985 23 1015 49
rect 1071 23 1101 49
rect 1157 23 1187 49
rect 1243 23 1273 49
rect 1329 23 1359 49
rect 1415 23 1445 49
rect 1501 23 1531 49
rect 1587 23 1617 49
rect 1673 23 1703 49
rect 1759 23 1789 49
rect 1845 23 1875 49
rect 1931 23 1961 49
rect 2017 23 2047 49
rect 2103 23 2133 49
rect 2189 23 2219 49
<< polycont >>
rect 60 285 94 319
rect 128 285 162 319
rect 196 285 230 319
rect 264 285 298 319
rect 376 281 410 315
rect 444 281 478 315
rect 512 281 546 315
rect 580 281 614 315
rect 648 281 682 315
rect 716 281 750 315
rect 784 281 818 315
rect 1026 285 1060 319
rect 1198 285 1232 319
rect 1370 285 1404 319
rect 1542 285 1576 319
rect 1714 285 1748 319
rect 1886 285 1920 319
rect 2058 285 2092 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 55 589 114 605
rect 55 555 71 589
rect 105 555 114 589
rect 55 510 114 555
rect 55 476 71 510
rect 105 476 114 510
rect 55 436 114 476
rect 148 572 200 649
rect 148 538 157 572
rect 191 538 200 572
rect 148 504 200 538
rect 148 470 157 504
rect 191 470 200 504
rect 148 454 200 470
rect 234 589 286 605
rect 234 555 243 589
rect 277 555 286 589
rect 234 510 286 555
rect 234 476 243 510
rect 277 476 286 510
rect 55 402 71 436
rect 105 420 114 436
rect 234 436 286 476
rect 320 572 381 649
rect 501 607 553 649
rect 320 538 333 572
rect 367 538 381 572
rect 320 504 381 538
rect 320 470 333 504
rect 367 470 381 504
rect 320 454 381 470
rect 418 589 467 605
rect 418 555 424 589
rect 458 555 467 589
rect 418 510 467 555
rect 418 476 424 510
rect 458 476 467 510
rect 234 420 243 436
rect 105 402 243 420
rect 277 420 286 436
rect 418 436 467 476
rect 277 402 384 420
rect 55 386 384 402
rect 19 319 314 352
rect 19 285 60 319
rect 94 285 128 319
rect 162 285 196 319
rect 230 285 264 319
rect 298 285 314 319
rect 19 283 314 285
rect 350 317 384 386
rect 418 402 424 436
rect 458 402 467 436
rect 501 573 510 607
rect 544 573 553 607
rect 673 607 725 649
rect 501 539 553 573
rect 501 505 510 539
rect 544 505 553 539
rect 501 471 553 505
rect 501 437 510 471
rect 544 437 553 471
rect 501 421 553 437
rect 587 589 639 605
rect 587 555 596 589
rect 630 555 639 589
rect 587 510 639 555
rect 587 476 596 510
rect 630 476 639 510
rect 587 436 639 476
rect 418 385 467 402
rect 587 402 596 436
rect 630 402 639 436
rect 673 573 682 607
rect 716 573 725 607
rect 845 607 897 649
rect 673 539 725 573
rect 673 505 682 539
rect 716 505 725 539
rect 673 471 725 505
rect 673 437 682 471
rect 716 437 725 471
rect 673 421 725 437
rect 759 589 811 605
rect 759 555 768 589
rect 802 555 811 589
rect 759 510 811 555
rect 759 476 768 510
rect 802 476 811 510
rect 759 436 811 476
rect 587 385 639 402
rect 759 402 768 436
rect 802 402 811 436
rect 845 573 854 607
rect 888 573 897 607
rect 845 539 897 573
rect 845 505 854 539
rect 888 505 897 539
rect 845 471 897 505
rect 845 437 854 471
rect 888 437 897 471
rect 845 421 897 437
rect 938 589 983 605
rect 938 555 940 589
rect 974 555 983 589
rect 938 510 983 555
rect 938 476 940 510
rect 974 476 983 510
rect 938 431 983 476
rect 759 385 811 402
rect 938 390 940 431
rect 974 390 983 431
rect 1017 599 1069 649
rect 1017 565 1026 599
rect 1060 565 1069 599
rect 1017 520 1069 565
rect 1017 486 1026 520
rect 1060 486 1069 520
rect 1017 441 1069 486
rect 1017 407 1026 441
rect 1060 407 1069 441
rect 1017 391 1069 407
rect 1103 589 1155 605
rect 1103 555 1112 589
rect 1146 555 1155 589
rect 1103 510 1155 555
rect 1103 476 1112 510
rect 1146 476 1155 510
rect 1103 431 1155 476
rect 418 351 904 385
rect 868 350 904 351
rect 350 315 834 317
rect 350 281 376 315
rect 410 281 444 315
rect 478 281 512 315
rect 546 281 580 315
rect 614 281 648 315
rect 682 281 716 315
rect 750 281 784 315
rect 818 281 834 315
rect 350 279 834 281
rect 868 316 870 350
rect 350 249 384 279
rect 55 215 384 249
rect 868 245 904 316
rect 55 187 114 215
rect 55 153 71 187
rect 105 153 114 187
rect 234 187 286 215
rect 55 113 114 153
rect 55 79 71 113
rect 105 79 114 113
rect 55 63 114 79
rect 148 165 200 181
rect 148 131 157 165
rect 191 131 200 165
rect 148 97 200 131
rect 148 63 157 97
rect 191 63 200 97
rect 234 153 243 187
rect 277 153 286 187
rect 418 211 904 245
rect 418 187 467 211
rect 234 113 286 153
rect 234 79 243 113
rect 277 79 286 113
rect 234 63 286 79
rect 320 165 374 181
rect 320 131 329 165
rect 363 131 374 165
rect 320 97 374 131
rect 320 63 329 97
rect 363 63 374 97
rect 418 153 424 187
rect 458 153 467 187
rect 587 187 639 211
rect 418 113 467 153
rect 418 79 424 113
rect 458 79 467 113
rect 418 63 467 79
rect 501 161 553 177
rect 501 127 510 161
rect 544 127 553 161
rect 501 93 553 127
rect 148 17 200 63
rect 320 17 374 63
rect 501 59 510 93
rect 544 59 553 93
rect 587 153 596 187
rect 630 153 639 187
rect 759 187 811 211
rect 587 113 639 153
rect 587 79 596 113
rect 630 79 639 113
rect 587 63 639 79
rect 673 161 725 177
rect 673 127 682 161
rect 716 127 725 161
rect 673 93 725 127
rect 501 17 553 59
rect 673 59 682 93
rect 716 59 725 93
rect 759 153 768 187
rect 802 153 811 187
rect 938 187 983 390
rect 1103 390 1112 431
rect 1146 390 1155 431
rect 1189 599 1241 649
rect 1189 565 1198 599
rect 1232 565 1241 599
rect 1189 520 1241 565
rect 1189 486 1198 520
rect 1232 486 1241 520
rect 1189 441 1241 486
rect 1189 407 1198 441
rect 1232 407 1241 441
rect 1189 391 1241 407
rect 1275 589 1327 605
rect 1275 555 1284 589
rect 1318 555 1327 589
rect 1275 510 1327 555
rect 1275 476 1284 510
rect 1318 476 1327 510
rect 1275 431 1327 476
rect 1017 350 1069 357
rect 1017 285 1026 350
rect 1060 285 1069 350
rect 1017 269 1069 285
rect 759 113 811 153
rect 759 79 768 113
rect 802 79 811 113
rect 759 63 811 79
rect 845 161 897 177
rect 845 127 854 161
rect 888 127 897 161
rect 845 93 897 127
rect 673 17 725 59
rect 845 59 854 93
rect 888 59 897 93
rect 938 153 940 187
rect 974 153 983 187
rect 938 113 983 153
rect 938 79 940 113
rect 974 79 983 113
rect 938 63 983 79
rect 1017 187 1069 216
rect 1017 153 1026 187
rect 1060 153 1069 187
rect 1017 113 1069 153
rect 1017 79 1026 113
rect 1060 79 1069 113
rect 845 17 897 59
rect 1017 17 1069 79
rect 1103 187 1155 390
rect 1275 390 1284 431
rect 1318 390 1327 431
rect 1361 599 1413 649
rect 1361 565 1370 599
rect 1404 565 1413 599
rect 1361 520 1413 565
rect 1361 486 1370 520
rect 1404 486 1413 520
rect 1361 441 1413 486
rect 1361 407 1370 441
rect 1404 407 1413 441
rect 1361 391 1413 407
rect 1447 589 1499 605
rect 1447 555 1456 589
rect 1490 555 1499 589
rect 1447 510 1499 555
rect 1447 476 1456 510
rect 1490 476 1499 510
rect 1447 431 1499 476
rect 1189 350 1241 357
rect 1189 285 1198 350
rect 1232 285 1241 350
rect 1189 269 1241 285
rect 1103 153 1112 187
rect 1146 153 1155 187
rect 1103 113 1155 153
rect 1103 79 1112 113
rect 1146 79 1155 113
rect 1103 63 1155 79
rect 1189 187 1241 216
rect 1189 153 1198 187
rect 1232 153 1241 187
rect 1189 113 1241 153
rect 1189 79 1198 113
rect 1232 79 1241 113
rect 1189 17 1241 79
rect 1275 187 1327 390
rect 1447 390 1456 431
rect 1490 390 1499 431
rect 1533 599 1585 649
rect 1533 565 1542 599
rect 1576 565 1585 599
rect 1533 520 1585 565
rect 1533 486 1542 520
rect 1576 486 1585 520
rect 1533 441 1585 486
rect 1533 407 1542 441
rect 1576 407 1585 441
rect 1533 391 1585 407
rect 1619 589 1671 605
rect 1619 555 1628 589
rect 1662 555 1671 589
rect 1619 510 1671 555
rect 1619 476 1628 510
rect 1662 476 1671 510
rect 1619 431 1671 476
rect 1361 350 1413 357
rect 1361 285 1370 350
rect 1404 285 1413 350
rect 1361 269 1413 285
rect 1275 153 1284 187
rect 1318 153 1327 187
rect 1275 113 1327 153
rect 1275 79 1284 113
rect 1318 79 1327 113
rect 1275 63 1327 79
rect 1361 187 1413 216
rect 1361 153 1370 187
rect 1404 153 1413 187
rect 1361 113 1413 153
rect 1361 79 1370 113
rect 1404 79 1413 113
rect 1361 17 1413 79
rect 1447 187 1499 390
rect 1619 390 1628 431
rect 1662 390 1671 431
rect 1705 599 1757 649
rect 1705 565 1714 599
rect 1748 565 1757 599
rect 1705 520 1757 565
rect 1705 486 1714 520
rect 1748 486 1757 520
rect 1705 441 1757 486
rect 1705 407 1714 441
rect 1748 407 1757 441
rect 1705 391 1757 407
rect 1791 589 1843 605
rect 1791 555 1800 589
rect 1834 555 1843 589
rect 1791 510 1843 555
rect 1791 476 1800 510
rect 1834 476 1843 510
rect 1791 431 1843 476
rect 1533 350 1585 357
rect 1533 285 1542 350
rect 1576 285 1585 350
rect 1533 269 1585 285
rect 1447 153 1456 187
rect 1490 153 1499 187
rect 1447 113 1499 153
rect 1447 79 1456 113
rect 1490 79 1499 113
rect 1447 63 1499 79
rect 1533 187 1585 216
rect 1533 153 1542 187
rect 1576 153 1585 187
rect 1533 113 1585 153
rect 1533 79 1542 113
rect 1576 79 1585 113
rect 1533 17 1585 79
rect 1619 187 1671 390
rect 1791 390 1800 431
rect 1834 390 1843 431
rect 1877 599 1929 649
rect 1877 565 1886 599
rect 1920 565 1929 599
rect 1877 520 1929 565
rect 1877 486 1886 520
rect 1920 486 1929 520
rect 1877 441 1929 486
rect 1877 407 1886 441
rect 1920 407 1929 441
rect 1877 391 1929 407
rect 1963 589 2015 605
rect 1963 555 1972 589
rect 2006 555 2015 589
rect 1963 510 2015 555
rect 1963 476 1972 510
rect 2006 476 2015 510
rect 1963 431 2015 476
rect 1705 350 1757 357
rect 1705 285 1714 350
rect 1748 285 1757 350
rect 1705 269 1757 285
rect 1619 153 1628 187
rect 1662 153 1671 187
rect 1619 113 1671 153
rect 1619 79 1628 113
rect 1662 79 1671 113
rect 1619 63 1671 79
rect 1705 187 1757 216
rect 1705 153 1714 187
rect 1748 153 1757 187
rect 1705 113 1757 153
rect 1705 79 1714 113
rect 1748 79 1757 113
rect 1705 17 1757 79
rect 1791 187 1843 390
rect 1963 390 1972 431
rect 2006 390 2015 431
rect 2049 599 2101 649
rect 2049 565 2058 599
rect 2092 565 2101 599
rect 2049 520 2101 565
rect 2049 486 2058 520
rect 2092 486 2101 520
rect 2049 441 2101 486
rect 2049 407 2058 441
rect 2092 407 2101 441
rect 2049 391 2101 407
rect 2135 589 2187 605
rect 2135 555 2144 589
rect 2178 555 2187 589
rect 2135 510 2187 555
rect 2135 476 2144 510
rect 2178 476 2187 510
rect 2135 431 2187 476
rect 1877 350 1929 357
rect 1877 285 1886 350
rect 1920 285 1929 350
rect 1877 269 1929 285
rect 1791 153 1800 187
rect 1834 153 1843 187
rect 1791 113 1843 153
rect 1791 79 1800 113
rect 1834 79 1843 113
rect 1791 63 1843 79
rect 1877 187 1929 216
rect 1877 153 1886 187
rect 1920 153 1929 187
rect 1877 113 1929 153
rect 1877 79 1886 113
rect 1920 79 1929 113
rect 1877 17 1929 79
rect 1963 187 2015 390
rect 2135 390 2144 431
rect 2178 390 2187 431
rect 2221 599 2280 649
rect 2221 565 2230 599
rect 2264 565 2280 599
rect 2221 520 2280 565
rect 2221 486 2230 520
rect 2264 486 2280 520
rect 2221 441 2280 486
rect 2221 407 2230 441
rect 2264 407 2280 441
rect 2221 391 2280 407
rect 2049 350 2101 357
rect 2049 285 2058 350
rect 2092 285 2101 350
rect 2049 269 2101 285
rect 1963 153 1972 187
rect 2006 153 2015 187
rect 1963 113 2015 153
rect 1963 79 1972 113
rect 2006 79 2015 113
rect 1963 63 2015 79
rect 2049 187 2101 216
rect 2049 153 2058 187
rect 2092 153 2101 187
rect 2049 113 2101 153
rect 2049 79 2058 113
rect 2092 79 2101 113
rect 2049 17 2101 79
rect 2135 187 2187 390
rect 2135 153 2144 187
rect 2178 153 2187 187
rect 2135 113 2187 153
rect 2135 79 2144 113
rect 2178 79 2187 113
rect 2135 63 2187 79
rect 2221 187 2280 216
rect 2221 153 2230 187
rect 2264 153 2280 187
rect 2221 113 2280 153
rect 2221 79 2230 113
rect 2264 79 2280 113
rect 2221 17 2280 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 940 397 974 424
rect 940 390 974 397
rect 870 316 904 350
rect 1112 397 1146 424
rect 1112 390 1146 397
rect 1026 319 1060 350
rect 1026 316 1060 319
rect 1284 397 1318 424
rect 1284 390 1318 397
rect 1198 319 1232 350
rect 1198 316 1232 319
rect 1456 397 1490 424
rect 1456 390 1490 397
rect 1370 319 1404 350
rect 1370 316 1404 319
rect 1628 397 1662 424
rect 1628 390 1662 397
rect 1542 319 1576 350
rect 1542 316 1576 319
rect 1800 397 1834 424
rect 1800 390 1834 397
rect 1714 319 1748 350
rect 1714 316 1748 319
rect 1972 397 2006 424
rect 1972 390 2006 397
rect 1886 319 1920 350
rect 1886 316 1920 319
rect 2144 397 2178 424
rect 2144 390 2178 397
rect 2058 319 2092 350
rect 2058 316 2092 319
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 928 424 2190 430
rect 928 390 940 424
rect 974 390 1112 424
rect 1146 390 1284 424
rect 1318 390 1456 424
rect 1490 390 1628 424
rect 1662 390 1800 424
rect 1834 390 1972 424
rect 2006 390 2144 424
rect 2178 390 2190 424
rect 928 384 2190 390
rect 858 350 2104 356
rect 858 316 870 350
rect 904 316 1026 350
rect 1060 316 1198 350
rect 1232 316 1370 350
rect 1404 316 1542 350
rect 1576 316 1714 350
rect 1748 316 1886 350
rect 1920 316 2058 350
rect 2092 316 2104 350
rect 858 310 2104 316
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
flabel pwell s 0 0 2304 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 2304 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 bufinv_16
flabel metal1 s 928 384 2190 430 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel metal1 s 0 617 2304 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 2304 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2304 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1612580
string GDS_START 1593036
<< end >>
