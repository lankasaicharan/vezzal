magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 70 241 438 243
rect 70 49 808 241
rect 0 0 864 49
<< scnmos >>
rect 149 49 179 217
rect 243 49 273 217
rect 329 49 359 217
rect 519 47 549 215
rect 605 47 635 215
rect 699 47 729 215
<< scpmoshvt >>
rect 149 367 179 619
rect 257 367 287 619
rect 335 367 365 619
rect 519 367 549 619
rect 591 367 621 619
rect 706 367 736 619
<< ndiff >>
rect 96 205 149 217
rect 96 171 104 205
rect 138 171 149 205
rect 96 101 149 171
rect 96 67 104 101
rect 138 67 149 101
rect 96 49 149 67
rect 179 167 243 217
rect 179 133 196 167
rect 230 133 243 167
rect 179 95 243 133
rect 179 61 196 95
rect 230 61 243 95
rect 179 49 243 61
rect 273 169 329 217
rect 273 135 284 169
rect 318 135 329 169
rect 273 49 329 135
rect 359 127 412 217
rect 359 93 370 127
rect 404 93 412 127
rect 359 49 412 93
rect 466 127 519 215
rect 466 93 474 127
rect 508 93 519 127
rect 466 47 519 93
rect 549 185 605 215
rect 549 151 560 185
rect 594 151 605 185
rect 549 101 605 151
rect 549 67 560 101
rect 594 67 605 101
rect 549 47 605 67
rect 635 187 699 215
rect 635 153 646 187
rect 680 153 699 187
rect 635 93 699 153
rect 635 59 646 93
rect 680 59 699 93
rect 635 47 699 59
rect 729 187 782 215
rect 729 153 740 187
rect 774 153 782 187
rect 729 101 782 153
rect 729 67 740 101
rect 774 67 782 101
rect 729 47 782 67
<< pdiff >>
rect 96 599 149 619
rect 96 565 104 599
rect 138 565 149 599
rect 96 515 149 565
rect 96 481 104 515
rect 138 481 149 515
rect 96 436 149 481
rect 96 402 104 436
rect 138 402 149 436
rect 96 367 149 402
rect 179 607 257 619
rect 179 573 201 607
rect 235 573 257 607
rect 179 492 257 573
rect 179 458 201 492
rect 235 458 257 492
rect 179 367 257 458
rect 287 367 335 619
rect 365 599 519 619
rect 365 565 376 599
rect 410 565 474 599
rect 508 565 519 599
rect 365 506 519 565
rect 365 472 376 506
rect 410 472 474 506
rect 508 472 519 506
rect 365 413 519 472
rect 365 379 376 413
rect 410 379 474 413
rect 508 379 519 413
rect 365 367 519 379
rect 549 367 591 619
rect 621 607 706 619
rect 621 573 644 607
rect 678 573 706 607
rect 621 525 706 573
rect 621 491 644 525
rect 678 491 706 525
rect 621 441 706 491
rect 621 407 644 441
rect 678 407 706 441
rect 621 367 706 407
rect 736 599 793 619
rect 736 565 747 599
rect 781 565 793 599
rect 736 504 793 565
rect 736 470 747 504
rect 781 470 793 504
rect 736 413 793 470
rect 736 379 747 413
rect 781 379 793 413
rect 736 367 793 379
<< ndiffc >>
rect 104 171 138 205
rect 104 67 138 101
rect 196 133 230 167
rect 196 61 230 95
rect 284 135 318 169
rect 370 93 404 127
rect 474 93 508 127
rect 560 151 594 185
rect 560 67 594 101
rect 646 153 680 187
rect 646 59 680 93
rect 740 153 774 187
rect 740 67 774 101
<< pdiffc >>
rect 104 565 138 599
rect 104 481 138 515
rect 104 402 138 436
rect 201 573 235 607
rect 201 458 235 492
rect 376 565 410 599
rect 474 565 508 599
rect 376 472 410 506
rect 474 472 508 506
rect 376 379 410 413
rect 474 379 508 413
rect 644 573 678 607
rect 644 491 678 525
rect 644 407 678 441
rect 747 565 781 599
rect 747 470 781 504
rect 747 379 781 413
<< poly >>
rect 149 619 179 645
rect 257 619 287 645
rect 335 619 365 645
rect 519 619 549 645
rect 591 619 621 645
rect 706 619 736 645
rect 149 335 179 367
rect 51 319 179 335
rect 51 285 67 319
rect 101 285 179 319
rect 257 308 287 367
rect 51 269 179 285
rect 149 217 179 269
rect 221 292 287 308
rect 335 305 365 367
rect 221 258 237 292
rect 271 258 287 292
rect 221 242 287 258
rect 329 289 397 305
rect 519 303 549 367
rect 329 255 347 289
rect 381 255 397 289
rect 243 217 273 242
rect 329 239 397 255
rect 461 287 549 303
rect 461 253 486 287
rect 520 253 549 287
rect 329 217 359 239
rect 461 237 549 253
rect 591 303 621 367
rect 706 303 736 367
rect 591 287 657 303
rect 591 253 607 287
rect 641 253 657 287
rect 591 237 657 253
rect 699 287 778 303
rect 699 253 717 287
rect 751 253 778 287
rect 699 237 778 253
rect 519 215 549 237
rect 605 215 635 237
rect 699 215 729 237
rect 149 23 179 49
rect 243 23 273 49
rect 329 23 359 49
rect 519 21 549 47
rect 605 21 635 47
rect 699 21 729 47
<< polycont >>
rect 67 285 101 319
rect 237 258 271 292
rect 347 255 381 289
rect 486 253 520 287
rect 607 253 641 287
rect 717 253 751 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 99 599 151 615
rect 99 565 104 599
rect 138 565 151 599
rect 99 515 151 565
rect 17 350 65 515
rect 99 481 104 515
rect 138 481 151 515
rect 99 436 151 481
rect 185 607 251 649
rect 185 573 201 607
rect 235 573 251 607
rect 185 492 251 573
rect 185 458 201 492
rect 235 458 251 492
rect 185 454 251 458
rect 360 599 526 615
rect 360 565 376 599
rect 410 565 474 599
rect 508 565 526 599
rect 360 506 526 565
rect 360 472 376 506
rect 410 472 474 506
rect 508 472 526 506
rect 99 402 104 436
rect 138 420 151 436
rect 360 420 526 472
rect 138 413 526 420
rect 138 402 376 413
rect 99 386 376 402
rect 17 319 113 350
rect 17 285 67 319
rect 101 285 113 319
rect 17 269 113 285
rect 17 151 65 269
rect 153 235 187 386
rect 360 379 376 386
rect 410 379 474 413
rect 508 379 526 413
rect 628 607 694 649
rect 628 573 644 607
rect 678 573 694 607
rect 628 525 694 573
rect 628 491 644 525
rect 678 491 694 525
rect 628 441 694 491
rect 628 407 644 441
rect 678 407 694 441
rect 731 599 847 615
rect 731 565 747 599
rect 781 565 847 599
rect 731 504 847 565
rect 731 470 747 504
rect 781 470 847 504
rect 731 413 847 470
rect 731 405 747 413
rect 360 373 526 379
rect 781 379 847 413
rect 221 292 277 350
rect 360 339 713 373
rect 747 339 847 379
rect 221 258 237 292
rect 271 258 277 292
rect 221 242 277 258
rect 313 289 381 305
rect 679 303 713 339
rect 313 255 347 289
rect 313 239 381 255
rect 415 287 555 303
rect 415 253 486 287
rect 520 253 555 287
rect 415 237 555 253
rect 591 287 645 303
rect 591 253 607 287
rect 641 253 645 287
rect 591 237 645 253
rect 679 287 751 303
rect 679 253 717 287
rect 679 237 751 253
rect 99 205 187 235
rect 99 171 104 205
rect 138 201 187 205
rect 785 203 847 339
rect 138 171 146 201
rect 99 101 146 171
rect 280 185 596 203
rect 280 169 560 185
rect 99 67 104 101
rect 138 67 146 101
rect 99 51 146 67
rect 180 133 196 167
rect 230 133 246 167
rect 180 95 246 133
rect 280 135 284 169
rect 318 135 320 169
rect 558 151 560 169
rect 594 151 596 185
rect 280 119 320 135
rect 354 127 420 135
rect 180 61 196 95
rect 230 85 246 95
rect 354 93 370 127
rect 404 93 420 127
rect 354 85 420 93
rect 230 61 420 85
rect 180 51 420 61
rect 458 127 524 135
rect 458 93 474 127
rect 508 93 524 127
rect 458 17 524 93
rect 558 101 596 151
rect 558 67 560 101
rect 594 67 596 101
rect 558 51 596 67
rect 630 187 696 203
rect 630 153 646 187
rect 680 153 696 187
rect 630 93 696 153
rect 630 59 646 93
rect 680 59 696 93
rect 630 17 696 59
rect 730 187 847 203
rect 730 153 740 187
rect 774 153 847 187
rect 730 101 847 153
rect 730 67 740 101
rect 774 67 847 101
rect 730 51 847 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221a_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4810038
string GDS_START 4801084
<< end >>
