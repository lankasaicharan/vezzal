magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
rect 563 299 731 331
<< pwell >>
rect 555 167 1093 211
rect 271 157 1093 167
rect 1 49 2015 157
rect 0 0 2016 49
<< scnmos >>
rect 84 47 114 131
rect 156 47 186 131
rect 354 57 384 141
rect 440 57 470 141
rect 654 101 684 185
rect 726 101 756 185
rect 885 101 915 185
rect 980 101 1010 185
rect 1082 47 1112 131
rect 1160 47 1190 131
rect 1384 47 1414 131
rect 1462 47 1492 131
rect 1570 47 1600 131
rect 1744 47 1774 131
rect 1830 47 1860 131
rect 1902 47 1932 131
<< scpmoshvt >>
rect 84 409 134 609
rect 320 411 370 611
rect 465 411 515 611
rect 710 419 760 619
rect 848 419 898 619
rect 946 419 996 619
rect 1160 419 1210 619
rect 1271 419 1321 619
rect 1383 419 1433 619
rect 1481 419 1531 619
rect 1642 419 1692 619
rect 1750 419 1800 619
rect 1858 419 1908 619
<< ndiff >>
rect 581 173 654 185
rect 27 111 84 131
rect 27 77 39 111
rect 73 77 84 111
rect 27 47 84 77
rect 114 47 156 131
rect 186 93 243 131
rect 186 59 197 93
rect 231 59 243 93
rect 186 47 243 59
rect 297 116 354 141
rect 297 82 309 116
rect 343 82 354 116
rect 297 57 354 82
rect 384 116 440 141
rect 384 82 395 116
rect 429 82 440 116
rect 384 57 440 82
rect 470 116 527 141
rect 470 82 481 116
rect 515 82 527 116
rect 581 139 593 173
rect 627 139 654 173
rect 581 101 654 139
rect 684 101 726 185
rect 756 160 885 185
rect 756 126 767 160
rect 801 126 885 160
rect 756 101 885 126
rect 915 101 980 185
rect 1010 173 1067 185
rect 1010 139 1021 173
rect 1055 139 1067 173
rect 1010 131 1067 139
rect 1010 101 1082 131
rect 470 57 527 82
rect 1032 47 1082 101
rect 1112 47 1160 131
rect 1190 93 1384 131
rect 1190 59 1323 93
rect 1357 59 1384 93
rect 1190 47 1384 59
rect 1414 47 1462 131
rect 1492 111 1570 131
rect 1492 77 1525 111
rect 1559 77 1570 111
rect 1492 47 1570 77
rect 1600 47 1744 131
rect 1774 106 1830 131
rect 1774 72 1785 106
rect 1819 72 1830 106
rect 1774 47 1830 72
rect 1860 47 1902 131
rect 1932 111 1989 131
rect 1932 77 1943 111
rect 1977 77 1989 111
rect 1932 47 1989 77
<< pdiff >>
rect 775 623 833 635
rect 775 619 787 623
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 191 609
rect 134 563 145 597
rect 179 563 191 597
rect 134 516 191 563
rect 134 482 145 516
rect 179 482 191 516
rect 134 409 191 482
rect 245 597 320 611
rect 245 563 257 597
rect 291 563 320 597
rect 245 527 320 563
rect 245 493 257 527
rect 291 493 320 527
rect 245 457 320 493
rect 245 423 257 457
rect 291 423 320 457
rect 245 411 320 423
rect 370 457 465 611
rect 370 423 397 457
rect 431 423 465 457
rect 370 411 465 423
rect 515 505 583 611
rect 515 471 537 505
rect 571 471 583 505
rect 515 411 583 471
rect 637 419 710 619
rect 760 589 787 619
rect 821 619 833 623
rect 821 589 848 619
rect 760 419 848 589
rect 898 419 946 619
rect 996 597 1160 619
rect 996 563 1007 597
rect 1041 563 1160 597
rect 996 469 1160 563
rect 996 435 1007 469
rect 1041 435 1160 469
rect 996 419 1160 435
rect 1210 419 1271 619
rect 1321 607 1383 619
rect 1321 573 1332 607
rect 1366 573 1383 607
rect 1321 508 1383 573
rect 1321 474 1332 508
rect 1366 474 1383 508
rect 1321 419 1383 474
rect 1433 419 1481 619
rect 1531 457 1642 619
rect 1531 423 1558 457
rect 1592 423 1642 457
rect 1531 419 1642 423
rect 1692 419 1750 619
rect 1800 596 1858 619
rect 1800 562 1813 596
rect 1847 562 1858 596
rect 1800 419 1858 562
rect 1908 597 1965 619
rect 1908 563 1919 597
rect 1953 563 1965 597
rect 1908 516 1965 563
rect 1908 482 1919 516
rect 1953 482 1965 516
rect 1908 419 1965 482
rect 637 381 695 419
rect 637 347 649 381
rect 683 347 695 381
rect 637 335 695 347
rect 1546 411 1604 419
<< ndiffc >>
rect 39 77 73 111
rect 197 59 231 93
rect 309 82 343 116
rect 395 82 429 116
rect 481 82 515 116
rect 593 139 627 173
rect 767 126 801 160
rect 1021 139 1055 173
rect 1323 59 1357 93
rect 1525 77 1559 111
rect 1785 72 1819 106
rect 1943 77 1977 111
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 482 179 516
rect 257 563 291 597
rect 257 493 291 527
rect 257 423 291 457
rect 397 423 431 457
rect 537 471 571 505
rect 787 589 821 623
rect 1007 563 1041 597
rect 1007 435 1041 469
rect 1332 573 1366 607
rect 1332 474 1366 508
rect 1558 423 1592 457
rect 1813 562 1847 596
rect 1919 563 1953 597
rect 1919 482 1953 516
rect 649 347 683 381
<< poly >>
rect 84 609 134 635
rect 320 611 370 637
rect 465 611 515 637
rect 710 619 760 645
rect 848 619 898 645
rect 946 619 996 645
rect 1160 619 1210 645
rect 1271 619 1321 645
rect 1383 619 1433 645
rect 1481 619 1531 645
rect 1642 619 1692 645
rect 1750 619 1800 645
rect 1858 619 1908 645
rect 84 252 134 409
rect 320 396 370 411
rect 320 366 417 396
rect 465 378 515 411
rect 206 344 272 360
rect 206 310 222 344
rect 256 324 272 344
rect 256 310 339 324
rect 206 294 339 310
rect 84 236 261 252
rect 84 222 211 236
rect 84 131 114 222
rect 195 202 211 222
rect 245 202 261 236
rect 195 186 261 202
rect 309 186 339 294
rect 387 264 417 366
rect 485 362 551 378
rect 485 328 501 362
rect 535 342 551 362
rect 535 328 605 342
rect 485 320 605 328
rect 710 320 760 419
rect 848 376 898 419
rect 485 312 760 320
rect 575 290 760 312
rect 804 360 898 376
rect 804 326 820 360
rect 854 326 898 360
rect 804 310 898 326
rect 946 383 996 419
rect 946 367 1043 383
rect 946 333 993 367
rect 1027 347 1043 367
rect 1160 352 1210 419
rect 1027 333 1112 347
rect 946 317 1112 333
rect 387 248 533 264
rect 387 234 483 248
rect 440 214 483 234
rect 517 214 533 248
rect 440 198 533 214
rect 654 230 684 290
rect 868 230 898 310
rect 974 259 1040 275
rect 654 200 756 230
rect 868 200 915 230
rect 974 225 990 259
rect 1024 225 1040 259
rect 974 209 1040 225
rect 195 176 225 186
rect 156 146 225 176
rect 309 156 384 186
rect 156 131 186 146
rect 354 141 384 156
rect 440 141 470 198
rect 654 185 684 200
rect 726 185 756 200
rect 885 185 915 200
rect 980 185 1010 209
rect 1082 131 1112 317
rect 1160 336 1229 352
rect 1160 302 1179 336
rect 1213 302 1229 336
rect 1160 286 1229 302
rect 1271 330 1321 419
rect 1383 330 1433 419
rect 1481 360 1531 419
rect 1642 387 1692 419
rect 1636 371 1702 387
rect 1481 330 1594 360
rect 1271 219 1301 330
rect 1383 282 1413 330
rect 1154 203 1301 219
rect 1348 266 1414 282
rect 1348 232 1364 266
rect 1398 232 1414 266
rect 1348 216 1414 232
rect 1456 266 1522 282
rect 1456 232 1472 266
rect 1506 232 1522 266
rect 1456 216 1522 232
rect 1564 219 1594 330
rect 1636 337 1652 371
rect 1686 337 1702 371
rect 1636 321 1702 337
rect 1750 300 1800 419
rect 1858 387 1908 419
rect 1858 371 1924 387
rect 1858 337 1874 371
rect 1908 337 1924 371
rect 1858 321 1924 337
rect 1744 284 1810 300
rect 1744 250 1760 284
rect 1794 250 1810 284
rect 1744 234 1810 250
rect 1154 169 1170 203
rect 1204 189 1301 203
rect 1204 169 1220 189
rect 1154 153 1220 169
rect 1160 131 1190 153
rect 1384 131 1414 216
rect 1462 131 1492 216
rect 1564 203 1694 219
rect 1564 189 1644 203
rect 1570 169 1644 189
rect 1678 169 1694 203
rect 1570 153 1694 169
rect 1570 131 1600 153
rect 1744 131 1774 234
rect 1858 176 1888 321
rect 1830 146 1932 176
rect 1830 131 1860 146
rect 1902 131 1932 146
rect 654 75 684 101
rect 726 75 756 101
rect 885 75 915 101
rect 980 75 1010 101
rect 84 21 114 47
rect 156 21 186 47
rect 354 31 384 57
rect 440 31 470 57
rect 1082 21 1112 47
rect 1160 21 1190 47
rect 1384 21 1414 47
rect 1462 21 1492 47
rect 1570 21 1600 47
rect 1744 21 1774 47
rect 1830 21 1860 47
rect 1902 21 1932 47
<< polycont >>
rect 222 310 256 344
rect 211 202 245 236
rect 501 328 535 362
rect 820 326 854 360
rect 993 333 1027 367
rect 483 214 517 248
rect 990 225 1024 259
rect 1179 302 1213 336
rect 1364 232 1398 266
rect 1472 232 1506 266
rect 1652 337 1686 371
rect 1874 337 1908 371
rect 1760 250 1794 284
rect 1170 169 1204 203
rect 1644 169 1678 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 526 89 563
rect 23 492 39 526
rect 73 492 89 526
rect 23 455 89 492
rect 129 597 195 649
rect 771 623 837 649
rect 129 563 145 597
rect 179 563 195 597
rect 129 516 195 563
rect 129 482 145 516
rect 179 482 195 516
rect 129 466 195 482
rect 241 597 657 613
rect 241 563 257 597
rect 291 579 657 597
rect 241 527 291 563
rect 241 493 257 527
rect 23 421 39 455
rect 73 421 89 455
rect 241 457 291 493
rect 241 430 257 457
rect 23 111 89 421
rect 125 423 257 430
rect 125 396 291 423
rect 327 509 501 543
rect 125 163 159 396
rect 327 360 361 509
rect 206 344 361 360
rect 206 310 222 344
rect 256 310 361 344
rect 206 294 361 310
rect 397 457 431 473
rect 397 252 431 423
rect 467 378 501 509
rect 537 505 587 543
rect 571 471 587 505
rect 623 537 657 579
rect 771 589 787 623
rect 821 589 837 623
rect 771 573 837 589
rect 991 597 1057 613
rect 991 563 1007 597
rect 1041 563 1057 597
rect 991 537 1057 563
rect 623 503 1057 537
rect 537 467 587 471
rect 537 433 753 467
rect 609 381 683 397
rect 467 362 551 378
rect 467 328 501 362
rect 535 328 551 362
rect 467 310 551 328
rect 609 347 649 381
rect 609 331 683 347
rect 609 264 643 331
rect 195 236 431 252
rect 195 202 211 236
rect 245 202 431 236
rect 195 199 431 202
rect 467 248 643 264
rect 719 259 753 433
rect 793 360 870 430
rect 793 326 820 360
rect 854 326 870 360
rect 793 310 870 326
rect 467 214 483 248
rect 517 214 643 248
rect 125 129 359 163
rect 23 77 39 111
rect 73 77 89 111
rect 293 116 359 129
rect 23 53 89 77
rect 181 59 197 93
rect 231 59 247 93
rect 181 17 247 59
rect 293 82 309 116
rect 343 82 359 116
rect 293 53 359 82
rect 395 116 429 199
rect 467 198 643 214
rect 577 173 643 198
rect 395 53 429 82
rect 465 116 531 145
rect 577 139 593 173
rect 627 139 643 173
rect 577 123 643 139
rect 679 225 871 259
rect 465 82 481 116
rect 515 87 531 116
rect 679 87 713 225
rect 515 82 713 87
rect 465 53 713 82
rect 751 160 801 189
rect 751 126 767 160
rect 751 17 801 126
rect 837 87 871 225
rect 907 173 941 503
rect 991 469 1057 503
rect 991 435 1007 469
rect 1041 435 1057 469
rect 1316 607 1382 649
rect 1316 573 1332 607
rect 1366 573 1382 607
rect 1316 508 1382 573
rect 1316 474 1332 508
rect 1366 474 1382 508
rect 1316 458 1382 474
rect 1418 579 1761 613
rect 991 419 1057 435
rect 1418 422 1452 579
rect 1093 388 1452 422
rect 1488 509 1670 543
rect 1093 383 1127 388
rect 977 367 1127 383
rect 977 333 993 367
rect 1027 349 1127 367
rect 1488 352 1522 509
rect 1027 333 1043 349
rect 977 317 1043 333
rect 1163 336 1229 352
rect 1163 302 1179 336
rect 1213 302 1229 336
rect 1163 289 1229 302
rect 1265 318 1522 352
rect 1265 289 1299 318
rect 1079 275 1299 289
rect 977 259 1299 275
rect 977 225 990 259
rect 1024 255 1299 259
rect 1348 266 1415 282
rect 1024 225 1113 255
rect 977 209 1113 225
rect 1348 232 1364 266
rect 1398 232 1415 266
rect 1154 203 1217 219
rect 1348 216 1415 232
rect 1456 266 1522 318
rect 1456 232 1472 266
rect 1506 232 1522 266
rect 1456 216 1522 232
rect 1558 457 1592 473
rect 907 139 1021 173
rect 1055 139 1071 173
rect 1154 169 1170 203
rect 1204 169 1217 203
rect 1558 180 1592 423
rect 1636 430 1670 509
rect 1727 500 1761 579
rect 1797 596 1863 649
rect 1797 562 1813 596
rect 1847 562 1863 596
rect 1797 536 1863 562
rect 1903 597 1994 613
rect 1903 563 1919 597
rect 1953 563 1994 597
rect 1903 516 1994 563
rect 1903 500 1919 516
rect 1727 482 1919 500
rect 1953 482 1994 516
rect 1727 466 1994 482
rect 1636 371 1924 430
rect 1636 337 1652 371
rect 1686 337 1874 371
rect 1908 337 1924 371
rect 1636 328 1924 337
rect 1657 284 1895 292
rect 1657 250 1760 284
rect 1794 250 1895 284
rect 1657 242 1895 250
rect 1960 206 1994 466
rect 1154 153 1217 169
rect 907 123 1071 139
rect 1253 146 1592 180
rect 1628 203 1994 206
rect 1628 169 1644 203
rect 1678 172 1994 203
rect 1678 169 1694 172
rect 1628 153 1694 169
rect 1253 87 1287 146
rect 1509 111 1592 146
rect 837 53 1287 87
rect 1323 93 1373 110
rect 1357 59 1373 93
rect 1323 17 1373 59
rect 1509 77 1525 111
rect 1559 77 1592 111
rect 1509 53 1592 77
rect 1769 106 1835 135
rect 1769 72 1785 106
rect 1819 72 1835 106
rect 1769 17 1835 72
rect 1927 111 1994 172
rect 1927 77 1943 111
rect 1977 77 1994 111
rect 1927 53 1994 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux4_lp
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 1663 390 1697 424 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 1759 390 1793 424 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 1855 390 1889 424 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 1183 168 1217 202 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1505652
string GDS_START 1491130
<< end >>
