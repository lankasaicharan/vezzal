magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 673 241 1151 263
rect 9 49 1151 241
rect 0 0 1152 49
<< scnmos >>
rect 88 47 118 215
rect 174 47 204 215
rect 260 47 290 215
rect 346 47 376 215
rect 432 47 462 215
rect 768 69 798 237
rect 854 69 884 237
rect 956 69 986 237
rect 1042 69 1072 237
<< scpmoshvt >>
rect 88 367 118 619
rect 354 367 384 619
rect 440 367 470 619
rect 526 367 556 619
rect 612 367 642 619
rect 768 367 798 619
rect 854 367 884 619
rect 956 367 986 619
rect 1042 367 1072 619
<< ndiff >>
rect 35 203 88 215
rect 35 169 43 203
rect 77 169 88 203
rect 35 101 88 169
rect 35 67 43 101
rect 77 67 88 101
rect 35 47 88 67
rect 118 207 174 215
rect 118 173 129 207
rect 163 173 174 207
rect 118 93 174 173
rect 118 59 129 93
rect 163 59 174 93
rect 118 47 174 59
rect 204 192 260 215
rect 204 158 215 192
rect 249 158 260 192
rect 204 101 260 158
rect 204 67 215 101
rect 249 67 260 101
rect 204 47 260 67
rect 290 133 346 215
rect 290 99 301 133
rect 335 99 346 133
rect 290 47 346 99
rect 376 192 432 215
rect 376 158 387 192
rect 421 158 432 192
rect 376 101 432 158
rect 376 67 387 101
rect 421 67 432 101
rect 376 47 432 67
rect 462 105 515 215
rect 699 225 768 237
rect 462 71 473 105
rect 507 71 515 105
rect 462 47 515 71
rect 699 191 707 225
rect 741 191 768 225
rect 699 157 768 191
rect 699 123 707 157
rect 741 123 768 157
rect 699 69 768 123
rect 798 179 854 237
rect 798 145 809 179
rect 843 145 854 179
rect 798 111 854 145
rect 798 77 809 111
rect 843 77 854 111
rect 798 69 854 77
rect 884 229 956 237
rect 884 195 909 229
rect 943 195 956 229
rect 884 157 956 195
rect 884 123 909 157
rect 943 123 956 157
rect 884 69 956 123
rect 986 227 1042 237
rect 986 193 997 227
rect 1031 193 1042 227
rect 986 111 1042 193
rect 986 77 997 111
rect 1031 77 1042 111
rect 986 69 1042 77
rect 1072 225 1125 237
rect 1072 191 1083 225
rect 1117 191 1125 225
rect 1072 115 1125 191
rect 1072 81 1083 115
rect 1117 81 1125 115
rect 1072 69 1125 81
<< pdiff >>
rect 35 599 88 619
rect 35 565 43 599
rect 77 565 88 599
rect 35 509 88 565
rect 35 475 43 509
rect 77 475 88 509
rect 35 413 88 475
rect 35 379 43 413
rect 77 379 88 413
rect 35 367 88 379
rect 118 607 171 619
rect 118 573 129 607
rect 163 573 171 607
rect 118 509 171 573
rect 118 475 129 509
rect 163 475 171 509
rect 118 413 171 475
rect 301 599 354 619
rect 301 565 309 599
rect 343 565 354 599
rect 301 509 354 565
rect 301 475 309 509
rect 343 475 354 509
rect 118 379 129 413
rect 163 379 171 413
rect 118 367 171 379
rect 301 413 354 475
rect 301 379 309 413
rect 343 379 354 413
rect 301 367 354 379
rect 384 607 440 619
rect 384 573 395 607
rect 429 573 440 607
rect 384 532 440 573
rect 384 498 395 532
rect 429 498 440 532
rect 384 453 440 498
rect 384 419 395 453
rect 429 419 440 453
rect 384 367 440 419
rect 470 599 526 619
rect 470 565 481 599
rect 515 565 526 599
rect 470 509 526 565
rect 470 475 481 509
rect 515 475 526 509
rect 470 413 526 475
rect 470 379 481 413
rect 515 379 526 413
rect 470 367 526 379
rect 556 607 612 619
rect 556 573 567 607
rect 601 573 612 607
rect 556 532 612 573
rect 556 498 567 532
rect 601 498 612 532
rect 556 455 612 498
rect 556 421 567 455
rect 601 421 612 455
rect 556 367 612 421
rect 642 599 768 619
rect 642 565 653 599
rect 687 565 723 599
rect 757 565 768 599
rect 642 517 768 565
rect 642 509 723 517
rect 642 475 653 509
rect 687 483 723 509
rect 757 483 768 517
rect 687 475 768 483
rect 642 434 768 475
rect 642 413 723 434
rect 642 379 653 413
rect 687 400 723 413
rect 757 400 768 434
rect 687 379 768 400
rect 642 367 768 379
rect 798 531 854 619
rect 798 497 809 531
rect 843 497 854 531
rect 798 436 854 497
rect 798 402 809 436
rect 843 402 854 436
rect 798 367 854 402
rect 884 599 956 619
rect 884 565 903 599
rect 937 565 956 599
rect 884 502 956 565
rect 884 468 903 502
rect 937 468 956 502
rect 884 367 956 468
rect 986 531 1042 619
rect 986 497 997 531
rect 1031 497 1042 531
rect 986 436 1042 497
rect 986 402 997 436
rect 1031 402 1042 436
rect 986 367 1042 402
rect 1072 599 1125 619
rect 1072 565 1083 599
rect 1117 565 1125 599
rect 1072 506 1125 565
rect 1072 472 1083 506
rect 1117 472 1125 506
rect 1072 413 1125 472
rect 1072 379 1083 413
rect 1117 379 1125 413
rect 1072 367 1125 379
<< ndiffc >>
rect 43 169 77 203
rect 43 67 77 101
rect 129 173 163 207
rect 129 59 163 93
rect 215 158 249 192
rect 215 67 249 101
rect 301 99 335 133
rect 387 158 421 192
rect 387 67 421 101
rect 473 71 507 105
rect 707 191 741 225
rect 707 123 741 157
rect 809 145 843 179
rect 809 77 843 111
rect 909 195 943 229
rect 909 123 943 157
rect 997 193 1031 227
rect 997 77 1031 111
rect 1083 191 1117 225
rect 1083 81 1117 115
<< pdiffc >>
rect 43 565 77 599
rect 43 475 77 509
rect 43 379 77 413
rect 129 573 163 607
rect 129 475 163 509
rect 309 565 343 599
rect 309 475 343 509
rect 129 379 163 413
rect 309 379 343 413
rect 395 573 429 607
rect 395 498 429 532
rect 395 419 429 453
rect 481 565 515 599
rect 481 475 515 509
rect 481 379 515 413
rect 567 573 601 607
rect 567 498 601 532
rect 567 421 601 455
rect 653 565 687 599
rect 723 565 757 599
rect 653 475 687 509
rect 723 483 757 517
rect 653 379 687 413
rect 723 400 757 434
rect 809 497 843 531
rect 809 402 843 436
rect 903 565 937 599
rect 903 468 937 502
rect 997 497 1031 531
rect 997 402 1031 436
rect 1083 565 1117 599
rect 1083 472 1117 506
rect 1083 379 1117 413
<< poly >>
rect 88 619 118 645
rect 354 619 384 645
rect 440 619 470 645
rect 526 619 556 645
rect 612 619 642 645
rect 768 619 798 645
rect 854 619 884 645
rect 956 619 986 645
rect 1042 619 1072 645
rect 203 433 269 449
rect 203 399 219 433
rect 253 399 269 433
rect 88 273 118 367
rect 203 365 269 399
rect 203 331 219 365
rect 253 345 269 365
rect 354 345 384 367
rect 440 345 470 367
rect 526 345 556 367
rect 612 345 642 367
rect 253 331 642 345
rect 768 335 798 367
rect 854 335 884 367
rect 956 335 986 367
rect 1042 335 1072 367
rect 203 315 642 331
rect 741 319 1072 335
rect 741 285 757 319
rect 791 285 825 319
rect 859 285 1072 319
rect 88 251 641 273
rect 741 269 1072 285
rect 88 237 591 251
rect 88 215 118 237
rect 174 215 204 237
rect 260 215 290 237
rect 346 215 376 237
rect 432 215 462 237
rect 575 217 591 237
rect 625 217 641 251
rect 768 237 798 269
rect 854 237 884 269
rect 956 237 986 269
rect 1042 237 1072 269
rect 575 201 641 217
rect 88 21 118 47
rect 174 21 204 47
rect 260 21 290 47
rect 346 21 376 47
rect 432 21 462 47
rect 768 43 798 69
rect 854 43 884 69
rect 956 43 986 69
rect 1042 43 1072 69
<< polycont >>
rect 219 399 253 433
rect 219 331 253 365
rect 757 285 791 319
rect 825 285 859 319
rect 591 217 625 251
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 27 599 86 615
rect 27 565 43 599
rect 77 565 86 599
rect 27 509 86 565
rect 27 475 43 509
rect 77 475 86 509
rect 27 413 86 475
rect 27 379 43 413
rect 77 379 86 413
rect 27 329 86 379
rect 120 607 179 649
rect 120 573 129 607
rect 163 573 179 607
rect 120 509 179 573
rect 120 475 129 509
rect 163 475 179 509
rect 120 413 179 475
rect 303 599 345 615
rect 303 565 309 599
rect 343 565 345 599
rect 303 509 345 565
rect 303 475 309 509
rect 343 475 345 509
rect 120 379 129 413
rect 163 379 179 413
rect 120 363 179 379
rect 213 433 269 449
rect 213 399 219 433
rect 253 399 269 433
rect 213 365 269 399
rect 213 331 219 365
rect 253 331 269 365
rect 303 413 345 475
rect 379 607 445 649
rect 379 573 395 607
rect 429 573 445 607
rect 379 532 445 573
rect 379 498 395 532
rect 429 498 445 532
rect 379 453 445 498
rect 379 419 395 453
rect 429 419 445 453
rect 479 599 517 615
rect 479 565 481 599
rect 515 565 517 599
rect 479 509 517 565
rect 479 475 481 509
rect 515 475 517 509
rect 303 379 309 413
rect 343 385 345 413
rect 479 413 517 475
rect 551 607 617 649
rect 551 573 567 607
rect 601 573 617 607
rect 551 532 617 573
rect 551 498 567 532
rect 601 498 617 532
rect 551 455 617 498
rect 551 421 567 455
rect 601 421 617 455
rect 651 599 1133 615
rect 651 565 653 599
rect 687 565 723 599
rect 757 581 903 599
rect 757 565 759 581
rect 651 517 759 565
rect 887 565 903 581
rect 937 581 1083 599
rect 937 565 953 581
rect 651 509 723 517
rect 651 475 653 509
rect 687 483 723 509
rect 757 483 759 517
rect 687 475 759 483
rect 651 434 759 475
rect 479 385 481 413
rect 343 379 481 385
rect 515 385 517 413
rect 651 413 723 434
rect 651 385 653 413
rect 515 379 653 385
rect 687 400 723 413
rect 757 400 759 434
rect 687 384 759 400
rect 793 531 853 547
rect 793 497 809 531
rect 843 497 853 531
rect 793 436 853 497
rect 887 502 953 565
rect 1079 565 1083 581
rect 1117 565 1133 599
rect 887 468 903 502
rect 937 468 953 502
rect 887 452 953 468
rect 987 531 1045 547
rect 987 497 997 531
rect 1031 497 1045 531
rect 793 402 809 436
rect 843 418 853 436
rect 987 436 1045 497
rect 987 418 997 436
rect 843 402 997 418
rect 1031 402 1045 436
rect 793 384 1045 402
rect 687 379 707 384
rect 303 351 707 379
rect 213 329 269 331
rect 27 284 269 329
rect 741 319 875 350
rect 27 203 86 284
rect 309 251 648 286
rect 741 285 757 319
rect 791 285 825 319
rect 859 285 875 319
rect 909 311 1045 384
rect 1079 506 1133 565
rect 1079 472 1083 506
rect 1117 472 1133 506
rect 1079 413 1133 472
rect 1079 379 1083 413
rect 1117 379 1133 413
rect 1079 363 1133 379
rect 909 277 1133 311
rect 909 251 959 277
rect 309 242 591 251
rect 27 169 43 203
rect 77 169 86 203
rect 27 101 86 169
rect 27 67 43 101
rect 77 67 86 101
rect 27 51 86 67
rect 120 207 172 223
rect 575 217 591 242
rect 625 217 648 251
rect 575 213 648 217
rect 691 229 959 251
rect 691 225 909 229
rect 120 173 129 207
rect 163 173 172 207
rect 120 93 172 173
rect 120 59 129 93
rect 163 59 172 93
rect 120 17 172 59
rect 206 192 541 208
rect 206 158 215 192
rect 249 174 387 192
rect 249 158 251 174
rect 206 101 251 158
rect 385 158 387 174
rect 421 179 541 192
rect 691 191 707 225
rect 741 217 909 225
rect 741 191 757 217
rect 421 158 638 179
rect 385 145 638 158
rect 206 67 215 101
rect 249 67 251 101
rect 206 51 251 67
rect 285 133 351 140
rect 285 99 301 133
rect 335 99 351 133
rect 285 17 351 99
rect 385 101 423 145
rect 385 67 387 101
rect 421 67 423 101
rect 385 51 423 67
rect 457 105 523 111
rect 457 71 473 105
rect 507 71 523 105
rect 457 17 523 71
rect 568 87 638 145
rect 691 157 757 191
rect 893 195 909 217
rect 943 195 959 229
rect 691 123 707 157
rect 741 123 757 157
rect 691 121 757 123
rect 793 145 809 179
rect 843 145 859 179
rect 793 111 859 145
rect 893 157 959 195
rect 893 123 909 157
rect 943 123 959 157
rect 993 227 1039 243
rect 993 193 997 227
rect 1031 193 1039 227
rect 793 87 809 111
rect 568 77 809 87
rect 843 87 859 111
rect 993 111 1039 193
rect 993 87 997 111
rect 843 77 997 87
rect 1031 77 1039 111
rect 568 53 1039 77
rect 1073 225 1133 277
rect 1073 191 1083 225
rect 1117 191 1133 225
rect 1073 115 1133 191
rect 1073 81 1083 115
rect 1117 81 1133 115
rect 1073 65 1133 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 einvp_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2841442
string GDS_START 2831826
<< end >>
