magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1288 -1260 2012 1741
use sky130_fd_pr__hvdfm1sd__example_55959141808233  sky130_fd_pr__hvdfm1sd__example_55959141808233_0
timestamp 1627201311
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180827  sky130_fd_pr__hvdfm1sd2__example_5595914180827_0
timestamp 1627201311
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180827  sky130_fd_pr__hvdfm1sd2__example_5595914180827_1
timestamp 1627201311
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180827  sky130_fd_pr__hvdfm1sd2__example_5595914180827_2
timestamp 1627201311
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180827  sky130_fd_pr__hvdfm1sd2__example_5595914180827_3
timestamp 1627201311
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd__example_55959141808240  sky130_fd_pr__dfm1sd__example_55959141808240_0
timestamp 1627201311
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 752 481 752 481 0 FreeSans 300 0 0 0 D
flabel comment s 596 481 596 481 0 FreeSans 300 0 0 0 S
flabel comment s 440 481 440 481 0 FreeSans 300 0 0 0 D
flabel comment s 284 481 284 481 0 FreeSans 300 0 0 0 S
flabel comment s 128 481 128 481 0 FreeSans 300 0 0 0 D
flabel comment s -28 481 -28 481 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 37234870
string GDS_START 37231882
<< end >>
