magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1778 1975
<< nwell >>
rect -38 331 518 704
<< pwell >>
rect 17 49 455 222
rect 0 0 480 49
<< scnmos >>
rect 100 112 130 196
rect 178 112 208 196
rect 264 112 294 196
rect 342 112 372 196
<< scpmoshvt >>
rect 84 374 134 574
rect 176 374 226 574
<< ndiff >>
rect 43 171 100 196
rect 43 137 55 171
rect 89 137 100 171
rect 43 112 100 137
rect 130 112 178 196
rect 208 171 264 196
rect 208 137 219 171
rect 253 137 264 171
rect 208 112 264 137
rect 294 112 342 196
rect 372 171 429 196
rect 372 137 383 171
rect 417 137 429 171
rect 372 112 429 137
<< pdiff >>
rect 27 566 84 574
rect 27 532 39 566
rect 73 532 84 566
rect 27 498 84 532
rect 27 464 39 498
rect 73 464 84 498
rect 27 430 84 464
rect 27 396 39 430
rect 73 396 84 430
rect 27 374 84 396
rect 134 374 176 574
rect 226 562 279 574
rect 226 528 237 562
rect 271 528 279 562
rect 226 494 279 528
rect 226 460 237 494
rect 271 460 279 494
rect 226 420 279 460
rect 226 386 237 420
rect 271 386 279 420
rect 226 374 279 386
<< ndiffc >>
rect 55 137 89 171
rect 219 137 253 171
rect 383 137 417 171
<< pdiffc >>
rect 39 532 73 566
rect 39 464 73 498
rect 39 396 73 430
rect 237 528 271 562
rect 237 460 271 494
rect 237 386 271 420
<< poly >>
rect 84 574 134 600
rect 176 574 226 600
rect 84 302 134 374
rect 176 359 226 374
rect 176 329 372 359
rect 64 286 134 302
rect 64 252 80 286
rect 114 266 134 286
rect 114 252 208 266
rect 64 236 208 252
rect 100 196 130 236
rect 178 196 208 236
rect 264 196 294 329
rect 342 302 372 329
rect 342 286 408 302
rect 342 252 358 286
rect 392 252 408 286
rect 342 236 408 252
rect 342 196 372 236
rect 100 86 130 112
rect 178 86 208 112
rect 264 86 294 112
rect 342 86 372 112
<< polycont >>
rect 80 252 114 286
rect 358 252 392 286
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 23 566 89 649
rect 23 532 39 566
rect 73 532 89 566
rect 23 498 89 532
rect 23 464 39 498
rect 73 464 89 498
rect 23 430 89 464
rect 23 396 39 430
rect 73 396 89 430
rect 203 562 279 578
rect 203 528 237 562
rect 271 528 279 562
rect 203 494 279 528
rect 203 460 237 494
rect 271 460 279 494
rect 203 420 279 460
rect 203 386 237 420
rect 271 386 279 420
rect 25 286 167 356
rect 25 252 80 286
rect 114 252 167 286
rect 25 236 167 252
rect 39 171 105 200
rect 39 137 55 171
rect 89 137 105 171
rect 39 17 105 137
rect 203 171 279 386
rect 313 286 455 578
rect 313 252 358 286
rect 392 252 455 286
rect 313 236 455 252
rect 203 137 219 171
rect 253 137 279 171
rect 203 88 279 137
rect 367 171 433 200
rect 367 137 383 171
rect 417 137 433 171
rect 367 17 433 137
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor2_lp2
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5289350
string GDS_START 5283282
<< end >>
