magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3046 1852
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 1 177 185 203
rect 735 177 1013 203
rect 1563 177 1747 203
rect 1 21 1747 177
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 174 47 204 151
rect 387 47 417 151
rect 503 47 533 151
rect 716 47 746 151
rect 811 47 841 177
rect 907 47 937 177
rect 1002 47 1032 151
rect 1215 47 1245 151
rect 1331 47 1361 151
rect 1544 47 1574 151
rect 1639 47 1669 177
<< scpmoshvt >>
rect 81 297 117 497
rect 186 333 222 497
rect 384 297 420 497
rect 500 297 536 497
rect 698 333 734 497
rect 803 297 839 497
rect 909 297 945 497
rect 1014 333 1050 497
rect 1212 297 1248 497
rect 1328 297 1364 497
rect 1526 333 1562 497
rect 1631 297 1667 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 151 159 177
rect 761 151 811 177
rect 109 47 174 151
rect 204 116 256 151
rect 204 82 214 116
rect 248 82 256 116
rect 204 47 256 82
rect 330 116 387 151
rect 330 82 338 116
rect 372 82 387 116
rect 330 47 387 82
rect 417 116 503 151
rect 417 82 443 116
rect 477 82 503 116
rect 417 47 503 82
rect 533 116 590 151
rect 533 82 548 116
rect 582 82 590 116
rect 533 47 590 82
rect 664 116 716 151
rect 664 82 672 116
rect 706 82 716 116
rect 664 47 716 82
rect 746 47 811 151
rect 841 161 907 177
rect 841 127 857 161
rect 891 127 907 161
rect 841 93 907 127
rect 841 59 857 93
rect 891 59 907 93
rect 841 47 907 59
rect 937 151 987 177
rect 1589 151 1639 177
rect 937 47 1002 151
rect 1032 116 1084 151
rect 1032 82 1042 116
rect 1076 82 1084 116
rect 1032 47 1084 82
rect 1158 116 1215 151
rect 1158 82 1166 116
rect 1200 82 1215 116
rect 1158 47 1215 82
rect 1245 116 1331 151
rect 1245 82 1271 116
rect 1305 82 1331 116
rect 1245 47 1331 82
rect 1361 116 1418 151
rect 1361 82 1376 116
rect 1410 82 1418 116
rect 1361 47 1418 82
rect 1492 116 1544 151
rect 1492 82 1500 116
rect 1534 82 1544 116
rect 1492 47 1544 82
rect 1574 47 1639 151
rect 1669 161 1721 177
rect 1669 127 1679 161
rect 1713 127 1721 161
rect 1669 93 1721 127
rect 1669 59 1679 93
rect 1713 59 1721 93
rect 1669 47 1721 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 333 186 497
rect 222 485 276 497
rect 222 451 234 485
rect 268 451 276 485
rect 222 417 276 451
rect 222 383 234 417
rect 268 383 276 417
rect 222 333 276 383
rect 330 479 384 497
rect 330 445 338 479
rect 372 445 384 479
rect 330 411 384 445
rect 330 377 338 411
rect 372 377 384 411
rect 330 343 384 377
rect 117 297 169 333
rect 330 309 338 343
rect 372 309 384 343
rect 330 297 384 309
rect 420 479 500 497
rect 420 445 443 479
rect 477 445 500 479
rect 420 411 500 445
rect 420 377 443 411
rect 477 377 500 411
rect 420 343 500 377
rect 420 309 443 343
rect 477 309 500 343
rect 420 297 500 309
rect 536 479 590 497
rect 536 445 548 479
rect 582 445 590 479
rect 536 411 590 445
rect 536 377 548 411
rect 582 377 590 411
rect 536 343 590 377
rect 536 309 548 343
rect 582 309 590 343
rect 644 485 698 497
rect 644 451 652 485
rect 686 451 698 485
rect 644 417 698 451
rect 644 383 652 417
rect 686 383 698 417
rect 644 333 698 383
rect 734 333 803 497
rect 536 297 590 309
rect 751 297 803 333
rect 839 485 909 497
rect 839 451 857 485
rect 891 451 909 485
rect 839 417 909 451
rect 839 383 857 417
rect 891 383 909 417
rect 839 349 909 383
rect 839 315 857 349
rect 891 315 909 349
rect 839 297 909 315
rect 945 333 1014 497
rect 1050 485 1104 497
rect 1050 451 1062 485
rect 1096 451 1104 485
rect 1050 417 1104 451
rect 1050 383 1062 417
rect 1096 383 1104 417
rect 1050 333 1104 383
rect 1158 479 1212 497
rect 1158 445 1166 479
rect 1200 445 1212 479
rect 1158 411 1212 445
rect 1158 377 1166 411
rect 1200 377 1212 411
rect 1158 343 1212 377
rect 945 297 997 333
rect 1158 309 1166 343
rect 1200 309 1212 343
rect 1158 297 1212 309
rect 1248 479 1328 497
rect 1248 445 1271 479
rect 1305 445 1328 479
rect 1248 411 1328 445
rect 1248 377 1271 411
rect 1305 377 1328 411
rect 1248 343 1328 377
rect 1248 309 1271 343
rect 1305 309 1328 343
rect 1248 297 1328 309
rect 1364 479 1418 497
rect 1364 445 1376 479
rect 1410 445 1418 479
rect 1364 411 1418 445
rect 1364 377 1376 411
rect 1410 377 1418 411
rect 1364 343 1418 377
rect 1364 309 1376 343
rect 1410 309 1418 343
rect 1472 485 1526 497
rect 1472 451 1480 485
rect 1514 451 1526 485
rect 1472 417 1526 451
rect 1472 383 1480 417
rect 1514 383 1526 417
rect 1472 333 1526 383
rect 1562 333 1631 497
rect 1364 297 1418 309
rect 1579 297 1631 333
rect 1667 485 1721 497
rect 1667 451 1679 485
rect 1713 451 1721 485
rect 1667 417 1721 451
rect 1667 383 1679 417
rect 1713 383 1721 417
rect 1667 349 1721 383
rect 1667 315 1679 349
rect 1713 315 1721 349
rect 1667 297 1721 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 214 82 248 116
rect 338 82 372 116
rect 443 82 477 116
rect 548 82 582 116
rect 672 82 706 116
rect 857 127 891 161
rect 857 59 891 93
rect 1042 82 1076 116
rect 1166 82 1200 116
rect 1271 82 1305 116
rect 1376 82 1410 116
rect 1500 82 1534 116
rect 1679 127 1713 161
rect 1679 59 1713 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 234 451 268 485
rect 234 383 268 417
rect 338 445 372 479
rect 338 377 372 411
rect 338 309 372 343
rect 443 445 477 479
rect 443 377 477 411
rect 443 309 477 343
rect 548 445 582 479
rect 548 377 582 411
rect 548 309 582 343
rect 652 451 686 485
rect 652 383 686 417
rect 857 451 891 485
rect 857 383 891 417
rect 857 315 891 349
rect 1062 451 1096 485
rect 1062 383 1096 417
rect 1166 445 1200 479
rect 1166 377 1200 411
rect 1166 309 1200 343
rect 1271 445 1305 479
rect 1271 377 1305 411
rect 1271 309 1305 343
rect 1376 445 1410 479
rect 1376 377 1410 411
rect 1376 309 1410 343
rect 1480 451 1514 485
rect 1480 383 1514 417
rect 1679 451 1713 485
rect 1679 383 1713 417
rect 1679 315 1713 349
<< poly >>
rect 81 497 117 523
rect 186 497 222 524
rect 384 497 420 523
rect 500 497 536 523
rect 698 497 734 524
rect 803 497 839 523
rect 909 497 945 523
rect 1014 497 1050 524
rect 1212 497 1248 523
rect 1328 497 1364 523
rect 1526 497 1562 524
rect 1631 497 1667 523
rect 81 282 117 297
rect 186 295 222 333
rect 184 285 298 295
rect 79 265 119 282
rect 184 265 248 285
rect 73 249 127 265
rect 73 215 83 249
rect 117 215 127 249
rect 232 251 248 265
rect 282 251 298 285
rect 384 282 420 297
rect 500 282 536 297
rect 698 295 734 333
rect 622 285 736 295
rect 232 241 298 251
rect 382 239 422 282
rect 73 199 127 215
rect 368 223 422 239
rect 79 177 109 199
rect 368 196 378 223
rect 174 189 378 196
rect 412 189 422 223
rect 174 173 422 189
rect 498 239 538 282
rect 622 251 638 285
rect 672 265 736 285
rect 803 282 839 297
rect 909 282 945 297
rect 1014 295 1050 333
rect 1012 285 1126 295
rect 801 265 841 282
rect 907 265 947 282
rect 1012 265 1076 285
rect 672 251 688 265
rect 622 241 688 251
rect 793 249 847 265
rect 498 223 552 239
rect 498 189 508 223
rect 542 196 552 223
rect 793 215 803 249
rect 837 215 847 249
rect 793 199 847 215
rect 901 249 955 265
rect 901 215 911 249
rect 945 215 955 249
rect 1060 251 1076 265
rect 1110 251 1126 285
rect 1212 282 1248 297
rect 1328 282 1364 297
rect 1526 295 1562 333
rect 1450 285 1564 295
rect 1060 241 1126 251
rect 1210 239 1250 282
rect 901 199 955 215
rect 1196 223 1250 239
rect 542 189 746 196
rect 498 173 746 189
rect 811 177 841 199
rect 907 177 937 199
rect 1196 196 1206 223
rect 1002 189 1206 196
rect 1240 189 1250 223
rect 174 166 417 173
rect 174 151 204 166
rect 387 151 417 166
rect 503 166 746 173
rect 503 151 533 166
rect 716 151 746 166
rect 1002 173 1250 189
rect 1326 239 1366 282
rect 1450 251 1466 285
rect 1500 265 1564 285
rect 1631 282 1667 297
rect 1629 265 1669 282
rect 1500 251 1516 265
rect 1450 241 1516 251
rect 1621 249 1675 265
rect 1326 223 1380 239
rect 1326 189 1336 223
rect 1370 196 1380 223
rect 1621 215 1631 249
rect 1665 215 1675 249
rect 1621 199 1675 215
rect 1370 189 1574 196
rect 1326 173 1574 189
rect 1639 177 1669 199
rect 1002 166 1245 173
rect 1002 151 1032 166
rect 1215 151 1245 166
rect 1331 166 1574 173
rect 1331 151 1361 166
rect 1544 151 1574 166
rect 79 21 109 47
rect 174 21 204 47
rect 387 21 417 47
rect 503 21 533 47
rect 716 21 746 47
rect 811 21 841 47
rect 907 21 937 47
rect 1002 21 1032 47
rect 1215 21 1245 47
rect 1331 21 1361 47
rect 1544 21 1574 47
rect 1639 21 1669 47
<< polycont >>
rect 83 215 117 249
rect 248 251 282 285
rect 378 189 412 223
rect 638 251 672 285
rect 508 189 542 223
rect 803 215 837 249
rect 911 215 945 249
rect 1076 251 1110 285
rect 1206 189 1240 223
rect 1466 251 1500 285
rect 1336 189 1370 223
rect 1631 215 1665 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 19 485 85 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 218 485 284 493
rect 218 451 234 485
rect 268 451 284 485
rect 218 417 284 451
rect 218 397 234 417
rect 19 349 85 383
rect 19 315 35 349
rect 69 315 85 349
rect 19 299 85 315
rect 180 391 234 397
rect 180 357 213 391
rect 268 383 284 417
rect 247 361 284 383
rect 322 479 388 493
rect 322 445 338 479
rect 372 445 388 479
rect 322 411 388 445
rect 322 377 338 411
rect 372 377 388 411
rect 247 357 259 361
rect 180 351 259 357
rect 67 249 146 265
rect 67 215 83 249
rect 117 215 146 249
rect 67 211 146 215
rect 26 161 78 177
rect 26 127 35 161
rect 69 127 78 161
rect 26 93 78 127
rect 26 59 35 93
rect 69 59 78 93
rect 112 125 146 211
rect 180 201 214 351
rect 322 343 388 377
rect 322 327 338 343
rect 292 309 338 327
rect 372 309 388 343
rect 292 301 388 309
rect 248 293 388 301
rect 433 479 493 527
rect 433 445 443 479
rect 477 445 493 479
rect 433 411 493 445
rect 433 377 443 411
rect 477 377 493 411
rect 433 343 493 377
rect 433 309 443 343
rect 477 309 493 343
rect 433 293 493 309
rect 532 479 598 493
rect 532 445 548 479
rect 582 445 598 479
rect 532 411 598 445
rect 532 377 548 411
rect 582 377 598 411
rect 532 343 598 377
rect 636 485 702 493
rect 636 451 652 485
rect 686 451 702 485
rect 636 417 702 451
rect 636 383 652 417
rect 686 397 702 417
rect 835 485 913 527
rect 835 451 857 485
rect 891 451 913 485
rect 835 417 913 451
rect 686 391 740 397
rect 636 361 673 383
rect 661 357 673 361
rect 707 357 740 391
rect 661 351 740 357
rect 532 309 548 343
rect 582 327 598 343
rect 582 309 628 327
rect 532 301 628 309
rect 532 293 672 301
rect 248 285 326 293
rect 282 251 326 285
rect 594 285 672 293
rect 248 235 326 251
rect 180 167 258 201
rect 112 79 167 125
rect 209 116 258 167
rect 292 151 326 235
rect 361 223 431 259
rect 361 189 378 223
rect 412 189 431 223
rect 489 223 559 259
rect 489 189 508 223
rect 542 189 559 223
rect 594 251 638 285
rect 594 235 672 251
rect 594 151 628 235
rect 706 201 740 351
rect 835 383 857 417
rect 891 383 913 417
rect 1046 485 1112 493
rect 1046 451 1062 485
rect 1096 451 1112 485
rect 1046 417 1112 451
rect 1046 397 1062 417
rect 835 349 913 383
rect 835 315 857 349
rect 891 315 913 349
rect 835 299 913 315
rect 1008 391 1062 397
rect 1008 357 1041 391
rect 1096 383 1112 417
rect 1075 361 1112 383
rect 1150 479 1216 493
rect 1150 445 1166 479
rect 1200 445 1216 479
rect 1150 411 1216 445
rect 1150 377 1166 411
rect 1200 377 1216 411
rect 1075 357 1087 361
rect 1008 351 1087 357
rect 292 117 380 151
rect 209 82 214 116
rect 248 82 258 116
rect 209 66 258 82
rect 330 116 380 117
rect 330 82 338 116
rect 372 82 380 116
rect 330 66 380 82
rect 427 116 493 132
rect 427 82 443 116
rect 477 82 493 116
rect 26 17 78 59
rect 427 17 493 82
rect 540 117 628 151
rect 662 167 740 201
rect 774 249 853 265
rect 774 215 803 249
rect 837 215 853 249
rect 774 211 853 215
rect 895 249 974 265
rect 895 215 911 249
rect 945 215 974 249
rect 895 211 974 215
rect 540 116 590 117
rect 540 82 548 116
rect 582 82 590 116
rect 540 66 590 82
rect 662 116 711 167
rect 774 125 808 211
rect 662 82 672 116
rect 706 82 711 116
rect 662 66 711 82
rect 753 79 808 125
rect 842 161 906 177
rect 842 127 857 161
rect 891 127 906 161
rect 842 93 906 127
rect 842 59 857 93
rect 891 59 906 93
rect 940 125 974 211
rect 1008 201 1042 351
rect 1150 343 1216 377
rect 1150 327 1166 343
rect 1120 309 1166 327
rect 1200 309 1216 343
rect 1120 301 1216 309
rect 1076 293 1216 301
rect 1255 479 1315 527
rect 1255 445 1271 479
rect 1305 445 1315 479
rect 1255 411 1315 445
rect 1255 377 1271 411
rect 1305 377 1315 411
rect 1255 343 1315 377
rect 1255 309 1271 343
rect 1305 309 1315 343
rect 1255 293 1315 309
rect 1360 479 1426 493
rect 1360 445 1376 479
rect 1410 445 1426 479
rect 1360 411 1426 445
rect 1360 377 1376 411
rect 1410 377 1426 411
rect 1360 343 1426 377
rect 1464 485 1530 493
rect 1464 451 1480 485
rect 1514 451 1530 485
rect 1464 417 1530 451
rect 1464 383 1480 417
rect 1514 397 1530 417
rect 1663 485 1729 527
rect 1663 451 1679 485
rect 1713 451 1729 485
rect 1663 417 1729 451
rect 1514 391 1568 397
rect 1464 361 1501 383
rect 1489 357 1501 361
rect 1535 357 1568 391
rect 1489 351 1568 357
rect 1360 309 1376 343
rect 1410 327 1426 343
rect 1410 309 1456 327
rect 1360 301 1456 309
rect 1360 293 1500 301
rect 1076 285 1154 293
rect 1110 251 1154 285
rect 1422 285 1500 293
rect 1076 235 1154 251
rect 1008 167 1086 201
rect 940 79 995 125
rect 1037 116 1086 167
rect 1120 151 1154 235
rect 1189 223 1259 259
rect 1189 189 1206 223
rect 1240 189 1259 223
rect 1317 223 1387 259
rect 1317 189 1336 223
rect 1370 189 1387 223
rect 1422 251 1466 285
rect 1422 235 1500 251
rect 1422 151 1456 235
rect 1534 201 1568 351
rect 1663 383 1679 417
rect 1713 383 1729 417
rect 1663 349 1729 383
rect 1663 315 1679 349
rect 1713 315 1729 349
rect 1663 299 1729 315
rect 1120 117 1208 151
rect 1037 82 1042 116
rect 1076 82 1086 116
rect 1037 66 1086 82
rect 1158 116 1208 117
rect 1158 82 1166 116
rect 1200 82 1208 116
rect 1158 66 1208 82
rect 1255 116 1321 132
rect 1255 82 1271 116
rect 1305 82 1321 116
rect 842 17 906 59
rect 1255 17 1321 82
rect 1368 117 1456 151
rect 1490 167 1568 201
rect 1602 249 1681 265
rect 1602 215 1631 249
rect 1665 215 1681 249
rect 1602 211 1681 215
rect 1368 116 1418 117
rect 1368 82 1376 116
rect 1410 82 1418 116
rect 1368 66 1418 82
rect 1490 116 1539 167
rect 1602 125 1636 211
rect 1490 82 1500 116
rect 1534 82 1539 116
rect 1490 66 1539 82
rect 1581 79 1636 125
rect 1670 161 1722 177
rect 1670 127 1679 161
rect 1713 127 1722 161
rect 1670 93 1722 127
rect 1670 59 1679 93
rect 1713 59 1722 93
rect 1670 17 1722 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 213 383 234 391
rect 234 383 247 391
rect 213 357 247 383
rect 673 383 686 391
rect 686 383 707 391
rect 673 357 707 383
rect 1041 383 1062 391
rect 1062 383 1075 391
rect 1041 357 1075 383
rect 1501 383 1514 391
rect 1514 383 1535 391
rect 1501 357 1535 383
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 201 391 259 397
rect 201 357 213 391
rect 247 388 259 391
rect 661 391 719 397
rect 661 388 673 391
rect 247 360 673 388
rect 247 357 259 360
rect 201 351 259 357
rect 661 357 673 360
rect 707 388 719 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 707 360 1041 388
rect 707 357 719 360
rect 661 351 719 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1489 391 1547 397
rect 1489 388 1501 391
rect 1075 360 1501 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1489 357 1501 360
rect 1535 357 1547 391
rect 1489 351 1547 357
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 S[0]
port 8 nsew signal input
flabel locali s 121 85 155 119 0 FreeSans 200 0 0 0 D[0]
port 4 nsew signal input
flabel locali s 765 85 799 119 0 FreeSans 200 180 0 0 D[1]
port 3 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 200 180 0 0 S[1]
port 7 nsew signal input
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 S[2]
port 6 nsew signal input
flabel locali s 949 85 983 119 0 FreeSans 200 0 0 0 D[2]
port 2 nsew signal input
flabel locali s 1593 85 1627 119 0 FreeSans 200 180 0 0 D[3]
port 1 nsew signal input
flabel locali s 1317 221 1351 255 0 FreeSans 200 180 0 0 S[3]
port 5 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 11 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 10 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 9 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 12 nsew power bidirectional
flabel metal1 s 213 357 247 391 0 FreeSans 200 0 0 0 Z
port 13 nsew signal output
rlabel comment s 0 0 0 0 4 muxb4to1_1
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1748 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 3051428
string GDS_START 3032294
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
