magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4562 1975
<< nwell >>
rect -38 331 3302 704
<< pwell >>
rect 1268 223 2153 235
rect 735 176 2153 223
rect 735 167 2406 176
rect 2839 167 3263 184
rect 735 157 3263 167
rect 25 49 3263 157
rect 0 0 3264 49
<< scnmos >>
rect 108 47 138 131
rect 186 47 216 131
rect 332 47 362 131
rect 410 47 440 131
rect 496 47 526 131
rect 574 47 604 131
rect 818 113 848 197
rect 890 113 920 197
rect 976 113 1006 197
rect 1048 113 1078 197
rect 1249 83 1279 167
rect 1351 125 1381 209
rect 1423 125 1453 209
rect 1699 125 1729 209
rect 1777 125 1807 209
rect 1885 125 1915 209
rect 1993 125 2023 209
rect 2142 66 2172 150
rect 2220 66 2250 150
rect 2293 66 2323 150
rect 2494 57 2524 141
rect 2566 57 2596 141
rect 2652 57 2682 141
rect 2724 57 2754 141
rect 2921 74 2951 158
rect 2993 74 3023 158
rect 3079 74 3109 158
rect 3151 74 3181 158
<< scpmoshvt >>
rect 84 409 134 609
rect 302 409 352 609
rect 408 409 458 609
rect 506 409 556 609
rect 612 409 662 609
rect 831 409 881 609
rect 937 409 987 609
rect 1151 419 1201 619
rect 1323 419 1373 619
rect 1429 419 1479 619
rect 1609 419 1659 619
rect 1715 419 1765 619
rect 1871 419 1921 619
rect 1969 419 2019 619
rect 2143 419 2193 619
rect 2257 419 2307 619
rect 2397 419 2447 619
rect 2614 400 2664 600
rect 2754 400 2804 600
rect 2972 374 3022 574
rect 3078 374 3128 574
<< ndiff >>
rect 761 179 818 197
rect 761 145 773 179
rect 807 145 818 179
rect 51 111 108 131
rect 51 77 63 111
rect 97 77 108 111
rect 51 47 108 77
rect 138 47 186 131
rect 216 106 332 131
rect 216 72 227 106
rect 261 72 332 106
rect 216 47 332 72
rect 362 47 410 131
rect 440 106 496 131
rect 440 72 451 106
rect 485 72 496 106
rect 440 47 496 72
rect 526 47 574 131
rect 604 96 661 131
rect 761 113 818 145
rect 848 113 890 197
rect 920 163 976 197
rect 920 129 931 163
rect 965 129 976 163
rect 920 113 976 129
rect 1006 113 1048 197
rect 1078 179 1135 197
rect 1078 145 1089 179
rect 1123 145 1135 179
rect 1294 184 1351 209
rect 1294 167 1306 184
rect 1078 113 1135 145
rect 1192 142 1249 167
rect 604 62 615 96
rect 649 62 661 96
rect 1192 108 1204 142
rect 1238 108 1249 142
rect 1192 83 1249 108
rect 1279 150 1306 167
rect 1340 150 1351 184
rect 1279 125 1351 150
rect 1381 125 1423 209
rect 1453 125 1525 209
rect 1642 180 1699 209
rect 1642 146 1654 180
rect 1688 146 1699 180
rect 1642 125 1699 146
rect 1729 125 1777 209
rect 1807 179 1885 209
rect 1807 145 1826 179
rect 1860 145 1885 179
rect 1807 125 1885 145
rect 1915 125 1993 209
rect 2023 197 2127 209
rect 2023 163 2081 197
rect 2115 163 2127 197
rect 2023 150 2127 163
rect 2023 125 2142 150
rect 1279 83 1329 125
rect 1468 123 1525 125
rect 1468 89 1479 123
rect 1513 89 1525 123
rect 2069 112 2142 125
rect 604 47 661 62
rect 1468 77 1525 89
rect 2069 78 2081 112
rect 2115 78 2142 112
rect 2069 66 2142 78
rect 2172 66 2220 150
rect 2250 66 2293 150
rect 2323 125 2380 150
rect 2323 91 2334 125
rect 2368 91 2380 125
rect 2323 66 2380 91
rect 2437 116 2494 141
rect 2437 82 2449 116
rect 2483 82 2494 116
rect 2437 57 2494 82
rect 2524 57 2566 141
rect 2596 116 2652 141
rect 2596 82 2607 116
rect 2641 82 2652 116
rect 2596 57 2652 82
rect 2682 57 2724 141
rect 2754 116 2811 141
rect 2754 82 2765 116
rect 2799 82 2811 116
rect 2754 57 2811 82
rect 2865 133 2921 158
rect 2865 99 2876 133
rect 2910 99 2921 133
rect 2865 74 2921 99
rect 2951 74 2993 158
rect 3023 133 3079 158
rect 3023 99 3034 133
rect 3068 99 3079 133
rect 3023 74 3079 99
rect 3109 74 3151 158
rect 3181 133 3237 158
rect 3181 99 3192 133
rect 3226 99 3237 133
rect 3181 74 3237 99
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 191 609
rect 134 563 145 597
rect 179 563 191 597
rect 134 526 191 563
rect 134 492 145 526
rect 179 492 191 526
rect 134 455 191 492
rect 134 421 145 455
rect 179 421 191 455
rect 134 409 191 421
rect 245 597 302 609
rect 245 563 257 597
rect 291 563 302 597
rect 245 526 302 563
rect 245 492 257 526
rect 291 492 302 526
rect 245 455 302 492
rect 245 421 257 455
rect 291 421 302 455
rect 245 409 302 421
rect 352 527 408 609
rect 352 493 363 527
rect 397 493 408 527
rect 352 455 408 493
rect 352 421 363 455
rect 397 421 408 455
rect 352 409 408 421
rect 458 409 506 609
rect 556 590 612 609
rect 556 556 567 590
rect 601 556 612 590
rect 556 409 612 556
rect 662 597 719 609
rect 662 563 673 597
rect 707 563 719 597
rect 662 514 719 563
rect 662 480 673 514
rect 707 480 719 514
rect 662 409 719 480
rect 774 597 831 609
rect 774 563 786 597
rect 820 563 831 597
rect 774 526 831 563
rect 774 492 786 526
rect 820 492 831 526
rect 774 455 831 492
rect 774 421 786 455
rect 820 421 831 455
rect 774 409 831 421
rect 881 597 937 609
rect 881 563 892 597
rect 926 563 937 597
rect 881 512 937 563
rect 881 478 892 512
rect 926 478 937 512
rect 881 409 937 478
rect 987 597 1042 609
rect 987 563 998 597
rect 1032 563 1042 597
rect 987 512 1042 563
rect 987 478 998 512
rect 1032 478 1042 512
rect 987 409 1042 478
rect 1096 496 1151 619
rect 1096 462 1106 496
rect 1140 462 1151 496
rect 1096 419 1151 462
rect 1201 496 1323 619
rect 1201 462 1278 496
rect 1312 462 1323 496
rect 1201 419 1323 462
rect 1373 419 1429 619
rect 1479 607 1609 619
rect 1479 573 1564 607
rect 1598 573 1609 607
rect 1479 419 1609 573
rect 1659 467 1715 619
rect 1659 433 1670 467
rect 1704 433 1715 467
rect 1659 419 1715 433
rect 1765 607 1871 619
rect 1765 573 1776 607
rect 1810 573 1871 607
rect 1765 419 1871 573
rect 1921 419 1969 619
rect 2019 597 2143 619
rect 2019 563 2057 597
rect 2091 563 2143 597
rect 2019 465 2143 563
rect 2019 431 2057 465
rect 2091 431 2143 465
rect 2019 419 2143 431
rect 2193 419 2257 619
rect 2307 611 2397 619
rect 2307 577 2318 611
rect 2352 577 2397 611
rect 2307 543 2397 577
rect 2307 509 2318 543
rect 2352 509 2397 543
rect 2307 419 2397 509
rect 2447 597 2504 619
rect 2447 563 2458 597
rect 2492 563 2504 597
rect 2447 465 2504 563
rect 2447 431 2458 465
rect 2492 431 2504 465
rect 2447 419 2504 431
rect 2558 527 2614 600
rect 2558 493 2569 527
rect 2603 493 2614 527
rect 2558 454 2614 493
rect 2558 420 2569 454
rect 2603 420 2614 454
rect 2558 400 2614 420
rect 2664 588 2754 600
rect 2664 554 2709 588
rect 2743 554 2754 588
rect 2664 517 2754 554
rect 2664 483 2709 517
rect 2743 483 2754 517
rect 2664 446 2754 483
rect 2664 412 2709 446
rect 2743 412 2754 446
rect 2664 400 2754 412
rect 2804 588 2861 600
rect 2804 554 2815 588
rect 2849 554 2861 588
rect 2804 517 2861 554
rect 2804 483 2815 517
rect 2849 483 2861 517
rect 2804 446 2861 483
rect 2804 412 2815 446
rect 2849 412 2861 446
rect 2804 400 2861 412
rect 2915 562 2972 574
rect 2915 528 2927 562
rect 2961 528 2972 562
rect 2915 491 2972 528
rect 2915 457 2927 491
rect 2961 457 2972 491
rect 2915 420 2972 457
rect 2915 386 2927 420
rect 2961 386 2972 420
rect 2915 374 2972 386
rect 3022 562 3078 574
rect 3022 528 3033 562
rect 3067 528 3078 562
rect 3022 491 3078 528
rect 3022 457 3033 491
rect 3067 457 3078 491
rect 3022 420 3078 457
rect 3022 386 3033 420
rect 3067 386 3078 420
rect 3022 374 3078 386
rect 3128 562 3185 574
rect 3128 528 3139 562
rect 3173 528 3185 562
rect 3128 491 3185 528
rect 3128 457 3139 491
rect 3173 457 3185 491
rect 3128 420 3185 457
rect 3128 386 3139 420
rect 3173 386 3185 420
rect 3128 374 3185 386
<< ndiffc >>
rect 773 145 807 179
rect 63 77 97 111
rect 227 72 261 106
rect 451 72 485 106
rect 931 129 965 163
rect 1089 145 1123 179
rect 615 62 649 96
rect 1204 108 1238 142
rect 1306 150 1340 184
rect 1654 146 1688 180
rect 1826 145 1860 179
rect 2081 163 2115 197
rect 1479 89 1513 123
rect 2081 78 2115 112
rect 2334 91 2368 125
rect 2449 82 2483 116
rect 2607 82 2641 116
rect 2765 82 2799 116
rect 2876 99 2910 133
rect 3034 99 3068 133
rect 3192 99 3226 133
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 492 179 526
rect 145 421 179 455
rect 257 563 291 597
rect 257 492 291 526
rect 257 421 291 455
rect 363 493 397 527
rect 363 421 397 455
rect 567 556 601 590
rect 673 563 707 597
rect 673 480 707 514
rect 786 563 820 597
rect 786 492 820 526
rect 786 421 820 455
rect 892 563 926 597
rect 892 478 926 512
rect 998 563 1032 597
rect 998 478 1032 512
rect 1106 462 1140 496
rect 1278 462 1312 496
rect 1564 573 1598 607
rect 1670 433 1704 467
rect 1776 573 1810 607
rect 2057 563 2091 597
rect 2057 431 2091 465
rect 2318 577 2352 611
rect 2318 509 2352 543
rect 2458 563 2492 597
rect 2458 431 2492 465
rect 2569 493 2603 527
rect 2569 420 2603 454
rect 2709 554 2743 588
rect 2709 483 2743 517
rect 2709 412 2743 446
rect 2815 554 2849 588
rect 2815 483 2849 517
rect 2815 412 2849 446
rect 2927 528 2961 562
rect 2927 457 2961 491
rect 2927 386 2961 420
rect 3033 528 3067 562
rect 3033 457 3067 491
rect 3033 386 3067 420
rect 3139 528 3173 562
rect 3139 457 3173 491
rect 3139 386 3173 420
<< poly >>
rect 84 609 134 635
rect 302 609 352 635
rect 408 609 458 635
rect 506 609 556 635
rect 612 609 662 635
rect 831 609 881 635
rect 937 609 987 635
rect 1151 619 1201 645
rect 1323 619 1373 645
rect 1429 619 1479 645
rect 1609 619 1659 645
rect 1715 619 1765 645
rect 1871 619 1921 645
rect 1969 619 2019 645
rect 2143 619 2193 645
rect 2257 619 2307 645
rect 2397 619 2447 645
rect 2614 600 2664 626
rect 2754 600 2804 626
rect 84 237 134 409
rect 302 351 352 409
rect 408 358 458 409
rect 506 358 556 409
rect 211 335 352 351
rect 211 301 227 335
rect 261 301 352 335
rect 211 285 352 301
rect 394 342 460 358
rect 394 308 410 342
rect 444 308 460 342
rect 394 292 460 308
rect 502 342 568 358
rect 502 308 518 342
rect 552 308 568 342
rect 84 221 252 237
rect 84 207 202 221
rect 108 131 138 207
rect 186 187 202 207
rect 236 187 252 221
rect 186 171 252 187
rect 316 176 346 285
rect 186 131 216 171
rect 316 146 362 176
rect 332 131 362 146
rect 410 131 440 292
rect 502 274 568 308
rect 502 240 518 274
rect 552 240 568 274
rect 502 224 568 240
rect 612 356 662 409
rect 831 356 881 409
rect 937 377 987 409
rect 937 361 1029 377
rect 612 340 738 356
rect 612 306 688 340
rect 722 306 738 340
rect 612 272 738 306
rect 612 238 688 272
rect 722 238 738 272
rect 502 176 532 224
rect 612 222 738 238
rect 818 340 895 356
rect 818 306 845 340
rect 879 306 895 340
rect 937 327 979 361
rect 1013 327 1029 361
rect 1151 356 1201 419
rect 1323 404 1373 419
rect 937 311 1029 327
rect 1135 340 1201 356
rect 818 263 895 306
rect 818 233 920 263
rect 616 176 646 222
rect 818 197 848 233
rect 890 197 920 233
rect 976 242 1006 311
rect 1135 306 1151 340
rect 1185 306 1201 340
rect 1135 290 1201 306
rect 1243 374 1373 404
rect 1243 242 1273 374
rect 1429 368 1479 419
rect 1609 381 1659 419
rect 1423 352 1553 368
rect 1315 310 1381 326
rect 1315 276 1331 310
rect 1365 276 1381 310
rect 1315 260 1381 276
rect 976 212 1273 242
rect 976 197 1006 212
rect 1048 197 1078 212
rect 496 146 532 176
rect 574 146 646 176
rect 496 131 526 146
rect 574 131 604 146
rect 1243 182 1279 212
rect 1351 209 1381 260
rect 1423 318 1503 352
rect 1537 318 1553 352
rect 1423 302 1553 318
rect 1601 365 1667 381
rect 1601 331 1617 365
rect 1651 331 1667 365
rect 1601 315 1667 331
rect 1423 209 1453 302
rect 1637 262 1667 315
rect 1715 376 1765 419
rect 1715 360 1813 376
rect 1871 374 1921 419
rect 1715 326 1763 360
rect 1797 326 1813 360
rect 1715 310 1813 326
rect 1855 358 1921 374
rect 1855 324 1871 358
rect 1905 324 1921 358
rect 1969 375 2019 419
rect 2143 387 2193 419
rect 1969 345 2101 375
rect 1637 232 1729 262
rect 1699 209 1729 232
rect 1777 209 1807 310
rect 1855 290 1921 324
rect 1855 256 1871 290
rect 1905 256 1921 290
rect 1855 240 1921 256
rect 1963 281 2029 297
rect 1963 247 1979 281
rect 2013 247 2029 281
rect 1885 209 1915 240
rect 1963 231 2029 247
rect 2071 273 2101 345
rect 2143 371 2209 387
rect 2257 377 2307 419
rect 2397 378 2447 419
rect 2972 574 3022 600
rect 3078 574 3128 600
rect 2143 337 2159 371
rect 2193 337 2209 371
rect 2143 321 2209 337
rect 2251 361 2355 377
rect 2251 327 2305 361
rect 2339 327 2355 361
rect 2251 293 2355 327
rect 2251 273 2305 293
rect 2071 243 2172 273
rect 1993 209 2023 231
rect 1249 167 1279 182
rect 818 87 848 113
rect 890 87 920 113
rect 976 87 1006 113
rect 1048 87 1078 113
rect 2142 150 2172 243
rect 2220 259 2305 273
rect 2339 259 2355 293
rect 2220 243 2355 259
rect 2397 362 2463 378
rect 2614 368 2664 400
rect 2397 328 2413 362
rect 2447 328 2463 362
rect 2397 312 2463 328
rect 2566 352 2664 368
rect 2566 318 2614 352
rect 2648 318 2664 352
rect 2220 150 2250 243
rect 2397 195 2427 312
rect 2566 284 2664 318
rect 2566 264 2614 284
rect 2293 165 2427 195
rect 2494 250 2614 264
rect 2648 264 2664 284
rect 2754 264 2804 400
rect 2648 250 2804 264
rect 2494 234 2804 250
rect 2293 150 2323 165
rect 1351 99 1381 125
rect 1423 99 1453 125
rect 1699 99 1729 125
rect 1777 99 1807 125
rect 1885 99 1915 125
rect 1993 99 2023 125
rect 1249 51 1279 83
rect 2494 141 2524 234
rect 2566 141 2596 234
rect 2724 203 2804 234
rect 2972 203 3022 374
rect 3078 332 3128 374
rect 3079 316 3145 332
rect 3079 282 3095 316
rect 3129 282 3145 316
rect 3079 248 3145 282
rect 3079 214 3095 248
rect 3129 228 3145 248
rect 3129 214 3181 228
rect 2724 186 3023 203
rect 2652 173 3023 186
rect 2652 156 2754 173
rect 2921 158 2951 173
rect 2993 158 3023 173
rect 3079 198 3181 214
rect 3079 158 3109 198
rect 3151 158 3181 198
rect 2652 141 2682 156
rect 2724 141 2754 156
rect 2142 51 2172 66
rect 108 21 138 47
rect 186 21 216 47
rect 332 21 362 47
rect 410 21 440 47
rect 496 21 526 47
rect 574 21 604 47
rect 1249 21 2172 51
rect 2220 40 2250 66
rect 2293 40 2323 66
rect 2494 31 2524 57
rect 2566 31 2596 57
rect 2652 31 2682 57
rect 2724 31 2754 57
rect 2921 48 2951 74
rect 2993 48 3023 74
rect 3079 48 3109 74
rect 3151 48 3181 74
<< polycont >>
rect 227 301 261 335
rect 410 308 444 342
rect 518 308 552 342
rect 202 187 236 221
rect 518 240 552 274
rect 688 306 722 340
rect 688 238 722 272
rect 845 306 879 340
rect 979 327 1013 361
rect 1151 306 1185 340
rect 1331 276 1365 310
rect 1503 318 1537 352
rect 1617 331 1651 365
rect 1763 326 1797 360
rect 1871 324 1905 358
rect 1871 256 1905 290
rect 1979 247 2013 281
rect 2159 337 2193 371
rect 2305 327 2339 361
rect 2305 259 2339 293
rect 2413 328 2447 362
rect 2614 318 2648 352
rect 2614 250 2648 284
rect 3095 282 3129 316
rect 3095 214 3129 248
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 526 89 563
rect 23 492 39 526
rect 73 492 89 526
rect 23 455 89 492
rect 23 421 39 455
rect 73 421 89 455
rect 23 351 89 421
rect 129 597 195 649
rect 129 563 145 597
rect 179 563 195 597
rect 129 526 195 563
rect 129 492 145 526
rect 179 492 195 526
rect 129 455 195 492
rect 129 421 145 455
rect 179 421 195 455
rect 129 405 195 421
rect 241 597 515 613
rect 241 563 257 597
rect 291 579 515 597
rect 291 563 307 579
rect 241 526 307 563
rect 241 492 257 526
rect 291 492 307 526
rect 241 455 307 492
rect 241 421 257 455
rect 291 421 307 455
rect 241 405 307 421
rect 347 527 413 543
rect 347 493 363 527
rect 397 493 413 527
rect 347 455 413 493
rect 481 498 515 579
rect 551 590 617 649
rect 551 556 567 590
rect 601 556 617 590
rect 551 534 617 556
rect 657 597 723 613
rect 657 563 673 597
rect 707 563 723 597
rect 657 514 723 563
rect 657 498 673 514
rect 481 480 673 498
rect 707 480 723 514
rect 481 464 723 480
rect 770 597 836 613
rect 770 563 786 597
rect 820 563 836 597
rect 770 526 836 563
rect 770 492 786 526
rect 820 492 836 526
rect 347 421 363 455
rect 397 428 413 455
rect 770 455 836 492
rect 876 597 942 649
rect 876 563 892 597
rect 926 563 942 597
rect 876 512 942 563
rect 876 478 892 512
rect 926 478 942 512
rect 876 462 942 478
rect 982 597 1512 613
rect 982 563 998 597
rect 1032 579 1512 597
rect 1032 563 1048 579
rect 982 512 1048 563
rect 982 478 998 512
rect 1032 478 1048 512
rect 982 462 1048 478
rect 1090 496 1156 543
rect 1090 462 1106 496
rect 1140 462 1156 496
rect 397 421 637 428
rect 347 394 637 421
rect 23 335 277 351
rect 23 301 227 335
rect 261 301 277 335
rect 23 285 277 301
rect 313 342 460 358
rect 313 308 410 342
rect 444 308 460 342
rect 313 292 460 308
rect 502 342 567 358
rect 502 308 518 342
rect 552 308 567 342
rect 23 111 113 285
rect 502 274 567 308
rect 502 256 518 274
rect 313 240 518 256
rect 552 240 567 274
rect 313 237 567 240
rect 186 222 567 237
rect 186 221 455 222
rect 186 187 202 221
rect 236 187 455 221
rect 186 171 455 187
rect 603 186 637 394
rect 770 421 786 455
rect 820 426 836 455
rect 1090 426 1156 462
rect 820 421 1028 426
rect 770 392 1028 421
rect 673 340 737 356
rect 673 306 688 340
rect 722 306 737 340
rect 673 272 737 306
rect 673 238 688 272
rect 722 238 737 272
rect 673 222 737 238
rect 773 201 807 392
rect 965 361 1028 392
rect 843 340 929 356
rect 843 306 845 340
rect 879 306 929 340
rect 965 327 979 361
rect 1013 327 1028 361
rect 965 311 1028 327
rect 1064 392 1156 426
rect 843 290 929 306
rect 1064 271 1098 392
rect 1192 356 1226 579
rect 1262 496 1328 543
rect 1478 537 1512 579
rect 1548 607 1614 649
rect 1548 573 1564 607
rect 1598 573 1614 607
rect 1760 607 1826 649
rect 1760 573 1776 607
rect 1810 573 1826 607
rect 2041 597 2107 613
rect 2041 563 2057 597
rect 2091 563 2107 597
rect 1478 503 1997 537
rect 1262 462 1278 496
rect 1312 462 1328 496
rect 1262 449 1328 462
rect 1262 415 1451 449
rect 1003 254 1098 271
rect 859 237 1098 254
rect 1134 340 1226 356
rect 1134 306 1151 340
rect 1185 326 1226 340
rect 1185 310 1381 326
rect 1185 306 1331 310
rect 1134 276 1331 306
rect 1365 276 1381 310
rect 1134 260 1381 276
rect 859 220 1037 237
rect 313 162 455 171
rect 491 152 735 186
rect 23 77 63 111
rect 97 77 113 111
rect 23 53 113 77
rect 211 106 277 135
rect 491 126 525 152
rect 211 72 227 106
rect 261 72 277 106
rect 211 17 277 72
rect 435 106 525 126
rect 435 72 451 106
rect 485 72 525 106
rect 435 53 525 72
rect 599 96 665 116
rect 599 62 615 96
rect 649 62 665 96
rect 599 17 665 62
rect 701 87 735 152
rect 773 179 823 201
rect 807 145 823 179
rect 773 123 823 145
rect 859 87 893 220
rect 701 53 893 87
rect 931 163 965 184
rect 931 17 965 129
rect 1003 87 1037 220
rect 1134 201 1168 260
rect 1073 179 1168 201
rect 1073 145 1089 179
rect 1123 145 1168 179
rect 1290 209 1356 213
rect 1417 209 1451 415
rect 1487 433 1670 467
rect 1704 433 1720 467
rect 1487 417 1720 433
rect 1487 352 1553 417
rect 1487 318 1503 352
rect 1537 318 1553 352
rect 1487 279 1553 318
rect 1601 365 1723 381
rect 1601 331 1617 365
rect 1651 331 1723 365
rect 1601 315 1723 331
rect 1487 245 1653 279
rect 1290 184 1583 209
rect 1073 123 1168 145
rect 1204 142 1254 171
rect 1238 108 1254 142
rect 1290 150 1306 184
rect 1340 175 1583 184
rect 1340 150 1356 175
rect 1290 121 1356 150
rect 1463 123 1513 139
rect 1204 87 1254 108
rect 1003 53 1254 87
rect 1463 89 1479 123
rect 1463 17 1513 89
rect 1549 87 1583 175
rect 1619 204 1653 245
rect 1689 274 1723 315
rect 1759 360 1813 376
rect 1759 350 1763 360
rect 1797 326 1813 360
rect 1793 316 1813 326
rect 1759 310 1813 316
rect 1855 358 1921 374
rect 1855 324 1871 358
rect 1905 324 1921 358
rect 1855 290 1921 324
rect 1855 274 1871 290
rect 1689 256 1871 274
rect 1905 256 1921 290
rect 1689 240 1921 256
rect 1963 355 1997 503
rect 2041 465 2107 563
rect 2302 611 2368 649
rect 2302 577 2318 611
rect 2352 577 2368 611
rect 2302 543 2368 577
rect 2302 509 2318 543
rect 2352 509 2368 543
rect 2302 493 2368 509
rect 2442 597 2673 613
rect 2442 563 2458 597
rect 2492 579 2673 597
rect 2041 431 2057 465
rect 2091 457 2107 465
rect 2442 465 2492 563
rect 2442 457 2458 465
rect 2091 431 2458 457
rect 2041 423 2492 431
rect 2041 415 2107 423
rect 2143 371 2196 387
rect 2143 355 2159 371
rect 1963 337 2159 355
rect 2193 337 2196 371
rect 1963 321 2196 337
rect 1963 281 2029 321
rect 1963 247 1979 281
rect 2013 247 2029 281
rect 1619 180 1704 204
rect 1619 146 1654 180
rect 1688 146 1704 180
rect 1619 123 1704 146
rect 1740 87 1774 240
rect 1963 231 2029 247
rect 2232 224 2266 423
rect 2442 415 2492 423
rect 2528 527 2603 543
rect 2528 493 2569 527
rect 2528 454 2603 493
rect 2528 420 2569 454
rect 2528 404 2603 420
rect 2302 361 2355 377
rect 2302 327 2305 361
rect 2339 327 2355 361
rect 2302 293 2355 327
rect 2397 362 2471 378
rect 2397 328 2413 362
rect 2447 350 2471 362
rect 2397 316 2431 328
rect 2465 316 2471 350
rect 2397 310 2471 316
rect 2302 259 2305 293
rect 2339 274 2355 293
rect 2528 274 2562 404
rect 2639 368 2673 579
rect 2709 588 2759 649
rect 2743 554 2759 588
rect 2709 517 2759 554
rect 2743 483 2759 517
rect 2709 446 2759 483
rect 2743 412 2759 446
rect 2709 396 2759 412
rect 2799 588 2849 604
rect 2799 554 2815 588
rect 2799 517 2849 554
rect 2799 483 2815 517
rect 2799 446 2849 483
rect 2799 412 2815 446
rect 2339 259 2562 274
rect 2302 240 2562 259
rect 2598 352 2673 368
rect 2799 356 2849 412
rect 2598 318 2614 352
rect 2648 318 2673 352
rect 2598 284 2673 318
rect 2598 250 2614 284
rect 2648 250 2673 284
rect 1549 53 1774 87
rect 1810 179 1876 204
rect 1810 145 1826 179
rect 1860 145 1876 179
rect 1810 17 1876 145
rect 2065 197 2266 224
rect 2065 163 2081 197
rect 2115 190 2266 197
rect 2115 163 2131 190
rect 2065 112 2131 163
rect 2065 78 2081 112
rect 2115 78 2131 112
rect 2065 62 2131 78
rect 2318 125 2384 154
rect 2318 91 2334 125
rect 2368 91 2384 125
rect 2318 17 2384 91
rect 2433 116 2499 240
rect 2598 234 2673 250
rect 2713 322 2849 356
rect 2892 562 2977 578
rect 2892 528 2927 562
rect 2961 528 2977 562
rect 2892 491 2977 528
rect 2892 457 2927 491
rect 2961 457 2977 491
rect 2892 420 2977 457
rect 2892 386 2927 420
rect 2961 386 2977 420
rect 2892 332 2977 386
rect 3017 562 3083 649
rect 3017 528 3033 562
rect 3067 528 3083 562
rect 3017 491 3083 528
rect 3017 457 3033 491
rect 3067 457 3083 491
rect 3017 420 3083 457
rect 3017 386 3033 420
rect 3067 386 3083 420
rect 3017 370 3083 386
rect 3123 562 3242 578
rect 3123 528 3139 562
rect 3173 528 3242 562
rect 3123 491 3242 528
rect 3123 457 3139 491
rect 3173 457 3242 491
rect 3123 420 3242 457
rect 3123 386 3139 420
rect 3173 386 3242 420
rect 3123 370 3242 386
rect 2713 145 2759 322
rect 2892 316 3145 332
rect 2892 298 3095 316
rect 2892 162 2926 298
rect 3079 282 3095 298
rect 3129 282 3145 316
rect 3079 248 3145 282
rect 3079 214 3095 248
rect 3129 214 3145 248
rect 3079 198 3145 214
rect 3208 162 3242 370
rect 2433 82 2449 116
rect 2483 82 2499 116
rect 2433 53 2499 82
rect 2591 116 2657 145
rect 2591 82 2607 116
rect 2641 82 2657 116
rect 2591 17 2657 82
rect 2713 116 2815 145
rect 2713 82 2765 116
rect 2799 82 2815 116
rect 2713 53 2815 82
rect 2860 133 2926 162
rect 2860 99 2876 133
rect 2910 99 2926 133
rect 2860 70 2926 99
rect 3018 133 3084 162
rect 3018 99 3034 133
rect 3068 99 3084 133
rect 3018 17 3084 99
rect 3176 133 3242 162
rect 3176 99 3192 133
rect 3226 99 3242 133
rect 3176 70 3242 99
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 1759 326 1763 350
rect 1763 326 1793 350
rect 1759 316 1793 326
rect 2431 328 2447 350
rect 2447 328 2465 350
rect 2431 316 2465 328
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
<< metal1 >>
rect 0 683 3264 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 0 617 3264 649
rect 1747 350 1805 356
rect 1747 316 1759 350
rect 1793 347 1805 350
rect 2419 350 2477 356
rect 2419 347 2431 350
rect 1793 319 2431 347
rect 1793 316 1805 319
rect 1747 310 1805 316
rect 2419 316 2431 319
rect 2465 316 2477 350
rect 2419 310 2477 316
rect 0 17 3264 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
rect 0 -49 3264 -17
<< labels >>
flabel pwell s 0 0 3264 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 3264 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfsbp_lp
flabel metal1 s 2431 316 2465 350 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel metal1 s 0 617 3264 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 3264 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2719 242 2753 276 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2719 316 2753 350 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3199 390 3233 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3199 464 3233 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3199 538 3233 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3264 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5593914
string GDS_START 5572226
<< end >>
