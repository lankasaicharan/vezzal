magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 564 235 858 241
rect 197 167 858 235
rect 1 49 858 167
rect 0 0 864 49
<< scnmos >>
rect 80 57 110 141
rect 276 125 306 209
rect 348 125 378 209
rect 420 125 450 209
rect 528 125 558 209
rect 643 47 673 215
rect 729 47 759 215
<< scpmoshvt >>
rect 106 375 136 459
rect 192 375 222 459
rect 278 375 308 459
rect 456 375 486 459
rect 551 375 581 459
rect 656 367 686 619
rect 742 367 772 619
<< ndiff >>
rect 27 116 80 141
rect 27 82 35 116
rect 69 82 80 116
rect 27 57 80 82
rect 110 116 163 141
rect 110 82 121 116
rect 155 82 163 116
rect 110 57 163 82
rect 590 209 643 215
rect 223 197 276 209
rect 223 163 231 197
rect 265 163 276 197
rect 223 125 276 163
rect 306 125 348 209
rect 378 125 420 209
rect 450 125 528 209
rect 558 125 643 209
rect 590 117 643 125
rect 590 83 598 117
rect 632 83 643 117
rect 590 47 643 83
rect 673 190 729 215
rect 673 156 684 190
rect 718 156 729 190
rect 673 101 729 156
rect 673 67 684 101
rect 718 67 729 101
rect 673 47 729 67
rect 759 202 832 215
rect 759 168 790 202
rect 824 168 832 202
rect 759 93 832 168
rect 759 59 770 93
rect 804 59 832 93
rect 759 47 832 59
<< pdiff >>
rect 603 607 656 619
rect 603 573 611 607
rect 645 573 656 607
rect 603 527 656 573
rect 603 493 611 527
rect 645 493 656 527
rect 603 459 656 493
rect 53 434 106 459
rect 53 400 61 434
rect 95 400 106 434
rect 53 375 106 400
rect 136 446 192 459
rect 136 412 147 446
rect 181 412 192 446
rect 136 375 192 412
rect 222 434 278 459
rect 222 400 233 434
rect 267 400 278 434
rect 222 375 278 400
rect 308 434 456 459
rect 308 400 319 434
rect 353 400 411 434
rect 445 400 456 434
rect 308 375 456 400
rect 486 434 551 459
rect 486 400 506 434
rect 540 400 551 434
rect 486 375 551 400
rect 581 444 656 459
rect 581 410 592 444
rect 626 410 656 444
rect 581 375 656 410
rect 603 367 656 375
rect 686 599 742 619
rect 686 565 697 599
rect 731 565 742 599
rect 686 504 742 565
rect 686 470 697 504
rect 731 470 742 504
rect 686 420 742 470
rect 686 386 697 420
rect 731 386 742 420
rect 686 367 742 386
rect 772 607 832 619
rect 772 573 783 607
rect 817 573 832 607
rect 772 511 832 573
rect 772 477 783 511
rect 817 477 832 511
rect 772 413 832 477
rect 772 379 790 413
rect 824 379 832 413
rect 772 367 832 379
<< ndiffc >>
rect 35 82 69 116
rect 121 82 155 116
rect 231 163 265 197
rect 598 83 632 117
rect 684 156 718 190
rect 684 67 718 101
rect 790 168 824 202
rect 770 59 804 93
<< pdiffc >>
rect 611 573 645 607
rect 611 493 645 527
rect 61 400 95 434
rect 147 412 181 446
rect 233 400 267 434
rect 319 400 353 434
rect 411 400 445 434
rect 506 400 540 434
rect 592 410 626 444
rect 697 565 731 599
rect 697 470 731 504
rect 697 386 731 420
rect 783 573 817 607
rect 783 477 817 511
rect 790 379 824 413
<< poly >>
rect 656 619 686 645
rect 742 619 772 645
rect 106 459 136 485
rect 192 459 222 485
rect 278 459 308 485
rect 456 459 486 485
rect 551 459 581 485
rect 106 297 136 375
rect 31 281 136 297
rect 31 247 47 281
rect 81 267 136 281
rect 81 247 110 267
rect 192 254 222 375
rect 278 343 308 375
rect 278 327 378 343
rect 278 293 317 327
rect 351 293 378 327
rect 456 308 486 375
rect 551 308 581 375
rect 656 308 686 367
rect 742 308 772 367
rect 278 277 378 293
rect 31 213 110 247
rect 31 179 47 213
rect 81 179 110 213
rect 31 163 110 179
rect 80 141 110 163
rect 178 224 222 254
rect 178 103 208 224
rect 276 209 306 235
rect 348 209 378 277
rect 420 292 486 308
rect 420 258 436 292
rect 470 258 486 292
rect 420 242 486 258
rect 528 292 594 308
rect 528 258 544 292
rect 578 258 594 292
rect 528 242 594 258
rect 636 292 772 308
rect 636 258 652 292
rect 686 258 772 292
rect 636 242 772 258
rect 420 209 450 242
rect 528 209 558 242
rect 643 215 673 242
rect 729 215 759 242
rect 276 103 306 125
rect 178 87 306 103
rect 348 99 378 125
rect 420 99 450 125
rect 528 99 558 125
rect 80 31 110 57
rect 178 53 201 87
rect 235 53 306 87
rect 178 37 306 53
rect 643 21 673 47
rect 729 21 759 47
<< polycont >>
rect 47 247 81 281
rect 317 293 351 327
rect 47 179 81 213
rect 436 258 470 292
rect 544 258 578 292
rect 652 258 686 292
rect 201 53 235 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 45 434 95 450
rect 45 400 61 434
rect 131 446 197 649
rect 131 412 147 446
rect 181 412 197 446
rect 131 407 197 412
rect 231 434 281 450
rect 45 373 95 400
rect 231 400 233 434
rect 267 400 281 434
rect 45 339 159 373
rect 17 281 85 297
rect 17 247 47 281
rect 81 247 85 281
rect 17 213 85 247
rect 17 179 47 213
rect 81 179 85 213
rect 17 163 85 179
rect 19 116 85 129
rect 19 82 35 116
rect 69 82 85 116
rect 19 17 85 82
rect 119 119 159 339
rect 231 201 281 400
rect 315 434 461 649
rect 576 607 661 649
rect 576 573 611 607
rect 645 573 661 607
rect 576 527 661 573
rect 576 493 611 527
rect 645 493 661 527
rect 315 400 319 434
rect 353 400 411 434
rect 445 400 461 434
rect 315 384 461 400
rect 504 434 542 450
rect 504 400 506 434
rect 540 400 542 434
rect 576 444 661 493
rect 576 410 592 444
rect 626 410 661 444
rect 695 599 740 615
rect 695 565 697 599
rect 731 565 740 599
rect 695 504 740 565
rect 695 470 697 504
rect 731 470 740 504
rect 695 420 740 470
rect 504 376 542 400
rect 695 386 697 420
rect 731 386 740 420
rect 777 607 840 649
rect 777 573 783 607
rect 817 573 840 607
rect 777 511 840 573
rect 777 477 783 511
rect 817 477 840 511
rect 777 413 840 477
rect 777 410 790 413
rect 695 376 740 386
rect 824 379 840 413
rect 315 327 367 350
rect 315 293 317 327
rect 351 293 367 327
rect 315 242 367 293
rect 401 292 470 350
rect 504 342 648 376
rect 695 342 756 376
rect 790 363 840 379
rect 614 308 648 342
rect 401 258 436 292
rect 401 235 470 258
rect 504 292 578 308
rect 504 258 544 292
rect 504 235 578 258
rect 614 292 686 308
rect 614 258 652 292
rect 614 242 686 258
rect 614 201 648 242
rect 720 208 756 342
rect 215 197 648 201
rect 215 163 231 197
rect 265 163 648 197
rect 215 159 648 163
rect 682 190 756 208
rect 682 156 684 190
rect 718 172 756 190
rect 790 202 840 219
rect 718 156 732 172
rect 119 116 251 119
rect 119 82 121 116
rect 155 87 251 116
rect 155 82 201 87
rect 119 53 201 82
rect 235 53 251 87
rect 119 51 251 53
rect 582 117 648 125
rect 582 83 598 117
rect 632 83 648 117
rect 582 17 648 83
rect 682 101 732 156
rect 824 168 840 202
rect 790 138 840 168
rect 682 67 684 101
rect 718 67 732 101
rect 682 51 732 67
rect 766 93 840 138
rect 766 59 770 93
rect 804 59 840 93
rect 766 17 840 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4b_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5361838
string GDS_START 5354064
<< end >>
