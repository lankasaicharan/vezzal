magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3698 1975
<< nwell >>
rect -38 331 2438 704
rect 1747 303 1959 331
<< pwell >>
rect 1951 241 2397 245
rect 65 161 739 233
rect 944 215 1339 235
rect 944 171 1511 215
rect 1751 171 2397 241
rect 944 161 2397 171
rect 65 49 2397 161
rect 0 0 2400 49
<< scnmos >>
rect 144 123 174 207
rect 230 123 260 207
rect 329 123 359 207
rect 453 123 483 207
rect 525 123 555 207
rect 611 123 641 207
rect 820 51 850 135
rect 1023 125 1053 209
rect 1113 125 1143 209
rect 1203 125 1233 209
rect 1398 61 1428 189
rect 1507 61 1537 145
rect 1640 61 1670 145
rect 1725 61 1755 145
rect 1830 47 1860 215
rect 2030 51 2060 219
rect 2116 51 2146 219
rect 2202 51 2232 219
rect 2288 51 2318 219
<< scpmoshvt >>
rect 180 491 210 619
rect 266 491 296 619
rect 338 491 368 619
rect 424 491 454 619
rect 518 491 548 619
rect 611 491 641 619
rect 855 481 885 609
rect 1045 463 1075 547
rect 1169 449 1199 533
rect 1241 449 1271 533
rect 1359 449 1389 617
rect 1445 449 1475 617
rect 1601 507 1631 591
rect 1673 507 1703 591
rect 1840 339 1870 591
rect 2030 367 2060 619
rect 2116 367 2146 619
rect 2202 367 2232 619
rect 2288 367 2318 619
<< ndiff >>
rect 91 177 144 207
rect 91 143 99 177
rect 133 143 144 177
rect 91 123 144 143
rect 174 182 230 207
rect 174 148 185 182
rect 219 148 230 182
rect 174 123 230 148
rect 260 123 329 207
rect 359 195 453 207
rect 359 161 389 195
rect 423 161 453 195
rect 359 123 453 161
rect 483 123 525 207
rect 555 169 611 207
rect 555 135 566 169
rect 600 135 611 169
rect 555 123 611 135
rect 641 195 713 207
rect 641 161 671 195
rect 705 161 713 195
rect 641 123 713 161
rect 970 183 1023 209
rect 970 149 978 183
rect 1012 149 1023 183
rect 767 107 820 135
rect 767 73 775 107
rect 809 73 820 107
rect 767 51 820 73
rect 850 103 903 135
rect 970 125 1023 149
rect 1053 183 1113 209
rect 1053 149 1068 183
rect 1102 149 1113 183
rect 1053 125 1113 149
rect 1143 125 1203 209
rect 1233 189 1313 209
rect 1233 125 1398 189
rect 850 69 861 103
rect 895 69 903 103
rect 850 51 903 69
rect 1255 75 1398 125
rect 1255 41 1267 75
rect 1301 61 1398 75
rect 1428 161 1485 189
rect 1428 127 1439 161
rect 1473 145 1485 161
rect 1777 187 1830 215
rect 1777 153 1785 187
rect 1819 153 1830 187
rect 1777 145 1830 153
rect 1473 127 1507 145
rect 1428 61 1507 127
rect 1537 119 1640 145
rect 1537 85 1595 119
rect 1629 85 1640 119
rect 1537 61 1640 85
rect 1670 61 1725 145
rect 1755 93 1830 145
rect 1755 61 1785 93
rect 1301 41 1313 61
rect 1255 33 1313 41
rect 1777 59 1785 61
rect 1819 59 1830 93
rect 1777 47 1830 59
rect 1860 185 1913 215
rect 1860 151 1871 185
rect 1905 151 1913 185
rect 1860 101 1913 151
rect 1860 67 1871 101
rect 1905 67 1913 101
rect 1860 47 1913 67
rect 1977 207 2030 219
rect 1977 173 1985 207
rect 2019 173 2030 207
rect 1977 97 2030 173
rect 1977 63 1985 97
rect 2019 63 2030 97
rect 1977 51 2030 63
rect 2060 205 2116 219
rect 2060 171 2071 205
rect 2105 171 2116 205
rect 2060 101 2116 171
rect 2060 67 2071 101
rect 2105 67 2116 101
rect 2060 51 2116 67
rect 2146 143 2202 219
rect 2146 109 2157 143
rect 2191 109 2202 143
rect 2146 51 2202 109
rect 2232 205 2288 219
rect 2232 171 2243 205
rect 2277 171 2288 205
rect 2232 101 2288 171
rect 2232 67 2243 101
rect 2277 67 2288 101
rect 2232 51 2288 67
rect 2318 143 2371 219
rect 2318 109 2329 143
rect 2363 109 2371 143
rect 2318 51 2371 109
<< pdiff >>
rect 127 573 180 619
rect 127 539 135 573
rect 169 539 180 573
rect 127 491 180 539
rect 210 578 266 619
rect 210 544 221 578
rect 255 544 266 578
rect 210 491 266 544
rect 296 491 338 619
rect 368 578 424 619
rect 368 544 379 578
rect 413 544 424 578
rect 368 491 424 544
rect 454 491 518 619
rect 548 582 611 619
rect 548 548 566 582
rect 600 548 611 582
rect 548 491 611 548
rect 641 607 694 619
rect 1286 631 1344 639
rect 641 573 652 607
rect 686 573 694 607
rect 641 539 694 573
rect 641 505 652 539
rect 686 505 694 539
rect 641 491 694 505
rect 748 578 855 609
rect 748 544 756 578
rect 790 544 855 578
rect 748 481 855 544
rect 885 529 938 609
rect 1286 597 1298 631
rect 1332 617 1344 631
rect 1332 597 1359 617
rect 885 495 896 529
rect 930 495 938 529
rect 885 481 938 495
rect 992 509 1045 547
rect 992 475 1000 509
rect 1034 475 1045 509
rect 992 463 1045 475
rect 1075 533 1147 547
rect 1286 533 1359 597
rect 1075 513 1169 533
rect 1075 479 1105 513
rect 1139 479 1169 513
rect 1075 463 1169 479
rect 1097 449 1169 463
rect 1199 449 1241 533
rect 1271 449 1359 533
rect 1389 491 1445 617
rect 1389 457 1400 491
rect 1434 457 1445 491
rect 1389 449 1445 457
rect 1475 591 1525 617
rect 1977 607 2030 619
rect 1475 566 1601 591
rect 1475 532 1556 566
rect 1590 532 1601 566
rect 1475 507 1601 532
rect 1631 507 1673 591
rect 1703 583 1840 591
rect 1703 566 1795 583
rect 1703 532 1714 566
rect 1748 549 1795 566
rect 1829 549 1840 583
rect 1748 532 1840 549
rect 1703 515 1840 532
rect 1703 507 1795 515
rect 1475 449 1525 507
rect 1783 481 1795 507
rect 1829 481 1840 515
rect 1783 339 1840 481
rect 1870 579 1923 591
rect 1870 545 1881 579
rect 1915 545 1923 579
rect 1870 484 1923 545
rect 1870 450 1881 484
rect 1915 450 1923 484
rect 1870 389 1923 450
rect 1870 355 1881 389
rect 1915 355 1923 389
rect 1977 573 1985 607
rect 2019 573 2030 607
rect 1977 512 2030 573
rect 1977 478 1985 512
rect 2019 478 2030 512
rect 1977 413 2030 478
rect 1977 379 1985 413
rect 2019 379 2030 413
rect 1977 367 2030 379
rect 2060 599 2116 619
rect 2060 565 2071 599
rect 2105 565 2116 599
rect 2060 512 2116 565
rect 2060 478 2071 512
rect 2105 478 2116 512
rect 2060 413 2116 478
rect 2060 379 2071 413
rect 2105 379 2116 413
rect 2060 367 2116 379
rect 2146 607 2202 619
rect 2146 573 2157 607
rect 2191 573 2202 607
rect 2146 519 2202 573
rect 2146 485 2157 519
rect 2191 485 2202 519
rect 2146 433 2202 485
rect 2146 399 2157 433
rect 2191 399 2202 433
rect 2146 367 2202 399
rect 2232 599 2288 619
rect 2232 565 2243 599
rect 2277 565 2288 599
rect 2232 512 2288 565
rect 2232 478 2243 512
rect 2277 478 2288 512
rect 2232 413 2288 478
rect 2232 379 2243 413
rect 2277 379 2288 413
rect 2232 367 2288 379
rect 2318 607 2371 619
rect 2318 573 2329 607
rect 2363 573 2371 607
rect 2318 530 2371 573
rect 2318 496 2329 530
rect 2363 496 2371 530
rect 2318 453 2371 496
rect 2318 419 2329 453
rect 2363 419 2371 453
rect 2318 367 2371 419
rect 1870 339 1923 355
<< ndiffc >>
rect 99 143 133 177
rect 185 148 219 182
rect 389 161 423 195
rect 566 135 600 169
rect 671 161 705 195
rect 978 149 1012 183
rect 775 73 809 107
rect 1068 149 1102 183
rect 861 69 895 103
rect 1267 41 1301 75
rect 1439 127 1473 161
rect 1785 153 1819 187
rect 1595 85 1629 119
rect 1785 59 1819 93
rect 1871 151 1905 185
rect 1871 67 1905 101
rect 1985 173 2019 207
rect 1985 63 2019 97
rect 2071 171 2105 205
rect 2071 67 2105 101
rect 2157 109 2191 143
rect 2243 171 2277 205
rect 2243 67 2277 101
rect 2329 109 2363 143
<< pdiffc >>
rect 135 539 169 573
rect 221 544 255 578
rect 379 544 413 578
rect 566 548 600 582
rect 652 573 686 607
rect 652 505 686 539
rect 756 544 790 578
rect 1298 597 1332 631
rect 896 495 930 529
rect 1000 475 1034 509
rect 1105 479 1139 513
rect 1400 457 1434 491
rect 1556 532 1590 566
rect 1714 532 1748 566
rect 1795 549 1829 583
rect 1795 481 1829 515
rect 1881 545 1915 579
rect 1881 450 1915 484
rect 1881 355 1915 389
rect 1985 573 2019 607
rect 1985 478 2019 512
rect 1985 379 2019 413
rect 2071 565 2105 599
rect 2071 478 2105 512
rect 2071 379 2105 413
rect 2157 573 2191 607
rect 2157 485 2191 519
rect 2157 399 2191 433
rect 2243 565 2277 599
rect 2243 478 2277 512
rect 2243 379 2277 413
rect 2329 573 2363 607
rect 2329 496 2363 530
rect 2329 419 2363 453
<< poly >>
rect 180 619 210 645
rect 266 619 296 645
rect 338 619 368 645
rect 424 619 454 645
rect 518 619 548 645
rect 611 619 641 645
rect 855 609 885 635
rect 180 453 210 491
rect 266 453 296 491
rect 80 423 296 453
rect 80 295 110 423
rect 188 365 254 381
rect 188 331 204 365
rect 238 345 254 365
rect 338 363 368 491
rect 424 459 454 491
rect 410 443 476 459
rect 410 409 426 443
rect 460 409 476 443
rect 410 393 476 409
rect 302 347 368 363
rect 238 331 260 345
rect 188 315 260 331
rect 80 279 146 295
rect 80 245 96 279
rect 130 259 146 279
rect 130 245 174 259
rect 80 229 174 245
rect 144 207 174 229
rect 230 207 260 315
rect 302 313 318 347
rect 352 313 368 347
rect 518 345 548 491
rect 611 376 641 491
rect 1359 617 1389 643
rect 1445 617 1475 643
rect 2030 619 2060 645
rect 2116 619 2146 645
rect 2202 619 2232 645
rect 2288 619 2318 645
rect 1045 547 1075 573
rect 855 459 885 481
rect 1169 533 1199 559
rect 1241 533 1271 559
rect 820 429 885 459
rect 1045 441 1075 463
rect 1601 591 1631 617
rect 1673 591 1703 617
rect 1840 591 1870 617
rect 611 360 701 376
rect 302 279 368 313
rect 489 329 555 345
rect 489 295 505 329
rect 539 295 555 329
rect 489 279 555 295
rect 302 245 318 279
rect 352 245 368 279
rect 302 229 368 245
rect 329 207 359 229
rect 453 207 483 233
rect 525 207 555 279
rect 611 326 651 360
rect 685 326 701 360
rect 611 292 701 326
rect 611 258 651 292
rect 685 258 701 292
rect 820 291 850 429
rect 934 411 1075 441
rect 934 381 964 411
rect 611 242 701 258
rect 784 275 850 291
rect 611 207 641 242
rect 784 241 800 275
rect 834 241 850 275
rect 898 365 964 381
rect 1169 369 1199 449
rect 898 331 914 365
rect 948 331 964 365
rect 898 297 964 331
rect 898 263 914 297
rect 948 263 964 297
rect 898 247 964 263
rect 1023 353 1199 369
rect 1023 319 1149 353
rect 1183 319 1199 353
rect 1023 303 1199 319
rect 1241 415 1271 449
rect 1241 399 1311 415
rect 1241 365 1261 399
rect 1295 365 1311 399
rect 1241 331 1311 365
rect 784 207 850 241
rect 1023 209 1053 303
rect 1241 297 1261 331
rect 1295 297 1311 331
rect 1241 281 1311 297
rect 1241 261 1271 281
rect 1359 277 1389 449
rect 1445 417 1475 449
rect 1445 401 1520 417
rect 1445 367 1470 401
rect 1504 367 1520 401
rect 1445 351 1520 367
rect 1601 309 1631 507
rect 1673 475 1703 507
rect 1673 459 1755 475
rect 1673 425 1701 459
rect 1735 425 1755 459
rect 1673 409 1755 425
rect 1539 279 1631 309
rect 1113 209 1143 235
rect 1203 231 1271 261
rect 1353 261 1428 277
rect 1203 209 1233 231
rect 1353 227 1369 261
rect 1403 227 1428 261
rect 1539 233 1569 279
rect 1353 211 1428 227
rect 784 173 800 207
rect 834 173 850 207
rect 784 157 850 173
rect 820 135 850 157
rect 144 55 174 123
rect 230 97 260 123
rect 329 97 359 123
rect 453 55 483 123
rect 525 97 555 123
rect 611 97 641 123
rect 144 25 483 55
rect 1398 189 1428 211
rect 1507 217 1575 233
rect 1023 99 1053 125
rect 1113 103 1143 125
rect 1095 87 1161 103
rect 1203 99 1233 125
rect 1095 53 1111 87
rect 1145 53 1161 87
rect 820 25 850 51
rect 1095 37 1161 53
rect 1507 183 1525 217
rect 1559 183 1575 217
rect 1507 167 1575 183
rect 1617 221 1683 237
rect 1617 187 1633 221
rect 1667 187 1683 221
rect 1617 171 1683 187
rect 1507 145 1537 167
rect 1640 145 1670 171
rect 1725 145 1755 409
rect 1840 303 1870 339
rect 2030 307 2060 367
rect 2116 307 2146 367
rect 2202 307 2232 367
rect 2288 307 2318 367
rect 1797 287 1870 303
rect 1797 253 1813 287
rect 1847 253 1870 287
rect 1797 237 1870 253
rect 1933 291 2318 307
rect 1933 257 1949 291
rect 1983 257 2017 291
rect 2051 257 2085 291
rect 2119 257 2153 291
rect 2187 257 2318 291
rect 1933 241 2318 257
rect 1830 215 1860 237
rect 2030 219 2060 241
rect 2116 219 2146 241
rect 2202 219 2232 241
rect 2288 219 2318 241
rect 1398 35 1428 61
rect 1507 35 1537 61
rect 1640 35 1670 61
rect 1725 35 1755 61
rect 1830 21 1860 47
rect 2030 25 2060 51
rect 2116 25 2146 51
rect 2202 25 2232 51
rect 2288 25 2318 51
<< polycont >>
rect 204 331 238 365
rect 426 409 460 443
rect 96 245 130 279
rect 318 313 352 347
rect 505 295 539 329
rect 318 245 352 279
rect 651 326 685 360
rect 651 258 685 292
rect 800 241 834 275
rect 914 331 948 365
rect 914 263 948 297
rect 1149 319 1183 353
rect 1261 365 1295 399
rect 1261 297 1295 331
rect 1470 367 1504 401
rect 1701 425 1735 459
rect 1369 227 1403 261
rect 800 173 834 207
rect 1111 53 1145 87
rect 1525 183 1559 217
rect 1633 187 1667 221
rect 1813 253 1847 287
rect 1949 257 1983 291
rect 2017 257 2051 291
rect 2085 257 2119 291
rect 2153 257 2187 291
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 26 573 171 589
rect 26 539 135 573
rect 169 539 171 573
rect 26 494 171 539
rect 205 578 271 649
rect 205 544 221 578
rect 255 544 271 578
rect 205 528 271 544
rect 363 578 530 594
rect 363 544 379 578
rect 413 544 530 578
rect 363 528 530 544
rect 564 582 602 649
rect 564 548 566 582
rect 600 548 602 582
rect 564 532 602 548
rect 636 607 702 615
rect 636 573 652 607
rect 686 573 702 607
rect 636 539 702 573
rect 496 498 530 528
rect 636 505 652 539
rect 686 505 702 539
rect 740 578 792 649
rect 1282 631 1348 649
rect 740 544 756 578
rect 790 544 792 578
rect 740 528 792 544
rect 826 579 1209 613
rect 1282 597 1298 631
rect 1332 597 1348 631
rect 1282 595 1348 597
rect 1699 583 1845 649
rect 1969 607 2028 649
rect 636 501 702 505
rect 26 460 462 494
rect 26 365 254 460
rect 410 443 462 460
rect 26 331 204 365
rect 238 331 254 365
rect 302 347 355 426
rect 410 409 426 443
rect 460 409 462 443
rect 496 464 511 498
rect 545 467 602 498
rect 668 494 702 501
rect 826 494 860 579
rect 1175 561 1209 579
rect 1554 566 1665 582
rect 545 464 615 467
rect 496 431 615 464
rect 668 460 860 494
rect 410 393 462 409
rect 26 193 62 331
rect 302 313 318 347
rect 352 313 355 347
rect 96 279 268 295
rect 130 245 268 279
rect 96 229 268 245
rect 302 279 355 313
rect 389 329 545 359
rect 389 295 505 329
rect 539 295 545 329
rect 389 279 545 295
rect 302 245 318 279
rect 352 245 355 279
rect 26 177 135 193
rect 26 143 99 177
rect 133 143 135 177
rect 26 127 135 143
rect 169 182 235 195
rect 169 148 185 182
rect 219 148 235 182
rect 169 17 235 148
rect 302 94 355 245
rect 581 243 615 431
rect 389 209 615 243
rect 651 360 739 424
rect 685 326 739 360
rect 651 292 739 326
rect 685 258 739 292
rect 651 238 739 258
rect 773 275 860 460
rect 773 241 800 275
rect 834 241 860 275
rect 389 195 427 209
rect 773 207 860 241
rect 773 204 800 207
rect 423 161 427 195
rect 655 195 800 204
rect 389 145 427 161
rect 550 169 616 175
rect 550 135 566 169
rect 600 135 616 169
rect 655 161 671 195
rect 705 173 800 195
rect 834 173 860 207
rect 705 161 860 173
rect 655 157 860 161
rect 894 529 950 545
rect 894 495 896 529
rect 930 495 950 529
rect 894 365 950 495
rect 894 331 914 365
rect 948 331 950 365
rect 894 297 950 331
rect 894 263 914 297
rect 948 263 950 297
rect 894 247 950 263
rect 984 509 1038 525
rect 984 498 1000 509
rect 984 464 991 498
rect 1034 475 1038 509
rect 1025 464 1038 475
rect 984 459 1038 464
rect 1072 513 1141 545
rect 1072 479 1105 513
rect 1139 479 1141 513
rect 550 17 616 135
rect 759 107 825 123
rect 894 119 933 247
rect 984 199 1030 459
rect 1072 445 1141 479
rect 1175 527 1520 561
rect 1072 261 1108 445
rect 1175 369 1209 527
rect 1384 491 1450 493
rect 1384 457 1400 491
rect 1434 457 1450 491
rect 1384 441 1450 457
rect 1384 415 1418 441
rect 1142 353 1209 369
rect 1142 319 1149 353
rect 1183 319 1209 353
rect 1142 303 1209 319
rect 1245 399 1418 415
rect 1486 407 1520 527
rect 1554 532 1556 566
rect 1590 532 1665 566
rect 1554 516 1665 532
rect 1699 566 1795 583
rect 1699 532 1714 566
rect 1748 549 1795 566
rect 1829 549 1845 583
rect 1748 532 1845 549
rect 1699 516 1845 532
rect 1245 365 1261 399
rect 1295 365 1418 399
rect 1454 401 1520 407
rect 1454 367 1470 401
rect 1504 367 1595 401
rect 1454 365 1595 367
rect 1245 331 1418 365
rect 1245 297 1261 331
rect 1295 297 1489 331
rect 1245 295 1489 297
rect 1072 227 1369 261
rect 1403 227 1419 261
rect 1072 224 1419 227
rect 967 183 1030 199
rect 967 149 978 183
rect 1012 149 1030 183
rect 967 133 1030 149
rect 1064 211 1419 224
rect 1064 183 1110 211
rect 1064 149 1068 183
rect 1102 149 1110 183
rect 1455 177 1489 295
rect 1561 303 1595 365
rect 1631 373 1665 516
rect 1779 515 1845 516
rect 1779 481 1795 515
rect 1829 481 1845 515
rect 1879 579 1919 595
rect 1879 545 1881 579
rect 1915 545 1919 579
rect 1879 484 1919 545
rect 1699 459 1745 475
rect 1699 425 1701 459
rect 1735 443 1745 459
rect 1879 450 1881 484
rect 1915 450 1919 484
rect 1879 443 1919 450
rect 1735 425 1919 443
rect 1699 409 1919 425
rect 1881 389 1919 409
rect 1631 339 1737 373
rect 1703 303 1737 339
rect 1915 355 1919 389
rect 1969 573 1985 607
rect 2019 573 2028 607
rect 1969 512 2028 573
rect 1969 478 1985 512
rect 2019 478 2028 512
rect 1969 413 2028 478
rect 1969 379 1985 413
rect 2019 379 2028 413
rect 1969 363 2028 379
rect 2062 599 2107 615
rect 2062 565 2071 599
rect 2105 565 2107 599
rect 2062 512 2107 565
rect 2062 478 2071 512
rect 2105 478 2107 512
rect 2062 413 2107 478
rect 2062 379 2071 413
rect 2105 379 2107 413
rect 2141 607 2207 649
rect 2141 573 2157 607
rect 2191 573 2207 607
rect 2141 519 2207 573
rect 2141 485 2157 519
rect 2191 485 2207 519
rect 2141 433 2207 485
rect 2141 399 2157 433
rect 2191 399 2207 433
rect 2241 599 2279 615
rect 2241 565 2243 599
rect 2277 565 2279 599
rect 2241 512 2279 565
rect 2241 478 2243 512
rect 2277 478 2279 512
rect 2241 413 2279 478
rect 2313 607 2379 649
rect 2313 573 2329 607
rect 2363 573 2379 607
rect 2313 530 2379 573
rect 2313 496 2329 530
rect 2363 496 2379 530
rect 2313 453 2379 496
rect 2313 419 2329 453
rect 2363 419 2379 453
rect 2062 365 2107 379
rect 2241 379 2243 413
rect 2277 385 2279 413
rect 2277 379 2382 385
rect 2241 365 2382 379
rect 1561 269 1667 303
rect 1064 133 1110 149
rect 1423 161 1489 177
rect 759 73 775 107
rect 809 73 825 107
rect 759 17 825 73
rect 859 103 933 119
rect 859 69 861 103
rect 895 99 933 103
rect 1144 111 1387 145
rect 1423 127 1439 161
rect 1473 127 1489 161
rect 1423 119 1489 127
rect 1523 217 1559 233
rect 1523 183 1525 217
rect 1144 99 1178 111
rect 895 87 1178 99
rect 895 69 1111 87
rect 859 53 1111 69
rect 1145 53 1178 87
rect 1353 85 1387 111
rect 1523 85 1559 183
rect 1595 221 1667 269
rect 1595 187 1633 221
rect 1595 171 1667 187
rect 1703 287 1847 303
rect 1703 253 1813 287
rect 1703 237 1847 253
rect 1881 297 1919 355
rect 2062 331 2382 365
rect 1881 291 2203 297
rect 1881 257 1949 291
rect 1983 257 2017 291
rect 2051 257 2085 291
rect 2119 257 2153 291
rect 2187 257 2203 291
rect 1703 135 1737 237
rect 859 51 1178 53
rect 1251 75 1317 77
rect 1251 41 1267 75
rect 1301 41 1317 75
rect 1353 51 1559 85
rect 1593 119 1737 135
rect 1593 85 1595 119
rect 1629 85 1737 119
rect 1593 69 1737 85
rect 1771 187 1835 203
rect 1881 201 1921 257
rect 2239 223 2382 331
rect 1771 153 1785 187
rect 1819 153 1835 187
rect 1771 93 1835 153
rect 1771 59 1785 93
rect 1819 59 1835 93
rect 1251 17 1317 41
rect 1771 17 1835 59
rect 1869 185 1921 201
rect 1869 151 1871 185
rect 1905 151 1921 185
rect 1869 101 1921 151
rect 1869 67 1871 101
rect 1905 67 1921 101
rect 1869 51 1921 67
rect 1969 207 2027 223
rect 1969 173 1985 207
rect 2019 173 2027 207
rect 1969 97 2027 173
rect 1969 63 1985 97
rect 2019 63 2027 97
rect 1969 17 2027 63
rect 2061 205 2382 223
rect 2061 171 2071 205
rect 2105 189 2243 205
rect 2105 171 2107 189
rect 2061 101 2107 171
rect 2241 171 2243 189
rect 2277 189 2382 205
rect 2277 171 2279 189
rect 2061 67 2071 101
rect 2105 67 2107 101
rect 2061 51 2107 67
rect 2141 143 2207 155
rect 2141 109 2157 143
rect 2191 109 2207 143
rect 2141 17 2207 109
rect 2241 101 2279 171
rect 2241 67 2243 101
rect 2277 67 2279 101
rect 2241 51 2279 67
rect 2313 143 2379 155
rect 2313 109 2329 143
rect 2363 109 2379 143
rect 2313 17 2379 109
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 511 464 545 498
rect 991 475 1000 498
rect 1000 475 1025 498
rect 991 464 1025 475
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 499 498 557 504
rect 499 464 511 498
rect 545 495 557 498
rect 979 498 1037 504
rect 979 495 991 498
rect 545 467 991 495
rect 545 464 557 467
rect 499 458 557 464
rect 979 464 991 467
rect 1025 464 1037 498
rect 979 458 1037 464
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< labels >>
flabel pwell s 0 0 2400 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2400 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfxtp_4
flabel metal1 s 0 617 2400 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2400 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2239 242 2273 276 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2335 242 2369 276 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2400 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4054852
string GDS_START 4036452
<< end >>
