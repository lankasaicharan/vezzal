magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 23 49 1605 241
rect 0 0 1632 49
<< scnmos >>
rect 102 47 132 215
rect 188 47 218 215
rect 274 47 304 215
rect 360 47 390 215
rect 446 47 476 215
rect 532 47 562 215
rect 618 47 648 215
rect 704 47 734 215
rect 790 47 820 215
rect 876 47 906 215
rect 976 47 1006 215
rect 1062 47 1092 215
rect 1148 47 1178 215
rect 1234 47 1264 215
rect 1394 47 1424 215
rect 1480 47 1510 215
<< scpmoshvt >>
rect 102 367 132 619
rect 188 367 218 619
rect 274 367 304 619
rect 360 367 390 619
rect 446 367 476 619
rect 532 367 562 619
rect 618 367 648 619
rect 704 367 734 619
rect 790 367 820 619
rect 876 367 906 619
rect 962 367 992 619
rect 1048 367 1078 619
rect 1188 367 1218 619
rect 1274 367 1304 619
rect 1406 367 1436 619
rect 1512 367 1542 619
<< ndiff >>
rect 49 165 102 215
rect 49 131 57 165
rect 91 131 102 165
rect 49 93 102 131
rect 49 59 57 93
rect 91 59 102 93
rect 49 47 102 59
rect 132 181 188 215
rect 132 147 143 181
rect 177 147 188 181
rect 132 101 188 147
rect 132 67 143 101
rect 177 67 188 101
rect 132 47 188 67
rect 218 105 274 215
rect 218 71 229 105
rect 263 71 274 105
rect 218 47 274 71
rect 304 181 360 215
rect 304 147 315 181
rect 349 147 360 181
rect 304 101 360 147
rect 304 67 315 101
rect 349 67 360 101
rect 304 47 360 67
rect 390 105 446 215
rect 390 71 401 105
rect 435 71 446 105
rect 390 47 446 71
rect 476 181 532 215
rect 476 147 487 181
rect 521 147 532 181
rect 476 101 532 147
rect 476 67 487 101
rect 521 67 532 101
rect 476 47 532 67
rect 562 105 618 215
rect 562 71 573 105
rect 607 71 618 105
rect 562 47 618 71
rect 648 203 704 215
rect 648 169 659 203
rect 693 169 704 203
rect 648 101 704 169
rect 648 67 659 101
rect 693 67 704 101
rect 648 47 704 67
rect 734 157 790 215
rect 734 123 745 157
rect 779 123 790 157
rect 734 89 790 123
rect 734 55 745 89
rect 779 55 790 89
rect 734 47 790 55
rect 820 203 876 215
rect 820 169 831 203
rect 865 169 876 203
rect 820 135 876 169
rect 820 101 831 135
rect 865 101 876 135
rect 820 47 876 101
rect 906 157 976 215
rect 906 123 926 157
rect 960 123 976 157
rect 906 89 976 123
rect 906 55 926 89
rect 960 55 976 89
rect 906 47 976 55
rect 1006 203 1062 215
rect 1006 169 1017 203
rect 1051 169 1062 203
rect 1006 101 1062 169
rect 1006 67 1017 101
rect 1051 67 1062 101
rect 1006 47 1062 67
rect 1092 190 1148 215
rect 1092 156 1103 190
rect 1137 156 1148 190
rect 1092 47 1148 156
rect 1178 93 1234 215
rect 1178 59 1189 93
rect 1223 59 1234 93
rect 1178 47 1234 59
rect 1264 190 1394 215
rect 1264 156 1275 190
rect 1309 156 1349 190
rect 1383 156 1394 190
rect 1264 47 1394 156
rect 1424 163 1480 215
rect 1424 129 1435 163
rect 1469 129 1480 163
rect 1424 91 1480 129
rect 1424 57 1435 91
rect 1469 57 1480 91
rect 1424 47 1480 57
rect 1510 165 1579 215
rect 1510 131 1537 165
rect 1571 131 1579 165
rect 1510 93 1579 131
rect 1510 59 1537 93
rect 1571 59 1579 93
rect 1510 47 1579 59
<< pdiff >>
rect 49 599 102 619
rect 49 565 57 599
rect 91 565 102 599
rect 49 507 102 565
rect 49 473 57 507
rect 91 473 102 507
rect 49 413 102 473
rect 49 379 57 413
rect 91 379 102 413
rect 49 367 102 379
rect 132 607 188 619
rect 132 573 143 607
rect 177 573 188 607
rect 132 536 188 573
rect 132 502 143 536
rect 177 502 188 536
rect 132 465 188 502
rect 132 431 143 465
rect 177 431 188 465
rect 132 367 188 431
rect 218 572 274 619
rect 218 538 229 572
rect 263 538 274 572
rect 218 367 274 538
rect 304 607 360 619
rect 304 573 315 607
rect 349 573 360 607
rect 304 504 360 573
rect 304 470 315 504
rect 349 470 360 504
rect 304 367 360 470
rect 390 572 446 619
rect 390 538 401 572
rect 435 538 446 572
rect 390 367 446 538
rect 476 611 532 619
rect 476 577 487 611
rect 521 577 532 611
rect 476 539 532 577
rect 476 505 487 539
rect 521 505 532 539
rect 476 465 532 505
rect 476 431 487 465
rect 521 431 532 465
rect 476 367 532 431
rect 562 527 618 619
rect 562 493 573 527
rect 607 493 618 527
rect 562 413 618 493
rect 562 379 573 413
rect 607 379 618 413
rect 562 367 618 379
rect 648 599 704 619
rect 648 565 659 599
rect 693 565 704 599
rect 648 529 704 565
rect 648 495 659 529
rect 693 495 704 529
rect 648 461 704 495
rect 648 427 659 461
rect 693 427 704 461
rect 648 367 704 427
rect 734 599 790 619
rect 734 565 745 599
rect 779 565 790 599
rect 734 529 790 565
rect 734 495 745 529
rect 779 495 790 529
rect 734 457 790 495
rect 734 423 745 457
rect 779 423 790 457
rect 734 367 790 423
rect 820 531 876 619
rect 820 497 831 531
rect 865 497 876 531
rect 820 457 876 497
rect 820 423 831 457
rect 865 423 876 457
rect 820 367 876 423
rect 906 599 962 619
rect 906 565 917 599
rect 951 565 962 599
rect 906 511 962 565
rect 906 477 917 511
rect 951 477 962 511
rect 906 367 962 477
rect 992 527 1048 619
rect 992 493 1003 527
rect 1037 493 1048 527
rect 992 457 1048 493
rect 992 423 1003 457
rect 1037 423 1048 457
rect 992 367 1048 423
rect 1078 600 1188 619
rect 1078 566 1143 600
rect 1177 566 1188 600
rect 1078 367 1188 566
rect 1218 445 1274 619
rect 1218 411 1229 445
rect 1263 411 1274 445
rect 1218 367 1274 411
rect 1304 600 1406 619
rect 1304 566 1327 600
rect 1361 566 1406 600
rect 1304 367 1406 566
rect 1436 527 1512 619
rect 1436 493 1467 527
rect 1501 493 1512 527
rect 1436 459 1512 493
rect 1436 425 1467 459
rect 1501 425 1512 459
rect 1436 367 1512 425
rect 1542 597 1604 619
rect 1542 563 1562 597
rect 1596 563 1604 597
rect 1542 529 1604 563
rect 1542 495 1562 529
rect 1596 495 1604 529
rect 1542 459 1604 495
rect 1542 425 1562 459
rect 1596 425 1604 459
rect 1542 367 1604 425
<< ndiffc >>
rect 57 131 91 165
rect 57 59 91 93
rect 143 147 177 181
rect 143 67 177 101
rect 229 71 263 105
rect 315 147 349 181
rect 315 67 349 101
rect 401 71 435 105
rect 487 147 521 181
rect 487 67 521 101
rect 573 71 607 105
rect 659 169 693 203
rect 659 67 693 101
rect 745 123 779 157
rect 745 55 779 89
rect 831 169 865 203
rect 831 101 865 135
rect 926 123 960 157
rect 926 55 960 89
rect 1017 169 1051 203
rect 1017 67 1051 101
rect 1103 156 1137 190
rect 1189 59 1223 93
rect 1275 156 1309 190
rect 1349 156 1383 190
rect 1435 129 1469 163
rect 1435 57 1469 91
rect 1537 131 1571 165
rect 1537 59 1571 93
<< pdiffc >>
rect 57 565 91 599
rect 57 473 91 507
rect 57 379 91 413
rect 143 573 177 607
rect 143 502 177 536
rect 143 431 177 465
rect 229 538 263 572
rect 315 573 349 607
rect 315 470 349 504
rect 401 538 435 572
rect 487 577 521 611
rect 487 505 521 539
rect 487 431 521 465
rect 573 493 607 527
rect 573 379 607 413
rect 659 565 693 599
rect 659 495 693 529
rect 659 427 693 461
rect 745 565 779 599
rect 745 495 779 529
rect 745 423 779 457
rect 831 497 865 531
rect 831 423 865 457
rect 917 565 951 599
rect 917 477 951 511
rect 1003 493 1037 527
rect 1003 423 1037 457
rect 1143 566 1177 600
rect 1229 411 1263 445
rect 1327 566 1361 600
rect 1467 493 1501 527
rect 1467 425 1501 459
rect 1562 563 1596 597
rect 1562 495 1596 529
rect 1562 425 1596 459
<< poly >>
rect 102 619 132 645
rect 188 619 218 645
rect 274 619 304 645
rect 360 619 390 645
rect 446 619 476 645
rect 532 619 562 645
rect 618 619 648 645
rect 704 619 734 645
rect 790 619 820 645
rect 876 619 906 645
rect 962 619 992 645
rect 1048 619 1078 645
rect 1188 619 1218 645
rect 1274 619 1304 645
rect 1406 619 1436 645
rect 1512 619 1542 645
rect 102 303 132 367
rect 66 287 132 303
rect 66 253 82 287
rect 116 253 132 287
rect 66 237 132 253
rect 102 215 132 237
rect 188 335 218 367
rect 274 335 304 367
rect 360 335 390 367
rect 446 335 476 367
rect 188 319 476 335
rect 188 285 204 319
rect 238 285 272 319
rect 306 285 340 319
rect 374 285 408 319
rect 442 285 476 319
rect 188 269 476 285
rect 188 215 218 269
rect 274 215 304 269
rect 360 215 390 269
rect 446 215 476 269
rect 532 317 562 367
rect 618 317 648 367
rect 704 317 734 367
rect 532 301 734 317
rect 532 267 548 301
rect 582 267 616 301
rect 650 267 684 301
rect 718 267 734 301
rect 532 251 734 267
rect 532 215 562 251
rect 618 215 648 251
rect 704 215 734 251
rect 790 345 820 367
rect 876 345 906 367
rect 962 345 992 367
rect 790 335 992 345
rect 1048 345 1078 367
rect 1188 345 1218 367
rect 1274 345 1304 367
rect 1406 345 1436 367
rect 790 319 1006 335
rect 790 285 815 319
rect 849 285 883 319
rect 917 285 951 319
rect 985 285 1006 319
rect 790 237 1006 285
rect 1048 315 1436 345
rect 1512 321 1542 367
rect 1048 303 1424 315
rect 1048 269 1064 303
rect 1098 269 1132 303
rect 1166 269 1200 303
rect 1234 269 1268 303
rect 1302 269 1336 303
rect 1370 269 1424 303
rect 1048 253 1424 269
rect 1478 305 1544 321
rect 1478 271 1494 305
rect 1528 271 1544 305
rect 1478 255 1544 271
rect 790 215 820 237
rect 876 215 906 237
rect 976 215 1006 237
rect 1062 215 1092 253
rect 1148 215 1178 253
rect 1234 215 1264 253
rect 1394 215 1424 253
rect 1480 215 1510 255
rect 102 21 132 47
rect 188 21 218 47
rect 274 21 304 47
rect 360 21 390 47
rect 446 21 476 47
rect 532 21 562 47
rect 618 21 648 47
rect 704 21 734 47
rect 790 21 820 47
rect 876 21 906 47
rect 976 21 1006 47
rect 1062 21 1092 47
rect 1148 21 1178 47
rect 1234 21 1264 47
rect 1394 21 1424 47
rect 1480 21 1510 47
<< polycont >>
rect 82 253 116 287
rect 204 285 238 319
rect 272 285 306 319
rect 340 285 374 319
rect 408 285 442 319
rect 548 267 582 301
rect 616 267 650 301
rect 684 267 718 301
rect 815 285 849 319
rect 883 285 917 319
rect 951 285 985 319
rect 1064 269 1098 303
rect 1132 269 1166 303
rect 1200 269 1234 303
rect 1268 269 1302 303
rect 1336 269 1370 303
rect 1494 271 1528 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 41 599 93 615
rect 41 565 57 599
rect 91 565 93 599
rect 41 507 93 565
rect 41 473 57 507
rect 91 473 93 507
rect 41 413 93 473
rect 127 607 193 615
rect 127 573 143 607
rect 177 573 193 607
rect 127 536 193 573
rect 127 502 143 536
rect 177 502 193 536
rect 227 572 265 649
rect 227 538 229 572
rect 263 538 265 572
rect 227 522 265 538
rect 299 607 365 615
rect 299 573 315 607
rect 349 573 365 607
rect 127 488 193 502
rect 299 504 365 573
rect 399 572 437 649
rect 399 538 401 572
rect 435 538 437 572
rect 399 522 437 538
rect 471 611 695 615
rect 471 577 487 611
rect 521 599 695 611
rect 521 577 659 599
rect 471 539 537 577
rect 649 565 659 577
rect 693 565 695 599
rect 299 488 315 504
rect 127 470 315 488
rect 349 488 365 504
rect 471 505 487 539
rect 521 505 537 539
rect 471 488 537 505
rect 349 470 537 488
rect 127 465 537 470
rect 127 431 143 465
rect 177 454 487 465
rect 177 431 193 454
rect 471 431 487 454
rect 521 431 537 465
rect 571 527 615 543
rect 571 493 573 527
rect 607 493 615 527
rect 41 379 57 413
rect 91 397 93 413
rect 229 397 435 420
rect 571 413 615 493
rect 571 397 573 413
rect 91 386 573 397
rect 91 379 263 386
rect 41 363 263 379
rect 401 379 573 386
rect 607 379 615 413
rect 649 529 695 565
rect 649 495 659 529
rect 693 495 695 529
rect 649 461 695 495
rect 649 427 659 461
rect 693 427 695 461
rect 649 411 695 427
rect 729 599 1105 615
rect 729 565 745 599
rect 779 581 917 599
rect 779 565 795 581
rect 729 529 795 565
rect 901 565 917 581
rect 951 579 1105 599
rect 951 565 967 579
rect 729 495 745 529
rect 779 495 795 529
rect 729 457 795 495
rect 729 423 745 457
rect 779 423 795 457
rect 401 375 615 379
rect 729 407 795 423
rect 829 531 867 547
rect 829 497 831 531
rect 865 497 867 531
rect 829 457 867 497
rect 901 511 967 565
rect 901 477 917 511
rect 951 477 967 511
rect 1001 527 1037 545
rect 1001 493 1003 527
rect 829 423 831 457
rect 865 443 867 457
rect 1001 457 1037 493
rect 1071 516 1105 579
rect 1139 600 1181 649
rect 1139 566 1143 600
rect 1177 566 1181 600
rect 1139 550 1181 566
rect 1311 600 1365 649
rect 1311 566 1327 600
rect 1361 566 1365 600
rect 1311 550 1365 566
rect 1399 597 1612 613
rect 1399 579 1562 597
rect 1399 516 1433 579
rect 1560 563 1562 579
rect 1596 563 1612 597
rect 1071 482 1433 516
rect 1467 527 1526 543
rect 1501 493 1526 527
rect 1001 443 1003 457
rect 865 423 1003 443
rect 1467 459 1526 493
rect 1037 445 1467 448
rect 1037 423 1229 445
rect 829 411 1229 423
rect 1263 425 1467 445
rect 1501 425 1526 459
rect 1263 411 1526 425
rect 829 407 1526 411
rect 1560 529 1612 563
rect 1560 495 1562 529
rect 1596 495 1612 529
rect 1560 459 1612 495
rect 1560 425 1562 459
rect 1596 425 1612 459
rect 1560 409 1612 425
rect 729 375 763 407
rect 401 363 763 375
rect 1492 375 1526 407
rect 297 319 367 352
rect 573 341 763 363
rect 797 339 1456 373
rect 1492 341 1615 375
rect 797 319 1001 339
rect 66 287 132 303
rect 66 253 82 287
rect 116 253 132 287
rect 188 285 204 319
rect 238 285 272 319
rect 306 285 340 319
rect 374 285 408 319
rect 442 285 458 319
rect 66 249 132 253
rect 492 267 548 301
rect 582 267 616 301
rect 650 267 684 301
rect 718 267 734 301
rect 492 265 734 267
rect 797 285 815 319
rect 849 285 883 319
rect 917 285 951 319
rect 985 285 1001 319
rect 1422 307 1456 339
rect 1422 305 1544 307
rect 797 265 1001 285
rect 1048 303 1386 305
rect 1048 269 1064 303
rect 1098 269 1132 303
rect 1166 269 1200 303
rect 1234 269 1268 303
rect 1302 269 1336 303
rect 1370 269 1386 303
rect 1422 271 1494 305
rect 1528 271 1544 305
rect 492 249 597 265
rect 66 215 597 249
rect 1087 240 1315 269
rect 1422 267 1544 271
rect 1578 233 1615 341
rect 655 203 1053 231
rect 1349 206 1615 233
rect 655 181 659 203
rect 41 165 93 181
rect 41 131 57 165
rect 91 131 93 165
rect 41 93 93 131
rect 41 59 57 93
rect 91 59 93 93
rect 41 17 93 59
rect 127 147 143 181
rect 177 147 315 181
rect 349 147 487 181
rect 521 169 659 181
rect 693 197 831 203
rect 693 169 695 197
rect 521 147 695 169
rect 865 197 1017 203
rect 865 169 876 197
rect 127 101 179 147
rect 127 67 143 101
rect 177 67 179 101
rect 127 51 179 67
rect 213 105 279 113
rect 213 71 229 105
rect 263 71 279 105
rect 213 17 279 71
rect 313 101 351 147
rect 313 67 315 101
rect 349 67 351 101
rect 313 51 351 67
rect 385 105 451 113
rect 385 71 401 105
rect 435 71 451 105
rect 385 17 451 71
rect 485 101 523 147
rect 485 67 487 101
rect 521 67 523 101
rect 485 51 523 67
rect 557 105 623 113
rect 557 71 573 105
rect 607 71 623 105
rect 557 17 623 71
rect 657 101 695 147
rect 657 67 659 101
rect 693 67 695 101
rect 657 51 695 67
rect 729 157 795 161
rect 729 123 745 157
rect 779 123 795 157
rect 729 89 795 123
rect 729 55 745 89
rect 779 55 795 89
rect 831 135 876 169
rect 1013 169 1017 197
rect 1051 169 1053 203
rect 865 101 876 135
rect 831 85 876 101
rect 910 157 976 161
rect 910 123 926 157
rect 960 123 976 157
rect 910 89 976 123
rect 729 17 795 55
rect 910 55 926 89
rect 960 55 976 89
rect 910 17 976 55
rect 1013 106 1053 169
rect 1093 199 1615 206
rect 1093 190 1385 199
rect 1093 156 1103 190
rect 1137 156 1275 190
rect 1309 156 1349 190
rect 1383 156 1385 190
rect 1093 140 1385 156
rect 1419 163 1485 165
rect 1419 129 1435 163
rect 1469 129 1485 163
rect 1419 106 1485 129
rect 1013 101 1485 106
rect 1013 67 1017 101
rect 1051 93 1485 101
rect 1051 67 1189 93
rect 1013 59 1189 67
rect 1223 91 1485 93
rect 1223 59 1435 91
rect 1013 57 1435 59
rect 1469 57 1485 91
rect 1013 51 1485 57
rect 1521 131 1537 165
rect 1571 131 1587 165
rect 1521 93 1587 131
rect 1521 59 1537 93
rect 1571 59 1587 93
rect 1521 17 1587 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o31ai_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1471 464 1505 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 260084
string GDS_START 247222
<< end >>
