magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 3506 1975
<< nwell >>
rect -38 335 2246 704
rect -38 332 645 335
rect 1384 332 2246 335
<< pwell >>
rect 499 274 603 283
rect 383 248 603 274
rect 187 237 603 248
rect 1072 237 1342 293
rect 187 229 1342 237
rect 2010 230 2207 268
rect 1908 229 2207 230
rect 187 184 2207 229
rect 7 49 2207 184
rect 0 0 2208 49
<< scpmos >>
rect 85 508 115 592
rect 175 508 205 592
rect 276 368 306 592
rect 477 368 507 592
rect 697 508 727 592
rect 787 508 817 592
rect 865 508 895 592
rect 967 508 997 592
rect 1161 392 1191 592
rect 1347 392 1377 592
rect 1517 508 1547 592
rect 1601 508 1631 592
rect 1709 508 1739 592
rect 1799 508 1829 592
rect 1993 424 2023 592
rect 2094 368 2124 592
<< nmoslvt >>
rect 90 74 120 158
rect 168 74 198 158
rect 270 74 300 222
rect 480 100 510 248
rect 684 127 714 211
rect 820 127 850 211
rect 892 127 922 211
rect 964 127 994 211
rect 1148 119 1178 267
rect 1236 119 1266 267
rect 1520 119 1550 203
rect 1598 119 1628 203
rect 1706 119 1736 203
rect 1784 119 1814 203
rect 1991 94 2021 204
rect 2093 94 2123 242
<< ndiff >>
rect 525 248 577 257
rect 213 158 270 222
rect 33 131 90 158
rect 33 97 45 131
rect 79 97 90 131
rect 33 74 90 97
rect 120 74 168 158
rect 198 133 270 158
rect 198 99 225 133
rect 259 99 270 133
rect 198 74 270 99
rect 300 202 355 222
rect 300 168 311 202
rect 345 168 355 202
rect 300 120 355 168
rect 300 86 311 120
rect 345 86 355 120
rect 300 74 355 86
rect 409 100 480 248
rect 510 245 577 248
rect 510 211 535 245
rect 569 211 577 245
rect 1098 211 1148 267
rect 510 100 577 211
rect 631 188 684 211
rect 631 154 639 188
rect 673 154 684 188
rect 631 127 684 154
rect 714 188 820 211
rect 714 154 775 188
rect 809 154 820 188
rect 714 127 820 154
rect 850 127 892 211
rect 922 127 964 211
rect 994 127 1148 211
rect 409 77 465 100
rect 409 43 420 77
rect 454 43 465 77
rect 409 31 465 43
rect 1009 124 1148 127
rect 1009 90 1021 124
rect 1055 119 1148 124
rect 1178 244 1236 267
rect 1178 210 1189 244
rect 1223 210 1236 244
rect 1178 169 1236 210
rect 1178 135 1189 169
rect 1223 135 1236 169
rect 1178 119 1236 135
rect 1266 203 1316 267
rect 2036 210 2093 242
rect 2036 204 2048 210
rect 1266 175 1520 203
rect 1266 141 1341 175
rect 1375 141 1475 175
rect 1509 141 1520 175
rect 1266 119 1520 141
rect 1550 119 1598 203
rect 1628 165 1706 203
rect 1628 131 1650 165
rect 1684 131 1706 165
rect 1628 119 1706 131
rect 1736 119 1784 203
rect 1814 170 1871 203
rect 1814 136 1825 170
rect 1859 136 1871 170
rect 1814 119 1871 136
rect 1934 166 1991 204
rect 1934 132 1946 166
rect 1980 132 1991 166
rect 1055 90 1067 119
rect 1009 78 1067 90
rect 1934 94 1991 132
rect 2021 176 2048 204
rect 2082 176 2093 210
rect 2021 138 2093 176
rect 2021 104 2048 138
rect 2082 104 2093 138
rect 2021 94 2093 104
rect 2123 214 2181 242
rect 2123 180 2134 214
rect 2168 180 2181 214
rect 2123 138 2181 180
rect 2123 104 2134 138
rect 2168 104 2181 138
rect 2123 94 2181 104
<< pdiff >>
rect 27 567 85 592
rect 27 533 38 567
rect 72 533 85 567
rect 27 508 85 533
rect 115 567 175 592
rect 115 533 128 567
rect 162 533 175 567
rect 115 508 175 533
rect 205 572 276 592
rect 205 538 228 572
rect 262 538 276 572
rect 205 508 276 538
rect 223 368 276 508
rect 306 421 364 592
rect 306 387 319 421
rect 353 387 364 421
rect 306 368 364 387
rect 418 581 477 592
rect 418 547 430 581
rect 464 547 477 581
rect 418 368 477 547
rect 507 413 584 592
rect 638 567 697 592
rect 638 533 650 567
rect 684 533 697 567
rect 638 508 697 533
rect 727 567 787 592
rect 727 533 740 567
rect 774 533 787 567
rect 727 508 787 533
rect 817 508 865 592
rect 895 567 967 592
rect 895 533 908 567
rect 942 533 967 567
rect 895 508 967 533
rect 997 567 1052 592
rect 997 533 1010 567
rect 1044 533 1052 567
rect 997 508 1052 533
rect 1106 580 1161 592
rect 1106 546 1114 580
rect 1148 546 1161 580
rect 1106 506 1161 546
rect 507 379 536 413
rect 570 379 584 413
rect 507 368 584 379
rect 1106 472 1114 506
rect 1148 472 1161 506
rect 1106 392 1161 472
rect 1191 580 1347 592
rect 1191 546 1205 580
rect 1239 546 1299 580
rect 1333 546 1347 580
rect 1191 512 1347 546
rect 1191 478 1205 512
rect 1239 478 1299 512
rect 1333 478 1347 512
rect 1191 444 1347 478
rect 1191 410 1205 444
rect 1239 410 1299 444
rect 1333 410 1347 444
rect 1191 392 1347 410
rect 1377 557 1517 592
rect 1377 523 1390 557
rect 1424 523 1470 557
rect 1504 523 1517 557
rect 1377 508 1517 523
rect 1547 508 1601 592
rect 1631 567 1709 592
rect 1631 533 1644 567
rect 1678 533 1709 567
rect 1631 508 1709 533
rect 1739 567 1799 592
rect 1739 533 1752 567
rect 1786 533 1799 567
rect 1739 508 1799 533
rect 1829 567 1884 592
rect 1829 533 1842 567
rect 1876 533 1884 567
rect 1829 508 1884 533
rect 1938 580 1993 592
rect 1938 546 1946 580
rect 1980 546 1993 580
rect 1377 392 1430 508
rect 1938 471 1993 546
rect 1938 437 1946 471
rect 1980 437 1993 471
rect 1938 424 1993 437
rect 2023 580 2094 592
rect 2023 546 2046 580
rect 2080 546 2094 580
rect 2023 470 2094 546
rect 2023 436 2046 470
rect 2080 436 2094 470
rect 2023 424 2094 436
rect 2041 368 2094 424
rect 2124 580 2181 592
rect 2124 546 2137 580
rect 2171 546 2181 580
rect 2124 497 2181 546
rect 2124 463 2137 497
rect 2171 463 2181 497
rect 2124 414 2181 463
rect 2124 380 2137 414
rect 2171 380 2181 414
rect 2124 368 2181 380
<< ndiffc >>
rect 45 97 79 131
rect 225 99 259 133
rect 311 168 345 202
rect 311 86 345 120
rect 535 211 569 245
rect 639 154 673 188
rect 775 154 809 188
rect 420 43 454 77
rect 1021 90 1055 124
rect 1189 210 1223 244
rect 1189 135 1223 169
rect 1341 141 1375 175
rect 1475 141 1509 175
rect 1650 131 1684 165
rect 1825 136 1859 170
rect 1946 132 1980 166
rect 2048 176 2082 210
rect 2048 104 2082 138
rect 2134 180 2168 214
rect 2134 104 2168 138
<< pdiffc >>
rect 38 533 72 567
rect 128 533 162 567
rect 228 538 262 572
rect 319 387 353 421
rect 430 547 464 581
rect 650 533 684 567
rect 740 533 774 567
rect 908 533 942 567
rect 1010 533 1044 567
rect 1114 546 1148 580
rect 536 379 570 413
rect 1114 472 1148 506
rect 1205 546 1239 580
rect 1299 546 1333 580
rect 1205 478 1239 512
rect 1299 478 1333 512
rect 1205 410 1239 444
rect 1299 410 1333 444
rect 1390 523 1424 557
rect 1470 523 1504 557
rect 1644 533 1678 567
rect 1752 533 1786 567
rect 1842 533 1876 567
rect 1946 546 1980 580
rect 1946 437 1980 471
rect 2046 546 2080 580
rect 2046 436 2080 470
rect 2137 546 2171 580
rect 2137 463 2171 497
rect 2137 380 2171 414
<< poly >>
rect 85 592 115 618
rect 175 592 205 618
rect 276 592 306 618
rect 477 592 507 618
rect 697 592 727 618
rect 787 592 817 618
rect 865 592 895 618
rect 967 592 997 618
rect 1161 592 1191 618
rect 1347 592 1377 618
rect 1517 592 1547 618
rect 1601 592 1631 618
rect 1709 592 1739 618
rect 1799 592 1829 618
rect 1993 592 2023 618
rect 2094 592 2124 618
rect 85 493 115 508
rect 175 493 205 508
rect 82 414 118 493
rect 57 384 118 414
rect 57 326 87 384
rect 172 336 208 493
rect 697 493 727 508
rect 787 493 817 508
rect 865 493 895 508
rect 967 493 997 508
rect 599 463 730 493
rect 276 353 306 368
rect 477 353 507 368
rect 21 310 87 326
rect 21 276 37 310
rect 71 276 87 310
rect 21 242 87 276
rect 162 320 228 336
rect 162 286 178 320
rect 212 286 228 320
rect 273 310 309 353
rect 474 336 510 353
rect 383 320 510 336
rect 162 270 228 286
rect 270 294 341 310
rect 21 208 37 242
rect 71 222 87 242
rect 71 208 120 222
rect 21 192 120 208
rect 90 158 120 192
rect 168 158 198 270
rect 270 260 291 294
rect 325 260 341 294
rect 383 286 399 320
rect 433 309 510 320
rect 599 309 629 463
rect 784 421 820 493
rect 677 418 820 421
rect 677 405 814 418
rect 677 371 693 405
rect 727 385 814 405
rect 727 371 743 385
rect 677 355 743 371
rect 862 370 898 493
rect 856 354 922 370
rect 856 320 872 354
rect 906 320 922 354
rect 433 286 792 309
rect 856 304 922 320
rect 383 279 792 286
rect 383 270 510 279
rect 270 244 341 260
rect 480 248 510 270
rect 270 222 300 244
rect 762 256 792 279
rect 684 211 714 237
rect 762 226 850 256
rect 820 211 850 226
rect 892 211 922 304
rect 964 360 1000 493
rect 1517 493 1547 508
rect 1601 493 1631 508
rect 1709 493 1739 508
rect 1799 493 1829 508
rect 1514 473 1547 493
rect 1462 457 1544 473
rect 1462 423 1478 457
rect 1512 423 1544 457
rect 1161 377 1191 392
rect 1347 377 1377 392
rect 1462 389 1544 423
rect 1158 360 1194 377
rect 964 344 1030 360
rect 964 310 980 344
rect 1014 310 1030 344
rect 964 294 1030 310
rect 1073 344 1194 360
rect 1073 310 1089 344
rect 1123 310 1194 344
rect 1073 294 1194 310
rect 1236 344 1302 360
rect 1236 310 1252 344
rect 1286 310 1302 344
rect 1236 294 1302 310
rect 964 211 994 294
rect 1148 267 1178 294
rect 1236 267 1266 294
rect 1344 291 1380 377
rect 1462 355 1478 389
rect 1512 355 1544 389
rect 1462 339 1544 355
rect 1598 467 1634 493
rect 1598 451 1664 467
rect 1598 417 1614 451
rect 1648 417 1664 451
rect 1598 401 1664 417
rect 1344 275 1484 291
rect 684 105 714 127
rect 90 48 120 74
rect 168 48 198 74
rect 270 48 300 74
rect 480 74 510 100
rect 607 89 741 105
rect 607 55 623 89
rect 657 55 691 89
rect 725 55 741 89
rect 607 39 741 55
rect 820 51 850 127
rect 892 101 922 127
rect 964 101 994 127
rect 1344 261 1366 275
rect 1350 241 1366 261
rect 1400 241 1434 275
rect 1468 255 1484 275
rect 1468 241 1550 255
rect 1350 225 1550 241
rect 1520 203 1550 225
rect 1598 203 1628 401
rect 1706 359 1742 493
rect 1796 409 1832 493
rect 1993 409 2023 424
rect 1796 379 2026 409
rect 1796 359 1850 379
rect 1676 343 1742 359
rect 1676 309 1692 343
rect 1726 309 1742 343
rect 1676 293 1742 309
rect 1784 343 1850 359
rect 2094 353 2124 368
rect 1784 309 1800 343
rect 1834 309 1850 343
rect 2091 330 2127 353
rect 1706 203 1736 293
rect 1784 275 1850 309
rect 1784 241 1800 275
rect 1834 255 1850 275
rect 2063 314 2129 330
rect 2063 280 2079 314
rect 2113 280 2129 314
rect 2063 264 2129 280
rect 1834 241 2021 255
rect 2093 242 2123 264
rect 1784 225 2021 241
rect 1784 203 1814 225
rect 1991 204 2021 225
rect 1148 93 1178 119
rect 1236 51 1266 119
rect 1520 93 1550 119
rect 1598 93 1628 119
rect 1706 93 1736 119
rect 1784 93 1814 119
rect 1991 68 2021 94
rect 2093 68 2123 94
rect 820 21 1266 51
<< polycont >>
rect 37 276 71 310
rect 178 286 212 320
rect 37 208 71 242
rect 291 260 325 294
rect 399 286 433 320
rect 693 371 727 405
rect 872 320 906 354
rect 1478 423 1512 457
rect 980 310 1014 344
rect 1089 310 1123 344
rect 1252 310 1286 344
rect 1478 355 1512 389
rect 1614 417 1648 451
rect 623 55 657 89
rect 691 55 725 89
rect 1366 241 1400 275
rect 1434 241 1468 275
rect 1692 309 1726 343
rect 1800 309 1834 343
rect 1800 241 1834 275
rect 2079 280 2113 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 22 567 88 649
rect 22 533 38 567
rect 72 533 88 567
rect 22 504 88 533
rect 128 567 178 596
rect 162 533 178 567
rect 128 470 178 533
rect 212 572 278 649
rect 212 538 228 572
rect 262 538 278 572
rect 212 531 278 538
rect 414 581 480 649
rect 414 547 430 581
rect 464 547 480 581
rect 414 531 480 547
rect 634 567 684 596
rect 634 533 650 567
rect 634 497 684 533
rect 724 567 811 596
rect 724 533 740 567
rect 774 533 811 567
rect 724 504 811 533
rect 892 567 958 649
rect 892 533 908 567
rect 942 533 958 567
rect 892 504 958 533
rect 994 567 1060 596
rect 994 533 1010 567
rect 1044 533 1060 567
rect 212 470 684 497
rect 108 463 684 470
rect 108 436 246 463
rect 21 310 74 430
rect 21 276 37 310
rect 71 276 74 310
rect 21 242 74 276
rect 21 208 37 242
rect 71 208 74 242
rect 21 192 74 208
rect 108 158 142 436
rect 303 421 433 429
rect 303 387 319 421
rect 353 387 433 421
rect 303 364 433 387
rect 176 350 257 356
rect 176 320 223 350
rect 176 286 178 320
rect 212 316 223 320
rect 212 286 257 316
rect 387 320 433 364
rect 176 270 257 286
rect 291 294 353 310
rect 325 260 353 294
rect 291 236 353 260
rect 387 286 399 320
rect 387 202 433 286
rect 295 168 311 202
rect 345 168 433 202
rect 29 131 142 158
rect 29 97 45 131
rect 79 97 142 131
rect 29 70 142 97
rect 209 133 259 162
rect 209 99 225 133
rect 209 17 259 99
rect 295 127 433 168
rect 467 161 501 463
rect 777 438 811 504
rect 994 438 1060 533
rect 1098 580 1164 649
rect 1098 546 1114 580
rect 1148 546 1164 580
rect 1098 506 1164 546
rect 1098 472 1114 506
rect 1148 472 1164 506
rect 1198 580 1340 596
rect 1198 546 1205 580
rect 1239 546 1299 580
rect 1333 546 1340 580
rect 1198 512 1340 546
rect 1198 478 1205 512
rect 1239 478 1299 512
rect 1333 478 1340 512
rect 1374 557 1520 573
rect 1374 523 1390 557
rect 1424 523 1470 557
rect 1504 541 1520 557
rect 1628 567 1694 649
rect 1504 523 1580 541
rect 1374 507 1580 523
rect 1198 444 1340 478
rect 535 421 588 429
rect 535 413 743 421
rect 535 379 536 413
rect 570 405 743 413
rect 570 379 693 405
rect 535 371 693 379
rect 727 371 743 405
rect 535 355 743 371
rect 777 404 1139 438
rect 1198 428 1205 444
rect 535 283 588 355
rect 535 249 741 283
rect 535 245 588 249
rect 569 211 588 245
rect 535 195 588 211
rect 623 188 673 215
rect 623 161 639 188
rect 467 154 639 161
rect 467 127 673 154
rect 295 120 361 127
rect 295 86 311 120
rect 345 86 361 120
rect 707 93 741 249
rect 777 215 811 404
rect 856 354 922 370
rect 856 320 872 354
rect 906 320 922 354
rect 856 304 922 320
rect 888 260 922 304
rect 964 350 1031 360
rect 964 344 991 350
rect 964 310 980 344
rect 1025 316 1031 350
rect 1014 310 1031 316
rect 964 294 1031 310
rect 1073 344 1139 404
rect 1073 310 1089 344
rect 1123 310 1139 344
rect 1073 294 1139 310
rect 1173 410 1205 428
rect 1239 410 1299 444
rect 1333 410 1340 444
rect 1173 394 1340 410
rect 1462 457 1512 473
rect 1462 423 1478 457
rect 1173 260 1207 394
rect 1462 389 1512 423
rect 1462 360 1478 389
rect 1241 355 1478 360
rect 1241 344 1512 355
rect 1241 310 1252 344
rect 1286 326 1512 344
rect 1286 310 1302 326
rect 1241 294 1302 310
rect 1350 275 1484 291
rect 888 244 1239 260
rect 1350 259 1366 275
rect 888 226 1189 244
rect 775 188 825 215
rect 1173 210 1189 226
rect 1223 210 1239 244
rect 809 154 825 188
rect 775 127 825 154
rect 859 158 1139 192
rect 859 93 893 158
rect 295 70 361 86
rect 404 77 470 93
rect 404 43 420 77
rect 454 43 470 77
rect 607 89 893 93
rect 607 55 623 89
rect 657 55 691 89
rect 725 55 893 89
rect 607 51 893 55
rect 1005 90 1021 124
rect 1055 90 1071 124
rect 404 17 470 43
rect 1005 17 1071 90
rect 1105 85 1139 158
rect 1173 169 1239 210
rect 1173 135 1189 169
rect 1223 135 1239 169
rect 1173 119 1239 135
rect 1273 241 1366 259
rect 1400 241 1434 275
rect 1468 241 1484 275
rect 1273 225 1484 241
rect 1546 259 1580 507
rect 1628 533 1644 567
rect 1678 533 1694 567
rect 1628 504 1694 533
rect 1736 567 1802 596
rect 1736 533 1752 567
rect 1786 533 1802 567
rect 1736 467 1802 533
rect 1842 567 1892 649
rect 1876 533 1892 567
rect 1842 504 1892 533
rect 1930 580 1996 596
rect 1930 546 1946 580
rect 1980 546 1996 580
rect 1930 471 1996 546
rect 1614 451 1810 467
rect 1930 461 1946 471
rect 1648 427 1810 451
rect 1980 437 1996 471
rect 1648 417 1912 427
rect 1614 393 1912 417
rect 1657 350 1742 359
rect 1657 316 1663 350
rect 1697 343 1742 350
rect 1657 309 1692 316
rect 1726 309 1742 343
rect 1657 293 1742 309
rect 1784 343 1844 359
rect 1784 309 1800 343
rect 1834 309 1844 343
rect 1784 275 1844 309
rect 1784 259 1800 275
rect 1546 241 1800 259
rect 1834 241 1844 275
rect 1546 225 1844 241
rect 1273 85 1307 225
rect 1546 191 1580 225
rect 1878 191 1912 393
rect 1341 175 1580 191
rect 1375 141 1475 175
rect 1509 141 1580 175
rect 1341 125 1580 141
rect 1623 165 1711 181
rect 1623 131 1650 165
rect 1684 131 1711 165
rect 1105 51 1307 85
rect 1623 17 1711 131
rect 1809 170 1912 191
rect 1809 136 1825 170
rect 1859 136 1912 170
rect 1809 115 1912 136
rect 1946 330 1996 437
rect 2030 580 2080 649
rect 2030 546 2046 580
rect 2030 470 2080 546
rect 2030 436 2046 470
rect 2030 420 2080 436
rect 2121 580 2191 596
rect 2121 546 2137 580
rect 2171 546 2191 580
rect 2121 497 2191 546
rect 2121 463 2137 497
rect 2171 463 2191 497
rect 2121 414 2191 463
rect 2121 380 2137 414
rect 2171 380 2191 414
rect 2121 364 2191 380
rect 1946 314 2123 330
rect 1946 280 2079 314
rect 2113 280 2123 314
rect 1946 264 2123 280
rect 1946 166 1996 264
rect 2157 230 2191 364
rect 1980 132 1996 166
rect 1946 106 1996 132
rect 2032 210 2082 226
rect 2032 176 2048 210
rect 2032 138 2082 176
rect 2032 104 2048 138
rect 2032 17 2082 104
rect 2118 214 2191 230
rect 2118 180 2134 214
rect 2168 180 2191 214
rect 2118 138 2191 180
rect 2118 104 2134 138
rect 2168 104 2191 138
rect 2118 88 2191 104
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 223 316 257 350
rect 991 344 1025 350
rect 991 316 1014 344
rect 1014 316 1025 344
rect 1663 343 1697 350
rect 1663 316 1692 343
rect 1692 316 1697 343
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 211 350 269 356
rect 211 316 223 350
rect 257 347 269 350
rect 979 350 1037 356
rect 979 347 991 350
rect 257 319 991 347
rect 257 316 269 319
rect 211 310 269 316
rect 979 316 991 319
rect 1025 347 1037 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1025 319 1663 347
rect 1025 316 1037 319
rect 979 310 1037 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfrtn_1
flabel comment s 983 39 983 39 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 223 316 257 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 2143 390 2177 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2143 464 2177 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2143 538 2177 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y R90
string GDS_END 3437588
string GDS_START 3420864
<< end >>
