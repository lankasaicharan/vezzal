magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3890 1975
<< nwell >>
rect -38 331 2630 704
rect 313 311 1196 331
rect 313 287 654 311
rect 960 305 1196 311
<< pwell >>
rect 1346 263 1541 281
rect 1206 235 1541 263
rect 920 229 1541 235
rect 444 195 1541 229
rect 12 167 1541 195
rect 1898 167 2322 237
rect 12 49 2591 167
rect 0 0 2592 49
<< scnmos >>
rect 95 85 125 169
rect 167 85 197 169
rect 267 85 297 169
rect 339 85 369 169
rect 425 85 455 169
rect 543 119 573 203
rect 615 119 645 203
rect 733 119 763 203
rect 805 119 835 203
rect 1019 125 1049 209
rect 1091 125 1121 209
rect 1309 153 1339 237
rect 1429 171 1459 255
rect 1626 57 1656 141
rect 1712 57 1742 141
rect 1784 57 1814 141
rect 1980 127 2010 211
rect 2052 127 2082 211
rect 2138 127 2168 211
rect 2210 127 2240 211
rect 2406 57 2436 141
rect 2478 57 2508 141
<< scpmoshvt >>
rect 83 403 133 603
rect 189 403 239 603
rect 405 323 455 523
rect 511 323 561 523
rect 728 347 778 547
rect 834 347 884 547
rect 1053 341 1103 541
rect 1289 419 1339 619
rect 1395 419 1445 619
rect 1507 419 1557 619
rect 1673 419 1723 619
rect 1906 367 1956 567
rect 2012 367 2062 567
rect 2458 409 2508 609
<< ndiff >>
rect 1372 243 1429 255
rect 1372 237 1384 243
rect 470 169 543 203
rect 38 144 95 169
rect 38 110 50 144
rect 84 110 95 144
rect 38 85 95 110
rect 125 85 167 169
rect 197 144 267 169
rect 197 110 222 144
rect 256 110 267 144
rect 197 85 267 110
rect 297 85 339 169
rect 369 144 425 169
rect 369 110 380 144
rect 414 110 425 144
rect 369 85 425 110
rect 455 161 543 169
rect 455 127 482 161
rect 516 127 543 161
rect 455 119 543 127
rect 573 119 615 203
rect 645 141 733 203
rect 645 119 672 141
rect 455 85 528 119
rect 660 107 672 119
rect 706 119 733 141
rect 763 119 805 203
rect 835 178 892 203
rect 835 144 846 178
rect 880 144 892 178
rect 835 119 892 144
rect 946 157 1019 209
rect 946 123 958 157
rect 992 125 1019 157
rect 1049 125 1091 209
rect 1121 184 1178 209
rect 1121 150 1132 184
rect 1166 150 1178 184
rect 1232 207 1309 237
rect 1232 173 1244 207
rect 1278 173 1309 207
rect 1232 153 1309 173
rect 1339 209 1384 237
rect 1418 209 1429 243
rect 1339 171 1429 209
rect 1459 217 1515 255
rect 1459 183 1470 217
rect 1504 183 1515 217
rect 1459 171 1515 183
rect 1339 153 1389 171
rect 1121 125 1178 150
rect 992 123 1004 125
rect 706 107 718 119
rect 660 95 718 107
rect 946 111 1004 123
rect 1924 186 1980 211
rect 1924 152 1935 186
rect 1969 152 1980 186
rect 1569 116 1626 141
rect 1569 82 1581 116
rect 1615 82 1626 116
rect 1569 57 1626 82
rect 1656 116 1712 141
rect 1656 82 1667 116
rect 1701 82 1712 116
rect 1656 57 1712 82
rect 1742 57 1784 141
rect 1814 116 1870 141
rect 1924 127 1980 152
rect 2010 127 2052 211
rect 2082 186 2138 211
rect 2082 152 2093 186
rect 2127 152 2138 186
rect 2082 127 2138 152
rect 2168 127 2210 211
rect 2240 186 2296 211
rect 2240 152 2251 186
rect 2285 152 2296 186
rect 2240 127 2296 152
rect 1814 82 1825 116
rect 1859 82 1870 116
rect 2350 116 2406 141
rect 1814 57 1870 82
rect 2350 82 2361 116
rect 2395 82 2406 116
rect 2350 57 2406 82
rect 2436 57 2478 141
rect 2508 116 2565 141
rect 2508 82 2519 116
rect 2553 82 2565 116
rect 2508 57 2565 82
<< pdiff >>
rect 27 591 83 603
rect 27 557 38 591
rect 72 557 83 591
rect 27 520 83 557
rect 27 486 38 520
rect 72 486 83 520
rect 27 449 83 486
rect 27 415 38 449
rect 72 415 83 449
rect 27 403 83 415
rect 133 590 189 603
rect 133 556 144 590
rect 178 556 189 590
rect 133 403 189 556
rect 239 449 295 603
rect 672 535 728 547
rect 239 415 250 449
rect 284 415 295 449
rect 239 403 295 415
rect 349 511 405 523
rect 349 477 360 511
rect 394 477 405 511
rect 349 323 405 477
rect 455 370 511 523
rect 455 336 466 370
rect 500 336 511 370
rect 455 323 511 336
rect 561 432 618 523
rect 561 398 572 432
rect 606 398 618 432
rect 561 323 618 398
rect 672 501 683 535
rect 717 501 728 535
rect 672 447 728 501
rect 672 413 683 447
rect 717 413 728 447
rect 672 347 728 413
rect 778 535 834 547
rect 778 501 789 535
rect 823 501 834 535
rect 778 447 834 501
rect 778 413 789 447
rect 823 413 834 447
rect 778 347 834 413
rect 884 535 941 547
rect 884 501 895 535
rect 929 501 941 535
rect 884 401 941 501
rect 884 367 895 401
rect 929 367 941 401
rect 884 347 941 367
rect 996 387 1053 541
rect 996 353 1008 387
rect 1042 353 1053 387
rect 996 341 1053 353
rect 1103 528 1160 541
rect 1103 494 1114 528
rect 1148 494 1160 528
rect 1103 341 1160 494
rect 1232 597 1289 619
rect 1232 563 1244 597
rect 1278 563 1289 597
rect 1232 465 1289 563
rect 1232 431 1244 465
rect 1278 431 1289 465
rect 1232 419 1289 431
rect 1339 597 1395 619
rect 1339 563 1350 597
rect 1384 563 1395 597
rect 1339 473 1395 563
rect 1339 439 1350 473
rect 1384 439 1395 473
rect 1339 419 1395 439
rect 1445 419 1507 619
rect 1557 607 1673 619
rect 1557 573 1575 607
rect 1609 573 1673 607
rect 1557 524 1673 573
rect 1557 490 1575 524
rect 1609 490 1673 524
rect 1557 419 1673 490
rect 1723 597 1780 619
rect 1723 563 1734 597
rect 1768 563 1780 597
rect 2401 597 2458 609
rect 1723 465 1780 563
rect 1723 431 1734 465
rect 1768 431 1780 465
rect 1723 419 1780 431
rect 1849 555 1906 567
rect 1849 521 1861 555
rect 1895 521 1906 555
rect 1849 484 1906 521
rect 1849 450 1861 484
rect 1895 450 1906 484
rect 1849 413 1906 450
rect 1849 379 1861 413
rect 1895 379 1906 413
rect 1849 367 1906 379
rect 1956 555 2012 567
rect 1956 521 1967 555
rect 2001 521 2012 555
rect 1956 484 2012 521
rect 1956 450 1967 484
rect 2001 450 2012 484
rect 1956 413 2012 450
rect 1956 379 1967 413
rect 2001 379 2012 413
rect 1956 367 2012 379
rect 2062 555 2119 567
rect 2062 521 2073 555
rect 2107 521 2119 555
rect 2062 484 2119 521
rect 2062 450 2073 484
rect 2107 450 2119 484
rect 2062 413 2119 450
rect 2062 379 2073 413
rect 2107 379 2119 413
rect 2401 563 2413 597
rect 2447 563 2458 597
rect 2401 473 2458 563
rect 2401 439 2413 473
rect 2447 439 2458 473
rect 2401 409 2458 439
rect 2508 597 2565 609
rect 2508 563 2519 597
rect 2553 563 2565 597
rect 2508 526 2565 563
rect 2508 492 2519 526
rect 2553 492 2565 526
rect 2508 455 2565 492
rect 2508 421 2519 455
rect 2553 421 2565 455
rect 2508 409 2565 421
rect 2062 367 2119 379
<< ndiffc >>
rect 50 110 84 144
rect 222 110 256 144
rect 380 110 414 144
rect 482 127 516 161
rect 672 107 706 141
rect 846 144 880 178
rect 958 123 992 157
rect 1132 150 1166 184
rect 1244 173 1278 207
rect 1384 209 1418 243
rect 1470 183 1504 217
rect 1935 152 1969 186
rect 1581 82 1615 116
rect 1667 82 1701 116
rect 2093 152 2127 186
rect 2251 152 2285 186
rect 1825 82 1859 116
rect 2361 82 2395 116
rect 2519 82 2553 116
<< pdiffc >>
rect 38 557 72 591
rect 38 486 72 520
rect 38 415 72 449
rect 144 556 178 590
rect 250 415 284 449
rect 360 477 394 511
rect 466 336 500 370
rect 572 398 606 432
rect 683 501 717 535
rect 683 413 717 447
rect 789 501 823 535
rect 789 413 823 447
rect 895 501 929 535
rect 895 367 929 401
rect 1008 353 1042 387
rect 1114 494 1148 528
rect 1244 563 1278 597
rect 1244 431 1278 465
rect 1350 563 1384 597
rect 1350 439 1384 473
rect 1575 573 1609 607
rect 1575 490 1609 524
rect 1734 563 1768 597
rect 1734 431 1768 465
rect 1861 521 1895 555
rect 1861 450 1895 484
rect 1861 379 1895 413
rect 1967 521 2001 555
rect 1967 450 2001 484
rect 1967 379 2001 413
rect 2073 521 2107 555
rect 2073 450 2107 484
rect 2073 379 2107 413
rect 2413 563 2447 597
rect 2413 439 2447 473
rect 2519 563 2553 597
rect 2519 492 2553 526
rect 2519 421 2553 455
<< poly >>
rect 83 603 133 629
rect 189 603 239 629
rect 397 615 1205 645
rect 1289 619 1339 645
rect 1395 619 1445 645
rect 1507 619 1557 645
rect 1673 619 1723 645
rect 397 605 463 615
rect 397 571 413 605
rect 447 571 463 605
rect 397 555 463 571
rect 405 523 455 555
rect 511 523 561 549
rect 728 547 778 573
rect 834 547 884 573
rect 83 257 133 403
rect 189 371 239 403
rect 189 355 297 371
rect 189 321 213 355
rect 247 321 297 355
rect 1053 541 1103 567
rect 728 332 778 347
rect 189 305 297 321
rect 95 241 197 257
rect 95 207 136 241
rect 170 207 197 241
rect 95 191 197 207
rect 95 169 125 191
rect 167 169 197 191
rect 267 249 297 305
rect 405 297 455 323
rect 267 219 369 249
rect 267 169 297 219
rect 339 169 369 219
rect 425 169 455 297
rect 511 248 561 323
rect 651 302 778 332
rect 834 315 884 347
rect 1053 326 1103 341
rect 1175 326 1205 615
rect 2458 609 2508 635
rect 1906 567 1956 593
rect 2012 567 2062 593
rect 1289 326 1339 419
rect 1395 387 1445 419
rect 1507 387 1557 419
rect 651 291 681 302
rect 615 275 681 291
rect 511 218 573 248
rect 543 203 573 218
rect 615 241 631 275
rect 665 241 681 275
rect 820 299 886 315
rect 820 265 836 299
rect 870 265 886 299
rect 1053 296 1339 326
rect 1387 371 1459 387
rect 1387 337 1403 371
rect 1437 337 1459 371
rect 1387 321 1459 337
rect 1507 371 1625 387
rect 1507 337 1575 371
rect 1609 337 1625 371
rect 1507 321 1625 337
rect 820 254 886 265
rect 1091 254 1121 296
rect 615 225 681 241
rect 615 203 645 225
rect 733 224 886 254
rect 1019 224 1121 254
rect 1309 237 1339 296
rect 1429 255 1459 321
rect 733 203 763 224
rect 805 203 835 224
rect 1019 209 1049 224
rect 1091 209 1121 224
rect 95 59 125 85
rect 167 59 197 85
rect 267 59 297 85
rect 339 59 369 85
rect 425 59 455 85
rect 543 51 573 119
rect 615 93 645 119
rect 1595 186 1625 321
rect 1673 368 1723 419
rect 1673 352 1742 368
rect 2458 377 2508 409
rect 1673 318 1689 352
rect 1723 318 1742 352
rect 1673 284 1742 318
rect 1673 250 1689 284
rect 1723 264 1742 284
rect 1906 317 1956 367
rect 2012 317 2062 367
rect 2401 361 2488 377
rect 2401 327 2417 361
rect 2451 327 2488 361
rect 1906 301 2353 317
rect 1906 267 1963 301
rect 1997 267 2031 301
rect 2065 267 2099 301
rect 2133 267 2167 301
rect 2201 267 2235 301
rect 2269 267 2303 301
rect 2337 267 2353 301
rect 1723 250 1814 264
rect 1906 251 2353 267
rect 2401 293 2488 327
rect 2401 259 2417 293
rect 2451 273 2488 293
rect 2451 259 2508 273
rect 1673 234 1814 250
rect 1309 127 1339 153
rect 733 93 763 119
rect 805 93 835 119
rect 1019 99 1049 125
rect 1091 99 1121 125
rect 1429 51 1459 171
rect 1595 156 1656 186
rect 1626 141 1656 156
rect 1712 141 1742 234
rect 1784 141 1814 234
rect 1980 211 2010 251
rect 2052 211 2082 251
rect 2138 211 2168 251
rect 2210 211 2240 251
rect 2401 243 2508 259
rect 2406 141 2436 243
rect 2478 141 2508 243
rect 1980 101 2010 127
rect 2052 101 2082 127
rect 2138 101 2168 127
rect 2210 101 2240 127
rect 543 21 1459 51
rect 1626 31 1656 57
rect 1712 31 1742 57
rect 1784 31 1814 57
rect 2406 31 2436 57
rect 2478 31 2508 57
<< polycont >>
rect 413 571 447 605
rect 213 321 247 355
rect 136 207 170 241
rect 631 241 665 275
rect 836 265 870 299
rect 1403 337 1437 371
rect 1575 337 1609 371
rect 1689 318 1723 352
rect 1689 250 1723 284
rect 2417 327 2451 361
rect 1963 267 1997 301
rect 2031 267 2065 301
rect 2099 267 2133 301
rect 2167 267 2201 301
rect 2235 267 2269 301
rect 2303 267 2337 301
rect 2417 259 2451 293
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 22 591 88 607
rect 22 557 38 591
rect 72 557 88 591
rect 22 520 88 557
rect 128 590 194 649
rect 128 556 144 590
rect 178 556 194 590
rect 128 555 194 556
rect 230 605 463 613
rect 230 571 413 605
rect 447 571 463 605
rect 230 555 463 571
rect 22 486 38 520
rect 72 519 88 520
rect 230 519 264 555
rect 667 535 733 551
rect 667 519 683 535
rect 72 486 264 519
rect 22 485 264 486
rect 344 511 683 519
rect 22 449 88 485
rect 344 477 360 511
rect 394 501 683 511
rect 717 501 733 535
rect 394 485 733 501
rect 394 477 410 485
rect 22 415 38 449
rect 72 415 88 449
rect 22 399 88 415
rect 234 415 250 449
rect 284 441 300 449
rect 556 441 622 449
rect 284 432 622 441
rect 284 415 572 432
rect 234 407 572 415
rect 22 144 84 399
rect 197 355 263 371
rect 197 321 213 355
rect 247 321 263 355
rect 197 305 263 321
rect 22 110 50 144
rect 22 81 84 110
rect 120 241 186 257
rect 120 207 136 241
rect 170 207 186 241
rect 120 88 186 207
rect 364 173 398 407
rect 556 398 572 407
rect 606 398 622 432
rect 556 397 622 398
rect 667 447 733 485
rect 667 413 683 447
rect 717 413 733 447
rect 667 397 733 413
rect 773 535 839 649
rect 773 501 789 535
rect 823 501 839 535
rect 773 447 839 501
rect 773 413 789 447
rect 823 413 839 447
rect 773 397 839 413
rect 879 535 956 551
rect 879 501 895 535
rect 929 501 956 535
rect 879 457 956 501
rect 1098 528 1164 649
rect 1098 494 1114 528
rect 1148 494 1164 528
rect 1098 493 1164 494
rect 1228 597 1294 613
rect 1228 563 1244 597
rect 1278 563 1294 597
rect 1228 465 1294 563
rect 1228 457 1244 465
rect 879 431 1244 457
rect 1278 431 1294 465
rect 879 423 1294 431
rect 1334 597 1400 613
rect 1334 563 1350 597
rect 1384 563 1400 597
rect 1334 473 1400 563
rect 1559 607 1625 649
rect 1559 573 1575 607
rect 1609 573 1625 607
rect 1559 524 1625 573
rect 1559 490 1575 524
rect 1609 490 1625 524
rect 1559 474 1625 490
rect 1718 597 1809 613
rect 1718 563 1734 597
rect 1768 563 1809 597
rect 1334 439 1350 473
rect 1384 457 1400 473
rect 1718 465 1809 563
rect 1384 439 1523 457
rect 1334 423 1523 439
rect 1718 438 1734 465
rect 879 401 956 423
rect 1228 415 1294 423
rect 450 370 516 371
rect 450 336 466 370
rect 500 361 516 370
rect 879 367 895 401
rect 929 367 956 401
rect 500 336 843 361
rect 879 351 956 367
rect 450 327 843 336
rect 450 319 532 327
rect 222 144 272 173
rect 256 110 272 144
rect 222 17 272 110
rect 364 144 430 173
rect 364 110 380 144
rect 414 110 430 144
rect 364 81 430 110
rect 466 161 532 319
rect 809 315 843 327
rect 809 299 886 315
rect 615 275 681 291
rect 615 241 631 275
rect 665 241 681 275
rect 809 265 836 299
rect 870 265 886 299
rect 809 263 886 265
rect 615 227 681 241
rect 922 227 956 351
rect 615 193 956 227
rect 992 353 1008 387
rect 1042 371 1058 387
rect 1387 371 1453 387
rect 1042 353 1403 371
rect 992 337 1403 353
rect 1437 337 1453 371
rect 466 127 482 161
rect 516 127 532 161
rect 830 178 896 193
rect 466 81 532 127
rect 656 141 722 157
rect 656 107 672 141
rect 706 107 722 141
rect 656 17 722 107
rect 830 144 846 178
rect 880 144 896 178
rect 830 87 896 144
rect 942 123 958 157
rect 992 123 1026 337
rect 1387 323 1453 337
rect 1062 267 1348 301
rect 1489 287 1523 423
rect 1559 431 1734 438
rect 1768 431 1809 465
rect 1559 404 1809 431
rect 1559 371 1625 404
rect 1559 337 1575 371
rect 1609 337 1625 371
rect 1559 323 1625 337
rect 1673 352 1739 368
rect 1673 318 1689 352
rect 1723 318 1739 352
rect 1673 287 1739 318
rect 1062 87 1096 267
rect 830 53 1096 87
rect 1132 184 1182 213
rect 1166 150 1182 184
rect 1132 17 1182 150
rect 1228 207 1278 231
rect 1228 173 1244 207
rect 1228 87 1278 173
rect 1314 157 1348 267
rect 1384 284 1739 287
rect 1384 253 1689 284
rect 1384 243 1418 253
rect 1673 250 1689 253
rect 1723 250 1739 284
rect 1673 234 1739 250
rect 1384 193 1418 209
rect 1454 183 1470 217
rect 1504 183 1520 217
rect 1454 157 1520 183
rect 1314 123 1520 157
rect 1775 145 1809 404
rect 1845 555 1911 578
rect 1845 521 1861 555
rect 1895 521 1911 555
rect 1845 484 1911 521
rect 1845 450 1861 484
rect 1895 450 1911 484
rect 1845 413 1911 450
rect 1845 379 1861 413
rect 1895 379 1911 413
rect 1845 215 1911 379
rect 1951 555 2017 649
rect 2397 597 2463 649
rect 1951 521 1967 555
rect 2001 521 2017 555
rect 1951 484 2017 521
rect 1951 450 1967 484
rect 2001 450 2017 484
rect 1951 413 2017 450
rect 1951 379 1967 413
rect 2001 379 2017 413
rect 1951 363 2017 379
rect 2057 555 2123 571
rect 2057 521 2073 555
rect 2107 521 2123 555
rect 2057 484 2123 521
rect 2057 450 2073 484
rect 2107 450 2123 484
rect 2057 413 2123 450
rect 2397 563 2413 597
rect 2447 563 2463 597
rect 2397 473 2463 563
rect 2397 439 2413 473
rect 2447 439 2463 473
rect 2397 423 2463 439
rect 2503 597 2569 613
rect 2503 563 2519 597
rect 2553 563 2569 597
rect 2503 526 2569 563
rect 2503 492 2519 526
rect 2553 492 2569 526
rect 2503 455 2569 492
rect 2057 379 2073 413
rect 2107 387 2123 413
rect 2503 421 2519 455
rect 2553 421 2569 455
rect 2107 379 2467 387
rect 2057 361 2467 379
rect 2057 353 2417 361
rect 2401 327 2417 353
rect 2451 327 2467 361
rect 1947 301 2353 317
rect 1947 267 1963 301
rect 1997 267 2031 301
rect 2065 267 2099 301
rect 2133 267 2167 301
rect 2201 267 2235 301
rect 2269 267 2303 301
rect 2337 267 2353 301
rect 1947 251 2353 267
rect 2401 293 2467 327
rect 2401 259 2417 293
rect 2451 259 2467 293
rect 1845 186 1985 215
rect 1845 181 1935 186
rect 1919 152 1935 181
rect 1969 152 1985 186
rect 1565 116 1631 145
rect 1565 87 1581 116
rect 1228 82 1581 87
rect 1615 82 1631 116
rect 1228 53 1631 82
rect 1667 116 1717 145
rect 1701 82 1717 116
rect 1667 17 1717 82
rect 1775 116 1875 145
rect 1919 123 1985 152
rect 1775 82 1825 116
rect 1859 87 1875 116
rect 2021 87 2055 251
rect 2401 243 2467 259
rect 2401 215 2435 243
rect 1859 82 2055 87
rect 1775 53 2055 82
rect 2093 186 2143 215
rect 2127 152 2143 186
rect 2093 17 2143 152
rect 2235 186 2435 215
rect 2235 152 2251 186
rect 2285 181 2435 186
rect 2285 152 2301 181
rect 2235 123 2301 152
rect 2345 116 2411 145
rect 2345 82 2361 116
rect 2395 82 2411 116
rect 2345 17 2411 82
rect 2503 116 2569 421
rect 2503 82 2519 116
rect 2553 82 2569 116
rect 2503 53 2569 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
flabel pwell s 0 0 2592 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 2592 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfxbp_lp
flabel metal1 s 0 617 2592 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 2592 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1855 390 1889 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1855 464 1889 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1855 538 1889 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2527 94 2561 128 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2527 168 2561 202 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2527 242 2561 276 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2527 316 2561 350 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2527 390 2561 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2527 464 2561 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2527 538 2561 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2592 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2524446
string GDS_START 2507084
<< end >>
