magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 3 49 1137 241
rect 0 0 1152 49
<< scnmos >>
rect 82 47 112 215
rect 168 47 198 215
rect 254 47 284 215
rect 340 47 370 215
rect 426 47 456 215
rect 512 47 542 215
rect 598 47 628 215
rect 684 47 714 215
rect 770 47 800 215
rect 856 47 886 215
rect 942 47 972 215
rect 1028 47 1058 215
<< scpmoshvt >>
rect 82 367 112 619
rect 168 367 198 619
rect 254 367 284 619
rect 340 367 370 619
rect 426 367 456 619
rect 512 367 542 619
rect 598 367 628 619
rect 684 367 714 619
rect 770 367 800 619
rect 856 367 886 619
rect 942 367 972 619
rect 1028 367 1058 619
<< ndiff >>
rect 29 192 82 215
rect 29 158 37 192
rect 71 158 82 192
rect 29 93 82 158
rect 29 59 37 93
rect 71 59 82 93
rect 29 47 82 59
rect 112 192 168 215
rect 112 158 123 192
rect 157 158 168 192
rect 112 101 168 158
rect 112 67 123 101
rect 157 67 168 101
rect 112 47 168 67
rect 198 131 254 215
rect 198 97 209 131
rect 243 97 254 131
rect 198 47 254 97
rect 284 192 340 215
rect 284 158 295 192
rect 329 158 340 192
rect 284 101 340 158
rect 284 67 295 101
rect 329 67 340 101
rect 284 47 340 67
rect 370 131 426 215
rect 370 97 381 131
rect 415 97 426 131
rect 370 47 426 97
rect 456 192 512 215
rect 456 158 467 192
rect 501 158 512 192
rect 456 101 512 158
rect 456 67 467 101
rect 501 67 512 101
rect 456 47 512 67
rect 542 95 598 215
rect 542 61 553 95
rect 587 61 598 95
rect 542 47 598 61
rect 628 175 684 215
rect 628 141 639 175
rect 673 141 684 175
rect 628 101 684 141
rect 628 67 639 101
rect 673 67 684 101
rect 628 47 684 67
rect 714 95 770 215
rect 714 61 725 95
rect 759 61 770 95
rect 714 47 770 61
rect 800 175 856 215
rect 800 141 811 175
rect 845 141 856 175
rect 800 101 856 141
rect 800 67 811 101
rect 845 67 856 101
rect 800 47 856 67
rect 886 95 942 215
rect 886 61 897 95
rect 931 61 942 95
rect 886 47 942 61
rect 972 175 1028 215
rect 972 141 983 175
rect 1017 141 1028 175
rect 972 101 1028 141
rect 972 67 983 101
rect 1017 67 1028 101
rect 972 47 1028 67
rect 1058 93 1111 215
rect 1058 59 1069 93
rect 1103 59 1111 93
rect 1058 47 1111 59
<< pdiff >>
rect 29 599 82 619
rect 29 565 37 599
rect 71 565 82 599
rect 29 513 82 565
rect 29 479 37 513
rect 71 479 82 513
rect 29 413 82 479
rect 29 379 37 413
rect 71 379 82 413
rect 29 367 82 379
rect 112 607 168 619
rect 112 573 123 607
rect 157 573 168 607
rect 112 531 168 573
rect 112 497 123 531
rect 157 497 168 531
rect 112 455 168 497
rect 112 421 123 455
rect 157 421 168 455
rect 112 367 168 421
rect 198 599 254 619
rect 198 565 209 599
rect 243 565 254 599
rect 198 513 254 565
rect 198 479 209 513
rect 243 479 254 513
rect 198 413 254 479
rect 198 379 209 413
rect 243 379 254 413
rect 198 367 254 379
rect 284 607 340 619
rect 284 573 295 607
rect 329 573 340 607
rect 284 531 340 573
rect 284 497 295 531
rect 329 497 340 531
rect 284 455 340 497
rect 284 421 295 455
rect 329 421 340 455
rect 284 367 340 421
rect 370 599 426 619
rect 370 565 381 599
rect 415 565 426 599
rect 370 513 426 565
rect 370 479 381 513
rect 415 479 426 513
rect 370 413 426 479
rect 370 379 381 413
rect 415 379 426 413
rect 370 367 426 379
rect 456 607 512 619
rect 456 573 467 607
rect 501 573 512 607
rect 456 526 512 573
rect 456 492 467 526
rect 501 492 512 526
rect 456 445 512 492
rect 456 411 467 445
rect 501 411 512 445
rect 456 367 512 411
rect 542 481 598 619
rect 542 447 553 481
rect 587 447 598 481
rect 542 413 598 447
rect 542 379 553 413
rect 587 379 598 413
rect 542 367 598 379
rect 628 585 684 619
rect 628 551 639 585
rect 673 551 684 585
rect 628 367 684 551
rect 714 425 770 619
rect 714 391 725 425
rect 759 391 770 425
rect 714 367 770 391
rect 800 585 856 619
rect 800 551 811 585
rect 845 551 856 585
rect 800 367 856 551
rect 886 413 942 619
rect 886 379 897 413
rect 931 379 942 413
rect 886 367 942 379
rect 972 585 1028 619
rect 972 551 983 585
rect 1017 551 1028 585
rect 972 367 1028 551
rect 1058 607 1115 619
rect 1058 573 1073 607
rect 1107 573 1115 607
rect 1058 539 1115 573
rect 1058 505 1073 539
rect 1107 505 1115 539
rect 1058 465 1115 505
rect 1058 431 1073 465
rect 1107 431 1115 465
rect 1058 367 1115 431
<< ndiffc >>
rect 37 158 71 192
rect 37 59 71 93
rect 123 158 157 192
rect 123 67 157 101
rect 209 97 243 131
rect 295 158 329 192
rect 295 67 329 101
rect 381 97 415 131
rect 467 158 501 192
rect 467 67 501 101
rect 553 61 587 95
rect 639 141 673 175
rect 639 67 673 101
rect 725 61 759 95
rect 811 141 845 175
rect 811 67 845 101
rect 897 61 931 95
rect 983 141 1017 175
rect 983 67 1017 101
rect 1069 59 1103 93
<< pdiffc >>
rect 37 565 71 599
rect 37 479 71 513
rect 37 379 71 413
rect 123 573 157 607
rect 123 497 157 531
rect 123 421 157 455
rect 209 565 243 599
rect 209 479 243 513
rect 209 379 243 413
rect 295 573 329 607
rect 295 497 329 531
rect 295 421 329 455
rect 381 565 415 599
rect 381 479 415 513
rect 381 379 415 413
rect 467 573 501 607
rect 467 492 501 526
rect 467 411 501 445
rect 553 447 587 481
rect 553 379 587 413
rect 639 551 673 585
rect 725 391 759 425
rect 811 551 845 585
rect 897 379 931 413
rect 983 551 1017 585
rect 1073 573 1107 607
rect 1073 505 1107 539
rect 1073 431 1107 465
<< poly >>
rect 82 619 112 645
rect 168 619 198 645
rect 254 619 284 645
rect 340 619 370 645
rect 426 619 456 645
rect 512 619 542 645
rect 598 619 628 645
rect 684 619 714 645
rect 770 619 800 645
rect 856 619 886 645
rect 942 619 972 645
rect 1028 619 1058 645
rect 82 303 112 367
rect 168 303 198 367
rect 254 303 284 367
rect 340 303 370 367
rect 32 287 370 303
rect 32 253 48 287
rect 82 253 116 287
rect 150 253 184 287
rect 218 253 252 287
rect 286 253 320 287
rect 354 253 370 287
rect 32 237 370 253
rect 82 215 112 237
rect 168 215 198 237
rect 254 215 284 237
rect 340 215 370 237
rect 426 303 456 367
rect 512 303 542 367
rect 598 303 628 367
rect 426 287 628 303
rect 426 253 442 287
rect 476 253 510 287
rect 544 253 578 287
rect 612 253 628 287
rect 426 237 628 253
rect 426 215 456 237
rect 512 215 542 237
rect 598 215 628 237
rect 684 335 714 367
rect 770 335 800 367
rect 856 335 886 367
rect 942 335 972 367
rect 684 319 972 335
rect 684 285 700 319
rect 734 285 768 319
rect 802 285 836 319
rect 870 285 904 319
rect 938 285 972 319
rect 1028 303 1058 367
rect 684 269 972 285
rect 684 215 714 269
rect 770 215 800 269
rect 856 215 886 269
rect 942 215 972 269
rect 1014 287 1080 303
rect 1014 253 1030 287
rect 1064 253 1080 287
rect 1014 237 1080 253
rect 1028 215 1058 237
rect 82 21 112 47
rect 168 21 198 47
rect 254 21 284 47
rect 340 21 370 47
rect 426 21 456 47
rect 512 21 542 47
rect 598 21 628 47
rect 684 21 714 47
rect 770 21 800 47
rect 856 21 886 47
rect 942 21 972 47
rect 1028 21 1058 47
<< polycont >>
rect 48 253 82 287
rect 116 253 150 287
rect 184 253 218 287
rect 252 253 286 287
rect 320 253 354 287
rect 442 253 476 287
rect 510 253 544 287
rect 578 253 612 287
rect 700 285 734 319
rect 768 285 802 319
rect 836 285 870 319
rect 904 285 938 319
rect 1030 253 1064 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 21 599 73 615
rect 21 565 37 599
rect 71 565 73 599
rect 21 513 73 565
rect 21 479 37 513
rect 71 479 73 513
rect 21 413 73 479
rect 107 607 173 649
rect 107 573 123 607
rect 157 573 173 607
rect 107 531 173 573
rect 107 497 123 531
rect 157 497 173 531
rect 107 455 173 497
rect 107 421 123 455
rect 157 421 173 455
rect 207 599 245 615
rect 207 565 209 599
rect 243 565 245 599
rect 207 513 245 565
rect 207 479 209 513
rect 243 479 245 513
rect 21 379 37 413
rect 71 379 73 413
rect 21 375 73 379
rect 207 413 245 479
rect 279 607 345 649
rect 279 573 295 607
rect 329 573 345 607
rect 279 531 345 573
rect 279 497 295 531
rect 329 497 345 531
rect 279 455 345 497
rect 279 421 295 455
rect 329 421 345 455
rect 379 599 417 615
rect 379 565 381 599
rect 415 565 417 599
rect 379 513 417 565
rect 379 479 381 513
rect 415 479 417 513
rect 207 379 209 413
rect 243 379 245 413
rect 207 375 245 379
rect 379 413 417 479
rect 379 379 381 413
rect 415 379 417 413
rect 451 607 1021 615
rect 451 573 467 607
rect 501 585 1021 607
rect 501 573 639 585
rect 451 551 639 573
rect 673 551 811 585
rect 845 551 983 585
rect 1017 551 1021 585
rect 451 535 1021 551
rect 1057 607 1123 615
rect 1057 573 1073 607
rect 1107 573 1123 607
rect 1057 539 1123 573
rect 451 526 517 535
rect 451 492 467 526
rect 501 492 517 526
rect 1057 505 1073 539
rect 1107 505 1123 539
rect 1057 499 1123 505
rect 451 445 517 492
rect 451 411 467 445
rect 501 411 517 445
rect 551 481 1123 499
rect 551 447 553 481
rect 587 465 1123 481
rect 587 447 603 465
rect 551 413 603 447
rect 1057 431 1073 465
rect 1107 431 1123 465
rect 379 375 417 379
rect 551 379 553 413
rect 587 379 603 413
rect 709 425 947 431
rect 709 391 725 425
rect 759 413 947 425
rect 759 391 897 413
rect 709 387 897 391
rect 551 375 603 379
rect 21 341 603 375
rect 881 379 897 387
rect 931 397 947 413
rect 931 379 1134 397
rect 881 363 1134 379
rect 684 329 847 353
rect 684 319 954 329
rect 19 287 370 303
rect 19 253 48 287
rect 82 253 116 287
rect 150 253 184 287
rect 218 253 252 287
rect 286 253 320 287
rect 354 253 370 287
rect 19 242 370 253
rect 404 287 650 303
rect 404 253 442 287
rect 476 253 510 287
rect 544 253 578 287
rect 612 253 650 287
rect 684 285 700 319
rect 734 285 768 319
rect 802 285 836 319
rect 870 285 904 319
rect 938 285 954 319
rect 684 283 954 285
rect 1014 287 1066 303
rect 404 249 650 253
rect 1014 253 1030 287
rect 1064 253 1066 287
rect 1014 249 1066 253
rect 404 242 1066 249
rect 607 215 1066 242
rect 21 192 81 208
rect 21 158 37 192
rect 71 158 81 192
rect 21 93 81 158
rect 21 59 37 93
rect 71 59 81 93
rect 21 17 81 59
rect 115 192 573 208
rect 115 158 123 192
rect 157 174 295 192
rect 157 158 159 174
rect 115 101 159 158
rect 293 158 295 174
rect 329 174 467 192
rect 329 158 331 174
rect 115 67 123 101
rect 157 67 159 101
rect 115 51 159 67
rect 193 131 259 140
rect 193 97 209 131
rect 243 97 259 131
rect 193 17 259 97
rect 293 101 331 158
rect 465 158 467 174
rect 501 179 573 192
rect 1100 179 1134 363
rect 501 175 1134 179
rect 501 158 639 175
rect 465 145 639 158
rect 293 67 295 101
rect 329 67 331 101
rect 293 51 331 67
rect 365 131 431 140
rect 365 97 381 131
rect 415 97 431 131
rect 365 17 431 97
rect 465 101 509 145
rect 623 141 639 145
rect 673 145 811 175
rect 673 141 689 145
rect 465 67 467 101
rect 501 67 509 101
rect 465 51 509 67
rect 543 95 589 111
rect 543 61 553 95
rect 587 61 589 95
rect 543 17 589 61
rect 623 101 689 141
rect 795 141 811 145
rect 845 145 983 175
rect 845 141 861 145
rect 623 67 639 101
rect 673 67 689 101
rect 623 51 689 67
rect 723 95 761 111
rect 723 61 725 95
rect 759 61 761 95
rect 723 17 761 61
rect 795 101 861 141
rect 967 141 983 145
rect 1017 145 1134 175
rect 1017 141 1033 145
rect 795 67 811 101
rect 845 67 861 101
rect 795 51 861 67
rect 895 95 933 111
rect 895 61 897 95
rect 931 61 933 95
rect 895 17 933 61
rect 967 101 1033 141
rect 967 67 983 101
rect 1017 67 1033 101
rect 967 51 1033 67
rect 1067 93 1119 111
rect 1067 59 1069 93
rect 1103 59 1119 93
rect 1067 17 1119 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor3_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2493482
string GDS_START 2483266
<< end >>
