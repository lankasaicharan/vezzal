magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 19 49 671 241
rect 0 0 672 49
<< scnmos >>
rect 98 47 128 215
rect 274 47 304 215
rect 360 47 390 215
rect 474 47 504 215
rect 562 47 592 215
<< scpmoshvt >>
rect 98 367 128 619
rect 195 367 225 619
rect 382 367 412 619
rect 468 367 498 619
rect 562 367 592 619
<< ndiff >>
rect 45 187 98 215
rect 45 153 53 187
rect 87 153 98 187
rect 45 103 98 153
rect 45 69 53 103
rect 87 69 98 103
rect 45 47 98 69
rect 128 125 274 215
rect 128 91 139 125
rect 173 91 229 125
rect 263 91 274 125
rect 128 47 274 91
rect 304 47 360 215
rect 390 47 474 215
rect 504 47 562 215
rect 592 201 645 215
rect 592 167 603 201
rect 637 167 645 201
rect 592 103 645 167
rect 592 69 603 103
rect 637 69 645 103
rect 592 47 645 69
<< pdiff >>
rect 45 599 98 619
rect 45 565 53 599
rect 87 565 98 599
rect 45 509 98 565
rect 45 475 53 509
rect 87 475 98 509
rect 45 413 98 475
rect 45 379 53 413
rect 87 379 98 413
rect 45 367 98 379
rect 128 599 195 619
rect 128 565 139 599
rect 173 565 195 599
rect 128 522 195 565
rect 128 488 139 522
rect 173 488 195 522
rect 128 441 195 488
rect 128 407 139 441
rect 173 407 195 441
rect 128 367 195 407
rect 225 607 382 619
rect 225 573 236 607
rect 270 573 337 607
rect 371 573 382 607
rect 225 514 382 573
rect 225 480 236 514
rect 270 492 382 514
rect 270 480 337 492
rect 225 458 337 480
rect 371 458 382 492
rect 225 367 382 458
rect 412 599 468 619
rect 412 565 423 599
rect 457 565 468 599
rect 412 509 468 565
rect 412 475 423 509
rect 457 475 468 509
rect 412 418 468 475
rect 412 384 423 418
rect 457 384 468 418
rect 412 367 468 384
rect 498 607 562 619
rect 498 573 513 607
rect 547 573 562 607
rect 498 492 562 573
rect 498 458 513 492
rect 547 458 562 492
rect 498 367 562 458
rect 592 599 645 619
rect 592 565 603 599
rect 637 565 645 599
rect 592 509 645 565
rect 592 475 603 509
rect 637 475 645 509
rect 592 418 645 475
rect 592 384 603 418
rect 637 384 645 418
rect 592 367 645 384
<< ndiffc >>
rect 53 153 87 187
rect 53 69 87 103
rect 139 91 173 125
rect 229 91 263 125
rect 603 167 637 201
rect 603 69 637 103
<< pdiffc >>
rect 53 565 87 599
rect 53 475 87 509
rect 53 379 87 413
rect 139 565 173 599
rect 139 488 173 522
rect 139 407 173 441
rect 236 573 270 607
rect 337 573 371 607
rect 236 480 270 514
rect 337 458 371 492
rect 423 565 457 599
rect 423 475 457 509
rect 423 384 457 418
rect 513 573 547 607
rect 513 458 547 492
rect 603 565 637 599
rect 603 475 637 509
rect 603 384 637 418
<< poly >>
rect 98 619 128 645
rect 195 619 225 645
rect 382 619 412 645
rect 468 619 498 645
rect 562 619 592 645
rect 98 303 128 367
rect 31 287 128 303
rect 31 253 47 287
rect 81 253 128 287
rect 31 237 128 253
rect 195 308 225 367
rect 382 308 412 367
rect 195 292 304 308
rect 195 258 211 292
rect 245 258 304 292
rect 195 242 304 258
rect 346 292 412 308
rect 468 303 498 367
rect 562 303 592 367
rect 346 258 362 292
rect 396 258 412 292
rect 346 242 412 258
rect 454 287 520 303
rect 454 253 470 287
rect 504 253 520 287
rect 98 215 128 237
rect 274 215 304 242
rect 360 215 390 242
rect 454 237 520 253
rect 562 287 634 303
rect 562 253 584 287
rect 618 253 634 287
rect 562 237 634 253
rect 474 215 504 237
rect 562 215 592 237
rect 98 21 128 47
rect 274 21 304 47
rect 360 21 390 47
rect 474 21 504 47
rect 562 21 592 47
<< polycont >>
rect 47 253 81 287
rect 211 258 245 292
rect 362 258 396 292
rect 470 253 504 287
rect 584 253 618 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 37 599 89 615
rect 37 565 53 599
rect 87 565 89 599
rect 37 509 89 565
rect 37 475 53 509
rect 87 475 89 509
rect 37 413 89 475
rect 37 379 53 413
rect 87 379 89 413
rect 123 599 181 615
rect 123 565 139 599
rect 173 565 181 599
rect 123 522 181 565
rect 123 488 139 522
rect 173 488 181 522
rect 123 441 181 488
rect 215 607 387 649
rect 215 573 236 607
rect 270 573 337 607
rect 371 573 387 607
rect 215 514 387 573
rect 215 480 236 514
rect 270 492 387 514
rect 270 480 337 492
rect 215 475 337 480
rect 291 458 337 475
rect 371 458 387 492
rect 291 453 387 458
rect 421 599 463 615
rect 421 565 423 599
rect 457 565 463 599
rect 421 509 463 565
rect 421 475 423 509
rect 457 475 463 509
rect 123 407 139 441
rect 173 419 257 441
rect 421 419 463 475
rect 497 607 563 649
rect 497 573 513 607
rect 547 573 563 607
rect 497 492 563 573
rect 497 458 513 492
rect 547 458 563 492
rect 497 452 563 458
rect 597 599 653 615
rect 597 565 603 599
rect 637 565 653 599
rect 597 509 653 565
rect 597 475 603 509
rect 637 475 653 509
rect 173 418 463 419
rect 597 418 653 475
rect 173 407 423 418
rect 223 385 423 407
rect 327 384 423 385
rect 457 384 603 418
rect 637 384 653 418
rect 37 373 89 379
rect 37 339 174 373
rect 17 287 81 303
rect 17 253 47 287
rect 17 237 81 253
rect 115 203 174 339
rect 208 292 271 350
rect 208 258 211 292
rect 245 258 271 292
rect 208 235 271 258
rect 305 292 412 350
rect 305 258 362 292
rect 396 258 412 292
rect 305 235 412 258
rect 454 287 550 350
rect 454 253 470 287
rect 504 253 550 287
rect 454 235 550 253
rect 584 287 655 350
rect 618 253 655 287
rect 584 237 655 253
rect 37 201 174 203
rect 37 187 603 201
rect 37 153 53 187
rect 87 167 603 187
rect 637 167 653 201
rect 87 153 89 167
rect 37 103 89 153
rect 37 69 53 103
rect 87 69 89 103
rect 37 53 89 69
rect 123 125 279 133
rect 123 91 139 125
rect 173 91 229 125
rect 263 91 279 125
rect 123 17 279 91
rect 587 103 653 167
rect 587 69 603 103
rect 637 69 653 103
rect 587 53 653 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a41oi_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1339194
string GDS_START 1332212
<< end >>
