magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 225 172 671 241
rect 2 49 671 172
rect 0 0 672 49
<< scnmos >>
rect 85 62 115 146
rect 304 47 334 215
rect 390 47 420 215
rect 476 47 506 215
rect 562 47 592 215
<< scpmoshvt >>
rect 85 367 115 495
rect 190 367 220 619
rect 276 367 306 619
rect 476 367 506 619
rect 562 367 592 619
<< ndiff >>
rect 251 203 304 215
rect 251 169 259 203
rect 293 169 304 203
rect 28 121 85 146
rect 28 87 36 121
rect 70 87 85 121
rect 28 62 85 87
rect 115 108 168 146
rect 115 74 126 108
rect 160 74 168 108
rect 115 62 168 74
rect 251 101 304 169
rect 251 67 259 101
rect 293 67 304 101
rect 251 47 304 67
rect 334 167 390 215
rect 334 133 345 167
rect 379 133 390 167
rect 334 93 390 133
rect 334 59 345 93
rect 379 59 390 93
rect 334 47 390 59
rect 420 203 476 215
rect 420 169 431 203
rect 465 169 476 203
rect 420 101 476 169
rect 420 67 431 101
rect 465 67 476 101
rect 420 47 476 67
rect 506 161 562 215
rect 506 127 517 161
rect 551 127 562 161
rect 506 47 562 127
rect 592 189 645 215
rect 592 155 603 189
rect 637 155 645 189
rect 592 101 645 155
rect 592 67 603 101
rect 637 67 645 101
rect 592 47 645 67
<< pdiff >>
rect 137 607 190 619
rect 137 573 145 607
rect 179 573 190 607
rect 137 522 190 573
rect 137 495 145 522
rect 32 481 85 495
rect 32 447 40 481
rect 74 447 85 481
rect 32 413 85 447
rect 32 379 40 413
rect 74 379 85 413
rect 32 367 85 379
rect 115 488 145 495
rect 179 488 190 522
rect 115 438 190 488
rect 115 404 136 438
rect 170 404 190 438
rect 115 367 190 404
rect 220 599 276 619
rect 220 565 231 599
rect 265 565 276 599
rect 220 526 276 565
rect 220 492 231 526
rect 265 492 276 526
rect 220 454 276 492
rect 220 420 231 454
rect 265 420 276 454
rect 220 367 276 420
rect 306 575 359 619
rect 306 541 317 575
rect 351 541 359 575
rect 306 367 359 541
rect 423 415 476 619
rect 423 381 431 415
rect 465 381 476 415
rect 423 367 476 381
rect 506 599 562 619
rect 506 565 517 599
rect 551 565 562 599
rect 506 529 562 565
rect 506 495 517 529
rect 551 495 562 529
rect 506 459 562 495
rect 506 425 517 459
rect 551 425 562 459
rect 506 367 562 425
rect 592 599 645 619
rect 592 565 603 599
rect 637 565 645 599
rect 592 507 645 565
rect 592 473 603 507
rect 637 473 645 507
rect 592 413 645 473
rect 592 379 603 413
rect 637 379 645 413
rect 592 367 645 379
<< ndiffc >>
rect 259 169 293 203
rect 36 87 70 121
rect 126 74 160 108
rect 259 67 293 101
rect 345 133 379 167
rect 345 59 379 93
rect 431 169 465 203
rect 431 67 465 101
rect 517 127 551 161
rect 603 155 637 189
rect 603 67 637 101
<< pdiffc >>
rect 145 573 179 607
rect 40 447 74 481
rect 40 379 74 413
rect 145 488 179 522
rect 136 404 170 438
rect 231 565 265 599
rect 231 492 265 526
rect 231 420 265 454
rect 317 541 351 575
rect 431 381 465 415
rect 517 565 551 599
rect 517 495 551 529
rect 517 425 551 459
rect 603 565 637 599
rect 603 473 637 507
rect 603 379 637 413
<< poly >>
rect 190 619 220 645
rect 276 619 306 645
rect 476 619 506 645
rect 562 619 592 645
rect 85 495 115 521
rect 85 345 115 367
rect 190 345 220 367
rect 276 345 306 367
rect 85 315 306 345
rect 85 286 160 315
rect 85 252 110 286
rect 144 252 160 286
rect 354 305 420 321
rect 354 271 370 305
rect 404 271 420 305
rect 354 267 420 271
rect 85 218 160 252
rect 85 184 110 218
rect 144 184 160 218
rect 304 237 420 267
rect 304 215 334 237
rect 390 215 420 237
rect 476 305 506 367
rect 562 305 592 367
rect 476 289 631 305
rect 476 275 581 289
rect 476 215 506 275
rect 562 255 581 275
rect 615 255 631 289
rect 562 239 631 255
rect 562 215 592 239
rect 85 168 160 184
rect 85 146 115 168
rect 85 36 115 62
rect 304 21 334 47
rect 390 21 420 47
rect 476 21 506 47
rect 562 21 592 47
<< polycont >>
rect 110 252 144 286
rect 370 271 404 305
rect 110 184 144 218
rect 581 255 615 289
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 120 607 186 649
rect 120 573 145 607
rect 179 573 186 607
rect 120 522 186 573
rect 20 481 86 497
rect 20 447 40 481
rect 74 447 86 481
rect 20 413 86 447
rect 20 379 40 413
rect 74 379 86 413
rect 120 488 145 522
rect 179 488 186 522
rect 120 438 186 488
rect 120 404 136 438
rect 170 404 186 438
rect 220 599 267 615
rect 220 565 231 599
rect 265 565 267 599
rect 220 526 267 565
rect 301 575 367 649
rect 301 541 317 575
rect 351 541 367 575
rect 301 533 367 541
rect 501 599 561 615
rect 501 565 517 599
rect 551 565 561 599
rect 220 492 231 526
rect 265 499 267 526
rect 501 529 561 565
rect 501 499 517 529
rect 265 495 517 499
rect 551 495 561 529
rect 265 492 561 495
rect 220 465 561 492
rect 220 454 281 465
rect 220 420 231 454
rect 265 420 281 454
rect 508 459 561 465
rect 220 404 281 420
rect 422 415 474 431
rect 20 370 86 379
rect 422 381 431 415
rect 465 381 474 415
rect 508 425 517 459
rect 551 425 561 459
rect 508 409 561 425
rect 595 599 653 615
rect 595 565 603 599
rect 637 565 653 599
rect 595 507 653 565
rect 595 473 603 507
rect 637 473 653 507
rect 595 413 653 473
rect 422 375 474 381
rect 595 379 603 413
rect 637 379 653 413
rect 595 375 653 379
rect 20 336 388 370
rect 422 341 653 375
rect 20 121 74 336
rect 354 307 388 336
rect 354 305 420 307
rect 110 286 189 302
rect 144 252 189 286
rect 354 271 370 305
rect 404 271 420 305
rect 354 269 420 271
rect 110 218 189 252
rect 144 184 189 218
rect 110 168 189 184
rect 243 203 465 235
rect 243 169 259 203
rect 293 201 431 203
rect 293 169 295 201
rect 20 87 36 121
rect 70 87 74 121
rect 20 71 74 87
rect 110 108 176 112
rect 110 74 126 108
rect 160 74 176 108
rect 110 17 176 74
rect 243 101 295 169
rect 429 169 431 201
rect 243 67 259 101
rect 293 67 295 101
rect 243 51 295 67
rect 329 133 345 167
rect 379 133 395 167
rect 329 93 395 133
rect 329 59 345 93
rect 379 59 395 93
rect 329 17 395 59
rect 429 101 465 169
rect 499 177 547 341
rect 581 289 655 305
rect 615 255 655 289
rect 581 239 655 255
rect 601 189 653 205
rect 499 161 567 177
rect 499 127 517 161
rect 551 127 567 161
rect 499 119 567 127
rect 601 155 603 189
rect 637 155 653 189
rect 429 67 431 101
rect 601 101 653 155
rect 601 85 603 101
rect 465 67 603 85
rect 637 67 653 101
rect 429 51 653 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 einvn_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4208680
string GDS_START 4202210
<< end >>
