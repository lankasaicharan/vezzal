magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1400 -1260 11646 1960
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_0
timestamp 1627201311
transform -1 0 -40 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_1
timestamp 1627201311
transform 1 0 314 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_2
timestamp 1627201311
transform 1 0 868 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_3
timestamp 1627201311
transform 1 0 1422 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_4
timestamp 1627201311
transform 1 0 1976 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_5
timestamp 1627201311
transform 1 0 2530 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_6
timestamp 1627201311
transform 1 0 3084 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_7
timestamp 1627201311
transform 1 0 3638 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_8
timestamp 1627201311
transform 1 0 4192 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_9
timestamp 1627201311
transform 1 0 4746 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_10
timestamp 1627201311
transform 1 0 5300 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_11
timestamp 1627201311
transform 1 0 5854 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_12
timestamp 1627201311
transform 1 0 6408 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_13
timestamp 1627201311
transform 1 0 6962 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_14
timestamp 1627201311
transform 1 0 7516 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_15
timestamp 1627201311
transform 1 0 8070 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_16
timestamp 1627201311
transform 1 0 8624 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_17
timestamp 1627201311
transform 1 0 9178 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_18
timestamp 1627201311
transform 1 0 9732 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_19
timestamp 1627201311
transform 1 0 10286 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 10386 675 10386 675 0 FreeSans 300 0 0 0 S
flabel comment s 10109 700 10109 700 0 FreeSans 300 0 0 0 D
flabel comment s 9832 675 9832 675 0 FreeSans 300 0 0 0 S
flabel comment s 9555 700 9555 700 0 FreeSans 300 0 0 0 D
flabel comment s 9278 675 9278 675 0 FreeSans 300 0 0 0 S
flabel comment s 9001 700 9001 700 0 FreeSans 300 0 0 0 D
flabel comment s 8724 675 8724 675 0 FreeSans 300 0 0 0 S
flabel comment s 8447 700 8447 700 0 FreeSans 300 0 0 0 D
flabel comment s 8170 675 8170 675 0 FreeSans 300 0 0 0 S
flabel comment s 7893 700 7893 700 0 FreeSans 300 0 0 0 D
flabel comment s 7616 675 7616 675 0 FreeSans 300 0 0 0 S
flabel comment s 7339 700 7339 700 0 FreeSans 300 0 0 0 D
flabel comment s 7062 675 7062 675 0 FreeSans 300 0 0 0 S
flabel comment s 6785 700 6785 700 0 FreeSans 300 0 0 0 D
flabel comment s 6508 675 6508 675 0 FreeSans 300 0 0 0 S
flabel comment s 6231 700 6231 700 0 FreeSans 300 0 0 0 D
flabel comment s 5954 675 5954 675 0 FreeSans 300 0 0 0 S
flabel comment s 5677 700 5677 700 0 FreeSans 300 0 0 0 D
flabel comment s 5400 675 5400 675 0 FreeSans 300 0 0 0 S
flabel comment s 5123 700 5123 700 0 FreeSans 300 0 0 0 D
flabel comment s 4846 675 4846 675 0 FreeSans 300 0 0 0 S
flabel comment s 4569 700 4569 700 0 FreeSans 300 0 0 0 D
flabel comment s 4292 675 4292 675 0 FreeSans 300 0 0 0 S
flabel comment s 4015 700 4015 700 0 FreeSans 300 0 0 0 D
flabel comment s 3738 675 3738 675 0 FreeSans 300 0 0 0 S
flabel comment s 3461 700 3461 700 0 FreeSans 300 0 0 0 D
flabel comment s 3184 675 3184 675 0 FreeSans 300 0 0 0 S
flabel comment s 2907 700 2907 700 0 FreeSans 300 0 0 0 D
flabel comment s 2630 675 2630 675 0 FreeSans 300 0 0 0 S
flabel comment s 2353 700 2353 700 0 FreeSans 300 0 0 0 D
flabel comment s 2076 675 2076 675 0 FreeSans 300 0 0 0 S
flabel comment s 1799 700 1799 700 0 FreeSans 300 0 0 0 D
flabel comment s 1522 675 1522 675 0 FreeSans 300 0 0 0 S
flabel comment s 1245 700 1245 700 0 FreeSans 300 0 0 0 D
flabel comment s 968 675 968 675 0 FreeSans 300 0 0 0 S
flabel comment s 691 700 691 700 0 FreeSans 300 0 0 0 D
flabel comment s 414 675 414 675 0 FreeSans 300 0 0 0 S
flabel comment s 137 700 137 700 0 FreeSans 300 0 0 0 D
flabel comment s -140 675 -140 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 15528204
string GDS_START 15508364
<< end >>
