magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 395 241 669 263
rect 4 49 669 241
rect 0 0 672 49
<< scnmos >>
rect 83 131 113 215
rect 188 47 218 215
rect 274 47 304 215
rect 474 69 504 237
rect 560 69 590 237
<< scpmoshvt >>
rect 83 367 113 495
rect 302 367 332 619
rect 388 367 418 619
rect 474 367 504 619
rect 560 367 590 619
<< ndiff >>
rect 421 225 474 237
rect 30 194 83 215
rect 30 160 38 194
rect 72 160 83 194
rect 30 131 83 160
rect 113 203 188 215
rect 113 169 124 203
rect 158 169 188 203
rect 113 131 188 169
rect 135 93 188 131
rect 135 59 143 93
rect 177 59 188 93
rect 135 47 188 59
rect 218 203 274 215
rect 218 169 229 203
rect 263 169 274 203
rect 218 101 274 169
rect 218 67 229 101
rect 263 67 274 101
rect 218 47 274 67
rect 304 179 357 215
rect 304 145 315 179
rect 349 145 357 179
rect 304 93 357 145
rect 304 59 315 93
rect 349 59 357 93
rect 421 191 429 225
rect 463 191 474 225
rect 421 115 474 191
rect 421 81 429 115
rect 463 81 474 115
rect 421 69 474 81
rect 504 229 560 237
rect 504 195 515 229
rect 549 195 560 229
rect 504 153 560 195
rect 504 119 515 153
rect 549 119 560 153
rect 504 69 560 119
rect 590 192 643 237
rect 590 158 601 192
rect 635 158 643 192
rect 590 115 643 158
rect 590 81 601 115
rect 635 81 643 115
rect 590 69 643 81
rect 304 47 357 59
<< pdiff >>
rect 249 599 302 619
rect 30 481 83 495
rect 30 447 38 481
rect 72 447 83 481
rect 30 413 83 447
rect 30 379 38 413
rect 72 379 83 413
rect 30 367 83 379
rect 113 483 166 495
rect 113 449 124 483
rect 158 449 166 483
rect 113 415 166 449
rect 113 381 124 415
rect 158 381 166 415
rect 113 367 166 381
rect 249 565 257 599
rect 291 565 302 599
rect 249 510 302 565
rect 249 476 257 510
rect 291 476 302 510
rect 249 413 302 476
rect 249 379 257 413
rect 291 379 302 413
rect 249 367 302 379
rect 332 611 388 619
rect 332 577 343 611
rect 377 577 388 611
rect 332 537 388 577
rect 332 503 343 537
rect 377 503 388 537
rect 332 457 388 503
rect 332 423 343 457
rect 377 423 388 457
rect 332 367 388 423
rect 418 599 474 619
rect 418 565 429 599
rect 463 565 474 599
rect 418 502 474 565
rect 418 468 429 502
rect 463 468 474 502
rect 418 409 474 468
rect 418 375 429 409
rect 463 375 474 409
rect 418 367 474 375
rect 504 536 560 619
rect 504 502 515 536
rect 549 502 560 536
rect 504 414 560 502
rect 504 380 515 414
rect 549 380 560 414
rect 504 367 560 380
rect 590 599 643 619
rect 590 565 601 599
rect 635 565 643 599
rect 590 517 643 565
rect 590 483 601 517
rect 635 483 643 517
rect 590 434 643 483
rect 590 400 601 434
rect 635 400 643 434
rect 590 367 643 400
<< ndiffc >>
rect 38 160 72 194
rect 124 169 158 203
rect 143 59 177 93
rect 229 169 263 203
rect 229 67 263 101
rect 315 145 349 179
rect 315 59 349 93
rect 429 191 463 225
rect 429 81 463 115
rect 515 195 549 229
rect 515 119 549 153
rect 601 158 635 192
rect 601 81 635 115
<< pdiffc >>
rect 38 447 72 481
rect 38 379 72 413
rect 124 449 158 483
rect 124 381 158 415
rect 257 565 291 599
rect 257 476 291 510
rect 257 379 291 413
rect 343 577 377 611
rect 343 503 377 537
rect 343 423 377 457
rect 429 565 463 599
rect 429 468 463 502
rect 429 375 463 409
rect 515 502 549 536
rect 515 380 549 414
rect 601 565 635 599
rect 601 483 635 517
rect 601 400 635 434
<< poly >>
rect 82 606 148 622
rect 302 619 332 645
rect 388 619 418 645
rect 474 619 504 645
rect 560 619 590 645
rect 82 572 98 606
rect 132 586 148 606
rect 132 572 218 586
rect 82 556 218 572
rect 83 495 113 556
rect 83 297 113 367
rect 188 297 218 556
rect 302 345 332 367
rect 388 345 418 367
rect 302 319 418 345
rect 302 315 368 319
rect 83 267 218 297
rect 352 285 368 315
rect 402 285 418 319
rect 352 269 418 285
rect 474 289 504 367
rect 560 325 590 367
rect 560 309 651 325
rect 560 289 601 309
rect 474 275 601 289
rect 635 275 651 309
rect 83 215 113 267
rect 188 237 304 267
rect 474 259 651 275
rect 474 237 504 259
rect 560 237 590 259
rect 188 215 218 237
rect 274 215 304 237
rect 83 105 113 131
rect 188 21 218 47
rect 274 21 304 47
rect 474 43 504 69
rect 560 43 590 69
<< polycont >>
rect 98 572 132 606
rect 368 285 402 319
rect 601 275 635 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 21 606 148 613
rect 21 572 98 606
rect 132 572 148 606
rect 21 533 148 572
rect 182 499 219 649
rect 22 481 80 497
rect 22 447 38 481
rect 72 447 80 481
rect 22 413 80 447
rect 22 379 38 413
rect 72 379 80 413
rect 22 319 80 379
rect 114 483 219 499
rect 114 449 124 483
rect 158 449 219 483
rect 114 415 219 449
rect 114 381 124 415
rect 158 381 219 415
rect 114 365 219 381
rect 253 599 293 615
rect 253 565 257 599
rect 291 565 293 599
rect 253 510 293 565
rect 253 476 257 510
rect 291 476 293 510
rect 253 413 293 476
rect 327 611 393 649
rect 327 577 343 611
rect 377 577 393 611
rect 327 537 393 577
rect 327 503 343 537
rect 377 503 393 537
rect 327 457 393 503
rect 327 423 343 457
rect 377 423 393 457
rect 427 599 651 615
rect 427 565 429 599
rect 463 581 601 599
rect 463 565 465 581
rect 427 502 465 565
rect 599 565 601 581
rect 635 565 651 599
rect 427 468 429 502
rect 463 468 465 502
rect 253 379 257 413
rect 291 389 293 413
rect 427 409 465 468
rect 427 389 429 409
rect 291 379 429 389
rect 253 375 429 379
rect 463 375 465 409
rect 253 355 465 375
rect 499 536 565 547
rect 499 502 515 536
rect 549 502 565 536
rect 499 414 565 502
rect 499 380 515 414
rect 549 380 565 414
rect 599 517 651 565
rect 599 483 601 517
rect 635 483 651 517
rect 599 434 651 483
rect 599 400 601 434
rect 635 400 651 434
rect 599 384 651 400
rect 22 285 368 319
rect 402 285 418 319
rect 22 194 74 285
rect 219 225 465 247
rect 22 160 38 194
rect 72 160 74 194
rect 22 144 74 160
rect 108 203 185 223
rect 108 169 124 203
rect 158 169 185 203
rect 108 93 185 169
rect 108 59 143 93
rect 177 59 185 93
rect 108 17 185 59
rect 219 213 429 225
rect 219 203 265 213
rect 219 169 229 203
rect 263 169 265 203
rect 413 191 429 213
rect 463 191 465 225
rect 219 101 265 169
rect 219 67 229 101
rect 263 67 265 101
rect 219 51 265 67
rect 299 145 315 179
rect 349 145 365 179
rect 299 93 365 145
rect 299 59 315 93
rect 349 59 365 93
rect 299 17 365 59
rect 413 115 465 191
rect 499 229 565 380
rect 599 309 651 350
rect 599 275 601 309
rect 635 275 651 309
rect 599 242 651 275
rect 499 195 515 229
rect 549 195 565 229
rect 499 153 565 195
rect 499 119 515 153
rect 549 119 565 153
rect 599 192 651 208
rect 599 158 601 192
rect 635 158 651 192
rect 413 81 429 115
rect 463 85 465 115
rect 599 115 651 158
rect 599 85 601 115
rect 463 81 601 85
rect 635 81 651 115
rect 413 51 651 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 einvp_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3023240
string GDS_START 3016202
<< end >>
