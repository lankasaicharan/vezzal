magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 332 1574 704
<< pwell >>
rect 645 258 1520 279
rect 638 248 1520 258
rect 9 49 1520 248
rect 0 0 1536 49
<< scpmos >>
rect 83 368 119 568
rect 199 368 235 592
rect 289 368 325 592
rect 385 368 421 592
rect 497 368 533 592
rect 607 392 643 592
rect 697 392 733 592
rect 804 392 840 592
rect 1006 392 1042 592
rect 1100 392 1136 592
rect 1190 392 1226 592
rect 1280 392 1316 592
rect 1370 392 1406 592
<< nmoslvt >>
rect 92 94 122 222
rect 203 74 233 222
rect 289 74 319 222
rect 417 74 447 222
rect 503 74 533 222
rect 721 125 751 253
rect 816 125 846 253
rect 934 125 964 253
rect 1020 125 1050 253
rect 1106 125 1136 253
rect 1192 125 1222 253
rect 1278 125 1308 253
rect 1408 125 1438 253
<< ndiff >>
rect 35 166 92 222
rect 35 132 47 166
rect 81 132 92 166
rect 35 94 92 132
rect 122 204 203 222
rect 122 170 133 204
rect 167 170 203 204
rect 122 136 203 170
rect 122 102 133 136
rect 167 102 203 136
rect 122 94 203 102
rect 153 74 203 94
rect 233 210 289 222
rect 233 176 244 210
rect 278 176 289 210
rect 233 120 289 176
rect 233 86 244 120
rect 278 86 289 120
rect 233 74 289 86
rect 319 146 417 222
rect 319 112 350 146
rect 384 112 417 146
rect 319 74 417 112
rect 447 210 503 222
rect 447 176 458 210
rect 492 176 503 210
rect 447 120 503 176
rect 447 86 458 120
rect 492 86 503 120
rect 447 74 503 86
rect 533 210 604 222
rect 533 176 558 210
rect 592 176 604 210
rect 533 120 604 176
rect 533 86 558 120
rect 592 86 604 120
rect 533 74 604 86
rect 671 232 721 253
rect 664 195 721 232
rect 664 161 676 195
rect 710 161 721 195
rect 664 125 721 161
rect 751 176 816 253
rect 751 142 766 176
rect 800 142 816 176
rect 751 125 816 142
rect 846 125 934 253
rect 964 173 1020 253
rect 964 139 975 173
rect 1009 139 1020 173
rect 964 125 1020 139
rect 1050 241 1106 253
rect 1050 207 1061 241
rect 1095 207 1106 241
rect 1050 171 1106 207
rect 1050 137 1061 171
rect 1095 137 1106 171
rect 1050 125 1106 137
rect 1136 173 1192 253
rect 1136 139 1147 173
rect 1181 139 1192 173
rect 1136 125 1192 139
rect 1222 239 1278 253
rect 1222 205 1233 239
rect 1267 205 1278 239
rect 1222 125 1278 205
rect 1308 171 1408 253
rect 1308 137 1341 171
rect 1375 137 1408 171
rect 1308 125 1408 137
rect 1438 173 1494 253
rect 1438 139 1449 173
rect 1483 139 1494 173
rect 1438 125 1494 139
rect 861 124 919 125
rect 861 90 873 124
rect 907 90 919 124
rect 861 78 919 90
<< pdiff >>
rect 134 580 199 592
rect 134 568 150 580
rect 27 556 83 568
rect 27 522 39 556
rect 73 522 83 556
rect 27 485 83 522
rect 27 451 39 485
rect 73 451 83 485
rect 27 414 83 451
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 546 150 568
rect 184 546 199 580
rect 119 368 199 546
rect 235 421 289 592
rect 235 387 245 421
rect 279 387 289 421
rect 235 368 289 387
rect 325 580 385 592
rect 325 546 338 580
rect 372 546 385 580
rect 325 368 385 546
rect 421 421 497 592
rect 421 387 431 421
rect 465 387 497 421
rect 421 368 497 387
rect 533 580 607 592
rect 533 546 544 580
rect 578 546 607 580
rect 533 392 607 546
rect 643 442 697 592
rect 643 408 653 442
rect 687 408 697 442
rect 643 392 697 408
rect 733 580 804 592
rect 733 546 760 580
rect 794 546 804 580
rect 733 392 804 546
rect 840 444 1006 592
rect 840 410 850 444
rect 884 410 962 444
rect 996 410 1006 444
rect 840 392 1006 410
rect 1042 580 1100 592
rect 1042 546 1054 580
rect 1088 546 1100 580
rect 1042 392 1100 546
rect 1136 441 1190 592
rect 1136 407 1146 441
rect 1180 407 1190 441
rect 1136 392 1190 407
rect 1226 580 1280 592
rect 1226 546 1236 580
rect 1270 546 1280 580
rect 1226 392 1280 546
rect 1316 444 1370 592
rect 1316 410 1326 444
rect 1360 410 1370 444
rect 1316 392 1370 410
rect 1406 580 1509 592
rect 1406 546 1439 580
rect 1473 546 1509 580
rect 1406 392 1509 546
rect 533 368 583 392
<< ndiffc >>
rect 47 132 81 166
rect 133 170 167 204
rect 133 102 167 136
rect 244 176 278 210
rect 244 86 278 120
rect 350 112 384 146
rect 458 176 492 210
rect 458 86 492 120
rect 558 176 592 210
rect 558 86 592 120
rect 676 161 710 195
rect 766 142 800 176
rect 975 139 1009 173
rect 1061 207 1095 241
rect 1061 137 1095 171
rect 1147 139 1181 173
rect 1233 205 1267 239
rect 1341 137 1375 171
rect 1449 139 1483 173
rect 873 90 907 124
<< pdiffc >>
rect 39 522 73 556
rect 39 451 73 485
rect 39 380 73 414
rect 150 546 184 580
rect 245 387 279 421
rect 338 546 372 580
rect 431 387 465 421
rect 544 546 578 580
rect 653 408 687 442
rect 760 546 794 580
rect 850 410 884 444
rect 962 410 996 444
rect 1054 546 1088 580
rect 1146 407 1180 441
rect 1236 546 1270 580
rect 1326 410 1360 444
rect 1439 546 1473 580
<< poly >>
rect 83 568 119 594
rect 199 592 235 618
rect 289 592 325 618
rect 385 592 421 618
rect 497 592 533 618
rect 607 592 643 618
rect 697 592 733 618
rect 804 592 840 618
rect 1006 592 1042 618
rect 1100 592 1136 618
rect 1190 592 1226 618
rect 1280 592 1316 618
rect 1370 592 1406 618
rect 83 310 119 368
rect 83 294 151 310
rect 199 294 235 368
rect 289 330 325 368
rect 385 330 421 368
rect 497 330 533 368
rect 607 336 643 392
rect 697 360 733 392
rect 804 360 840 392
rect 697 344 950 360
rect 1006 347 1042 392
rect 289 314 533 330
rect 289 294 313 314
rect 83 260 101 294
rect 135 260 151 294
rect 83 244 151 260
rect 203 280 313 294
rect 347 280 381 314
rect 415 280 449 314
rect 483 280 533 314
rect 203 264 533 280
rect 583 320 649 336
rect 697 330 832 344
rect 583 286 599 320
rect 633 286 649 320
rect 583 270 649 286
rect 816 310 832 330
rect 866 310 900 344
rect 934 310 950 344
rect 816 299 950 310
rect 92 222 122 244
rect 203 222 233 264
rect 289 222 319 264
rect 417 222 447 264
rect 503 222 533 264
rect 92 68 122 94
rect 203 48 233 74
rect 289 48 319 74
rect 417 48 447 74
rect 503 48 533 74
rect 619 51 649 270
rect 721 253 751 279
rect 816 269 964 299
rect 816 253 846 269
rect 934 253 964 269
rect 1012 298 1042 347
rect 1012 268 1050 298
rect 1100 279 1136 392
rect 1190 360 1226 392
rect 1280 360 1316 392
rect 1190 344 1316 360
rect 1190 324 1266 344
rect 1020 253 1050 268
rect 1106 253 1136 279
rect 1192 310 1266 324
rect 1300 310 1316 344
rect 1192 294 1316 310
rect 1370 360 1406 392
rect 1370 344 1438 360
rect 1370 310 1386 344
rect 1420 310 1438 344
rect 1370 294 1438 310
rect 1192 253 1222 294
rect 1278 253 1308 294
rect 1408 253 1438 294
rect 721 51 751 125
rect 816 99 846 125
rect 934 99 964 125
rect 1020 51 1050 125
rect 619 21 1050 51
rect 1106 51 1136 125
rect 1192 99 1222 125
rect 1278 99 1308 125
rect 1408 51 1438 125
rect 1106 21 1438 51
<< polycont >>
rect 101 260 135 294
rect 313 280 347 314
rect 381 280 415 314
rect 449 280 483 314
rect 599 286 633 320
rect 832 310 866 344
rect 900 310 934 344
rect 1266 310 1300 344
rect 1386 310 1420 344
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 130 580 205 649
rect 17 556 89 572
rect 17 522 39 556
rect 73 522 89 556
rect 130 546 150 580
rect 184 546 205 580
rect 319 580 391 649
rect 319 546 338 580
rect 372 546 391 580
rect 527 580 596 649
rect 527 546 544 580
rect 578 546 596 580
rect 744 580 810 649
rect 744 546 760 580
rect 794 546 810 580
rect 1036 580 1106 649
rect 1036 546 1054 580
rect 1088 546 1106 580
rect 1220 580 1286 649
rect 1220 546 1236 580
rect 1270 546 1286 580
rect 1400 580 1513 649
rect 1400 546 1439 580
rect 1473 546 1513 580
rect 17 512 89 522
rect 17 485 1504 512
rect 17 451 39 485
rect 73 478 1504 485
rect 73 451 89 478
rect 17 414 89 451
rect 17 380 39 414
rect 73 380 89 414
rect 17 364 89 380
rect 217 421 481 444
rect 217 387 245 421
rect 279 387 431 421
rect 465 387 481 421
rect 217 364 481 387
rect 515 442 850 444
rect 515 408 653 442
rect 687 410 850 442
rect 884 410 962 444
rect 996 441 1326 444
rect 996 410 1146 441
rect 687 408 1146 410
rect 515 407 1146 408
rect 1180 410 1326 441
rect 1360 410 1376 444
rect 1180 407 1376 410
rect 515 394 1376 407
rect 515 390 703 394
rect 17 204 51 364
rect 85 294 167 310
rect 85 260 101 294
rect 135 260 167 294
rect 85 238 167 260
rect 217 230 263 364
rect 515 330 549 390
rect 1130 388 1216 394
rect 297 314 549 330
rect 297 280 313 314
rect 347 280 381 314
rect 415 280 449 314
rect 483 280 549 314
rect 297 264 549 280
rect 583 320 649 356
rect 583 286 599 320
rect 633 286 649 320
rect 793 344 1031 360
rect 793 310 832 344
rect 866 310 900 344
rect 934 310 1031 344
rect 793 294 1031 310
rect 583 270 649 286
rect 1182 260 1216 388
rect 1250 344 1335 360
rect 1250 310 1266 344
rect 1300 310 1335 344
rect 1250 294 1335 310
rect 1369 344 1436 360
rect 1369 310 1386 344
rect 1420 310 1436 344
rect 1369 294 1436 310
rect 1301 260 1335 294
rect 1470 260 1504 478
rect 692 241 1095 260
rect 692 236 1061 241
rect 217 210 508 230
rect 660 226 1061 236
rect 17 166 81 204
rect 17 132 47 166
rect 17 90 81 132
rect 117 170 133 204
rect 167 170 183 204
rect 117 136 183 170
rect 117 102 133 136
rect 167 102 183 136
rect 117 17 183 102
rect 217 176 244 210
rect 278 196 458 210
rect 278 176 294 196
rect 217 120 294 176
rect 442 176 458 196
rect 492 176 508 210
rect 217 86 244 120
rect 278 86 294 120
rect 217 70 294 86
rect 334 146 400 162
rect 334 112 350 146
rect 384 112 400 146
rect 334 17 400 112
rect 442 120 508 176
rect 442 86 458 120
rect 492 86 508 120
rect 442 70 508 86
rect 542 210 608 226
rect 542 176 558 210
rect 592 176 608 210
rect 542 120 608 176
rect 660 195 726 226
rect 660 161 676 195
rect 710 161 726 195
rect 1182 239 1267 260
rect 1182 226 1233 239
rect 660 121 726 161
rect 762 176 1025 192
rect 762 142 766 176
rect 800 173 1025 176
rect 800 158 975 173
rect 800 142 821 158
rect 762 126 821 142
rect 959 139 975 158
rect 1009 139 1025 173
rect 542 86 558 120
rect 592 86 608 120
rect 542 17 608 86
rect 857 90 873 124
rect 907 90 923 124
rect 959 121 1025 139
rect 1061 171 1095 207
rect 1216 205 1233 226
rect 1301 226 1504 260
rect 857 17 923 90
rect 1061 85 1095 137
rect 1131 173 1181 192
rect 1216 187 1267 205
rect 1131 139 1147 173
rect 1325 171 1391 187
rect 1325 153 1341 171
rect 1181 139 1341 153
rect 1131 137 1341 139
rect 1375 137 1391 171
rect 1131 119 1391 137
rect 1433 173 1499 192
rect 1433 139 1449 173
rect 1483 139 1499 173
rect 1433 85 1499 139
rect 1061 51 1499 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4b_4
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 3223778
string GDS_START 3212952
<< end >>
