magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 4946 1975
<< nwell >>
rect -38 332 3686 704
<< pwell >>
rect 662 235 1026 272
rect 1447 235 1978 261
rect 2743 248 2931 290
rect 662 229 1978 235
rect 6 218 1978 229
rect 6 192 2073 218
rect 2346 192 3647 248
rect 6 49 3647 192
rect 0 0 3648 49
<< scpmos >>
rect 83 464 119 592
rect 173 464 209 592
rect 251 464 287 592
rect 341 464 377 592
rect 543 464 579 592
rect 745 368 781 592
rect 835 368 871 592
rect 1037 464 1073 548
rect 1121 464 1157 548
rect 1228 464 1264 592
rect 1559 424 1595 592
rect 1643 424 1679 592
rect 1751 424 1787 592
rect 1953 424 1989 592
rect 2031 424 2067 592
rect 2138 508 2174 592
rect 2216 508 2252 592
rect 2421 392 2457 592
rect 2523 392 2559 592
rect 2607 392 2643 592
rect 2809 399 2845 527
rect 3045 368 3081 592
rect 3135 368 3171 592
rect 3334 384 3370 584
rect 3439 368 3475 592
rect 3529 368 3565 592
<< nmoslvt >>
rect 89 119 119 203
rect 167 119 197 203
rect 333 119 363 203
rect 411 119 441 203
rect 547 119 577 203
rect 745 98 775 246
rect 913 98 943 246
rect 1155 125 1185 209
rect 1227 125 1257 209
rect 1318 125 1348 209
rect 1565 125 1595 235
rect 1651 125 1681 235
rect 1772 125 1802 235
rect 1872 125 1902 235
rect 1967 82 1997 192
rect 2217 82 2247 166
rect 2295 82 2325 166
rect 2422 74 2452 222
rect 2526 74 2556 222
rect 2612 74 2642 222
rect 2825 180 2855 264
rect 3031 74 3061 222
rect 3117 74 3147 222
rect 3329 94 3359 222
rect 3449 74 3479 222
rect 3535 74 3565 222
<< ndiff >>
rect 688 234 745 246
rect 32 170 89 203
rect 32 136 44 170
rect 78 136 89 170
rect 32 119 89 136
rect 119 119 167 203
rect 197 175 333 203
rect 197 141 208 175
rect 242 141 288 175
rect 322 141 333 175
rect 197 119 333 141
rect 363 119 411 203
rect 441 169 547 203
rect 441 135 452 169
rect 486 135 547 169
rect 441 119 547 135
rect 577 180 634 203
rect 577 146 588 180
rect 622 146 634 180
rect 577 119 634 146
rect 688 200 700 234
rect 734 200 745 234
rect 688 98 745 200
rect 775 98 913 246
rect 943 237 1000 246
rect 943 203 954 237
rect 988 203 1000 237
rect 943 169 1000 203
rect 943 135 954 169
rect 988 135 1000 169
rect 943 98 1000 135
rect 1078 125 1155 209
rect 1185 125 1227 209
rect 1257 184 1318 209
rect 1257 150 1273 184
rect 1307 150 1318 184
rect 1257 125 1318 150
rect 1348 179 1419 209
rect 1348 145 1373 179
rect 1407 145 1419 179
rect 1348 125 1419 145
rect 1473 125 1565 235
rect 1595 189 1651 235
rect 1595 155 1606 189
rect 1640 155 1651 189
rect 1595 125 1651 155
rect 1681 171 1772 235
rect 1681 137 1716 171
rect 1750 137 1772 171
rect 1681 125 1772 137
rect 1802 171 1872 235
rect 1802 137 1827 171
rect 1861 137 1872 171
rect 1802 125 1872 137
rect 1902 192 1952 235
rect 1902 125 1967 192
rect 1078 118 1140 125
rect 790 82 848 98
rect 790 48 802 82
rect 836 48 848 82
rect 790 36 848 48
rect 1078 84 1092 118
rect 1126 84 1140 118
rect 1078 72 1140 84
rect 1473 119 1550 125
rect 1473 85 1494 119
rect 1528 85 1550 119
rect 1473 73 1550 85
rect 1917 82 1967 125
rect 1997 166 2047 192
rect 2769 251 2825 264
rect 2372 166 2422 222
rect 1997 154 2217 166
rect 1997 120 2008 154
rect 2042 120 2090 154
rect 2124 120 2172 154
rect 2206 120 2217 154
rect 1997 82 2217 120
rect 2247 82 2295 166
rect 2325 86 2422 166
rect 2325 82 2356 86
rect 2340 52 2356 82
rect 2390 74 2422 86
rect 2452 120 2526 222
rect 2452 86 2472 120
rect 2506 86 2526 120
rect 2452 74 2526 86
rect 2556 172 2612 222
rect 2556 138 2567 172
rect 2601 138 2612 172
rect 2556 74 2612 138
rect 2642 99 2715 222
rect 2769 217 2780 251
rect 2814 217 2825 251
rect 2769 180 2825 217
rect 2855 222 2905 264
rect 2855 210 3031 222
rect 2855 180 2986 210
rect 2978 176 2986 180
rect 3020 176 3031 210
rect 2642 74 2669 99
rect 2390 52 2407 74
rect 2340 40 2407 52
rect 2657 65 2669 74
rect 2703 65 2715 99
rect 2978 120 3031 176
rect 2978 86 2986 120
rect 3020 86 3031 120
rect 2978 74 3031 86
rect 3061 210 3117 222
rect 3061 176 3072 210
rect 3106 176 3117 210
rect 3061 120 3117 176
rect 3061 86 3072 120
rect 3106 86 3117 120
rect 3061 74 3117 86
rect 3147 210 3209 222
rect 3147 176 3158 210
rect 3192 176 3209 210
rect 3147 120 3209 176
rect 3147 86 3158 120
rect 3192 86 3209 120
rect 3272 214 3329 222
rect 3272 180 3284 214
rect 3318 180 3329 214
rect 3272 146 3329 180
rect 3272 112 3284 146
rect 3318 112 3329 146
rect 3272 94 3329 112
rect 3359 194 3449 222
rect 3359 160 3390 194
rect 3424 160 3449 194
rect 3359 120 3449 160
rect 3359 94 3390 120
rect 3147 74 3209 86
rect 2657 53 2715 65
rect 3378 86 3390 94
rect 3424 86 3449 120
rect 3378 74 3449 86
rect 3479 194 3535 222
rect 3479 160 3490 194
rect 3524 160 3535 194
rect 3479 120 3535 160
rect 3479 86 3490 120
rect 3524 86 3535 120
rect 3479 74 3535 86
rect 3565 210 3621 222
rect 3565 176 3576 210
rect 3610 176 3621 210
rect 3565 120 3621 176
rect 3565 86 3576 120
rect 3610 86 3621 120
rect 3565 74 3621 86
<< pdiff >>
rect 2860 619 3030 631
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 511 83 546
rect 27 477 39 511
rect 73 477 83 511
rect 27 464 83 477
rect 119 579 173 592
rect 119 545 129 579
rect 163 545 173 579
rect 119 464 173 545
rect 209 464 251 592
rect 287 520 341 592
rect 287 486 297 520
rect 331 486 341 520
rect 287 464 341 486
rect 377 580 433 592
rect 377 546 387 580
rect 421 546 433 580
rect 377 510 433 546
rect 377 476 387 510
rect 421 476 433 510
rect 377 464 433 476
rect 487 580 543 592
rect 487 546 499 580
rect 533 546 543 580
rect 487 510 543 546
rect 487 476 499 510
rect 533 476 543 510
rect 487 464 543 476
rect 579 580 635 592
rect 579 546 589 580
rect 623 546 635 580
rect 579 510 635 546
rect 579 476 589 510
rect 623 476 635 510
rect 579 464 635 476
rect 689 580 745 592
rect 689 546 701 580
rect 735 546 745 580
rect 689 510 745 546
rect 689 476 701 510
rect 735 476 745 510
rect 689 440 745 476
rect 689 406 701 440
rect 735 406 745 440
rect 689 368 745 406
rect 781 580 835 592
rect 781 546 791 580
rect 825 546 835 580
rect 781 502 835 546
rect 781 468 791 502
rect 825 468 835 502
rect 781 368 835 468
rect 871 580 927 592
rect 871 546 881 580
rect 915 546 927 580
rect 1172 548 1228 592
rect 871 499 927 546
rect 871 465 881 499
rect 915 465 927 499
rect 871 418 927 465
rect 981 528 1037 548
rect 981 494 993 528
rect 1027 494 1037 528
rect 981 464 1037 494
rect 1073 464 1121 548
rect 1157 520 1228 548
rect 1157 486 1184 520
rect 1218 486 1228 520
rect 1157 464 1228 486
rect 1264 520 1330 592
rect 1264 486 1284 520
rect 1318 486 1330 520
rect 1264 464 1330 486
rect 1384 580 1559 592
rect 1384 546 1396 580
rect 1430 546 1515 580
rect 1549 546 1559 580
rect 871 384 881 418
rect 915 384 927 418
rect 871 368 927 384
rect 1384 424 1559 546
rect 1595 424 1643 592
rect 1679 543 1751 592
rect 1679 509 1689 543
rect 1723 509 1751 543
rect 1679 424 1751 509
rect 1787 580 1843 592
rect 1787 546 1797 580
rect 1831 546 1843 580
rect 1787 470 1843 546
rect 1787 436 1797 470
rect 1831 436 1843 470
rect 1787 424 1843 436
rect 1897 580 1953 592
rect 1897 546 1909 580
rect 1943 546 1953 580
rect 1897 508 1953 546
rect 1897 474 1909 508
rect 1943 474 1953 508
rect 1897 424 1953 474
rect 1989 424 2031 592
rect 2067 580 2138 592
rect 2067 546 2077 580
rect 2111 546 2138 580
rect 2067 508 2138 546
rect 2174 508 2216 592
rect 2252 575 2308 592
rect 2252 541 2262 575
rect 2296 541 2308 575
rect 2252 508 2308 541
rect 2365 580 2421 592
rect 2365 546 2377 580
rect 2411 546 2421 580
rect 2067 470 2123 508
rect 2067 436 2077 470
rect 2111 436 2123 470
rect 2067 424 2123 436
rect 2365 502 2421 546
rect 2365 468 2377 502
rect 2411 468 2421 502
rect 2365 392 2421 468
rect 2457 575 2523 592
rect 2457 541 2477 575
rect 2511 541 2523 575
rect 2457 392 2523 541
rect 2559 392 2607 592
rect 2643 580 2699 592
rect 2643 546 2653 580
rect 2687 546 2699 580
rect 2860 585 2872 619
rect 2906 585 2984 619
rect 3018 592 3030 619
rect 3018 585 3045 592
rect 2643 462 2699 546
rect 2860 529 3045 585
rect 2860 527 2984 529
rect 2643 428 2653 462
rect 2687 428 2699 462
rect 2643 392 2699 428
rect 2753 451 2809 527
rect 2753 417 2765 451
rect 2799 417 2809 451
rect 2753 399 2809 417
rect 2845 495 2984 527
rect 3018 495 3045 529
rect 2845 447 3045 495
rect 2845 413 2984 447
rect 3018 413 3045 447
rect 2845 399 3045 413
rect 2995 368 3045 399
rect 3081 580 3135 592
rect 3081 546 3091 580
rect 3125 546 3135 580
rect 3081 497 3135 546
rect 3081 463 3091 497
rect 3125 463 3135 497
rect 3081 414 3135 463
rect 3081 380 3091 414
rect 3125 380 3135 414
rect 3081 368 3135 380
rect 3171 580 3225 592
rect 3385 584 3439 592
rect 3171 546 3181 580
rect 3215 546 3225 580
rect 3171 510 3225 546
rect 3171 476 3181 510
rect 3215 476 3225 510
rect 3171 440 3225 476
rect 3171 406 3181 440
rect 3215 406 3225 440
rect 3171 368 3225 406
rect 3279 572 3334 584
rect 3279 538 3290 572
rect 3324 538 3334 572
rect 3279 501 3334 538
rect 3279 467 3290 501
rect 3324 467 3334 501
rect 3279 430 3334 467
rect 3279 396 3290 430
rect 3324 396 3334 430
rect 3279 384 3334 396
rect 3370 576 3439 584
rect 3370 542 3395 576
rect 3429 542 3439 576
rect 3370 498 3439 542
rect 3370 464 3395 498
rect 3429 464 3439 498
rect 3370 426 3439 464
rect 3370 392 3395 426
rect 3429 392 3439 426
rect 3370 384 3439 392
rect 3389 368 3439 384
rect 3475 580 3529 592
rect 3475 546 3485 580
rect 3519 546 3529 580
rect 3475 497 3529 546
rect 3475 463 3485 497
rect 3519 463 3529 497
rect 3475 414 3529 463
rect 3475 380 3485 414
rect 3519 380 3529 414
rect 3475 368 3529 380
rect 3565 580 3621 592
rect 3565 546 3575 580
rect 3609 546 3621 580
rect 3565 497 3621 546
rect 3565 463 3575 497
rect 3609 463 3621 497
rect 3565 414 3621 463
rect 3565 380 3575 414
rect 3609 380 3621 414
rect 3565 368 3621 380
<< ndiffc >>
rect 44 136 78 170
rect 208 141 242 175
rect 288 141 322 175
rect 452 135 486 169
rect 588 146 622 180
rect 700 200 734 234
rect 954 203 988 237
rect 954 135 988 169
rect 1273 150 1307 184
rect 1373 145 1407 179
rect 1606 155 1640 189
rect 1716 137 1750 171
rect 1827 137 1861 171
rect 802 48 836 82
rect 1092 84 1126 118
rect 1494 85 1528 119
rect 2008 120 2042 154
rect 2090 120 2124 154
rect 2172 120 2206 154
rect 2356 52 2390 86
rect 2472 86 2506 120
rect 2567 138 2601 172
rect 2780 217 2814 251
rect 2986 176 3020 210
rect 2669 65 2703 99
rect 2986 86 3020 120
rect 3072 176 3106 210
rect 3072 86 3106 120
rect 3158 176 3192 210
rect 3158 86 3192 120
rect 3284 180 3318 214
rect 3284 112 3318 146
rect 3390 160 3424 194
rect 3390 86 3424 120
rect 3490 160 3524 194
rect 3490 86 3524 120
rect 3576 176 3610 210
rect 3576 86 3610 120
<< pdiffc >>
rect 39 546 73 580
rect 39 477 73 511
rect 129 545 163 579
rect 297 486 331 520
rect 387 546 421 580
rect 387 476 421 510
rect 499 546 533 580
rect 499 476 533 510
rect 589 546 623 580
rect 589 476 623 510
rect 701 546 735 580
rect 701 476 735 510
rect 701 406 735 440
rect 791 546 825 580
rect 791 468 825 502
rect 881 546 915 580
rect 881 465 915 499
rect 993 494 1027 528
rect 1184 486 1218 520
rect 1284 486 1318 520
rect 1396 546 1430 580
rect 1515 546 1549 580
rect 881 384 915 418
rect 1689 509 1723 543
rect 1797 546 1831 580
rect 1797 436 1831 470
rect 1909 546 1943 580
rect 1909 474 1943 508
rect 2077 546 2111 580
rect 2262 541 2296 575
rect 2377 546 2411 580
rect 2077 436 2111 470
rect 2377 468 2411 502
rect 2477 541 2511 575
rect 2653 546 2687 580
rect 2872 585 2906 619
rect 2984 585 3018 619
rect 2653 428 2687 462
rect 2765 417 2799 451
rect 2984 495 3018 529
rect 2984 413 3018 447
rect 3091 546 3125 580
rect 3091 463 3125 497
rect 3091 380 3125 414
rect 3181 546 3215 580
rect 3181 476 3215 510
rect 3181 406 3215 440
rect 3290 538 3324 572
rect 3290 467 3324 501
rect 3290 396 3324 430
rect 3395 542 3429 576
rect 3395 464 3429 498
rect 3395 392 3429 426
rect 3485 546 3519 580
rect 3485 463 3519 497
rect 3485 380 3519 414
rect 3575 546 3609 580
rect 3575 463 3609 497
rect 3575 380 3609 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 251 592 287 618
rect 341 592 377 618
rect 543 592 579 618
rect 745 592 781 618
rect 835 592 871 618
rect 1228 592 1264 618
rect 1559 592 1595 618
rect 1643 592 1679 618
rect 1751 592 1787 618
rect 1953 592 1989 618
rect 2031 592 2067 618
rect 2138 592 2174 618
rect 2216 592 2252 618
rect 2421 592 2457 618
rect 2523 592 2559 618
rect 2607 592 2643 618
rect 83 427 119 464
rect 44 411 119 427
rect 44 377 60 411
rect 94 377 119 411
rect 44 343 119 377
rect 173 359 209 464
rect 251 437 287 464
rect 341 440 377 464
rect 543 440 579 464
rect 251 407 299 437
rect 341 410 441 440
rect 543 410 665 440
rect 44 309 60 343
rect 94 309 119 343
rect 44 275 119 309
rect 44 241 60 275
rect 94 241 119 275
rect 44 225 119 241
rect 161 343 227 359
rect 161 309 177 343
rect 211 309 227 343
rect 161 275 227 309
rect 269 358 299 407
rect 411 362 441 410
rect 269 342 363 358
rect 269 308 313 342
rect 347 308 363 342
rect 269 292 363 308
rect 161 241 177 275
rect 211 241 227 275
rect 161 225 227 241
rect 89 203 119 225
rect 167 203 197 225
rect 333 203 363 292
rect 411 346 587 362
rect 411 332 537 346
rect 411 203 441 332
rect 521 312 537 332
rect 571 312 587 346
rect 521 296 587 312
rect 635 248 665 410
rect 1037 548 1073 574
rect 1121 548 1157 574
rect 1037 432 1073 464
rect 1007 416 1073 432
rect 1007 382 1023 416
rect 1057 382 1073 416
rect 745 336 781 368
rect 713 320 781 336
rect 835 334 871 368
rect 1007 366 1073 382
rect 1121 368 1157 464
rect 1228 449 1264 464
rect 1227 419 1264 449
rect 713 286 729 320
rect 763 286 781 320
rect 713 270 781 286
rect 823 318 943 334
rect 823 284 839 318
rect 873 284 943 318
rect 547 218 665 248
rect 745 246 775 270
rect 823 268 943 284
rect 913 246 943 268
rect 1041 254 1071 366
rect 1119 352 1185 368
rect 1119 318 1135 352
rect 1169 318 1185 352
rect 1119 302 1185 318
rect 547 203 577 218
rect 89 93 119 119
rect 167 51 197 119
rect 333 93 363 119
rect 411 93 441 119
rect 547 51 577 119
rect 1041 224 1185 254
rect 1155 209 1185 224
rect 1227 209 1257 419
rect 1407 375 1473 391
rect 1299 355 1365 371
rect 1299 321 1315 355
rect 1349 321 1365 355
rect 1299 305 1365 321
rect 1407 341 1423 375
rect 1457 341 1473 375
rect 1407 307 1473 341
rect 1318 209 1348 305
rect 1407 273 1423 307
rect 1457 287 1473 307
rect 1559 287 1595 424
rect 1457 273 1595 287
rect 1407 257 1595 273
rect 1643 391 1679 424
rect 1643 375 1709 391
rect 1643 341 1659 375
rect 1693 341 1709 375
rect 1643 307 1709 341
rect 1643 273 1659 307
rect 1693 273 1709 307
rect 1751 356 1787 424
rect 1953 382 1989 424
rect 1872 366 1989 382
rect 1751 340 1824 356
rect 1751 306 1774 340
rect 1808 306 1824 340
rect 1751 290 1824 306
rect 1872 332 1939 366
rect 1973 332 1989 366
rect 1872 316 1989 332
rect 2031 351 2067 424
rect 2138 399 2174 508
rect 2216 476 2252 508
rect 2216 460 2282 476
rect 2216 426 2232 460
rect 2266 440 2282 460
rect 2266 426 2349 440
rect 2216 410 2349 426
rect 2031 335 2097 351
rect 1643 257 1709 273
rect 1565 235 1595 257
rect 1651 235 1681 257
rect 1772 235 1802 290
rect 1872 235 1902 316
rect 2031 301 2047 335
rect 2081 301 2097 335
rect 2031 285 2097 301
rect 2139 237 2169 399
rect 2211 303 2277 319
rect 2211 269 2227 303
rect 2261 269 2277 303
rect 2211 253 2277 269
rect 1967 207 2169 237
rect 1967 192 1997 207
rect 745 72 775 98
rect 167 21 577 51
rect 913 51 943 98
rect 1155 99 1185 125
rect 1227 51 1257 125
rect 1318 99 1348 125
rect 1565 99 1595 125
rect 1651 99 1681 125
rect 1772 99 1802 125
rect 1872 99 1902 125
rect 2217 166 2247 253
rect 2319 211 2349 410
rect 3045 592 3081 618
rect 3135 592 3171 618
rect 2809 527 2845 553
rect 2421 310 2457 392
rect 2523 310 2559 392
rect 2607 360 2643 392
rect 2809 367 2845 399
rect 3334 584 3370 610
rect 3439 592 3475 618
rect 3529 592 3565 618
rect 2607 344 2673 360
rect 2607 310 2623 344
rect 2657 310 2673 344
rect 2391 294 2457 310
rect 2391 260 2407 294
rect 2441 260 2457 294
rect 2391 244 2457 260
rect 2499 294 2565 310
rect 2607 294 2673 310
rect 2789 351 2855 367
rect 2789 317 2805 351
rect 2839 317 2855 351
rect 2789 301 2855 317
rect 2499 260 2515 294
rect 2549 260 2565 294
rect 2499 244 2565 260
rect 2422 222 2452 244
rect 2526 222 2556 244
rect 2612 222 2642 294
rect 2825 264 2855 301
rect 2897 336 2963 352
rect 2897 302 2913 336
rect 2947 329 2963 336
rect 3045 329 3081 368
rect 3135 329 3171 368
rect 3334 330 3370 384
rect 3334 329 3365 330
rect 2947 302 3365 329
rect 3439 310 3475 368
rect 3529 310 3565 368
rect 2897 286 3365 302
rect 3031 270 3365 286
rect 3407 294 3565 310
rect 2295 181 2349 211
rect 2295 166 2325 181
rect 1967 51 1997 82
rect 2217 56 2247 82
rect 2295 56 2325 82
rect 913 21 1997 51
rect 3031 222 3061 270
rect 3117 222 3147 270
rect 3329 222 3359 270
rect 3407 260 3423 294
rect 3457 260 3565 294
rect 3407 244 3565 260
rect 3449 222 3479 244
rect 3535 222 3565 244
rect 2825 154 2855 180
rect 2422 48 2452 74
rect 2526 48 2556 74
rect 2612 48 2642 74
rect 3031 48 3061 74
rect 3117 48 3147 74
rect 3329 68 3359 94
rect 3449 48 3479 74
rect 3535 48 3565 74
<< polycont >>
rect 60 377 94 411
rect 60 309 94 343
rect 60 241 94 275
rect 177 309 211 343
rect 313 308 347 342
rect 177 241 211 275
rect 537 312 571 346
rect 1023 382 1057 416
rect 729 286 763 320
rect 839 284 873 318
rect 1135 318 1169 352
rect 1315 321 1349 355
rect 1423 341 1457 375
rect 1423 273 1457 307
rect 1659 341 1693 375
rect 1659 273 1693 307
rect 1774 306 1808 340
rect 1939 332 1973 366
rect 2232 426 2266 460
rect 2047 301 2081 335
rect 2227 269 2261 303
rect 2623 310 2657 344
rect 2407 260 2441 294
rect 2805 317 2839 351
rect 2515 260 2549 294
rect 2913 302 2947 336
rect 3423 260 3457 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3648 683
rect 23 580 73 596
rect 23 546 39 580
rect 23 511 73 546
rect 113 579 179 649
rect 113 545 129 579
rect 163 545 179 579
rect 113 529 179 545
rect 213 581 437 615
rect 23 477 39 511
rect 213 495 247 581
rect 371 580 437 581
rect 73 477 247 495
rect 23 461 247 477
rect 281 520 331 547
rect 281 486 297 520
rect 281 460 331 486
rect 371 546 387 580
rect 421 546 437 580
rect 371 510 437 546
rect 371 476 387 510
rect 421 476 437 510
rect 371 460 437 476
rect 483 580 549 649
rect 483 546 499 580
rect 533 546 549 580
rect 483 510 549 546
rect 483 476 499 510
rect 533 476 549 510
rect 483 460 549 476
rect 589 580 639 596
rect 623 546 639 580
rect 589 510 639 546
rect 623 476 639 510
rect 25 411 110 427
rect 25 377 60 411
rect 94 377 110 411
rect 297 426 331 460
rect 297 392 431 426
rect 25 343 110 377
rect 25 309 60 343
rect 94 309 110 343
rect 25 275 110 309
rect 25 241 60 275
rect 94 241 110 275
rect 25 225 110 241
rect 161 343 263 359
rect 161 309 177 343
rect 211 309 263 343
rect 161 275 263 309
rect 297 342 363 358
rect 297 308 313 342
rect 347 308 363 342
rect 297 292 363 308
rect 161 241 177 275
rect 211 241 263 275
rect 397 258 431 392
rect 589 362 639 476
rect 685 580 735 596
rect 685 546 701 580
rect 685 510 735 546
rect 685 476 701 510
rect 685 440 735 476
rect 775 580 841 649
rect 775 546 791 580
rect 825 546 841 580
rect 775 502 841 546
rect 775 468 791 502
rect 825 468 841 502
rect 775 458 841 468
rect 881 580 957 596
rect 915 546 957 580
rect 881 499 957 546
rect 915 465 957 499
rect 993 528 1043 649
rect 1027 494 1043 528
rect 993 470 1043 494
rect 1077 581 1565 615
rect 685 406 701 440
rect 735 406 847 424
rect 685 390 847 406
rect 521 346 639 362
rect 521 312 537 346
rect 571 312 639 346
rect 521 296 639 312
rect 161 225 263 241
rect 297 224 554 258
rect 297 191 338 224
rect 28 170 94 191
rect 28 136 44 170
rect 78 136 94 170
rect 28 17 94 136
rect 192 175 338 191
rect 192 141 208 175
rect 242 141 288 175
rect 322 141 338 175
rect 192 125 338 141
rect 436 169 486 190
rect 436 135 452 169
rect 436 17 486 135
rect 520 85 554 224
rect 588 180 639 296
rect 697 320 779 356
rect 697 286 729 320
rect 763 286 779 320
rect 697 270 779 286
rect 813 334 847 390
rect 881 418 957 465
rect 1077 436 1111 581
rect 1380 580 1565 581
rect 915 384 957 418
rect 881 368 957 384
rect 813 318 889 334
rect 813 284 839 318
rect 873 284 889 318
rect 813 268 889 284
rect 923 270 957 368
rect 1007 416 1111 436
rect 1007 382 1023 416
rect 1057 402 1111 416
rect 1168 520 1234 547
rect 1168 486 1184 520
rect 1218 486 1234 520
rect 1168 442 1234 486
rect 1268 520 1334 547
rect 1380 546 1396 580
rect 1430 546 1515 580
rect 1549 546 1609 580
rect 1268 486 1284 520
rect 1318 510 1334 520
rect 1318 486 1541 510
rect 1268 476 1541 486
rect 1168 408 1473 442
rect 1057 382 1073 402
rect 1007 366 1073 382
rect 1407 375 1473 408
rect 1299 368 1365 371
rect 1119 355 1365 368
rect 1119 352 1315 355
rect 1119 318 1135 352
rect 1169 321 1315 352
rect 1349 321 1365 355
rect 1169 318 1365 321
rect 1119 305 1365 318
rect 1407 341 1423 375
rect 1457 341 1473 375
rect 1407 307 1473 341
rect 1119 276 1223 305
rect 1119 270 1183 276
rect 813 234 847 268
rect 923 242 1183 270
rect 1217 242 1223 276
rect 1407 273 1423 307
rect 1457 273 1473 307
rect 1407 271 1473 273
rect 923 237 1223 242
rect 923 236 954 237
rect 684 200 700 234
rect 734 200 847 234
rect 938 203 954 236
rect 988 236 1223 237
rect 1257 237 1473 271
rect 622 146 639 180
rect 938 169 988 203
rect 588 119 639 146
rect 673 132 904 166
rect 673 85 707 132
rect 520 51 707 85
rect 786 82 836 98
rect 786 48 802 82
rect 870 85 904 132
rect 938 135 954 169
rect 938 119 988 135
rect 1022 168 1223 202
rect 1022 85 1056 168
rect 870 51 1056 85
rect 1090 118 1144 134
rect 1090 84 1092 118
rect 1126 84 1144 118
rect 786 17 836 48
rect 1090 17 1144 84
rect 1189 87 1223 168
rect 1257 184 1323 237
rect 1507 203 1541 476
rect 1257 150 1273 184
rect 1307 150 1323 184
rect 1257 121 1323 150
rect 1357 179 1541 203
rect 1575 459 1609 546
rect 1673 543 1739 649
rect 1673 509 1689 543
rect 1723 509 1739 543
rect 1673 493 1739 509
rect 1781 580 1847 596
rect 1781 546 1797 580
rect 1831 546 1847 580
rect 1781 470 1847 546
rect 1781 459 1797 470
rect 1575 436 1797 459
rect 1831 436 1847 470
rect 1893 580 1959 649
rect 1893 546 1909 580
rect 1943 546 1959 580
rect 1893 508 1959 546
rect 1893 474 1909 508
rect 1943 474 1959 508
rect 1893 458 1959 474
rect 2061 580 2127 596
rect 2061 546 2077 580
rect 2111 546 2127 580
rect 2061 470 2127 546
rect 2246 575 2312 649
rect 2246 541 2262 575
rect 2296 541 2312 575
rect 2246 520 2312 541
rect 2361 580 2427 596
rect 2361 546 2377 580
rect 2411 546 2427 580
rect 2361 502 2427 546
rect 2461 575 2527 649
rect 2856 619 3034 649
rect 2461 541 2477 575
rect 2511 541 2527 575
rect 2461 520 2527 541
rect 2637 580 2687 596
rect 2637 546 2653 580
rect 2856 585 2872 619
rect 2906 585 2984 619
rect 3018 585 3034 619
rect 2856 569 3034 585
rect 2637 535 2687 546
rect 2361 486 2377 502
rect 1575 425 1847 436
rect 1575 223 1609 425
rect 1781 424 1847 425
rect 2061 436 2077 470
rect 2111 454 2127 470
rect 2216 468 2377 486
rect 2411 486 2427 502
rect 2637 501 2931 535
rect 2637 486 2687 501
rect 2411 468 2687 486
rect 2216 462 2687 468
rect 2216 460 2653 462
rect 2111 436 2182 454
rect 1643 375 1724 391
rect 1781 390 1989 424
rect 2061 420 2182 436
rect 1643 341 1659 375
rect 1693 341 1724 375
rect 1923 366 1989 390
rect 1643 307 1724 341
rect 1643 273 1659 307
rect 1693 273 1724 307
rect 1758 350 1889 356
rect 1758 340 1855 350
rect 1758 306 1774 340
rect 1808 316 1855 340
rect 1923 332 1939 366
rect 1973 332 1989 366
rect 2148 384 2182 420
rect 2216 426 2232 460
rect 2266 452 2653 460
rect 2266 426 2282 452
rect 2216 418 2282 426
rect 2637 428 2653 452
rect 2316 384 2533 418
rect 2637 412 2687 428
rect 2721 451 2815 467
rect 2721 417 2765 451
rect 2799 417 2815 451
rect 1923 316 1989 332
rect 2031 335 2097 351
rect 2148 350 2350 384
rect 2499 378 2533 384
rect 2721 401 2815 417
rect 1808 306 1889 316
rect 1758 290 1889 306
rect 2031 301 2047 335
rect 2081 316 2097 335
rect 2081 303 2277 316
rect 2081 301 2227 303
rect 1643 257 1724 273
rect 1690 256 1724 257
rect 2031 276 2227 301
rect 1575 189 1656 223
rect 1690 222 1945 256
rect 2031 242 2047 276
rect 2081 269 2227 276
rect 2261 269 2277 303
rect 2081 256 2277 269
rect 2081 242 2097 256
rect 2031 236 2097 242
rect 2311 222 2345 350
rect 2391 316 2431 350
rect 2499 344 2673 378
rect 2391 294 2465 316
rect 2607 310 2623 344
rect 2657 310 2673 344
rect 2391 260 2407 294
rect 2441 260 2465 294
rect 2391 236 2465 260
rect 2499 294 2565 310
rect 2607 294 2673 310
rect 2499 260 2515 294
rect 2549 260 2565 294
rect 2721 267 2755 401
rect 2789 351 2855 367
rect 2789 317 2805 351
rect 2839 317 2855 351
rect 2789 301 2855 317
rect 2897 352 2931 501
rect 2965 529 3034 569
rect 2965 495 2984 529
rect 3018 495 3034 529
rect 2965 447 3034 495
rect 2965 413 2984 447
rect 3018 413 3034 447
rect 2965 390 3034 413
rect 3075 580 3125 596
rect 3075 546 3091 580
rect 3075 497 3125 546
rect 3075 463 3091 497
rect 3075 414 3125 463
rect 3075 380 3091 414
rect 3165 580 3231 649
rect 3165 546 3181 580
rect 3215 546 3231 580
rect 3165 510 3231 546
rect 3165 476 3181 510
rect 3215 476 3231 510
rect 3165 440 3231 476
rect 3165 406 3181 440
rect 3215 406 3231 440
rect 3165 390 3231 406
rect 3268 572 3340 588
rect 3268 538 3290 572
rect 3324 538 3340 572
rect 3268 501 3340 538
rect 3268 467 3290 501
rect 3324 467 3340 501
rect 3268 430 3340 467
rect 3268 396 3290 430
rect 3324 396 3340 430
rect 3075 356 3125 380
rect 2897 336 2963 352
rect 2897 302 2913 336
rect 2947 302 2963 336
rect 2897 286 2963 302
rect 3075 310 3143 356
rect 3268 310 3340 396
rect 3379 576 3445 649
rect 3379 542 3395 576
rect 3429 542 3445 576
rect 3379 498 3445 542
rect 3379 464 3395 498
rect 3429 464 3445 498
rect 3379 426 3445 464
rect 3379 392 3395 426
rect 3429 392 3445 426
rect 3379 364 3445 392
rect 3479 580 3541 596
rect 3479 546 3485 580
rect 3519 546 3541 580
rect 3479 497 3541 546
rect 3479 463 3485 497
rect 3519 463 3541 497
rect 3479 414 3541 463
rect 3479 380 3485 414
rect 3519 380 3541 414
rect 3479 364 3541 380
rect 3575 580 3625 649
rect 3609 546 3625 580
rect 3575 497 3625 546
rect 3609 463 3625 497
rect 3575 414 3625 463
rect 3609 380 3625 414
rect 3575 364 3625 380
rect 2721 260 2830 267
rect 2499 251 2830 260
rect 1357 145 1373 179
rect 1407 169 1541 179
rect 1407 145 1423 169
rect 1357 87 1423 145
rect 1590 155 1606 189
rect 1640 155 1656 189
rect 1189 53 1423 87
rect 1469 119 1554 135
rect 1590 121 1656 155
rect 1690 171 1777 187
rect 1690 137 1716 171
rect 1750 137 1777 171
rect 1690 121 1777 137
rect 1811 171 1877 188
rect 1811 137 1827 171
rect 1861 137 1877 171
rect 1469 85 1494 119
rect 1528 87 1554 119
rect 1690 87 1724 121
rect 1528 85 1724 87
rect 1469 53 1724 85
rect 1811 17 1877 137
rect 1911 86 1945 222
rect 2188 188 2345 222
rect 2499 226 2780 251
rect 2499 188 2533 226
rect 2721 217 2780 226
rect 2814 217 2830 251
rect 2721 201 2830 217
rect 2897 201 2931 286
rect 3075 244 3122 310
rect 2188 170 2222 188
rect 1992 154 2222 170
rect 2379 154 2533 188
rect 2567 172 2617 192
rect 1992 120 2008 154
rect 2042 120 2090 154
rect 2124 120 2172 154
rect 2206 120 2222 154
rect 2268 120 2413 154
rect 2601 167 2617 172
rect 2864 167 2931 201
rect 2965 210 3022 226
rect 2965 176 2986 210
rect 3020 176 3022 210
rect 2601 138 2898 167
rect 2567 133 2898 138
rect 2268 86 2302 120
rect 2447 86 2472 120
rect 2506 86 2531 120
rect 2567 119 2617 133
rect 2965 120 3022 176
rect 1911 52 2302 86
rect 2336 52 2356 86
rect 2390 52 2411 86
rect 2336 17 2411 52
rect 2447 85 2531 86
rect 2653 85 2669 99
rect 2447 65 2669 85
rect 2703 65 2719 99
rect 2447 51 2719 65
rect 2965 86 2986 120
rect 3020 86 3022 120
rect 2965 17 3022 86
rect 3056 210 3122 244
rect 3268 294 3473 310
rect 3268 260 3423 294
rect 3457 260 3473 294
rect 3268 244 3473 260
rect 3056 176 3072 210
rect 3106 176 3122 210
rect 3056 120 3122 176
rect 3056 86 3072 120
rect 3106 86 3122 120
rect 3056 70 3122 86
rect 3156 210 3222 226
rect 3156 176 3158 210
rect 3192 176 3222 210
rect 3156 120 3222 176
rect 3156 86 3158 120
rect 3192 86 3222 120
rect 3268 214 3334 244
rect 3268 180 3284 214
rect 3318 180 3334 214
rect 3507 210 3541 364
rect 3268 146 3334 180
rect 3268 112 3284 146
rect 3318 112 3334 146
rect 3268 108 3334 112
rect 3374 194 3440 210
rect 3374 160 3390 194
rect 3424 160 3440 194
rect 3374 120 3440 160
rect 3156 17 3222 86
rect 3374 86 3390 120
rect 3424 86 3440 120
rect 3374 17 3440 86
rect 3474 194 3541 210
rect 3474 160 3490 194
rect 3524 160 3541 194
rect 3474 120 3541 160
rect 3474 86 3490 120
rect 3524 86 3541 120
rect 3474 70 3541 86
rect 3576 210 3626 226
rect 3610 176 3626 210
rect 3576 120 3626 176
rect 3610 86 3626 120
rect 3576 17 3626 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3648 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 3583 649 3617 683
rect 1183 242 1217 276
rect 1855 316 1889 350
rect 2047 242 2081 276
rect 2431 316 2465 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
<< metal1 >>
rect 0 683 3648 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3648 683
rect 0 617 3648 649
rect 1843 350 1901 356
rect 1843 316 1855 350
rect 1889 347 1901 350
rect 2419 350 2477 356
rect 2419 347 2431 350
rect 1889 319 2431 347
rect 1889 316 1901 319
rect 1843 310 1901 316
rect 2419 316 2431 319
rect 2465 316 2477 350
rect 2419 310 2477 316
rect 1171 276 1229 282
rect 1171 242 1183 276
rect 1217 273 1229 276
rect 2035 276 2093 282
rect 2035 273 2047 276
rect 1217 245 2047 273
rect 1217 242 1229 245
rect 1171 236 1229 242
rect 2035 242 2047 245
rect 2081 242 2093 276
rect 2035 236 2093 242
rect 0 17 3648 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3648 17
rect 0 -49 3648 -17
<< labels >>
flabel pwell s 0 0 3648 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 3648 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfbbn_2
flabel metal1 s 2431 316 2465 350 0 FreeSans 340 0 0 0 SET_B
port 6 nsew signal input
flabel metal1 s 0 617 3648 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 3648 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 3103 316 3137 350 0 FreeSans 340 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 3487 390 3521 424 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 2815 316 2849 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3648 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 1787922
string GDS_START 1762592
<< end >>
