magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1265 -1309 2225 2641
<< nwell >>
rect -5 997 965 1370
rect -5 -38 965 335
<< pwell >>
rect 5 912 91 921
rect 869 912 955 921
rect 5 692 955 912
rect 5 420 357 692
rect 5 411 91 420
rect 869 411 955 692
<< scnmos >>
rect 246 718 276 886
rect 318 718 348 886
rect 404 718 434 886
rect 476 718 506 886
rect 682 718 712 886
rect 754 718 784 886
rect 176 446 206 530
rect 248 446 278 530
<< scpmoshvt >>
rect 246 1085 276 1285
rect 318 1085 348 1285
rect 404 1085 434 1285
rect 476 1085 506 1285
rect 682 1085 712 1285
rect 754 1085 784 1285
rect 176 47 206 247
rect 248 47 278 247
<< ndiff >>
rect 193 874 246 886
rect 193 840 201 874
rect 235 840 246 874
rect 193 767 246 840
rect 193 733 201 767
rect 235 733 246 767
rect 193 718 246 733
rect 276 718 318 886
rect 348 878 404 886
rect 348 844 359 878
rect 393 844 404 878
rect 348 760 404 844
rect 348 726 359 760
rect 393 726 404 760
rect 348 718 404 726
rect 434 718 476 886
rect 506 872 563 886
rect 506 838 517 872
rect 551 838 563 872
rect 506 760 563 838
rect 506 726 517 760
rect 551 726 563 760
rect 506 718 563 726
rect 625 846 682 886
rect 625 812 637 846
rect 671 812 682 846
rect 625 760 682 812
rect 625 726 637 760
rect 671 726 682 760
rect 625 718 682 726
rect 712 718 754 886
rect 784 874 837 886
rect 784 840 795 874
rect 829 840 837 874
rect 784 764 837 840
rect 784 730 795 764
rect 829 730 837 764
rect 784 718 837 730
rect 123 505 176 530
rect 123 471 131 505
rect 165 471 176 505
rect 123 446 176 471
rect 206 446 248 530
rect 278 505 331 530
rect 278 471 289 505
rect 323 471 331 505
rect 278 446 331 471
<< pdiff >>
rect 193 1273 246 1285
rect 193 1239 201 1273
rect 235 1239 246 1273
rect 193 1199 246 1239
rect 193 1165 201 1199
rect 235 1165 246 1199
rect 193 1131 246 1165
rect 193 1097 201 1131
rect 235 1097 246 1131
rect 193 1085 246 1097
rect 276 1085 318 1285
rect 348 1277 404 1285
rect 348 1243 359 1277
rect 393 1243 404 1277
rect 348 1173 404 1243
rect 348 1139 359 1173
rect 393 1139 404 1173
rect 348 1085 404 1139
rect 434 1085 476 1285
rect 506 1277 563 1285
rect 506 1243 517 1277
rect 551 1243 563 1277
rect 506 1195 563 1243
rect 506 1161 517 1195
rect 551 1161 563 1195
rect 506 1127 563 1161
rect 506 1093 517 1127
rect 551 1093 563 1127
rect 506 1085 563 1093
rect 625 1277 682 1285
rect 625 1243 637 1277
rect 671 1243 682 1277
rect 625 1202 682 1243
rect 625 1168 637 1202
rect 671 1168 682 1202
rect 625 1134 682 1168
rect 625 1100 637 1134
rect 671 1100 682 1134
rect 625 1085 682 1100
rect 712 1085 754 1285
rect 784 1273 837 1285
rect 784 1239 795 1273
rect 829 1239 837 1273
rect 784 1202 837 1239
rect 784 1168 795 1202
rect 829 1168 837 1202
rect 784 1131 837 1168
rect 784 1097 795 1131
rect 829 1097 837 1131
rect 784 1085 837 1097
rect 123 235 176 247
rect 123 201 131 235
rect 165 201 176 235
rect 123 164 176 201
rect 123 130 131 164
rect 165 130 176 164
rect 123 93 176 130
rect 123 59 131 93
rect 165 59 176 93
rect 123 47 176 59
rect 206 47 248 247
rect 278 235 331 247
rect 278 201 289 235
rect 323 201 331 235
rect 278 164 331 201
rect 278 130 289 164
rect 323 130 331 164
rect 278 93 331 130
rect 278 59 289 93
rect 323 59 331 93
rect 278 47 331 59
<< ndiffc >>
rect 201 840 235 874
rect 201 733 235 767
rect 359 844 393 878
rect 359 726 393 760
rect 517 838 551 872
rect 517 726 551 760
rect 637 812 671 846
rect 637 726 671 760
rect 795 840 829 874
rect 795 730 829 764
rect 131 471 165 505
rect 289 471 323 505
<< pdiffc >>
rect 201 1239 235 1273
rect 201 1165 235 1199
rect 201 1097 235 1131
rect 359 1243 393 1277
rect 359 1139 393 1173
rect 517 1243 551 1277
rect 517 1161 551 1195
rect 517 1093 551 1127
rect 637 1243 671 1277
rect 637 1168 671 1202
rect 637 1100 671 1134
rect 795 1239 829 1273
rect 795 1168 829 1202
rect 795 1097 829 1131
rect 131 201 165 235
rect 131 130 165 164
rect 131 59 165 93
rect 289 201 323 235
rect 289 130 323 164
rect 289 59 323 93
<< psubdiff >>
rect 31 871 65 895
rect 31 788 65 837
rect 31 730 65 754
rect 895 871 929 895
rect 895 788 929 837
rect 895 730 929 754
rect 31 578 65 602
rect 31 495 65 544
rect 895 578 929 602
rect 31 437 65 461
rect 895 495 929 544
rect 895 437 929 461
<< nsubdiff >>
rect 31 1244 65 1268
rect 31 1157 65 1210
rect 31 1099 65 1123
rect 895 1244 929 1268
rect 895 1157 929 1210
rect 895 1099 929 1123
rect 31 209 65 233
rect 31 122 65 175
rect 31 64 65 88
rect 895 209 929 233
rect 895 122 929 175
rect 895 64 929 88
<< psubdiffcont >>
rect 31 837 65 871
rect 31 754 65 788
rect 895 837 929 871
rect 895 754 929 788
rect 31 544 65 578
rect 895 544 929 578
rect 31 461 65 495
rect 895 461 929 495
<< nsubdiffcont >>
rect 31 1210 65 1244
rect 31 1123 65 1157
rect 895 1210 929 1244
rect 895 1123 929 1157
rect 31 175 65 209
rect 31 88 65 122
rect 895 175 929 209
rect 895 88 929 122
<< poly >>
rect 246 1285 276 1311
rect 318 1285 348 1311
rect 404 1285 434 1311
rect 476 1285 506 1311
rect 682 1285 712 1311
rect 754 1285 784 1311
rect 246 1053 276 1085
rect 318 1053 348 1085
rect 404 1070 434 1085
rect 476 1070 506 1085
rect 404 1053 636 1070
rect 246 1037 348 1053
rect 246 1003 286 1037
rect 320 1003 348 1037
rect 246 987 348 1003
rect 390 1040 636 1053
rect 390 1037 456 1040
rect 390 1003 406 1037
rect 440 1003 456 1037
rect 390 987 456 1003
rect 606 1017 636 1040
rect 682 1017 712 1085
rect 754 1017 784 1085
rect 498 982 564 998
rect 606 987 784 1017
rect 498 948 514 982
rect 548 948 564 982
rect 498 938 564 948
rect 404 932 564 938
rect 246 886 276 912
rect 318 886 348 912
rect 404 908 528 932
rect 404 886 434 908
rect 476 886 506 908
rect 682 886 712 987
rect 754 886 784 987
rect 246 618 276 718
rect 318 618 348 718
rect 404 692 434 718
rect 476 692 506 718
rect 682 692 712 718
rect 754 692 784 718
rect 246 602 382 618
rect 246 598 264 602
rect 248 568 264 598
rect 298 568 332 602
rect 366 568 382 602
rect 176 530 206 556
rect 248 552 382 568
rect 248 530 278 552
rect 176 426 206 446
rect 248 426 278 446
rect 117 408 278 426
rect 117 374 133 408
rect 167 374 201 408
rect 235 374 278 408
rect 117 358 278 374
rect 176 247 206 358
rect 248 247 278 358
rect 176 21 206 47
rect 248 21 278 47
<< polycont >>
rect 286 1003 320 1037
rect 406 1003 440 1037
rect 514 948 548 982
rect 264 568 298 602
rect 332 568 366 602
rect 133 374 167 408
rect 201 374 235 408
<< locali >>
rect 0 1315 31 1349
rect 65 1315 127 1349
rect 161 1315 223 1349
rect 257 1315 319 1349
rect 353 1315 415 1349
rect 449 1315 511 1349
rect 545 1315 607 1349
rect 641 1315 703 1349
rect 737 1315 799 1349
rect 833 1315 895 1349
rect 929 1315 960 1349
rect 18 1244 78 1279
rect 18 1210 31 1244
rect 65 1210 78 1244
rect 18 1157 78 1210
rect 18 1123 31 1157
rect 65 1123 78 1157
rect 18 1044 78 1123
rect 185 1273 255 1281
rect 185 1239 201 1273
rect 235 1239 255 1273
rect 185 1199 255 1239
rect 185 1165 201 1199
rect 235 1165 255 1199
rect 185 1131 255 1165
rect 343 1277 409 1315
rect 343 1243 359 1277
rect 393 1243 409 1277
rect 343 1173 409 1243
rect 343 1139 359 1173
rect 393 1139 409 1173
rect 501 1277 567 1279
rect 501 1243 517 1277
rect 551 1243 567 1277
rect 501 1195 567 1243
rect 501 1161 517 1195
rect 551 1161 567 1195
rect 185 1097 201 1131
rect 235 1097 255 1131
rect 501 1127 567 1161
rect 501 1105 517 1127
rect 185 1087 255 1097
rect 302 1093 517 1105
rect 551 1093 567 1127
rect 621 1277 687 1315
rect 621 1243 637 1277
rect 671 1243 687 1277
rect 621 1202 687 1243
rect 621 1168 637 1202
rect 671 1168 687 1202
rect 621 1134 687 1168
rect 621 1100 637 1134
rect 671 1100 687 1134
rect 779 1273 845 1281
rect 779 1239 795 1273
rect 829 1239 845 1273
rect 779 1202 845 1239
rect 779 1168 795 1202
rect 829 1168 845 1202
rect 779 1131 845 1168
rect 185 964 236 1087
rect 302 1071 567 1093
rect 302 1053 336 1071
rect 270 1037 336 1053
rect 533 1066 567 1071
rect 779 1097 795 1131
rect 829 1097 845 1131
rect 270 1003 286 1037
rect 320 1003 336 1037
rect 270 998 336 1003
rect 374 1003 406 1037
rect 440 1003 456 1037
rect 533 1032 632 1066
rect 374 1002 456 1003
rect 374 964 408 1002
rect 490 982 564 998
rect 490 968 514 982
rect 18 871 78 954
rect 18 837 31 871
rect 65 837 78 871
rect 18 788 78 837
rect 18 754 31 788
rect 65 754 78 788
rect 18 683 78 754
rect 185 930 408 964
rect 442 948 514 968
rect 548 948 564 982
rect 185 874 241 930
rect 442 922 519 948
rect 442 896 476 922
rect 598 914 632 1032
rect 185 840 201 874
rect 235 840 241 874
rect 185 767 241 840
rect 185 733 201 767
rect 235 733 241 767
rect 185 717 241 733
rect 343 878 399 896
rect 343 844 359 878
rect 393 844 399 878
rect 343 760 399 844
rect 343 726 359 760
rect 393 726 399 760
rect 343 683 399 726
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 399 683
rect 433 862 476 896
rect 553 888 632 914
rect 510 880 632 888
rect 510 872 587 880
rect 18 578 78 649
rect 18 544 31 578
rect 65 544 78 578
rect 18 495 78 544
rect 18 461 31 495
rect 65 461 78 495
rect 115 505 181 649
rect 115 471 131 505
rect 165 471 181 505
rect 115 461 181 471
rect 215 602 382 615
rect 215 568 264 602
rect 298 568 332 602
rect 366 568 382 602
rect 215 555 382 568
rect 18 378 78 461
rect 215 427 249 555
rect 433 521 467 862
rect 510 838 517 872
rect 551 838 587 872
rect 779 874 845 1097
rect 882 1244 942 1279
rect 882 1210 895 1244
rect 929 1210 942 1244
rect 882 1157 942 1210
rect 882 1123 895 1157
rect 929 1123 942 1157
rect 882 1044 942 1123
rect 510 828 587 838
rect 501 760 587 828
rect 501 726 517 760
rect 551 726 587 760
rect 501 717 587 726
rect 621 812 637 846
rect 671 812 687 846
rect 621 760 687 812
rect 621 726 637 760
rect 671 726 687 760
rect 621 683 687 726
rect 779 840 795 874
rect 829 840 845 874
rect 779 764 845 840
rect 779 730 795 764
rect 829 730 845 764
rect 779 717 845 730
rect 882 871 942 954
rect 882 837 895 871
rect 929 837 942 871
rect 882 788 942 837
rect 882 754 895 788
rect 929 754 942 788
rect 882 683 942 754
rect 501 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 117 408 249 427
rect 117 374 133 408
rect 167 374 201 408
rect 235 374 249 408
rect 117 306 249 374
rect 283 505 467 521
rect 283 471 289 505
rect 323 487 467 505
rect 882 578 942 649
rect 882 544 895 578
rect 929 544 942 578
rect 882 495 942 544
rect 323 471 343 487
rect 18 209 78 288
rect 283 272 343 471
rect 882 461 895 495
rect 929 461 942 495
rect 882 378 942 461
rect 273 235 343 272
rect 18 175 31 209
rect 65 175 78 209
rect 18 122 78 175
rect 18 88 31 122
rect 65 88 78 122
rect 18 53 78 88
rect 115 201 131 235
rect 165 201 181 235
rect 115 164 181 201
rect 115 130 131 164
rect 165 130 181 164
rect 115 93 181 130
rect 115 59 131 93
rect 165 59 181 93
rect 115 17 181 59
rect 273 201 289 235
rect 323 201 343 235
rect 273 164 343 201
rect 273 130 289 164
rect 323 130 343 164
rect 273 93 343 130
rect 273 59 289 93
rect 323 59 343 93
rect 273 53 343 59
rect 882 209 942 288
rect 882 175 895 209
rect 929 175 942 209
rect 882 122 942 175
rect 882 88 895 122
rect 929 88 942 122
rect 882 53 942 88
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 1315 65 1349
rect 127 1315 161 1349
rect 223 1315 257 1349
rect 319 1315 353 1349
rect 415 1315 449 1349
rect 511 1315 545 1349
rect 607 1315 641 1349
rect 703 1315 737 1349
rect 799 1315 833 1349
rect 895 1315 929 1349
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 1349 960 1381
rect 0 1315 31 1349
rect 65 1315 127 1349
rect 161 1315 223 1349
rect 257 1315 319 1349
rect 353 1315 415 1349
rect 449 1315 511 1349
rect 545 1315 607 1349
rect 641 1315 703 1349
rect 737 1315 799 1349
rect 833 1315 895 1349
rect 929 1315 960 1349
rect 0 1283 960 1315
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel locali s 799 760 833 794 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 799 834 833 868 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 799 1130 833 1164 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 799 1056 833 1090 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 799 982 833 1016 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 799 908 833 942 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 128 316 162 350 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 31 1204 65 1238 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
flabel locali s 31 1130 65 1164 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
flabel locali s 895 94 929 128 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 895 1204 929 1238 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
flabel locali s 895 1130 929 1164 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
flabel locali s 895 1056 929 1090 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 31 1056 65 1090 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
rlabel comment s 0 0 0 0 4 lsbuf_lp
flabel metal1 s 0 0 960 49 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 1283 960 1332 0 FreeSans 200 0 0 0 DESTPWR
port 2 nsew power bidirectional
flabel metal1 s 0 617 960 715 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 1332
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 474048
string GDS_START 460884
<< end >>
