magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
rect 261 309 1089 331
rect 764 307 1089 309
<< pwell >>
rect 1397 211 2017 241
rect 272 183 382 211
rect 836 183 2017 211
rect 272 167 2017 183
rect 1 49 2017 167
rect 0 0 2112 49
<< scnmos >>
rect 84 57 114 141
rect 156 57 186 141
rect 378 73 408 157
rect 450 73 480 157
rect 536 73 566 157
rect 608 73 638 157
rect 942 101 972 185
rect 1028 101 1058 185
rect 1106 101 1136 185
rect 1208 101 1238 185
rect 1480 47 1510 215
rect 1558 47 1588 215
rect 1827 47 1857 215
rect 1899 47 1929 215
<< scpmoshvt >>
rect 84 470 114 598
rect 156 470 186 598
rect 354 345 384 473
rect 456 345 486 473
rect 587 345 617 473
rect 659 345 689 473
rect 857 343 887 471
rect 966 343 996 427
rect 1164 387 1194 515
rect 1273 387 1303 471
rect 1477 367 1507 619
rect 1563 367 1593 619
rect 1635 367 1665 619
rect 1721 367 1751 619
rect 1919 367 1949 619
rect 1997 367 2027 619
<< ndiff >>
rect 298 173 356 185
rect 27 116 84 141
rect 27 82 39 116
rect 73 82 84 116
rect 27 57 84 82
rect 114 57 156 141
rect 186 116 243 141
rect 186 82 197 116
rect 231 82 243 116
rect 186 57 243 82
rect 298 139 310 173
rect 344 157 356 173
rect 862 160 942 185
rect 344 139 378 157
rect 298 73 378 139
rect 408 73 450 157
rect 480 123 536 157
rect 480 89 491 123
rect 525 89 536 123
rect 480 73 536 89
rect 566 73 608 157
rect 638 123 695 157
rect 638 89 649 123
rect 683 89 695 123
rect 862 126 874 160
rect 908 126 942 160
rect 862 101 942 126
rect 972 173 1028 185
rect 972 139 983 173
rect 1017 139 1028 173
rect 972 101 1028 139
rect 1058 101 1106 185
rect 1136 147 1208 185
rect 1136 113 1147 147
rect 1181 113 1208 147
rect 1136 101 1208 113
rect 1238 160 1295 185
rect 1238 126 1249 160
rect 1283 126 1295 160
rect 1238 101 1295 126
rect 638 73 695 89
rect 1423 125 1480 215
rect 1423 91 1435 125
rect 1469 91 1480 125
rect 1423 47 1480 91
rect 1510 47 1558 215
rect 1588 93 1827 215
rect 1588 59 1599 93
rect 1633 59 1827 93
rect 1588 47 1827 59
rect 1857 47 1899 215
rect 1929 203 1991 215
rect 1929 169 1945 203
rect 1979 169 1991 203
rect 1929 103 1991 169
rect 1929 69 1945 103
rect 1979 69 1991 103
rect 1929 47 1991 69
<< pdiff >>
rect 27 586 84 598
rect 27 552 39 586
rect 73 552 84 586
rect 27 516 84 552
rect 27 482 39 516
rect 73 482 84 516
rect 27 470 84 482
rect 114 470 156 598
rect 186 586 243 598
rect 186 552 197 586
rect 231 552 243 586
rect 186 516 243 552
rect 186 482 197 516
rect 231 482 243 516
rect 186 470 243 482
rect 297 461 354 473
rect 297 427 309 461
rect 343 427 354 461
rect 297 391 354 427
rect 297 357 309 391
rect 343 357 354 391
rect 297 345 354 357
rect 384 345 456 473
rect 486 449 587 473
rect 486 415 497 449
rect 531 415 587 449
rect 486 345 587 415
rect 617 345 659 473
rect 689 461 746 473
rect 689 427 700 461
rect 734 427 746 461
rect 689 391 746 427
rect 689 357 700 391
rect 734 357 746 391
rect 689 345 746 357
rect 800 430 857 471
rect 800 396 812 430
rect 846 396 857 430
rect 800 343 857 396
rect 887 427 944 471
rect 1420 597 1477 619
rect 1420 563 1432 597
rect 1466 563 1477 597
rect 1107 477 1164 515
rect 1107 443 1119 477
rect 1153 443 1164 477
rect 887 407 966 427
rect 887 373 898 407
rect 932 373 966 407
rect 887 343 966 373
rect 996 402 1053 427
rect 996 368 1007 402
rect 1041 368 1053 402
rect 1107 387 1164 443
rect 1194 481 1251 515
rect 1420 505 1477 563
rect 1194 447 1205 481
rect 1239 471 1251 481
rect 1420 471 1432 505
rect 1466 471 1477 505
rect 1239 447 1273 471
rect 1194 387 1273 447
rect 1303 446 1360 471
rect 1303 412 1314 446
rect 1348 412 1360 446
rect 1303 387 1360 412
rect 1420 413 1477 471
rect 996 343 1053 368
rect 1420 379 1432 413
rect 1466 379 1477 413
rect 1420 367 1477 379
rect 1507 596 1563 619
rect 1507 562 1518 596
rect 1552 562 1563 596
rect 1507 367 1563 562
rect 1593 367 1635 619
rect 1665 413 1721 619
rect 1665 379 1676 413
rect 1710 379 1721 413
rect 1665 367 1721 379
rect 1751 597 1808 619
rect 1751 563 1762 597
rect 1796 563 1808 597
rect 1751 483 1808 563
rect 1751 449 1762 483
rect 1796 449 1808 483
rect 1751 367 1808 449
rect 1862 607 1919 619
rect 1862 573 1874 607
rect 1908 573 1919 607
rect 1862 483 1919 573
rect 1862 449 1874 483
rect 1908 449 1919 483
rect 1862 367 1919 449
rect 1949 367 1997 619
rect 2027 597 2084 619
rect 2027 563 2038 597
rect 2072 563 2084 597
rect 2027 505 2084 563
rect 2027 471 2038 505
rect 2072 471 2084 505
rect 2027 413 2084 471
rect 2027 379 2038 413
rect 2072 379 2084 413
rect 2027 367 2084 379
<< ndiffc >>
rect 39 82 73 116
rect 197 82 231 116
rect 310 139 344 173
rect 491 89 525 123
rect 649 89 683 123
rect 874 126 908 160
rect 983 139 1017 173
rect 1147 113 1181 147
rect 1249 126 1283 160
rect 1435 91 1469 125
rect 1599 59 1633 93
rect 1945 169 1979 203
rect 1945 69 1979 103
<< pdiffc >>
rect 39 552 73 586
rect 39 482 73 516
rect 197 552 231 586
rect 197 482 231 516
rect 309 427 343 461
rect 309 357 343 391
rect 497 415 531 449
rect 700 427 734 461
rect 700 357 734 391
rect 812 396 846 430
rect 1432 563 1466 597
rect 1119 443 1153 477
rect 898 373 932 407
rect 1007 368 1041 402
rect 1205 447 1239 481
rect 1432 471 1466 505
rect 1314 412 1348 446
rect 1432 379 1466 413
rect 1518 562 1552 596
rect 1676 379 1710 413
rect 1762 563 1796 597
rect 1762 449 1796 483
rect 1874 573 1908 607
rect 1874 449 1908 483
rect 2038 563 2072 597
rect 2038 471 2072 505
rect 2038 379 2072 413
<< poly >>
rect 84 598 114 624
rect 156 598 186 624
rect 1477 619 1507 645
rect 1563 619 1593 645
rect 1635 619 1665 645
rect 1721 619 1751 645
rect 1919 619 1949 645
rect 1997 619 2027 645
rect 294 597 360 613
rect 294 563 310 597
rect 344 577 360 597
rect 1087 597 1194 613
rect 344 563 996 577
rect 294 547 996 563
rect 1087 563 1103 597
rect 1137 563 1194 597
rect 1087 547 1194 563
rect 354 473 384 499
rect 456 473 486 499
rect 587 473 617 499
rect 659 473 689 499
rect 84 370 114 470
rect 156 370 186 470
rect 84 354 186 370
rect 84 320 100 354
rect 134 320 186 354
rect 857 471 887 497
rect 84 286 186 320
rect 84 252 100 286
rect 134 252 186 286
rect 84 236 186 252
rect 84 141 114 236
rect 156 141 186 236
rect 354 313 384 345
rect 456 313 486 345
rect 354 297 486 313
rect 354 263 412 297
rect 446 263 486 297
rect 587 323 617 345
rect 659 323 689 345
rect 966 427 996 547
rect 1164 515 1194 547
rect 1273 471 1303 497
rect 587 293 689 323
rect 587 282 638 293
rect 354 229 486 263
rect 354 200 412 229
rect 378 195 412 200
rect 446 195 486 229
rect 528 266 638 282
rect 528 232 544 266
rect 578 232 638 266
rect 528 216 638 232
rect 378 179 486 195
rect 378 157 408 179
rect 450 157 480 179
rect 536 157 566 216
rect 608 157 638 216
rect 686 237 752 245
rect 857 237 887 343
rect 966 321 996 343
rect 966 291 1058 321
rect 1164 315 1194 387
rect 686 229 972 237
rect 686 195 702 229
rect 736 207 972 229
rect 736 195 752 207
rect 686 179 752 195
rect 942 185 972 207
rect 1028 185 1058 291
rect 1106 285 1194 315
rect 1106 185 1136 285
rect 1273 237 1303 387
rect 1477 303 1507 367
rect 1563 335 1593 367
rect 1635 335 1665 367
rect 1558 319 1665 335
rect 1721 325 1751 367
rect 1919 345 1949 367
rect 1444 287 1510 303
rect 1444 253 1460 287
rect 1494 253 1510 287
rect 1444 237 1510 253
rect 1208 207 1365 237
rect 1480 215 1510 237
rect 1558 285 1574 319
rect 1608 305 1665 319
rect 1713 309 1779 325
rect 1608 285 1624 305
rect 1558 269 1624 285
rect 1713 275 1729 309
rect 1763 275 1779 309
rect 1899 315 1949 345
rect 1899 303 1929 315
rect 1558 215 1588 269
rect 1713 259 1779 275
rect 1827 287 1929 303
rect 1827 253 1843 287
rect 1877 267 1929 287
rect 1997 267 2027 367
rect 1877 253 2027 267
rect 1827 237 2027 253
rect 1827 215 1857 237
rect 1899 215 1929 237
rect 1208 185 1238 207
rect 1335 187 1365 207
rect 1335 171 1401 187
rect 1335 137 1351 171
rect 1385 137 1401 171
rect 1335 103 1401 137
rect 942 75 972 101
rect 1028 75 1058 101
rect 1106 75 1136 101
rect 1208 75 1238 101
rect 84 31 114 57
rect 156 31 186 57
rect 378 47 408 73
rect 450 47 480 73
rect 536 47 566 73
rect 608 47 638 73
rect 1335 69 1351 103
rect 1385 69 1401 103
rect 1335 53 1401 69
rect 1480 21 1510 47
rect 1558 21 1588 47
rect 1827 21 1857 47
rect 1899 21 1929 47
<< polycont >>
rect 310 563 344 597
rect 1103 563 1137 597
rect 100 320 134 354
rect 100 252 134 286
rect 412 263 446 297
rect 412 195 446 229
rect 544 232 578 266
rect 702 195 736 229
rect 1460 253 1494 287
rect 1574 285 1608 319
rect 1729 275 1763 309
rect 1843 253 1877 287
rect 1351 137 1385 171
rect 1351 69 1385 103
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 23 586 89 649
rect 23 552 39 586
rect 73 552 89 586
rect 23 516 89 552
rect 23 482 39 516
rect 73 482 89 516
rect 23 466 89 482
rect 181 586 247 602
rect 181 552 197 586
rect 231 552 247 586
rect 181 516 247 552
rect 181 482 197 516
rect 231 482 247 516
rect 181 466 247 482
rect 25 354 167 430
rect 25 320 100 354
rect 134 320 167 354
rect 25 286 167 320
rect 25 252 100 286
rect 134 252 167 286
rect 25 236 167 252
rect 213 145 247 466
rect 23 116 89 145
rect 23 82 39 116
rect 73 82 89 116
rect 23 17 89 82
rect 181 116 247 145
rect 293 597 360 613
rect 293 563 310 597
rect 344 563 360 597
rect 293 461 360 563
rect 293 427 309 461
rect 343 427 360 461
rect 293 391 360 427
rect 293 357 309 391
rect 343 357 360 391
rect 481 449 547 649
rect 481 415 497 449
rect 531 415 547 449
rect 481 388 547 415
rect 700 597 1153 613
rect 700 563 1103 597
rect 1137 563 1153 597
rect 700 547 1153 563
rect 700 461 750 547
rect 734 427 750 461
rect 700 391 750 427
rect 293 173 360 357
rect 734 357 750 391
rect 293 139 310 173
rect 344 139 360 173
rect 293 123 360 139
rect 396 318 664 352
rect 396 297 462 318
rect 396 263 412 297
rect 446 263 462 297
rect 396 229 462 263
rect 396 195 412 229
rect 446 195 462 229
rect 505 266 594 282
rect 505 232 544 266
rect 578 232 594 266
rect 505 216 594 232
rect 630 245 664 318
rect 700 315 750 357
rect 796 477 1153 511
rect 796 430 862 477
rect 1103 443 1119 477
rect 796 396 812 430
rect 846 396 862 430
rect 796 351 862 396
rect 898 407 948 441
rect 932 373 948 407
rect 700 281 822 315
rect 630 229 752 245
rect 396 179 462 195
rect 630 195 702 229
rect 736 195 752 229
rect 630 179 752 195
rect 181 82 197 116
rect 231 87 247 116
rect 396 87 430 179
rect 788 143 822 281
rect 898 303 948 373
rect 991 402 1057 431
rect 1103 409 1153 443
rect 1189 481 1255 649
rect 1189 447 1205 481
rect 1239 447 1255 481
rect 1416 597 1482 613
rect 1416 563 1432 597
rect 1466 563 1482 597
rect 1416 505 1482 563
rect 1518 596 1568 649
rect 1552 562 1568 596
rect 1518 535 1568 562
rect 1762 597 1812 613
rect 1796 563 1812 597
rect 1189 409 1255 447
rect 1298 446 1364 475
rect 1298 412 1314 446
rect 1348 412 1364 446
rect 991 368 1007 402
rect 1041 373 1057 402
rect 1298 373 1364 412
rect 1041 368 1364 373
rect 991 339 1364 368
rect 1416 471 1432 505
rect 1466 499 1482 505
rect 1762 499 1812 563
rect 1466 483 1812 499
rect 1466 471 1762 483
rect 1416 465 1762 471
rect 1416 413 1482 465
rect 1796 449 1812 483
rect 1762 433 1812 449
rect 1858 607 1924 649
rect 1858 573 1874 607
rect 1908 573 1924 607
rect 1858 483 1924 573
rect 1858 449 1874 483
rect 1908 449 1924 483
rect 1858 433 1924 449
rect 2022 597 2088 613
rect 2022 563 2038 597
rect 2072 563 2088 597
rect 2022 505 2088 563
rect 2022 471 2038 505
rect 2072 471 2088 505
rect 1416 379 1432 413
rect 1466 379 1482 413
rect 1416 363 1482 379
rect 1660 413 1726 429
rect 1660 379 1676 413
rect 1710 397 1726 413
rect 2022 413 2088 471
rect 1710 379 1849 397
rect 1660 363 1849 379
rect 1558 319 1624 356
rect 898 287 1510 303
rect 898 269 1460 287
rect 231 82 430 87
rect 181 53 430 82
rect 475 123 541 143
rect 475 89 491 123
rect 525 89 541 123
rect 475 17 541 89
rect 633 123 822 143
rect 633 89 649 123
rect 683 109 822 123
rect 858 160 924 189
rect 858 126 874 160
rect 908 126 924 160
rect 683 89 699 109
rect 633 69 699 89
rect 858 87 924 126
rect 967 173 1017 269
rect 1444 253 1460 269
rect 1494 253 1510 287
rect 1558 285 1574 319
rect 1608 285 1624 319
rect 1558 269 1624 285
rect 1713 309 1779 325
rect 1713 275 1729 309
rect 1763 275 1779 309
rect 1444 233 1510 253
rect 1713 233 1779 275
rect 967 139 983 173
rect 967 123 1017 139
rect 1053 199 1299 233
rect 1444 199 1779 233
rect 1815 303 1849 363
rect 2022 379 2038 413
rect 2072 379 2088 413
rect 1815 287 1893 303
rect 1815 253 1843 287
rect 1877 253 1893 287
rect 1815 237 1893 253
rect 1053 87 1087 199
rect 858 53 1087 87
rect 1131 147 1197 163
rect 1131 113 1147 147
rect 1181 113 1197 147
rect 1131 17 1197 113
rect 1233 160 1299 199
rect 1233 126 1249 160
rect 1283 126 1299 160
rect 1233 97 1299 126
rect 1335 171 1401 187
rect 1335 137 1351 171
rect 1385 163 1401 171
rect 1815 163 1849 237
rect 2022 219 2088 379
rect 1385 137 1849 163
rect 1335 129 1849 137
rect 1929 203 2088 219
rect 1929 169 1945 203
rect 1979 169 2088 203
rect 1335 125 1485 129
rect 1335 103 1435 125
rect 1335 69 1351 103
rect 1385 91 1435 103
rect 1469 91 1485 125
rect 1929 103 2088 169
rect 1385 69 1485 91
rect 1335 53 1485 69
rect 1583 59 1599 93
rect 1633 59 1649 93
rect 1583 17 1649 59
rect 1929 69 1945 103
rect 1979 69 2088 103
rect 1929 53 2088 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrtp_lp
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 2047 94 2081 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 168 2081 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 464 2081 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 538 2081 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1897908
string GDS_START 1883634
<< end >>
