magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3966 1852
<< nwell >>
rect -38 261 2706 582
<< pwell >>
rect 1 21 2651 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 277 47 307 177
rect 371 47 401 177
rect 475 47 505 177
rect 559 47 589 177
rect 653 47 683 177
rect 747 47 777 177
rect 841 47 871 177
rect 935 47 965 177
rect 1039 47 1069 177
rect 1123 47 1153 177
rect 1217 47 1247 177
rect 1311 47 1341 177
rect 1405 47 1435 177
rect 1499 47 1529 177
rect 1593 47 1623 177
rect 1687 47 1717 177
rect 1781 47 1811 177
rect 1875 47 1905 177
rect 1969 47 1999 177
rect 2063 47 2093 177
rect 2157 47 2187 177
rect 2251 47 2281 177
rect 2345 47 2375 177
rect 2439 47 2469 177
rect 2543 47 2573 177
<< scpmoshvt >>
rect 81 297 117 497
rect 279 297 315 497
rect 373 297 409 497
rect 467 297 503 497
rect 561 297 597 497
rect 655 297 691 497
rect 749 297 785 497
rect 843 297 879 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1125 297 1161 497
rect 1219 297 1255 497
rect 1313 297 1349 497
rect 1407 297 1443 497
rect 1501 297 1537 497
rect 1595 297 1631 497
rect 1689 297 1725 497
rect 1783 297 1819 497
rect 1877 297 1913 497
rect 1971 297 2007 497
rect 2065 297 2101 497
rect 2159 297 2195 497
rect 2253 297 2289 497
rect 2347 297 2383 497
rect 2441 297 2477 497
rect 2535 297 2571 497
<< ndiff >>
rect 27 165 89 177
rect 27 131 35 165
rect 69 131 89 165
rect 27 97 89 131
rect 27 63 35 97
rect 69 63 89 97
rect 27 47 89 63
rect 119 165 171 177
rect 119 131 129 165
rect 163 131 171 165
rect 119 97 171 131
rect 119 63 129 97
rect 163 63 171 97
rect 119 47 171 63
rect 225 165 277 177
rect 225 131 233 165
rect 267 131 277 165
rect 225 97 277 131
rect 225 63 233 97
rect 267 63 277 97
rect 225 47 277 63
rect 307 97 371 177
rect 307 63 327 97
rect 361 63 371 97
rect 307 47 371 63
rect 401 165 475 177
rect 401 131 421 165
rect 455 131 475 165
rect 401 97 475 131
rect 401 63 421 97
rect 455 63 475 97
rect 401 47 475 63
rect 505 97 559 177
rect 505 63 515 97
rect 549 63 559 97
rect 505 47 559 63
rect 589 165 653 177
rect 589 131 609 165
rect 643 131 653 165
rect 589 97 653 131
rect 589 63 609 97
rect 643 63 653 97
rect 589 47 653 63
rect 683 97 747 177
rect 683 63 703 97
rect 737 63 747 97
rect 683 47 747 63
rect 777 165 841 177
rect 777 131 797 165
rect 831 131 841 165
rect 777 97 841 131
rect 777 63 797 97
rect 831 63 841 97
rect 777 47 841 63
rect 871 97 935 177
rect 871 63 891 97
rect 925 63 935 97
rect 871 47 935 63
rect 965 165 1039 177
rect 965 131 985 165
rect 1019 131 1039 165
rect 965 97 1039 131
rect 965 63 985 97
rect 1019 63 1039 97
rect 965 47 1039 63
rect 1069 97 1123 177
rect 1069 63 1079 97
rect 1113 63 1123 97
rect 1069 47 1123 63
rect 1153 165 1217 177
rect 1153 131 1173 165
rect 1207 131 1217 165
rect 1153 97 1217 131
rect 1153 63 1173 97
rect 1207 63 1217 97
rect 1153 47 1217 63
rect 1247 97 1311 177
rect 1247 63 1267 97
rect 1301 63 1311 97
rect 1247 47 1311 63
rect 1341 165 1405 177
rect 1341 131 1361 165
rect 1395 131 1405 165
rect 1341 97 1405 131
rect 1341 63 1361 97
rect 1395 63 1405 97
rect 1341 47 1405 63
rect 1435 97 1499 177
rect 1435 63 1455 97
rect 1489 63 1499 97
rect 1435 47 1499 63
rect 1529 165 1593 177
rect 1529 131 1549 165
rect 1583 131 1593 165
rect 1529 97 1593 131
rect 1529 63 1549 97
rect 1583 63 1593 97
rect 1529 47 1593 63
rect 1623 97 1687 177
rect 1623 63 1643 97
rect 1677 63 1687 97
rect 1623 47 1687 63
rect 1717 165 1781 177
rect 1717 131 1737 165
rect 1771 131 1781 165
rect 1717 97 1781 131
rect 1717 63 1737 97
rect 1771 63 1781 97
rect 1717 47 1781 63
rect 1811 97 1875 177
rect 1811 63 1831 97
rect 1865 63 1875 97
rect 1811 47 1875 63
rect 1905 165 1969 177
rect 1905 131 1925 165
rect 1959 131 1969 165
rect 1905 97 1969 131
rect 1905 63 1925 97
rect 1959 63 1969 97
rect 1905 47 1969 63
rect 1999 97 2063 177
rect 1999 63 2019 97
rect 2053 63 2063 97
rect 1999 47 2063 63
rect 2093 165 2157 177
rect 2093 131 2113 165
rect 2147 131 2157 165
rect 2093 97 2157 131
rect 2093 63 2113 97
rect 2147 63 2157 97
rect 2093 47 2157 63
rect 2187 97 2251 177
rect 2187 63 2207 97
rect 2241 63 2251 97
rect 2187 47 2251 63
rect 2281 165 2345 177
rect 2281 131 2301 165
rect 2335 131 2345 165
rect 2281 97 2345 131
rect 2281 63 2301 97
rect 2335 63 2345 97
rect 2281 47 2345 63
rect 2375 97 2439 177
rect 2375 63 2395 97
rect 2429 63 2439 97
rect 2375 47 2439 63
rect 2469 165 2543 177
rect 2469 131 2489 165
rect 2523 131 2543 165
rect 2469 97 2543 131
rect 2469 63 2489 97
rect 2523 63 2543 97
rect 2469 47 2543 63
rect 2573 97 2625 177
rect 2573 63 2583 97
rect 2617 63 2625 97
rect 2573 47 2625 63
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 479 171 497
rect 117 445 129 479
rect 163 445 171 479
rect 117 411 171 445
rect 117 377 129 411
rect 163 377 171 411
rect 117 343 171 377
rect 117 309 129 343
rect 163 309 171 343
rect 117 297 171 309
rect 225 479 279 497
rect 225 445 233 479
rect 267 445 279 479
rect 225 411 279 445
rect 225 377 233 411
rect 267 377 279 411
rect 225 343 279 377
rect 225 309 233 343
rect 267 309 279 343
rect 225 297 279 309
rect 315 485 373 497
rect 315 451 327 485
rect 361 451 373 485
rect 315 417 373 451
rect 315 383 327 417
rect 361 383 373 417
rect 315 297 373 383
rect 409 479 467 497
rect 409 445 421 479
rect 455 445 467 479
rect 409 411 467 445
rect 409 377 421 411
rect 455 377 467 411
rect 409 343 467 377
rect 409 309 421 343
rect 455 309 467 343
rect 409 297 467 309
rect 503 485 561 497
rect 503 451 515 485
rect 549 451 561 485
rect 503 417 561 451
rect 503 383 515 417
rect 549 383 561 417
rect 503 297 561 383
rect 597 479 655 497
rect 597 445 609 479
rect 643 445 655 479
rect 597 411 655 445
rect 597 377 609 411
rect 643 377 655 411
rect 597 343 655 377
rect 597 309 609 343
rect 643 309 655 343
rect 597 297 655 309
rect 691 485 749 497
rect 691 451 703 485
rect 737 451 749 485
rect 691 417 749 451
rect 691 383 703 417
rect 737 383 749 417
rect 691 297 749 383
rect 785 479 843 497
rect 785 445 797 479
rect 831 445 843 479
rect 785 411 843 445
rect 785 377 797 411
rect 831 377 843 411
rect 785 343 843 377
rect 785 309 797 343
rect 831 309 843 343
rect 785 297 843 309
rect 879 485 937 497
rect 879 451 891 485
rect 925 451 937 485
rect 879 417 937 451
rect 879 383 891 417
rect 925 383 937 417
rect 879 297 937 383
rect 973 479 1031 497
rect 973 445 985 479
rect 1019 445 1031 479
rect 973 411 1031 445
rect 973 377 985 411
rect 1019 377 1031 411
rect 973 343 1031 377
rect 973 309 985 343
rect 1019 309 1031 343
rect 973 297 1031 309
rect 1067 485 1125 497
rect 1067 451 1079 485
rect 1113 451 1125 485
rect 1067 417 1125 451
rect 1067 383 1079 417
rect 1113 383 1125 417
rect 1067 297 1125 383
rect 1161 479 1219 497
rect 1161 445 1173 479
rect 1207 445 1219 479
rect 1161 411 1219 445
rect 1161 377 1173 411
rect 1207 377 1219 411
rect 1161 343 1219 377
rect 1161 309 1173 343
rect 1207 309 1219 343
rect 1161 297 1219 309
rect 1255 485 1313 497
rect 1255 451 1267 485
rect 1301 451 1313 485
rect 1255 417 1313 451
rect 1255 383 1267 417
rect 1301 383 1313 417
rect 1255 297 1313 383
rect 1349 479 1407 497
rect 1349 445 1361 479
rect 1395 445 1407 479
rect 1349 411 1407 445
rect 1349 377 1361 411
rect 1395 377 1407 411
rect 1349 343 1407 377
rect 1349 309 1361 343
rect 1395 309 1407 343
rect 1349 297 1407 309
rect 1443 485 1501 497
rect 1443 451 1455 485
rect 1489 451 1501 485
rect 1443 417 1501 451
rect 1443 383 1455 417
rect 1489 383 1501 417
rect 1443 297 1501 383
rect 1537 479 1595 497
rect 1537 445 1549 479
rect 1583 445 1595 479
rect 1537 411 1595 445
rect 1537 377 1549 411
rect 1583 377 1595 411
rect 1537 343 1595 377
rect 1537 309 1549 343
rect 1583 309 1595 343
rect 1537 297 1595 309
rect 1631 485 1689 497
rect 1631 451 1643 485
rect 1677 451 1689 485
rect 1631 417 1689 451
rect 1631 383 1643 417
rect 1677 383 1689 417
rect 1631 297 1689 383
rect 1725 479 1783 497
rect 1725 445 1737 479
rect 1771 445 1783 479
rect 1725 411 1783 445
rect 1725 377 1737 411
rect 1771 377 1783 411
rect 1725 343 1783 377
rect 1725 309 1737 343
rect 1771 309 1783 343
rect 1725 297 1783 309
rect 1819 485 1877 497
rect 1819 451 1831 485
rect 1865 451 1877 485
rect 1819 417 1877 451
rect 1819 383 1831 417
rect 1865 383 1877 417
rect 1819 297 1877 383
rect 1913 479 1971 497
rect 1913 445 1925 479
rect 1959 445 1971 479
rect 1913 411 1971 445
rect 1913 377 1925 411
rect 1959 377 1971 411
rect 1913 343 1971 377
rect 1913 309 1925 343
rect 1959 309 1971 343
rect 1913 297 1971 309
rect 2007 485 2065 497
rect 2007 451 2019 485
rect 2053 451 2065 485
rect 2007 417 2065 451
rect 2007 383 2019 417
rect 2053 383 2065 417
rect 2007 297 2065 383
rect 2101 479 2159 497
rect 2101 445 2113 479
rect 2147 445 2159 479
rect 2101 411 2159 445
rect 2101 377 2113 411
rect 2147 377 2159 411
rect 2101 343 2159 377
rect 2101 309 2113 343
rect 2147 309 2159 343
rect 2101 297 2159 309
rect 2195 485 2253 497
rect 2195 451 2207 485
rect 2241 451 2253 485
rect 2195 417 2253 451
rect 2195 383 2207 417
rect 2241 383 2253 417
rect 2195 297 2253 383
rect 2289 479 2347 497
rect 2289 445 2301 479
rect 2335 445 2347 479
rect 2289 411 2347 445
rect 2289 377 2301 411
rect 2335 377 2347 411
rect 2289 343 2347 377
rect 2289 309 2301 343
rect 2335 309 2347 343
rect 2289 297 2347 309
rect 2383 485 2441 497
rect 2383 451 2395 485
rect 2429 451 2441 485
rect 2383 417 2441 451
rect 2383 383 2395 417
rect 2429 383 2441 417
rect 2383 297 2441 383
rect 2477 479 2535 497
rect 2477 445 2489 479
rect 2523 445 2535 479
rect 2477 411 2535 445
rect 2477 377 2489 411
rect 2523 377 2535 411
rect 2477 343 2535 377
rect 2477 309 2489 343
rect 2523 309 2535 343
rect 2477 297 2535 309
rect 2571 485 2625 497
rect 2571 451 2583 485
rect 2617 451 2625 485
rect 2571 417 2625 451
rect 2571 383 2583 417
rect 2617 383 2625 417
rect 2571 297 2625 383
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 129 131 163 165
rect 129 63 163 97
rect 233 131 267 165
rect 233 63 267 97
rect 327 63 361 97
rect 421 131 455 165
rect 421 63 455 97
rect 515 63 549 97
rect 609 131 643 165
rect 609 63 643 97
rect 703 63 737 97
rect 797 131 831 165
rect 797 63 831 97
rect 891 63 925 97
rect 985 131 1019 165
rect 985 63 1019 97
rect 1079 63 1113 97
rect 1173 131 1207 165
rect 1173 63 1207 97
rect 1267 63 1301 97
rect 1361 131 1395 165
rect 1361 63 1395 97
rect 1455 63 1489 97
rect 1549 131 1583 165
rect 1549 63 1583 97
rect 1643 63 1677 97
rect 1737 131 1771 165
rect 1737 63 1771 97
rect 1831 63 1865 97
rect 1925 131 1959 165
rect 1925 63 1959 97
rect 2019 63 2053 97
rect 2113 131 2147 165
rect 2113 63 2147 97
rect 2207 63 2241 97
rect 2301 131 2335 165
rect 2301 63 2335 97
rect 2395 63 2429 97
rect 2489 131 2523 165
rect 2489 63 2523 97
rect 2583 63 2617 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 445 163 479
rect 129 377 163 411
rect 129 309 163 343
rect 233 445 267 479
rect 233 377 267 411
rect 233 309 267 343
rect 327 451 361 485
rect 327 383 361 417
rect 421 445 455 479
rect 421 377 455 411
rect 421 309 455 343
rect 515 451 549 485
rect 515 383 549 417
rect 609 445 643 479
rect 609 377 643 411
rect 609 309 643 343
rect 703 451 737 485
rect 703 383 737 417
rect 797 445 831 479
rect 797 377 831 411
rect 797 309 831 343
rect 891 451 925 485
rect 891 383 925 417
rect 985 445 1019 479
rect 985 377 1019 411
rect 985 309 1019 343
rect 1079 451 1113 485
rect 1079 383 1113 417
rect 1173 445 1207 479
rect 1173 377 1207 411
rect 1173 309 1207 343
rect 1267 451 1301 485
rect 1267 383 1301 417
rect 1361 445 1395 479
rect 1361 377 1395 411
rect 1361 309 1395 343
rect 1455 451 1489 485
rect 1455 383 1489 417
rect 1549 445 1583 479
rect 1549 377 1583 411
rect 1549 309 1583 343
rect 1643 451 1677 485
rect 1643 383 1677 417
rect 1737 445 1771 479
rect 1737 377 1771 411
rect 1737 309 1771 343
rect 1831 451 1865 485
rect 1831 383 1865 417
rect 1925 445 1959 479
rect 1925 377 1959 411
rect 1925 309 1959 343
rect 2019 451 2053 485
rect 2019 383 2053 417
rect 2113 445 2147 479
rect 2113 377 2147 411
rect 2113 309 2147 343
rect 2207 451 2241 485
rect 2207 383 2241 417
rect 2301 445 2335 479
rect 2301 377 2335 411
rect 2301 309 2335 343
rect 2395 451 2429 485
rect 2395 383 2429 417
rect 2489 445 2523 479
rect 2489 377 2523 411
rect 2489 309 2523 343
rect 2583 451 2617 485
rect 2583 383 2617 417
<< poly >>
rect 81 497 117 523
rect 279 497 315 523
rect 373 497 409 523
rect 467 497 503 523
rect 561 497 597 523
rect 655 497 691 523
rect 749 497 785 523
rect 843 497 879 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1125 497 1161 523
rect 1219 497 1255 523
rect 1313 497 1349 523
rect 1407 497 1443 523
rect 1501 497 1537 523
rect 1595 497 1631 523
rect 1689 497 1725 523
rect 1783 497 1819 523
rect 1877 497 1913 523
rect 1971 497 2007 523
rect 2065 497 2101 523
rect 2159 497 2195 523
rect 2253 497 2289 523
rect 2347 497 2383 523
rect 2441 497 2477 523
rect 2535 497 2571 523
rect 81 282 117 297
rect 279 282 315 297
rect 373 282 409 297
rect 467 282 503 297
rect 561 282 597 297
rect 655 282 691 297
rect 749 282 785 297
rect 843 282 879 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1125 282 1161 297
rect 1219 282 1255 297
rect 1313 282 1349 297
rect 1407 282 1443 297
rect 1501 282 1537 297
rect 1595 282 1631 297
rect 1689 282 1725 297
rect 1783 282 1819 297
rect 1877 282 1913 297
rect 1971 282 2007 297
rect 2065 282 2101 297
rect 2159 282 2195 297
rect 2253 282 2289 297
rect 2347 282 2383 297
rect 2441 282 2477 297
rect 2535 282 2571 297
rect 79 265 119 282
rect 22 249 119 265
rect 22 215 38 249
rect 72 215 119 249
rect 22 199 119 215
rect 89 177 119 199
rect 277 259 317 282
rect 371 259 411 282
rect 465 259 505 282
rect 277 249 505 259
rect 277 215 327 249
rect 361 215 395 249
rect 429 215 505 249
rect 277 205 505 215
rect 277 177 307 205
rect 371 177 401 205
rect 475 177 505 205
rect 559 259 599 282
rect 653 259 693 282
rect 747 259 787 282
rect 841 259 881 282
rect 935 259 975 282
rect 1029 259 1069 282
rect 559 249 1069 259
rect 559 215 583 249
rect 617 215 661 249
rect 695 215 739 249
rect 773 215 817 249
rect 851 215 895 249
rect 929 215 963 249
rect 997 215 1069 249
rect 559 205 1069 215
rect 559 177 589 205
rect 653 177 683 205
rect 747 177 777 205
rect 841 177 871 205
rect 935 177 965 205
rect 1039 177 1069 205
rect 1123 259 1163 282
rect 1217 259 1257 282
rect 1311 259 1351 282
rect 1405 259 1445 282
rect 1499 259 1539 282
rect 1593 259 1633 282
rect 1687 259 1727 282
rect 1781 259 1821 282
rect 1875 259 1915 282
rect 1969 259 2009 282
rect 2063 259 2103 282
rect 2157 259 2197 282
rect 2251 259 2291 282
rect 2345 259 2385 282
rect 2439 259 2479 282
rect 2533 259 2573 282
rect 1123 249 2573 259
rect 1123 215 1143 249
rect 1177 215 1221 249
rect 1255 215 1299 249
rect 1333 215 1377 249
rect 1411 215 1455 249
rect 1489 215 1523 249
rect 1557 215 1601 249
rect 1635 215 1679 249
rect 1713 215 1757 249
rect 1791 215 1835 249
rect 1869 215 1903 249
rect 1937 215 1981 249
rect 2015 215 2059 249
rect 2093 215 2137 249
rect 2171 215 2215 249
rect 2249 215 2293 249
rect 2327 215 2361 249
rect 2395 215 2439 249
rect 2473 215 2573 249
rect 1123 205 2573 215
rect 1123 177 1153 205
rect 1217 177 1247 205
rect 1311 177 1341 205
rect 1405 177 1435 205
rect 1499 177 1529 205
rect 1593 177 1623 205
rect 1687 177 1717 205
rect 1781 177 1811 205
rect 1875 177 1905 205
rect 1969 177 1999 205
rect 2063 177 2093 205
rect 2157 177 2187 205
rect 2251 177 2281 205
rect 2345 177 2375 205
rect 2439 177 2469 205
rect 2543 177 2573 205
rect 89 21 119 47
rect 277 21 307 47
rect 371 21 401 47
rect 475 21 505 47
rect 559 21 589 47
rect 653 21 683 47
rect 747 21 777 47
rect 841 21 871 47
rect 935 21 965 47
rect 1039 21 1069 47
rect 1123 21 1153 47
rect 1217 21 1247 47
rect 1311 21 1341 47
rect 1405 21 1435 47
rect 1499 21 1529 47
rect 1593 21 1623 47
rect 1687 21 1717 47
rect 1781 21 1811 47
rect 1875 21 1905 47
rect 1969 21 1999 47
rect 2063 21 2093 47
rect 2157 21 2187 47
rect 2251 21 2281 47
rect 2345 21 2375 47
rect 2439 21 2469 47
rect 2543 21 2573 47
<< polycont >>
rect 38 215 72 249
rect 327 215 361 249
rect 395 215 429 249
rect 583 215 617 249
rect 661 215 695 249
rect 739 215 773 249
rect 817 215 851 249
rect 895 215 929 249
rect 963 215 997 249
rect 1143 215 1177 249
rect 1221 215 1255 249
rect 1299 215 1333 249
rect 1377 215 1411 249
rect 1455 215 1489 249
rect 1523 215 1557 249
rect 1601 215 1635 249
rect 1679 215 1713 249
rect 1757 215 1791 249
rect 1835 215 1869 249
rect 1903 215 1937 249
rect 1981 215 2015 249
rect 2059 215 2093 249
rect 2137 215 2171 249
rect 2215 215 2249 249
rect 2293 215 2327 249
rect 2361 215 2395 249
rect 2439 215 2473 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 35 485 69 527
rect 35 417 69 451
rect 35 349 69 383
rect 35 289 69 315
rect 103 479 179 493
rect 103 445 129 479
rect 163 445 179 479
rect 103 411 179 445
rect 103 377 129 411
rect 163 377 179 411
rect 103 343 179 377
rect 103 309 129 343
rect 163 309 179 343
rect 103 289 179 309
rect 217 479 283 493
rect 217 445 233 479
rect 267 445 283 479
rect 217 411 283 445
rect 217 377 233 411
rect 267 377 283 411
rect 217 343 283 377
rect 327 485 361 527
rect 327 417 361 451
rect 327 357 361 383
rect 395 479 471 493
rect 395 445 421 479
rect 455 445 471 479
rect 395 411 471 445
rect 395 377 421 411
rect 455 377 471 411
rect 217 309 233 343
rect 267 323 283 343
rect 395 343 471 377
rect 515 485 549 527
rect 515 417 549 451
rect 515 357 549 383
rect 583 479 659 493
rect 583 445 609 479
rect 643 445 659 479
rect 583 411 659 445
rect 583 377 609 411
rect 643 377 659 411
rect 395 323 421 343
rect 267 309 421 323
rect 455 323 471 343
rect 583 343 659 377
rect 703 485 737 527
rect 703 417 737 451
rect 703 367 737 383
rect 771 479 847 493
rect 771 445 797 479
rect 831 445 847 479
rect 771 411 847 445
rect 771 377 797 411
rect 831 377 847 411
rect 455 309 549 323
rect 217 289 549 309
rect 583 309 609 343
rect 643 323 659 343
rect 771 343 847 377
rect 891 485 925 527
rect 891 417 925 451
rect 891 367 925 383
rect 959 479 1035 493
rect 959 445 985 479
rect 1019 445 1035 479
rect 959 411 1035 445
rect 959 377 985 411
rect 1019 377 1035 411
rect 771 323 797 343
rect 643 309 797 323
rect 831 323 847 343
rect 959 343 1035 377
rect 1079 485 1113 527
rect 1079 417 1113 451
rect 1079 367 1113 383
rect 1147 479 1223 493
rect 1147 445 1173 479
rect 1207 445 1223 479
rect 1147 411 1223 445
rect 1147 377 1173 411
rect 1207 377 1223 411
rect 959 323 985 343
rect 831 309 985 323
rect 1019 323 1035 343
rect 1147 343 1223 377
rect 1267 485 1301 527
rect 1267 417 1301 451
rect 1267 367 1301 383
rect 1335 479 1411 493
rect 1335 445 1361 479
rect 1395 445 1411 479
rect 1335 411 1411 445
rect 1335 377 1361 411
rect 1395 377 1411 411
rect 1019 309 1113 323
rect 583 289 1113 309
rect 1147 309 1173 343
rect 1207 323 1223 343
rect 1335 343 1411 377
rect 1455 485 1489 527
rect 1455 417 1489 451
rect 1455 367 1489 383
rect 1523 479 1599 493
rect 1523 445 1549 479
rect 1583 445 1599 479
rect 1523 411 1599 445
rect 1523 377 1549 411
rect 1583 377 1599 411
rect 1335 323 1361 343
rect 1207 309 1361 323
rect 1395 323 1411 343
rect 1523 343 1599 377
rect 1643 485 1677 527
rect 1643 417 1677 451
rect 1643 367 1677 383
rect 1711 479 1787 493
rect 1711 445 1737 479
rect 1771 445 1787 479
rect 1711 411 1787 445
rect 1711 377 1737 411
rect 1771 377 1787 411
rect 1523 323 1549 343
rect 1395 309 1549 323
rect 1583 323 1599 343
rect 1711 343 1787 377
rect 1831 485 1865 527
rect 1831 417 1865 451
rect 1831 367 1865 383
rect 1899 479 1975 493
rect 1899 445 1925 479
rect 1959 445 1975 479
rect 1899 411 1975 445
rect 1899 377 1925 411
rect 1959 377 1975 411
rect 1711 323 1737 343
rect 1583 309 1737 323
rect 1771 323 1787 343
rect 1899 343 1975 377
rect 2019 485 2053 527
rect 2019 417 2053 451
rect 2019 367 2053 383
rect 2087 479 2163 493
rect 2087 445 2113 479
rect 2147 445 2163 479
rect 2087 411 2163 445
rect 2087 377 2113 411
rect 2147 377 2163 411
rect 1899 323 1925 343
rect 1771 309 1925 323
rect 1959 323 1975 343
rect 2087 343 2163 377
rect 2207 485 2241 527
rect 2207 417 2241 451
rect 2207 367 2241 383
rect 2275 479 2351 493
rect 2275 445 2301 479
rect 2335 445 2351 479
rect 2275 411 2351 445
rect 2275 377 2301 411
rect 2335 377 2351 411
rect 2087 323 2113 343
rect 1959 309 2113 323
rect 2147 323 2163 343
rect 2275 343 2351 377
rect 2395 485 2429 527
rect 2395 417 2429 451
rect 2395 367 2429 383
rect 2463 479 2539 493
rect 2463 445 2489 479
rect 2523 445 2539 479
rect 2463 411 2539 445
rect 2463 377 2489 411
rect 2523 377 2539 411
rect 2275 323 2301 343
rect 2147 309 2301 323
rect 2335 323 2351 343
rect 2463 343 2539 377
rect 2583 485 2617 527
rect 2583 417 2617 451
rect 2583 367 2617 383
rect 2463 323 2489 343
rect 2335 309 2489 323
rect 2523 323 2539 343
rect 2523 309 2644 323
rect 1147 289 2644 309
rect 132 255 179 289
rect 515 255 549 289
rect 1078 255 1113 289
rect 22 249 88 255
rect 22 215 38 249
rect 72 215 88 249
rect 132 249 471 255
rect 132 215 327 249
rect 361 215 395 249
rect 429 215 471 249
rect 515 249 1027 255
rect 515 215 583 249
rect 617 215 661 249
rect 695 215 739 249
rect 773 215 817 249
rect 851 215 895 249
rect 929 215 963 249
rect 997 215 1027 249
rect 1078 249 2540 255
rect 1078 215 1143 249
rect 1177 215 1221 249
rect 1255 215 1299 249
rect 1333 215 1377 249
rect 1411 215 1455 249
rect 1489 215 1523 249
rect 1557 215 1601 249
rect 1635 215 1679 249
rect 1713 215 1757 249
rect 1791 215 1835 249
rect 1869 215 1903 249
rect 1937 215 1981 249
rect 2015 215 2059 249
rect 2093 215 2137 249
rect 2171 215 2215 249
rect 2249 215 2293 249
rect 2327 215 2361 249
rect 2395 215 2439 249
rect 2473 215 2540 249
rect 132 181 179 215
rect 515 181 549 215
rect 1078 181 1113 215
rect 2584 181 2644 289
rect 35 165 69 181
rect 35 97 69 131
rect 35 17 69 63
rect 103 165 179 181
rect 103 131 129 165
rect 163 131 179 165
rect 103 97 179 131
rect 103 63 129 97
rect 163 63 179 97
rect 103 52 179 63
rect 217 165 549 181
rect 217 131 233 165
rect 267 147 421 165
rect 267 131 283 147
rect 217 97 283 131
rect 395 131 421 147
rect 455 147 549 165
rect 583 165 1113 181
rect 455 131 471 147
rect 217 63 233 97
rect 267 63 283 97
rect 217 52 283 63
rect 327 97 361 113
rect 327 17 361 63
rect 395 97 471 131
rect 583 131 609 165
rect 643 147 797 165
rect 643 131 659 147
rect 395 63 421 97
rect 455 63 471 97
rect 395 52 471 63
rect 515 97 549 113
rect 515 17 549 63
rect 583 97 659 131
rect 771 131 797 147
rect 831 147 985 165
rect 831 131 847 147
rect 583 63 609 97
rect 643 63 659 97
rect 583 52 659 63
rect 703 97 737 113
rect 703 17 737 63
rect 771 97 847 131
rect 959 131 985 147
rect 1019 147 1113 165
rect 1147 165 2644 181
rect 1019 131 1035 147
rect 771 63 797 97
rect 831 63 847 97
rect 771 52 847 63
rect 891 97 925 113
rect 891 17 925 63
rect 959 97 1035 131
rect 1147 131 1173 165
rect 1207 147 1361 165
rect 1207 131 1223 147
rect 959 63 985 97
rect 1019 63 1035 97
rect 959 52 1035 63
rect 1079 97 1113 113
rect 1079 17 1113 63
rect 1147 97 1223 131
rect 1335 131 1361 147
rect 1395 147 1549 165
rect 1395 131 1411 147
rect 1147 63 1173 97
rect 1207 63 1223 97
rect 1147 52 1223 63
rect 1267 97 1301 113
rect 1147 51 1207 52
rect 1267 17 1301 63
rect 1335 97 1411 131
rect 1523 131 1549 147
rect 1583 147 1737 165
rect 1583 131 1599 147
rect 1335 63 1361 97
rect 1395 63 1411 97
rect 1335 52 1411 63
rect 1455 97 1489 113
rect 1361 51 1395 52
rect 1455 17 1489 63
rect 1523 97 1599 131
rect 1711 131 1737 147
rect 1771 147 1925 165
rect 1771 131 1787 147
rect 1523 63 1549 97
rect 1583 63 1599 97
rect 1523 52 1599 63
rect 1643 97 1677 113
rect 1549 51 1583 52
rect 1643 17 1677 63
rect 1711 97 1787 131
rect 1899 131 1925 147
rect 1959 147 2113 165
rect 1959 131 1975 147
rect 1711 63 1737 97
rect 1771 63 1787 97
rect 1711 52 1787 63
rect 1831 97 1865 113
rect 1831 17 1865 63
rect 1899 97 1975 131
rect 2087 131 2113 147
rect 2147 147 2301 165
rect 2147 131 2163 147
rect 1899 63 1925 97
rect 1959 63 1975 97
rect 1899 52 1975 63
rect 2019 97 2053 113
rect 2019 17 2053 63
rect 2087 97 2163 131
rect 2275 131 2301 147
rect 2335 147 2489 165
rect 2335 131 2351 147
rect 2087 63 2113 97
rect 2147 63 2163 97
rect 2087 52 2163 63
rect 2207 97 2241 113
rect 2207 17 2241 63
rect 2275 97 2351 131
rect 2463 131 2489 147
rect 2523 147 2644 165
rect 2523 131 2539 147
rect 2275 63 2301 97
rect 2335 63 2351 97
rect 2275 52 2351 63
rect 2395 97 2429 113
rect 2395 17 2429 63
rect 2463 97 2539 131
rect 2463 63 2489 97
rect 2523 63 2539 97
rect 2463 52 2539 63
rect 2583 97 2617 113
rect 2583 17 2617 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
<< metal1 >>
rect 0 561 2668 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 0 496 2668 527
rect 0 17 2668 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
rect 0 -48 2668 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 2594 221 2628 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 2594 289 2628 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 bufbuf_16
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2668 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1977410
string GDS_START 1957960
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
