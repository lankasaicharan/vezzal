magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
<< pwell >>
rect 53 163 1086 247
rect 53 49 1191 163
rect 0 0 1248 49
<< scnmos >>
rect 132 137 162 221
rect 240 53 270 221
rect 338 53 368 221
rect 442 53 472 221
rect 528 53 558 221
rect 668 53 698 221
rect 754 53 784 221
rect 864 53 894 221
rect 950 53 980 221
rect 1082 53 1112 137
<< scpmoshvt >>
rect 132 367 162 451
rect 240 367 270 619
rect 330 367 360 619
rect 420 367 450 619
rect 528 367 558 619
rect 719 367 749 619
rect 805 367 835 619
rect 891 367 921 619
rect 977 367 1007 619
rect 1082 367 1112 451
<< ndiff >>
rect 79 196 132 221
rect 79 162 87 196
rect 121 162 132 196
rect 79 137 132 162
rect 162 192 240 221
rect 162 158 175 192
rect 209 158 240 192
rect 162 137 240 158
rect 187 99 240 137
rect 187 65 195 99
rect 229 65 240 99
rect 187 53 240 65
rect 270 206 338 221
rect 270 172 289 206
rect 323 172 338 206
rect 270 101 338 172
rect 270 67 288 101
rect 322 67 338 101
rect 270 53 338 67
rect 368 163 442 221
rect 368 129 389 163
rect 423 129 442 163
rect 368 95 442 129
rect 368 61 389 95
rect 423 61 442 95
rect 368 53 442 61
rect 472 209 528 221
rect 472 175 483 209
rect 517 175 528 209
rect 472 101 528 175
rect 472 67 483 101
rect 517 67 528 101
rect 472 53 528 67
rect 558 73 668 221
rect 558 53 592 73
rect 580 39 592 53
rect 626 53 668 73
rect 698 213 754 221
rect 698 179 709 213
rect 743 179 754 213
rect 698 53 754 179
rect 784 73 864 221
rect 784 53 807 73
rect 626 39 638 53
rect 580 31 638 39
rect 799 39 807 53
rect 841 53 864 73
rect 894 213 950 221
rect 894 179 905 213
rect 939 179 950 213
rect 894 53 950 179
rect 980 137 1060 221
rect 980 73 1082 137
rect 980 53 1014 73
rect 841 39 849 53
rect 799 27 849 39
rect 1002 39 1014 53
rect 1048 53 1082 73
rect 1112 112 1165 137
rect 1112 78 1123 112
rect 1157 78 1165 112
rect 1112 53 1165 78
rect 1048 39 1060 53
rect 1002 31 1060 39
<< pdiff >>
rect 187 607 240 619
rect 187 573 195 607
rect 229 573 240 607
rect 187 496 240 573
rect 187 462 195 496
rect 229 462 240 496
rect 187 451 240 462
rect 79 426 132 451
rect 79 392 87 426
rect 121 392 132 426
rect 79 367 132 392
rect 162 367 240 451
rect 270 367 330 619
rect 360 367 420 619
rect 450 367 528 619
rect 558 599 611 619
rect 558 565 569 599
rect 603 565 611 599
rect 558 505 611 565
rect 558 471 569 505
rect 603 471 611 505
rect 558 413 611 471
rect 558 379 569 413
rect 603 379 611 413
rect 558 367 611 379
rect 666 607 719 619
rect 666 573 674 607
rect 708 573 719 607
rect 666 529 719 573
rect 666 495 674 529
rect 708 495 719 529
rect 666 453 719 495
rect 666 419 674 453
rect 708 419 719 453
rect 666 367 719 419
rect 749 599 805 619
rect 749 565 760 599
rect 794 565 805 599
rect 749 502 805 565
rect 749 468 760 502
rect 794 468 805 502
rect 749 413 805 468
rect 749 379 760 413
rect 794 379 805 413
rect 749 367 805 379
rect 835 607 891 619
rect 835 573 846 607
rect 880 573 891 607
rect 835 528 891 573
rect 835 494 846 528
rect 880 494 891 528
rect 835 451 891 494
rect 835 417 846 451
rect 880 417 891 451
rect 835 367 891 417
rect 921 599 977 619
rect 921 565 932 599
rect 966 565 977 599
rect 921 502 977 565
rect 921 468 932 502
rect 966 468 977 502
rect 921 413 977 468
rect 921 379 932 413
rect 966 379 977 413
rect 921 367 977 379
rect 1007 607 1060 619
rect 1007 573 1018 607
rect 1052 573 1060 607
rect 1007 528 1060 573
rect 1007 494 1018 528
rect 1052 494 1060 528
rect 1007 451 1060 494
rect 1007 417 1018 451
rect 1052 417 1082 451
rect 1007 367 1082 417
rect 1112 426 1165 451
rect 1112 392 1123 426
rect 1157 392 1165 426
rect 1112 367 1165 392
<< ndiffc >>
rect 87 162 121 196
rect 175 158 209 192
rect 195 65 229 99
rect 289 172 323 206
rect 288 67 322 101
rect 389 129 423 163
rect 389 61 423 95
rect 483 175 517 209
rect 483 67 517 101
rect 592 39 626 73
rect 709 179 743 213
rect 807 39 841 73
rect 905 179 939 213
rect 1014 39 1048 73
rect 1123 78 1157 112
<< pdiffc >>
rect 195 573 229 607
rect 195 462 229 496
rect 87 392 121 426
rect 569 565 603 599
rect 569 471 603 505
rect 569 379 603 413
rect 674 573 708 607
rect 674 495 708 529
rect 674 419 708 453
rect 760 565 794 599
rect 760 468 794 502
rect 760 379 794 413
rect 846 573 880 607
rect 846 494 880 528
rect 846 417 880 451
rect 932 565 966 599
rect 932 468 966 502
rect 932 379 966 413
rect 1018 573 1052 607
rect 1018 494 1052 528
rect 1018 417 1052 451
rect 1123 392 1157 426
<< poly >>
rect 240 619 270 645
rect 330 619 360 645
rect 420 619 450 645
rect 528 619 558 645
rect 719 619 749 645
rect 805 619 835 645
rect 891 619 921 645
rect 977 619 1007 645
rect 132 451 162 477
rect 1082 451 1112 477
rect 132 309 162 367
rect 240 309 270 367
rect 330 335 360 367
rect 420 335 450 367
rect 21 293 162 309
rect 21 259 37 293
rect 71 259 162 293
rect 21 243 162 259
rect 204 293 270 309
rect 204 259 220 293
rect 254 259 270 293
rect 312 319 378 335
rect 312 285 328 319
rect 362 285 378 319
rect 312 269 378 285
rect 420 319 486 335
rect 420 285 436 319
rect 470 285 486 319
rect 420 269 486 285
rect 528 309 558 367
rect 719 331 749 367
rect 805 331 835 367
rect 891 331 921 367
rect 977 331 1007 367
rect 674 315 1007 331
rect 528 293 626 309
rect 674 295 690 315
rect 204 243 270 259
rect 132 221 162 243
rect 240 221 270 243
rect 338 221 368 269
rect 442 221 472 269
rect 528 259 576 293
rect 610 259 626 293
rect 528 243 626 259
rect 668 281 690 295
rect 724 281 758 315
rect 792 281 826 315
rect 860 281 894 315
rect 928 301 1007 315
rect 1082 325 1112 367
rect 1082 309 1227 325
rect 928 281 980 301
rect 668 265 980 281
rect 528 221 558 243
rect 668 221 698 265
rect 754 221 784 265
rect 864 221 894 265
rect 950 221 980 265
rect 1082 275 1177 309
rect 1211 275 1227 309
rect 1082 241 1227 275
rect 132 111 162 137
rect 240 27 270 53
rect 338 27 368 53
rect 442 27 472 53
rect 528 27 558 53
rect 668 27 698 53
rect 754 27 784 53
rect 1082 207 1177 241
rect 1211 207 1227 241
rect 1082 191 1227 207
rect 1082 137 1112 191
rect 864 27 894 53
rect 950 27 980 53
rect 1082 27 1112 53
<< polycont >>
rect 37 259 71 293
rect 220 259 254 293
rect 328 285 362 319
rect 436 285 470 319
rect 576 259 610 293
rect 690 281 724 315
rect 758 281 792 315
rect 826 281 860 315
rect 894 281 928 315
rect 1177 275 1211 309
rect 1177 207 1211 241
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 179 607 245 649
rect 179 573 195 607
rect 229 573 245 607
rect 179 496 245 573
rect 179 462 195 496
rect 229 462 245 496
rect 179 453 245 462
rect 553 599 619 615
rect 553 565 569 599
rect 603 565 619 599
rect 553 505 619 565
rect 553 471 569 505
rect 603 471 619 505
rect 71 426 137 442
rect 71 392 87 426
rect 121 419 137 426
rect 121 392 470 419
rect 71 385 470 392
rect 553 413 619 471
rect 658 607 724 649
rect 658 573 674 607
rect 708 573 724 607
rect 658 529 724 573
rect 658 495 674 529
rect 708 495 724 529
rect 658 453 724 495
rect 658 419 674 453
rect 708 419 724 453
rect 758 599 796 615
rect 758 565 760 599
rect 794 565 796 599
rect 758 502 796 565
rect 758 468 760 502
rect 794 468 796 502
rect 553 385 569 413
rect 71 384 141 385
rect 17 293 73 350
rect 17 259 37 293
rect 71 259 73 293
rect 17 242 73 259
rect 107 208 141 384
rect 204 293 271 351
rect 204 259 220 293
rect 254 259 271 293
rect 305 319 378 351
rect 305 285 328 319
rect 362 285 378 319
rect 305 269 378 285
rect 420 319 470 385
rect 420 285 436 319
rect 420 269 470 285
rect 506 379 569 385
rect 603 385 619 413
rect 758 413 796 468
rect 830 607 896 649
rect 830 573 846 607
rect 880 573 896 607
rect 830 528 896 573
rect 830 494 846 528
rect 880 494 896 528
rect 830 451 896 494
rect 830 417 846 451
rect 880 417 896 451
rect 930 599 968 615
rect 930 565 932 599
rect 966 565 968 599
rect 930 502 968 565
rect 930 468 932 502
rect 966 468 968 502
rect 603 379 708 385
rect 506 351 708 379
rect 204 242 271 259
rect 506 233 540 351
rect 660 315 708 351
rect 758 379 760 413
rect 794 383 796 413
rect 930 413 968 468
rect 1002 607 1068 649
rect 1002 573 1018 607
rect 1052 573 1068 607
rect 1002 528 1068 573
rect 1002 494 1018 528
rect 1052 494 1068 528
rect 1002 451 1068 494
rect 1002 417 1018 451
rect 1052 417 1068 451
rect 1102 426 1173 442
rect 930 383 932 413
rect 794 379 932 383
rect 966 383 968 413
rect 1102 392 1123 426
rect 1157 392 1173 426
rect 1102 384 1173 392
rect 966 379 1045 383
rect 758 349 1045 379
rect 305 209 540 233
rect 305 208 483 209
rect 71 196 141 208
rect 71 162 87 196
rect 121 162 141 196
rect 71 146 141 162
rect 175 192 239 208
rect 209 158 239 192
rect 175 99 239 158
rect 175 65 195 99
rect 229 65 239 99
rect 175 17 239 65
rect 273 206 483 208
rect 273 172 289 206
rect 323 199 483 206
rect 323 172 339 199
rect 273 101 339 172
rect 473 175 483 199
rect 517 175 540 209
rect 273 67 288 101
rect 322 67 339 101
rect 273 51 339 67
rect 373 129 389 163
rect 423 129 439 163
rect 373 95 439 129
rect 373 61 389 95
rect 423 61 439 95
rect 373 17 439 61
rect 473 101 540 175
rect 574 293 626 309
rect 574 259 576 293
rect 610 259 626 293
rect 660 281 690 315
rect 724 281 758 315
rect 792 281 826 315
rect 860 281 894 315
rect 928 281 944 315
rect 660 265 944 281
rect 574 145 626 259
rect 978 229 1045 349
rect 693 213 1045 229
rect 693 179 709 213
rect 743 179 905 213
rect 939 179 1045 213
rect 1102 145 1141 384
rect 1175 309 1231 350
rect 1175 275 1177 309
rect 1211 275 1231 309
rect 1175 241 1231 275
rect 1175 207 1177 241
rect 1211 207 1231 241
rect 1175 191 1231 207
rect 574 143 1141 145
rect 574 112 1173 143
rect 574 111 1123 112
rect 473 67 483 101
rect 517 67 540 101
rect 1107 78 1123 111
rect 1157 78 1173 112
rect 473 51 540 67
rect 576 73 642 77
rect 576 39 592 73
rect 626 39 642 73
rect 576 17 642 39
rect 791 73 857 77
rect 791 39 807 73
rect 841 39 857 73
rect 791 17 857 39
rect 998 73 1064 77
rect 998 39 1014 73
rect 1048 39 1064 73
rect 1107 62 1173 78
rect 998 17 1064 39
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or4bb_4
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6796874
string GDS_START 6787062
<< end >>
