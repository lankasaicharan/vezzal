magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 1 228 211 248
rect 1 49 863 228
rect 0 0 864 49
<< scnmos >>
rect 84 74 114 222
rect 296 74 326 202
rect 396 74 426 202
rect 510 74 540 202
rect 608 74 638 202
rect 750 74 780 202
<< scpmoshvt >>
rect 86 368 116 592
rect 306 397 336 565
rect 413 368 443 592
rect 497 368 527 592
rect 611 368 641 592
rect 725 368 755 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 184 185 222
rect 114 150 125 184
rect 159 150 185 184
rect 114 116 185 150
rect 114 82 125 116
rect 159 82 185 116
rect 114 74 185 82
rect 239 190 296 202
rect 239 156 251 190
rect 285 156 296 190
rect 239 120 296 156
rect 239 86 251 120
rect 285 86 296 120
rect 239 74 296 86
rect 326 188 396 202
rect 326 154 351 188
rect 385 154 396 188
rect 326 120 396 154
rect 326 86 351 120
rect 385 86 396 120
rect 326 74 396 86
rect 426 120 510 202
rect 426 86 451 120
rect 485 86 510 120
rect 426 74 510 86
rect 540 188 608 202
rect 540 154 551 188
rect 585 154 608 188
rect 540 120 608 154
rect 540 86 551 120
rect 585 86 608 120
rect 540 74 608 86
rect 638 120 750 202
rect 638 86 671 120
rect 705 86 750 120
rect 638 74 750 86
rect 780 190 837 202
rect 780 156 791 190
rect 825 156 837 190
rect 780 120 837 156
rect 780 86 791 120
rect 825 86 837 120
rect 780 74 837 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 508 86 546
rect 27 474 39 508
rect 73 474 86 508
rect 27 368 86 474
rect 116 580 273 592
rect 116 546 139 580
rect 173 546 225 580
rect 259 565 273 580
rect 354 565 413 592
rect 259 546 306 565
rect 116 492 306 546
rect 116 458 139 492
rect 173 458 258 492
rect 292 458 306 492
rect 116 397 306 458
rect 336 553 413 565
rect 336 519 366 553
rect 400 519 413 553
rect 336 443 413 519
rect 336 409 366 443
rect 400 409 413 443
rect 336 397 413 409
rect 116 368 169 397
rect 360 368 413 397
rect 443 368 497 592
rect 527 368 611 592
rect 641 368 725 592
rect 755 580 837 592
rect 755 546 768 580
rect 802 546 837 580
rect 755 498 837 546
rect 755 464 768 498
rect 802 464 837 498
rect 755 368 837 464
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 150 159 184
rect 125 82 159 116
rect 251 156 285 190
rect 251 86 285 120
rect 351 154 385 188
rect 351 86 385 120
rect 451 86 485 120
rect 551 154 585 188
rect 551 86 585 120
rect 671 86 705 120
rect 791 156 825 190
rect 791 86 825 120
<< pdiffc >>
rect 39 546 73 580
rect 39 474 73 508
rect 139 546 173 580
rect 225 546 259 580
rect 139 458 173 492
rect 258 458 292 492
rect 366 519 400 553
rect 366 409 400 443
rect 768 546 802 580
rect 768 464 802 498
<< poly >>
rect 86 592 116 618
rect 413 592 443 618
rect 497 592 527 618
rect 611 592 641 618
rect 725 592 755 618
rect 306 565 336 591
rect 306 382 336 397
rect 86 353 116 368
rect 83 336 119 353
rect 250 352 339 382
rect 413 353 443 368
rect 497 353 527 368
rect 611 353 641 368
rect 725 353 755 368
rect 250 340 326 352
rect 83 320 157 336
rect 83 286 107 320
rect 141 286 157 320
rect 250 306 266 340
rect 300 306 326 340
rect 250 290 326 306
rect 410 304 446 353
rect 83 270 157 286
rect 84 222 114 270
rect 296 202 326 290
rect 374 288 446 304
rect 374 254 390 288
rect 424 274 446 288
rect 494 310 530 353
rect 608 326 644 353
rect 722 336 758 353
rect 608 310 674 326
rect 494 294 560 310
rect 424 254 440 274
rect 374 238 440 254
rect 494 260 510 294
rect 544 260 560 294
rect 494 244 560 260
rect 608 276 624 310
rect 658 276 674 310
rect 608 260 674 276
rect 722 320 788 336
rect 722 286 738 320
rect 772 286 788 320
rect 722 270 788 286
rect 396 202 426 238
rect 510 202 540 244
rect 608 202 638 260
rect 750 202 780 270
rect 84 48 114 74
rect 296 48 326 74
rect 396 48 426 74
rect 510 48 540 74
rect 608 48 638 74
rect 750 48 780 74
<< polycont >>
rect 107 286 141 320
rect 266 306 300 340
rect 390 254 424 288
rect 510 260 544 294
rect 624 276 658 310
rect 738 286 772 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 508 89 546
rect 23 474 39 508
rect 73 474 89 508
rect 23 458 89 474
rect 123 580 308 649
rect 123 546 139 580
rect 173 546 225 580
rect 259 546 308 580
rect 752 580 841 649
rect 123 492 308 546
rect 123 458 139 492
rect 173 458 258 492
rect 292 458 308 492
rect 350 553 416 569
rect 350 519 366 553
rect 400 519 416 553
rect 23 226 57 458
rect 350 443 416 519
rect 350 424 366 443
rect 91 409 366 424
rect 400 409 416 443
rect 91 390 416 409
rect 91 320 157 390
rect 91 286 107 320
rect 141 286 157 320
rect 217 340 316 356
rect 217 306 266 340
rect 300 306 316 340
rect 217 290 316 306
rect 91 270 157 286
rect 123 256 157 270
rect 374 288 455 356
rect 23 210 75 226
rect 123 222 301 256
rect 374 254 390 288
rect 424 254 455 288
rect 374 238 455 254
rect 494 294 560 578
rect 494 260 510 294
rect 544 260 560 294
rect 601 310 674 578
rect 752 546 768 580
rect 802 546 841 580
rect 752 498 841 546
rect 752 464 768 498
rect 802 464 841 498
rect 601 276 624 310
rect 658 276 674 310
rect 601 260 674 276
rect 722 320 839 430
rect 722 286 738 320
rect 772 286 839 320
rect 722 270 839 286
rect 494 244 560 260
rect 23 176 39 210
rect 73 176 75 210
rect 235 190 301 222
rect 775 204 841 206
rect 23 120 75 176
rect 23 86 39 120
rect 73 86 75 120
rect 23 70 75 86
rect 109 184 189 188
rect 109 150 125 184
rect 159 150 189 184
rect 109 116 189 150
rect 109 82 125 116
rect 159 82 189 116
rect 109 17 189 82
rect 235 156 251 190
rect 285 156 301 190
rect 235 120 301 156
rect 235 86 251 120
rect 285 86 301 120
rect 235 70 301 86
rect 335 190 841 204
rect 335 188 791 190
rect 335 154 351 188
rect 385 170 551 188
rect 385 154 401 170
rect 335 120 401 154
rect 535 154 551 170
rect 585 170 791 188
rect 585 154 601 170
rect 335 86 351 120
rect 385 86 401 120
rect 335 70 401 86
rect 435 120 501 136
rect 435 86 451 120
rect 485 86 501 120
rect 435 17 501 86
rect 535 120 601 154
rect 775 156 791 170
rect 825 156 841 190
rect 535 86 551 120
rect 585 86 601 120
rect 535 70 601 86
rect 635 120 741 136
rect 635 86 671 120
rect 705 86 741 120
rect 635 17 741 86
rect 775 120 841 156
rect 775 86 791 120
rect 825 86 841 120
rect 775 70 841 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o41a_1
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 440794
string GDS_START 432522
<< end >>
