magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 331 1478 704
<< pwell >>
rect 5 49 1435 241
rect 0 0 1440 49
<< scnmos >>
rect 84 47 114 215
rect 170 47 200 215
rect 256 47 286 215
rect 342 47 372 215
rect 436 47 466 215
rect 522 47 552 215
rect 676 47 706 215
rect 763 47 793 215
rect 880 47 910 215
rect 966 47 996 215
rect 1064 47 1094 215
rect 1150 47 1180 215
rect 1236 47 1266 215
rect 1322 47 1352 215
<< scpmoshvt >>
rect 84 367 114 619
rect 170 367 200 619
rect 256 367 286 619
rect 350 367 380 619
rect 436 367 466 619
rect 522 367 552 619
rect 712 367 742 619
rect 798 367 828 619
rect 884 367 914 619
rect 970 367 1000 619
rect 1069 367 1099 619
rect 1157 367 1187 619
rect 1243 367 1273 619
rect 1329 367 1359 619
<< ndiff >>
rect 31 203 84 215
rect 31 169 39 203
rect 73 169 84 203
rect 31 93 84 169
rect 31 59 39 93
rect 73 59 84 93
rect 31 47 84 59
rect 114 203 170 215
rect 114 169 125 203
rect 159 169 170 203
rect 114 101 170 169
rect 114 67 125 101
rect 159 67 170 101
rect 114 47 170 67
rect 200 169 256 215
rect 200 135 211 169
rect 245 135 256 169
rect 200 47 256 135
rect 286 172 342 215
rect 286 138 297 172
rect 331 138 342 172
rect 286 93 342 138
rect 286 59 297 93
rect 331 59 342 93
rect 286 47 342 59
rect 372 163 436 215
rect 372 129 387 163
rect 421 129 436 163
rect 372 93 436 129
rect 372 59 387 93
rect 421 59 436 93
rect 372 47 436 59
rect 466 203 522 215
rect 466 169 477 203
rect 511 169 522 203
rect 466 101 522 169
rect 466 67 477 101
rect 511 67 522 101
rect 466 47 522 67
rect 552 104 676 215
rect 552 70 563 104
rect 597 70 631 104
rect 665 70 676 104
rect 552 47 676 70
rect 706 173 763 215
rect 706 139 717 173
rect 751 139 763 173
rect 706 101 763 139
rect 706 67 717 101
rect 751 67 763 101
rect 706 47 763 67
rect 793 95 880 215
rect 793 61 819 95
rect 853 61 880 95
rect 793 47 880 61
rect 910 172 966 215
rect 910 138 921 172
rect 955 138 966 172
rect 910 101 966 138
rect 910 67 921 101
rect 955 67 966 101
rect 910 47 966 67
rect 996 161 1064 215
rect 996 127 1011 161
rect 1045 127 1064 161
rect 996 93 1064 127
rect 996 59 1011 93
rect 1045 59 1064 93
rect 996 47 1064 59
rect 1094 203 1150 215
rect 1094 169 1105 203
rect 1139 169 1150 203
rect 1094 101 1150 169
rect 1094 67 1105 101
rect 1139 67 1150 101
rect 1094 47 1150 67
rect 1180 173 1236 215
rect 1180 139 1191 173
rect 1225 139 1236 173
rect 1180 89 1236 139
rect 1180 55 1191 89
rect 1225 55 1236 89
rect 1180 47 1236 55
rect 1266 203 1322 215
rect 1266 169 1277 203
rect 1311 169 1322 203
rect 1266 101 1322 169
rect 1266 67 1277 101
rect 1311 67 1322 101
rect 1266 47 1322 67
rect 1352 179 1409 215
rect 1352 145 1363 179
rect 1397 145 1409 179
rect 1352 89 1409 145
rect 1352 55 1363 89
rect 1397 55 1409 89
rect 1352 47 1409 55
<< pdiff >>
rect 27 599 84 619
rect 27 565 35 599
rect 69 565 84 599
rect 27 507 84 565
rect 27 473 35 507
rect 69 473 84 507
rect 27 413 84 473
rect 27 379 35 413
rect 69 379 84 413
rect 27 367 84 379
rect 114 568 170 619
rect 114 534 125 568
rect 159 534 170 568
rect 114 367 170 534
rect 200 599 256 619
rect 200 565 211 599
rect 245 565 256 599
rect 200 510 256 565
rect 200 476 211 510
rect 245 476 256 510
rect 200 367 256 476
rect 286 568 350 619
rect 286 534 301 568
rect 335 534 350 568
rect 286 367 350 534
rect 380 599 436 619
rect 380 565 391 599
rect 425 565 436 599
rect 380 507 436 565
rect 380 473 391 507
rect 425 473 436 507
rect 380 413 436 473
rect 380 379 391 413
rect 425 379 436 413
rect 380 367 436 379
rect 466 531 522 619
rect 466 497 477 531
rect 511 497 522 531
rect 466 413 522 497
rect 466 379 477 413
rect 511 379 522 413
rect 466 367 522 379
rect 552 607 605 619
rect 552 573 563 607
rect 597 573 605 607
rect 552 524 605 573
rect 552 490 563 524
rect 597 490 605 524
rect 552 367 605 490
rect 659 572 712 619
rect 659 538 667 572
rect 701 538 712 572
rect 659 367 712 538
rect 742 584 798 619
rect 742 550 753 584
rect 787 550 798 584
rect 742 367 798 550
rect 828 424 884 619
rect 828 390 839 424
rect 873 390 884 424
rect 828 367 884 390
rect 914 584 970 619
rect 914 550 925 584
rect 959 550 970 584
rect 914 367 970 550
rect 1000 572 1069 619
rect 1000 538 1020 572
rect 1054 538 1069 572
rect 1000 367 1069 538
rect 1099 599 1157 619
rect 1099 565 1112 599
rect 1146 565 1157 599
rect 1099 508 1157 565
rect 1099 474 1112 508
rect 1146 474 1157 508
rect 1099 409 1157 474
rect 1099 375 1112 409
rect 1146 375 1157 409
rect 1099 367 1157 375
rect 1187 607 1243 619
rect 1187 573 1198 607
rect 1232 573 1243 607
rect 1187 539 1243 573
rect 1187 505 1198 539
rect 1232 505 1243 539
rect 1187 469 1243 505
rect 1187 435 1198 469
rect 1232 435 1243 469
rect 1187 367 1243 435
rect 1273 599 1329 619
rect 1273 565 1284 599
rect 1318 565 1329 599
rect 1273 508 1329 565
rect 1273 474 1284 508
rect 1318 474 1329 508
rect 1273 409 1329 474
rect 1273 375 1284 409
rect 1318 375 1329 409
rect 1273 367 1329 375
rect 1359 607 1412 619
rect 1359 573 1370 607
rect 1404 573 1412 607
rect 1359 539 1412 573
rect 1359 505 1370 539
rect 1404 505 1412 539
rect 1359 469 1412 505
rect 1359 435 1370 469
rect 1404 435 1412 469
rect 1359 367 1412 435
<< ndiffc >>
rect 39 169 73 203
rect 39 59 73 93
rect 125 169 159 203
rect 125 67 159 101
rect 211 135 245 169
rect 297 138 331 172
rect 297 59 331 93
rect 387 129 421 163
rect 387 59 421 93
rect 477 169 511 203
rect 477 67 511 101
rect 563 70 597 104
rect 631 70 665 104
rect 717 139 751 173
rect 717 67 751 101
rect 819 61 853 95
rect 921 138 955 172
rect 921 67 955 101
rect 1011 127 1045 161
rect 1011 59 1045 93
rect 1105 169 1139 203
rect 1105 67 1139 101
rect 1191 139 1225 173
rect 1191 55 1225 89
rect 1277 169 1311 203
rect 1277 67 1311 101
rect 1363 145 1397 179
rect 1363 55 1397 89
<< pdiffc >>
rect 35 565 69 599
rect 35 473 69 507
rect 35 379 69 413
rect 125 534 159 568
rect 211 565 245 599
rect 211 476 245 510
rect 301 534 335 568
rect 391 565 425 599
rect 391 473 425 507
rect 391 379 425 413
rect 477 497 511 531
rect 477 379 511 413
rect 563 573 597 607
rect 563 490 597 524
rect 667 538 701 572
rect 753 550 787 584
rect 839 390 873 424
rect 925 550 959 584
rect 1020 538 1054 572
rect 1112 565 1146 599
rect 1112 474 1146 508
rect 1112 375 1146 409
rect 1198 573 1232 607
rect 1198 505 1232 539
rect 1198 435 1232 469
rect 1284 565 1318 599
rect 1284 474 1318 508
rect 1284 375 1318 409
rect 1370 573 1404 607
rect 1370 505 1404 539
rect 1370 435 1404 469
<< poly >>
rect 84 619 114 645
rect 170 619 200 645
rect 256 619 286 645
rect 350 619 380 645
rect 436 619 466 645
rect 522 619 552 645
rect 712 619 742 645
rect 798 619 828 645
rect 884 619 914 645
rect 970 619 1000 645
rect 1069 619 1099 645
rect 1157 619 1187 645
rect 1243 619 1273 645
rect 1329 619 1359 645
rect 84 335 114 367
rect 48 319 114 335
rect 48 285 64 319
rect 98 285 114 319
rect 48 269 114 285
rect 84 215 114 269
rect 170 335 200 367
rect 256 335 286 367
rect 350 335 380 367
rect 170 319 286 335
rect 170 285 195 319
rect 229 285 286 319
rect 170 269 286 285
rect 328 319 394 335
rect 328 285 344 319
rect 378 285 394 319
rect 328 269 394 285
rect 436 285 466 367
rect 522 321 552 367
rect 712 345 742 367
rect 522 305 601 321
rect 522 285 551 305
rect 436 271 551 285
rect 585 271 601 305
rect 685 315 742 345
rect 798 333 828 367
rect 884 333 914 367
rect 793 317 914 333
rect 685 303 715 315
rect 170 215 200 269
rect 256 215 286 269
rect 342 215 372 269
rect 436 255 601 271
rect 649 287 715 303
rect 436 215 466 255
rect 522 215 552 255
rect 649 253 665 287
rect 699 253 715 287
rect 793 283 809 317
rect 843 303 914 317
rect 970 303 1000 367
rect 1069 331 1099 367
rect 1157 331 1187 367
rect 1243 331 1273 367
rect 1329 331 1359 367
rect 1069 315 1359 331
rect 843 283 910 303
rect 793 267 910 283
rect 649 237 715 253
rect 763 237 910 267
rect 956 287 1022 303
rect 1069 295 1085 315
rect 956 253 972 287
rect 1006 253 1022 287
rect 956 237 1022 253
rect 1064 281 1085 295
rect 1119 281 1153 315
rect 1187 281 1221 315
rect 1255 281 1289 315
rect 1323 281 1359 315
rect 1064 265 1359 281
rect 676 215 706 237
rect 763 215 793 237
rect 880 215 910 237
rect 966 215 996 237
rect 1064 215 1094 265
rect 1150 215 1180 265
rect 1236 215 1266 265
rect 1322 215 1352 265
rect 84 21 114 47
rect 170 21 200 47
rect 256 21 286 47
rect 342 21 372 47
rect 436 21 466 47
rect 522 21 552 47
rect 676 21 706 47
rect 763 21 793 47
rect 880 21 910 47
rect 966 21 996 47
rect 1064 21 1094 47
rect 1150 21 1180 47
rect 1236 21 1266 47
rect 1322 21 1352 47
<< polycont >>
rect 64 285 98 319
rect 195 285 229 319
rect 344 285 378 319
rect 551 271 585 305
rect 665 253 699 287
rect 809 283 843 317
rect 972 253 1006 287
rect 1085 281 1119 315
rect 1153 281 1187 315
rect 1221 281 1255 315
rect 1289 281 1323 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 19 599 75 615
rect 19 565 35 599
rect 69 565 75 599
rect 19 507 75 565
rect 109 568 175 649
rect 109 534 125 568
rect 159 534 175 568
rect 109 526 175 534
rect 209 599 251 615
rect 209 565 211 599
rect 245 565 251 599
rect 19 473 35 507
rect 69 492 75 507
rect 209 510 251 565
rect 285 568 351 649
rect 285 534 301 568
rect 335 534 351 568
rect 285 526 351 534
rect 387 607 613 615
rect 387 599 563 607
rect 387 565 391 599
rect 425 581 563 599
rect 425 565 435 581
rect 209 492 211 510
rect 69 476 211 492
rect 245 492 251 510
rect 387 507 435 565
rect 547 573 563 581
rect 597 573 613 607
rect 387 492 391 507
rect 245 476 391 492
rect 69 473 391 476
rect 425 473 435 507
rect 19 458 435 473
rect 19 413 75 458
rect 19 379 35 413
rect 69 379 75 413
rect 19 363 75 379
rect 109 390 327 424
rect 109 329 143 390
rect 48 319 143 329
rect 48 285 64 319
rect 98 285 143 319
rect 48 269 143 285
rect 179 319 259 356
rect 179 285 195 319
rect 229 285 259 319
rect 179 281 259 285
rect 293 329 327 390
rect 387 413 435 458
rect 387 379 391 413
rect 425 379 435 413
rect 387 363 435 379
rect 469 531 513 547
rect 469 497 477 531
rect 511 497 513 531
rect 469 454 513 497
rect 547 524 613 573
rect 651 572 717 649
rect 651 538 667 572
rect 701 538 717 572
rect 651 530 717 538
rect 751 584 970 600
rect 751 550 753 584
rect 787 550 925 584
rect 959 550 970 584
rect 751 534 970 550
rect 1004 572 1070 649
rect 1004 538 1020 572
rect 1054 538 1070 572
rect 1004 530 1070 538
rect 1110 599 1148 615
rect 1110 565 1112 599
rect 1146 565 1148 599
rect 547 490 563 524
rect 597 490 613 524
rect 1110 508 1148 565
rect 547 488 613 490
rect 647 462 1076 496
rect 647 454 681 462
rect 469 420 681 454
rect 715 424 889 428
rect 469 413 513 420
rect 469 379 477 413
rect 511 379 513 413
rect 715 390 839 424
rect 873 390 889 424
rect 715 386 889 390
rect 293 319 394 329
rect 293 285 344 319
rect 378 285 394 319
rect 293 281 394 285
rect 469 247 513 379
rect 23 203 80 219
rect 23 169 39 203
rect 73 169 80 203
rect 23 93 80 169
rect 23 59 39 93
rect 73 59 80 93
rect 23 17 80 59
rect 114 203 170 219
rect 114 169 125 203
rect 159 169 170 203
rect 114 101 170 169
rect 204 213 513 247
rect 204 169 247 213
rect 473 203 513 213
rect 204 135 211 169
rect 245 135 247 169
rect 204 119 247 135
rect 281 172 347 179
rect 281 138 297 172
rect 331 138 347 172
rect 114 67 125 101
rect 159 85 170 101
rect 281 93 347 138
rect 281 85 297 93
rect 159 67 297 85
rect 114 59 297 67
rect 331 59 347 93
rect 114 51 347 59
rect 381 163 437 179
rect 381 129 387 163
rect 421 129 437 163
rect 381 93 437 129
rect 381 59 387 93
rect 421 59 437 93
rect 381 17 437 59
rect 473 169 477 203
rect 511 169 513 203
rect 473 101 513 169
rect 551 352 749 386
rect 551 305 585 352
rect 793 317 859 350
rect 551 179 585 271
rect 649 253 665 287
rect 699 253 715 287
rect 793 283 809 317
rect 843 283 859 317
rect 1042 317 1076 462
rect 1110 474 1112 508
rect 1146 474 1148 508
rect 1110 409 1148 474
rect 1182 607 1248 649
rect 1182 573 1198 607
rect 1232 573 1248 607
rect 1182 539 1248 573
rect 1182 505 1198 539
rect 1232 505 1248 539
rect 1182 469 1248 505
rect 1182 435 1198 469
rect 1232 435 1248 469
rect 1182 419 1248 435
rect 1282 599 1326 615
rect 1282 565 1284 599
rect 1318 565 1326 599
rect 1282 508 1326 565
rect 1282 474 1284 508
rect 1318 474 1326 508
rect 1110 375 1112 409
rect 1146 385 1148 409
rect 1282 409 1326 474
rect 1360 607 1420 649
rect 1360 573 1370 607
rect 1404 573 1420 607
rect 1360 539 1420 573
rect 1360 505 1370 539
rect 1404 505 1420 539
rect 1360 469 1420 505
rect 1360 435 1370 469
rect 1404 435 1420 469
rect 1360 419 1420 435
rect 1282 385 1284 409
rect 1146 375 1284 385
rect 1318 385 1326 409
rect 1318 375 1409 385
rect 1110 351 1409 375
rect 1042 315 1339 317
rect 895 287 1008 303
rect 649 247 715 253
rect 895 253 972 287
rect 1006 253 1008 287
rect 1042 281 1085 315
rect 1119 281 1153 315
rect 1187 281 1221 315
rect 1255 281 1289 315
rect 1323 281 1339 315
rect 895 247 1008 253
rect 1375 247 1409 351
rect 649 213 1008 247
rect 1095 213 1409 247
rect 1095 203 1141 213
rect 551 173 971 179
rect 551 145 717 173
rect 715 139 717 145
rect 751 172 971 173
rect 751 145 921 172
rect 751 139 767 145
rect 473 67 477 101
rect 511 67 513 101
rect 473 51 513 67
rect 547 104 681 111
rect 547 70 563 104
rect 597 70 631 104
rect 665 70 681 104
rect 547 17 681 70
rect 715 101 767 139
rect 905 138 921 145
rect 955 138 971 172
rect 715 67 717 101
rect 751 67 767 101
rect 715 51 767 67
rect 803 95 869 111
rect 803 61 819 95
rect 853 61 869 95
rect 803 17 869 61
rect 905 101 971 138
rect 905 67 921 101
rect 955 67 971 101
rect 905 51 971 67
rect 1005 161 1061 177
rect 1005 127 1011 161
rect 1045 127 1061 161
rect 1005 93 1061 127
rect 1005 59 1011 93
rect 1045 59 1061 93
rect 1005 17 1061 59
rect 1095 169 1105 203
rect 1139 169 1141 203
rect 1275 203 1313 213
rect 1095 101 1141 169
rect 1095 67 1105 101
rect 1139 67 1141 101
rect 1095 51 1141 67
rect 1175 139 1191 173
rect 1225 139 1241 173
rect 1175 89 1241 139
rect 1175 55 1191 89
rect 1225 55 1241 89
rect 1175 17 1241 55
rect 1275 169 1277 203
rect 1311 169 1313 203
rect 1275 101 1313 169
rect 1275 67 1277 101
rect 1311 67 1313 101
rect 1275 51 1313 67
rect 1347 145 1363 179
rect 1397 145 1413 179
rect 1347 89 1413 145
rect 1347 55 1363 89
rect 1397 55 1413 89
rect 1347 17 1413 55
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2bb2o_4
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6017308
string GDS_START 6005574
<< end >>
