magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 288 248 671 259
rect 1 49 671 248
rect 0 0 672 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 273 368 309 592
rect 364 368 400 592
rect 463 368 499 592
rect 553 368 589 592
<< nmoslvt >>
rect 81 74 111 222
rect 167 74 197 222
rect 253 74 283 222
rect 364 85 394 233
rect 450 85 480 233
rect 561 85 591 233
<< ndiff >>
rect 314 222 364 233
rect 27 196 81 222
rect 27 162 36 196
rect 70 162 81 196
rect 27 120 81 162
rect 27 86 36 120
rect 70 86 81 120
rect 27 74 81 86
rect 111 116 167 222
rect 111 82 122 116
rect 156 82 167 116
rect 111 74 167 82
rect 197 184 253 222
rect 197 150 208 184
rect 242 150 253 184
rect 197 116 253 150
rect 197 82 208 116
rect 242 82 253 116
rect 197 74 253 82
rect 283 85 364 222
rect 394 221 450 233
rect 394 187 405 221
rect 439 187 450 221
rect 394 85 450 187
rect 480 85 561 233
rect 591 221 645 233
rect 591 187 602 221
rect 636 187 645 221
rect 591 131 645 187
rect 591 97 602 131
rect 636 97 645 131
rect 591 85 645 97
rect 283 74 307 85
rect 298 51 307 74
rect 341 51 349 85
rect 298 39 349 51
rect 495 51 503 85
rect 537 51 546 85
rect 495 39 546 51
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 497 173 546
rect 119 463 129 497
rect 163 463 173 497
rect 119 414 173 463
rect 119 380 129 414
rect 163 380 173 414
rect 119 368 173 380
rect 209 576 273 592
rect 209 542 229 576
rect 263 542 273 576
rect 209 368 273 542
rect 309 580 364 592
rect 309 546 319 580
rect 353 546 364 580
rect 309 499 364 546
rect 309 465 319 499
rect 353 465 364 499
rect 309 368 364 465
rect 400 576 463 592
rect 400 542 419 576
rect 453 542 463 576
rect 400 368 463 542
rect 499 580 553 592
rect 499 546 509 580
rect 543 546 553 580
rect 499 492 553 546
rect 499 458 509 492
rect 543 458 553 492
rect 499 368 553 458
rect 589 580 645 592
rect 589 546 599 580
rect 633 546 645 580
rect 589 497 645 546
rect 589 463 599 497
rect 633 463 645 497
rect 589 414 645 463
rect 589 380 599 414
rect 633 380 645 414
rect 589 368 645 380
<< ndiffc >>
rect 36 162 70 196
rect 36 86 70 120
rect 122 82 156 116
rect 208 150 242 184
rect 208 82 242 116
rect 405 187 439 221
rect 602 187 636 221
rect 602 97 636 131
rect 307 51 341 85
rect 503 51 537 85
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 229 542 263 576
rect 319 546 353 580
rect 319 465 353 499
rect 419 542 453 576
rect 509 546 543 580
rect 509 458 543 492
rect 599 546 633 580
rect 599 463 633 497
rect 599 380 633 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 273 592 309 618
rect 364 592 400 618
rect 463 592 499 618
rect 553 592 589 618
rect 83 310 119 368
rect 173 310 209 368
rect 273 336 309 368
rect 364 336 400 368
rect 463 336 499 368
rect 253 320 319 336
rect 81 294 203 310
rect 81 260 97 294
rect 131 260 203 294
rect 81 244 203 260
rect 253 286 269 320
rect 303 286 319 320
rect 253 270 319 286
rect 364 320 499 336
rect 553 330 589 368
rect 364 286 409 320
rect 443 286 499 320
rect 364 270 499 286
rect 547 314 613 330
rect 547 280 563 314
rect 597 280 613 314
rect 81 222 111 244
rect 167 222 197 244
rect 253 222 283 270
rect 364 233 394 270
rect 450 233 480 270
rect 547 264 613 280
rect 561 233 591 264
rect 81 48 111 74
rect 167 48 197 74
rect 253 48 283 74
rect 364 59 394 85
rect 450 59 480 85
rect 561 59 591 85
<< polycont >>
rect 97 260 131 294
rect 269 286 303 320
rect 409 286 443 320
rect 563 280 597 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 497 179 546
rect 213 576 263 649
rect 213 542 229 576
rect 213 526 263 542
rect 303 580 369 596
rect 303 546 319 580
rect 353 546 369 580
rect 113 463 129 497
rect 163 492 179 497
rect 303 499 369 546
rect 403 576 469 649
rect 403 542 419 576
rect 453 542 469 576
rect 403 526 469 542
rect 505 580 559 596
rect 505 546 509 580
rect 543 546 559 580
rect 303 492 319 499
rect 163 465 319 492
rect 353 492 369 499
rect 505 492 559 546
rect 353 465 509 492
rect 163 463 509 465
rect 113 458 509 463
rect 543 458 559 492
rect 599 580 649 649
rect 633 546 649 580
rect 599 497 649 546
rect 633 463 649 497
rect 113 414 219 458
rect 113 380 129 414
rect 163 380 219 414
rect 113 364 219 380
rect 25 294 147 310
rect 25 260 97 294
rect 131 260 147 294
rect 25 236 147 260
rect 185 252 219 364
rect 285 390 565 424
rect 285 336 359 390
rect 253 320 359 336
rect 253 286 269 320
rect 303 310 359 320
rect 393 320 459 356
rect 303 286 319 310
rect 393 286 409 320
rect 443 286 459 320
rect 531 330 565 390
rect 599 414 649 463
rect 633 380 649 414
rect 599 364 649 380
rect 531 314 613 330
rect 531 280 563 314
rect 597 280 613 314
rect 531 264 613 280
rect 185 221 455 252
rect 185 218 405 221
rect 20 196 86 202
rect 20 162 36 196
rect 70 184 86 196
rect 389 187 405 218
rect 439 187 455 221
rect 586 221 652 230
rect 586 187 602 221
rect 636 187 652 221
rect 70 162 208 184
rect 20 150 208 162
rect 242 153 274 184
rect 586 153 652 187
rect 242 150 652 153
rect 20 120 70 150
rect 20 86 36 120
rect 208 131 652 150
rect 208 119 602 131
rect 208 116 242 119
rect 20 70 70 86
rect 106 82 122 116
rect 156 82 172 116
rect 106 17 172 82
rect 589 97 602 119
rect 636 97 652 131
rect 208 66 242 82
rect 291 51 307 85
rect 341 51 503 85
rect 537 51 553 85
rect 589 81 652 97
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand3_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 286964
string GDS_START 280528
<< end >>
