magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2126 1852
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 793 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 185 47 215 177
rect 287 93 317 177
rect 495 47 525 177
rect 591 47 621 177
rect 675 47 705 177
<< scpmoshvt >>
rect 81 297 117 497
rect 177 297 213 497
rect 289 297 325 381
rect 487 297 523 497
rect 583 297 619 497
rect 677 297 713 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 165 185 177
rect 109 131 130 165
rect 164 131 185 165
rect 109 97 185 131
rect 109 63 130 97
rect 164 63 185 97
rect 109 47 185 63
rect 215 157 287 177
rect 215 123 230 157
rect 264 123 287 157
rect 215 93 287 123
rect 317 165 379 177
rect 317 131 337 165
rect 371 131 379 165
rect 317 93 379 131
rect 433 93 495 177
rect 215 89 272 93
rect 215 55 226 89
rect 260 55 272 89
rect 215 47 272 55
rect 433 59 441 93
rect 475 59 495 93
rect 433 47 495 59
rect 525 163 591 177
rect 525 129 538 163
rect 572 129 591 163
rect 525 47 591 129
rect 621 47 675 177
rect 705 165 767 177
rect 705 131 725 165
rect 759 131 767 165
rect 705 47 767 131
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 297 81 451
rect 117 469 177 497
rect 117 435 130 469
rect 164 435 177 469
rect 117 401 177 435
rect 117 367 130 401
rect 164 367 177 401
rect 117 297 177 367
rect 213 489 302 497
rect 213 455 244 489
rect 278 455 302 489
rect 213 435 302 455
rect 433 439 487 497
rect 213 381 272 435
rect 433 405 441 439
rect 475 405 487 439
rect 213 297 289 381
rect 325 345 379 381
rect 325 311 337 345
rect 371 311 379 345
rect 325 297 379 311
rect 433 371 487 405
rect 433 337 441 371
rect 475 337 487 371
rect 433 297 487 337
rect 523 485 583 497
rect 523 451 535 485
rect 569 451 583 485
rect 523 417 583 451
rect 523 383 535 417
rect 569 383 583 417
rect 523 297 583 383
rect 619 489 677 497
rect 619 455 631 489
rect 665 455 677 489
rect 619 297 677 455
rect 713 485 767 497
rect 713 451 725 485
rect 759 451 767 485
rect 713 417 767 451
rect 713 383 725 417
rect 759 383 767 417
rect 713 297 767 383
<< ndiffc >>
rect 35 59 69 93
rect 130 131 164 165
rect 130 63 164 97
rect 230 123 264 157
rect 337 131 371 165
rect 226 55 260 89
rect 441 59 475 93
rect 538 129 572 163
rect 725 131 759 165
<< pdiffc >>
rect 35 451 69 485
rect 130 435 164 469
rect 130 367 164 401
rect 244 455 278 489
rect 441 405 475 439
rect 337 311 371 345
rect 441 337 475 371
rect 535 451 569 485
rect 535 383 569 417
rect 631 455 665 489
rect 725 451 759 485
rect 725 383 759 417
<< poly >>
rect 81 497 117 523
rect 177 497 213 523
rect 487 497 523 523
rect 583 497 619 523
rect 677 497 713 523
rect 289 381 325 407
rect 81 282 117 297
rect 177 282 213 297
rect 289 282 325 297
rect 487 282 523 297
rect 583 282 619 297
rect 677 282 713 297
rect 79 259 119 282
rect 175 259 215 282
rect 79 249 215 259
rect 79 215 140 249
rect 174 215 215 249
rect 79 205 215 215
rect 79 177 109 205
rect 185 177 215 205
rect 287 265 327 282
rect 485 265 525 282
rect 581 265 621 282
rect 287 249 341 265
rect 287 215 297 249
rect 331 215 341 249
rect 287 199 341 215
rect 421 249 525 265
rect 421 215 431 249
rect 465 215 525 249
rect 287 177 317 199
rect 421 198 525 215
rect 567 249 621 265
rect 567 215 577 249
rect 611 215 621 249
rect 567 199 621 215
rect 495 177 525 198
rect 591 177 621 199
rect 675 265 715 282
rect 675 249 729 265
rect 675 215 685 249
rect 719 215 729 249
rect 675 199 729 215
rect 675 177 705 199
rect 287 67 317 93
rect 79 21 109 47
rect 185 21 215 47
rect 495 21 525 47
rect 591 21 621 47
rect 675 21 705 47
<< polycont >>
rect 140 215 174 249
rect 297 215 331 249
rect 431 215 465 249
rect 577 215 611 249
rect 685 215 719 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 485 85 527
rect 228 489 294 527
rect 18 451 35 485
rect 69 451 85 485
rect 129 469 180 485
rect 129 435 130 469
rect 164 435 180 469
rect 228 455 244 489
rect 278 455 294 489
rect 129 401 180 435
rect 425 439 475 493
rect 425 421 441 439
rect 22 367 130 401
rect 164 367 180 401
rect 243 405 441 421
rect 243 379 475 405
rect 22 177 76 367
rect 243 333 277 379
rect 441 371 475 379
rect 124 299 277 333
rect 311 311 337 345
rect 371 311 407 345
rect 124 249 190 299
rect 373 265 407 311
rect 509 485 585 493
rect 509 451 535 485
rect 569 451 585 485
rect 509 417 585 451
rect 631 489 665 527
rect 631 437 665 455
rect 699 485 775 493
rect 699 451 725 485
rect 759 451 775 485
rect 509 383 535 417
rect 569 403 585 417
rect 699 417 775 451
rect 699 403 725 417
rect 569 383 725 403
rect 759 383 775 417
rect 509 369 775 383
rect 441 335 475 337
rect 441 301 543 335
rect 124 215 140 249
rect 174 215 190 249
rect 245 249 339 265
rect 245 215 297 249
rect 331 215 339 249
rect 245 199 339 215
rect 373 249 465 265
rect 373 215 431 249
rect 373 199 465 215
rect 22 165 180 177
rect 373 165 407 199
rect 22 143 130 165
rect 104 131 130 143
rect 164 131 180 165
rect 18 93 69 109
rect 18 59 35 93
rect 104 97 180 131
rect 104 63 130 97
rect 164 63 180 97
rect 214 123 230 157
rect 264 123 280 157
rect 321 131 337 165
rect 371 131 407 165
rect 499 165 543 301
rect 577 249 617 323
rect 611 215 617 249
rect 577 199 617 215
rect 675 249 733 323
rect 675 215 685 249
rect 719 215 733 249
rect 675 199 733 215
rect 499 163 588 165
rect 499 129 538 163
rect 572 129 588 163
rect 499 127 588 129
rect 699 131 725 165
rect 759 131 775 165
rect 214 89 280 123
rect 18 17 69 59
rect 214 55 226 89
rect 260 55 280 89
rect 214 17 280 55
rect 425 59 441 93
rect 475 59 491 93
rect 425 17 491 59
rect 699 17 775 131
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 245 199 339 265 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 684 221 718 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 30 357 64 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 582 289 616 323 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21bo_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1603388
string GDS_START 1596804
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
