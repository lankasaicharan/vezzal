magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3230 1852
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 201 1533 203
rect 1 23 1910 201
rect 1 21 309 23
rect 797 21 1007 23
rect 1448 21 1910 23
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 183 47 213 177
rect 298 93 328 177
rect 541 49 571 177
rect 629 49 659 177
rect 901 47 931 177
rect 1097 49 1127 177
rect 1258 49 1288 133
rect 1417 49 1447 177
rect 1556 47 1586 167
rect 1667 47 1697 175
rect 1751 47 1781 175
<< scpmoshvt >>
rect 81 297 117 497
rect 179 297 215 497
rect 300 297 336 425
rect 520 325 556 493
rect 627 297 663 465
rect 849 297 885 497
rect 1089 297 1125 465
rect 1250 297 1286 425
rect 1419 329 1455 457
rect 1548 329 1584 497
rect 1659 297 1695 497
rect 1753 297 1789 497
<< ndiff >>
rect 27 129 79 177
rect 27 95 35 129
rect 69 95 79 129
rect 27 47 79 95
rect 109 129 183 177
rect 109 95 133 129
rect 167 95 183 129
rect 109 47 183 95
rect 213 93 298 177
rect 328 169 423 177
rect 328 135 377 169
rect 411 135 423 169
rect 328 93 423 135
rect 477 165 541 177
rect 477 131 487 165
rect 521 131 541 165
rect 213 89 283 93
rect 213 55 231 89
rect 265 55 283 89
rect 213 47 283 55
rect 477 49 541 131
rect 571 91 629 177
rect 571 57 583 91
rect 617 57 629 91
rect 571 49 629 57
rect 659 91 739 177
rect 659 57 693 91
rect 727 57 739 91
rect 659 49 739 57
rect 823 157 901 177
rect 823 123 837 157
rect 871 123 901 157
rect 823 89 901 123
rect 823 55 837 89
rect 871 55 901 89
rect 823 47 901 55
rect 931 165 983 177
rect 931 131 941 165
rect 975 131 983 165
rect 931 124 983 131
rect 931 47 981 124
rect 1037 104 1097 177
rect 1035 97 1097 104
rect 1035 63 1043 97
rect 1077 63 1097 97
rect 1035 49 1097 63
rect 1127 133 1227 177
rect 1313 169 1417 177
rect 1313 135 1359 169
rect 1393 135 1417 169
rect 1313 133 1417 135
rect 1127 126 1258 133
rect 1127 92 1137 126
rect 1171 92 1258 126
rect 1127 49 1258 92
rect 1288 49 1417 133
rect 1447 167 1507 177
rect 1607 167 1667 175
rect 1447 93 1556 167
rect 1447 59 1469 93
rect 1503 59 1556 93
rect 1447 49 1556 59
rect 1474 47 1556 49
rect 1586 142 1667 167
rect 1586 108 1613 142
rect 1647 108 1667 142
rect 1586 47 1667 108
rect 1697 97 1751 175
rect 1697 63 1707 97
rect 1741 63 1751 97
rect 1697 47 1751 63
rect 1781 101 1884 175
rect 1781 67 1837 101
rect 1871 67 1884 101
rect 1781 47 1884 67
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 477 179 497
rect 117 443 133 477
rect 167 443 179 477
rect 117 409 179 443
rect 117 375 133 409
rect 167 375 179 409
rect 117 341 179 375
rect 117 307 133 341
rect 167 307 179 341
rect 117 297 179 307
rect 215 477 283 497
rect 215 443 236 477
rect 270 443 283 477
rect 215 425 283 443
rect 215 297 300 425
rect 336 341 394 425
rect 336 307 348 341
rect 382 307 394 341
rect 453 413 520 493
rect 453 379 474 413
rect 508 379 520 413
rect 453 325 520 379
rect 556 481 610 493
rect 556 447 568 481
rect 602 465 610 481
rect 795 481 849 497
rect 602 447 627 465
rect 556 325 627 447
rect 336 297 394 307
rect 575 297 627 325
rect 663 423 741 465
rect 795 447 803 481
rect 837 447 849 481
rect 795 435 849 447
rect 663 339 742 423
rect 663 305 696 339
rect 730 305 742 339
rect 663 297 742 305
rect 796 297 849 435
rect 885 343 949 497
rect 1488 489 1548 497
rect 885 309 897 343
rect 931 309 949 343
rect 885 297 949 309
rect 1003 405 1089 465
rect 1003 371 1011 405
rect 1045 371 1089 405
rect 1003 297 1089 371
rect 1125 425 1226 465
rect 1488 457 1500 489
rect 1348 425 1419 457
rect 1125 409 1250 425
rect 1125 375 1177 409
rect 1211 375 1250 409
rect 1125 341 1250 375
rect 1125 307 1177 341
rect 1211 307 1250 341
rect 1125 297 1250 307
rect 1286 390 1419 425
rect 1286 356 1359 390
rect 1393 356 1419 390
rect 1286 329 1419 356
rect 1455 455 1500 457
rect 1534 455 1548 489
rect 1455 329 1548 455
rect 1584 341 1659 497
rect 1584 329 1613 341
rect 1286 297 1383 329
rect 1601 307 1613 329
rect 1647 307 1659 341
rect 1601 297 1659 307
rect 1695 489 1753 497
rect 1695 455 1707 489
rect 1741 455 1753 489
rect 1695 297 1753 455
rect 1789 477 1884 497
rect 1789 443 1838 477
rect 1872 443 1884 477
rect 1789 409 1884 443
rect 1789 375 1839 409
rect 1873 375 1884 409
rect 1789 297 1884 375
<< ndiffc >>
rect 35 95 69 129
rect 133 95 167 129
rect 377 135 411 169
rect 487 131 521 165
rect 231 55 265 89
rect 583 57 617 91
rect 693 57 727 91
rect 837 123 871 157
rect 837 55 871 89
rect 941 131 975 165
rect 1043 63 1077 97
rect 1359 135 1393 169
rect 1137 92 1171 126
rect 1469 59 1503 93
rect 1613 108 1647 142
rect 1707 63 1741 97
rect 1837 67 1871 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 133 443 167 477
rect 133 375 167 409
rect 133 307 167 341
rect 236 443 270 477
rect 348 307 382 341
rect 474 379 508 413
rect 568 447 602 481
rect 803 447 837 481
rect 696 305 730 339
rect 897 309 931 343
rect 1011 371 1045 405
rect 1177 375 1211 409
rect 1177 307 1211 341
rect 1359 356 1393 390
rect 1500 455 1534 489
rect 1613 307 1647 341
rect 1707 455 1741 489
rect 1838 443 1872 477
rect 1839 375 1873 409
<< poly >>
rect 81 497 117 523
rect 179 497 215 523
rect 520 493 556 519
rect 298 451 338 483
rect 300 425 336 451
rect 627 465 663 504
rect 849 497 885 523
rect 520 310 556 325
rect 81 282 117 297
rect 179 282 215 297
rect 300 282 336 297
rect 79 265 119 282
rect 177 265 217 282
rect 298 265 338 282
rect 518 271 558 310
rect 1087 493 1457 523
rect 1548 497 1584 523
rect 1659 497 1695 523
rect 1753 497 1789 523
rect 1087 491 1127 493
rect 1089 465 1125 491
rect 1417 483 1457 493
rect 1419 457 1455 483
rect 1250 425 1286 451
rect 1419 314 1455 329
rect 1548 314 1584 329
rect 627 282 663 297
rect 849 282 885 297
rect 1089 282 1125 297
rect 1250 282 1286 297
rect 518 265 571 271
rect 625 265 665 282
rect 79 249 256 265
rect 79 215 212 249
rect 246 215 256 249
rect 79 199 256 215
rect 298 249 571 265
rect 298 215 488 249
rect 522 215 571 249
rect 298 199 571 215
rect 613 249 677 265
rect 613 215 623 249
rect 657 215 677 249
rect 847 247 887 282
rect 1087 247 1127 282
rect 1248 265 1288 282
rect 847 217 1127 247
rect 613 199 677 215
rect 79 177 109 199
rect 183 177 213 199
rect 298 177 328 199
rect 541 177 571 199
rect 629 177 659 199
rect 901 177 931 217
rect 1097 177 1127 217
rect 1169 249 1288 265
rect 1169 215 1179 249
rect 1213 215 1288 249
rect 1169 199 1288 215
rect 298 67 328 93
rect 79 21 109 47
rect 183 21 213 47
rect 541 21 571 49
rect 629 21 659 49
rect 1258 133 1288 199
rect 1417 265 1457 314
rect 1417 249 1481 265
rect 1546 255 1586 314
rect 1659 282 1695 297
rect 1753 282 1789 297
rect 1657 265 1697 282
rect 1417 215 1427 249
rect 1461 215 1481 249
rect 1417 199 1481 215
rect 1523 239 1586 255
rect 1523 205 1533 239
rect 1567 205 1586 239
rect 1417 177 1447 199
rect 1523 189 1586 205
rect 1629 249 1697 265
rect 1629 215 1639 249
rect 1673 215 1697 249
rect 1629 199 1697 215
rect 1556 167 1586 189
rect 1667 175 1697 199
rect 1751 265 1791 282
rect 1751 249 1839 265
rect 1751 215 1785 249
rect 1819 215 1839 249
rect 1751 199 1839 215
rect 1751 175 1781 199
rect 901 21 931 47
rect 1097 21 1127 49
rect 1258 23 1288 49
rect 1417 21 1447 49
rect 1556 21 1586 47
rect 1667 21 1697 47
rect 1751 21 1781 47
<< polycont >>
rect 212 215 246 249
rect 488 215 522 249
rect 623 215 657 249
rect 1179 215 1213 249
rect 1427 215 1461 249
rect 1533 205 1567 239
rect 1639 215 1673 249
rect 1785 215 1819 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 17 485 75 527
rect 17 451 35 485
rect 69 451 75 485
rect 17 417 75 451
rect 17 383 35 417
rect 69 383 75 417
rect 17 349 75 383
rect 17 315 35 349
rect 69 315 75 349
rect 17 298 75 315
rect 109 477 173 493
rect 109 443 133 477
rect 167 443 173 477
rect 209 477 286 527
rect 787 481 853 527
rect 1691 489 1758 527
rect 209 443 236 477
rect 270 443 286 477
rect 322 447 568 481
rect 602 447 636 481
rect 787 447 803 481
rect 837 447 853 481
rect 940 455 1500 489
rect 1534 455 1599 489
rect 1691 455 1707 489
rect 1741 455 1758 489
rect 1838 477 1897 493
rect 109 409 173 443
rect 322 409 366 447
rect 940 413 974 455
rect 109 375 133 409
rect 167 375 173 409
rect 109 341 173 375
rect 109 307 133 341
rect 167 307 173 341
rect 17 129 75 147
rect 17 95 35 129
rect 69 95 75 129
rect 17 17 75 95
rect 109 129 173 307
rect 209 375 366 409
rect 434 379 474 413
rect 508 379 974 413
rect 1011 405 1045 421
rect 209 249 253 375
rect 299 307 348 341
rect 382 307 636 341
rect 209 215 212 249
rect 246 215 253 249
rect 209 173 253 215
rect 209 139 343 173
rect 109 95 133 129
rect 167 95 173 129
rect 109 70 173 95
rect 207 89 265 105
rect 207 55 231 89
rect 207 17 265 55
rect 299 85 343 139
rect 377 169 411 307
rect 602 265 636 307
rect 680 305 696 339
rect 730 323 757 339
rect 701 289 723 305
rect 701 275 757 289
rect 445 249 568 265
rect 445 215 488 249
rect 522 215 568 249
rect 602 249 667 265
rect 602 215 623 249
rect 657 215 667 249
rect 602 199 667 215
rect 377 119 411 135
rect 471 165 547 181
rect 471 131 487 165
rect 521 159 547 165
rect 701 159 735 275
rect 791 241 825 379
rect 871 309 897 343
rect 931 309 975 343
rect 871 289 975 309
rect 521 131 735 159
rect 471 125 735 131
rect 769 207 825 241
rect 769 91 803 207
rect 917 187 975 289
rect 536 85 583 91
rect 299 57 583 85
rect 617 57 633 91
rect 677 57 693 91
rect 727 57 803 91
rect 837 157 871 173
rect 837 89 871 123
rect 299 51 633 57
rect 951 165 975 187
rect 917 131 941 153
rect 917 83 975 131
rect 1011 119 1045 371
rect 1079 178 1113 455
rect 1872 443 1897 477
rect 1838 421 1897 443
rect 1359 409 1897 421
rect 1159 375 1177 409
rect 1211 375 1242 409
rect 1159 341 1242 375
rect 1159 307 1177 341
rect 1211 323 1242 341
rect 1359 390 1839 409
rect 1393 387 1839 390
rect 1790 375 1839 387
rect 1873 375 1897 409
rect 1211 307 1213 323
rect 1159 289 1213 307
rect 1247 289 1325 323
rect 1162 249 1247 254
rect 1162 215 1179 249
rect 1213 215 1247 249
rect 1162 199 1247 215
rect 1205 187 1247 199
rect 1079 165 1131 178
rect 1079 144 1171 165
rect 1087 131 1171 144
rect 1137 126 1171 131
rect 1205 153 1213 187
rect 1205 126 1247 153
rect 1011 85 1019 119
rect 837 17 871 55
rect 1011 63 1043 85
rect 1077 63 1093 97
rect 1137 64 1171 92
rect 1291 85 1325 289
rect 1359 169 1393 356
rect 1427 289 1553 323
rect 1597 307 1613 341
rect 1647 307 1807 341
rect 1597 299 1807 307
rect 1427 249 1471 289
rect 1773 265 1807 299
rect 1461 215 1471 249
rect 1427 199 1471 215
rect 1505 239 1567 255
rect 1505 205 1533 239
rect 1611 249 1739 265
rect 1611 215 1639 249
rect 1673 215 1739 249
rect 1773 249 1829 265
rect 1773 215 1785 249
rect 1819 215 1829 249
rect 1505 189 1567 205
rect 1773 199 1829 215
rect 1505 187 1546 189
rect 1505 153 1509 187
rect 1543 153 1546 187
rect 1773 181 1807 199
rect 1505 146 1546 153
rect 1613 150 1807 181
rect 1605 147 1807 150
rect 1359 119 1393 135
rect 1605 142 1663 147
rect 1605 119 1613 142
rect 1427 85 1469 93
rect 1011 53 1093 63
rect 1291 59 1469 85
rect 1503 59 1530 93
rect 1605 85 1611 119
rect 1647 108 1663 142
rect 1863 117 1897 375
rect 1645 85 1663 108
rect 1605 59 1663 85
rect 1707 97 1741 113
rect 1291 51 1530 59
rect 1707 17 1741 63
rect 1837 101 1897 117
rect 1871 67 1897 101
rect 1837 51 1897 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 723 305 730 323
rect 730 305 757 323
rect 723 289 757 305
rect 917 165 951 187
rect 917 153 941 165
rect 941 153 951 165
rect 1213 289 1247 323
rect 1213 153 1247 187
rect 1019 97 1053 119
rect 1019 85 1043 97
rect 1043 85 1053 97
rect 1509 153 1543 187
rect 1611 108 1613 119
rect 1613 108 1645 119
rect 1611 85 1645 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 711 323 769 329
rect 711 289 723 323
rect 757 320 769 323
rect 1201 323 1259 329
rect 1201 320 1213 323
rect 757 292 1213 320
rect 757 289 769 292
rect 711 283 769 289
rect 1201 289 1213 292
rect 1247 289 1259 323
rect 1201 283 1259 289
rect 905 187 963 193
rect 905 153 917 187
rect 951 184 963 187
rect 1201 187 1259 193
rect 1201 184 1213 187
rect 951 156 1213 184
rect 951 153 963 156
rect 905 147 963 153
rect 1201 153 1213 156
rect 1247 184 1259 187
rect 1497 187 1555 193
rect 1497 184 1509 187
rect 1247 156 1509 184
rect 1247 153 1259 156
rect 1201 147 1259 153
rect 1497 153 1509 156
rect 1543 153 1555 187
rect 1497 147 1555 153
rect 1007 119 1065 125
rect 1007 85 1019 119
rect 1053 116 1065 119
rect 1599 119 1657 125
rect 1599 116 1611 119
rect 1053 88 1611 116
rect 1053 85 1065 88
rect 1007 79 1065 85
rect 1599 85 1611 88
rect 1645 85 1657 119
rect 1599 79 1657 85
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 131 357 165 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1500 289 1534 323 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 488 221 522 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1686 221 1720 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xnor3_2
flabel comment s 0 544 0 544 3 FreeSans 200 0 0 0 HHNEC
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1263666
string GDS_START 1250874
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
