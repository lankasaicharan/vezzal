magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 1 49 964 157
rect 0 0 1056 49
<< scnmos >>
rect 80 47 110 131
rect 166 47 196 131
rect 252 47 282 131
rect 338 47 368 131
rect 424 47 454 131
rect 510 47 540 131
rect 596 47 626 131
rect 682 47 712 131
rect 768 47 798 131
rect 854 47 884 131
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 252 367 282 619
rect 338 367 368 619
rect 424 367 454 619
rect 510 367 540 619
rect 596 367 626 619
rect 682 367 712 619
rect 768 367 798 619
rect 854 367 884 619
<< ndiff >>
rect 27 106 80 131
rect 27 72 35 106
rect 69 72 80 106
rect 27 47 80 72
rect 110 106 166 131
rect 110 72 121 106
rect 155 72 166 106
rect 110 47 166 72
rect 196 106 252 131
rect 196 72 207 106
rect 241 72 252 106
rect 196 47 252 72
rect 282 106 338 131
rect 282 72 293 106
rect 327 72 338 106
rect 282 47 338 72
rect 368 97 424 131
rect 368 63 379 97
rect 413 63 424 97
rect 368 47 424 63
rect 454 106 510 131
rect 454 72 465 106
rect 499 72 510 106
rect 454 47 510 72
rect 540 97 596 131
rect 540 63 551 97
rect 585 63 596 97
rect 540 47 596 63
rect 626 106 682 131
rect 626 72 637 106
rect 671 72 682 106
rect 626 47 682 72
rect 712 97 768 131
rect 712 63 723 97
rect 757 63 768 97
rect 712 47 768 63
rect 798 106 854 131
rect 798 72 809 106
rect 843 72 854 106
rect 798 47 854 72
rect 884 97 938 131
rect 884 63 896 97
rect 930 63 938 97
rect 884 47 938 63
<< pdiff >>
rect 27 595 80 619
rect 27 561 35 595
rect 69 561 80 595
rect 27 511 80 561
rect 27 477 35 511
rect 69 477 80 511
rect 27 425 80 477
rect 27 391 35 425
rect 69 391 80 425
rect 27 367 80 391
rect 110 595 166 619
rect 110 561 121 595
rect 155 561 166 595
rect 110 511 166 561
rect 110 477 121 511
rect 155 477 166 511
rect 110 425 166 477
rect 110 391 121 425
rect 155 391 166 425
rect 110 367 166 391
rect 196 595 252 619
rect 196 561 207 595
rect 241 561 252 595
rect 196 511 252 561
rect 196 477 207 511
rect 241 477 252 511
rect 196 425 252 477
rect 196 391 207 425
rect 241 391 252 425
rect 196 367 252 391
rect 282 595 338 619
rect 282 561 293 595
rect 327 561 338 595
rect 282 511 338 561
rect 282 477 293 511
rect 327 477 338 511
rect 282 425 338 477
rect 282 391 293 425
rect 327 391 338 425
rect 282 367 338 391
rect 368 599 424 619
rect 368 565 379 599
rect 413 565 424 599
rect 368 531 424 565
rect 368 497 379 531
rect 413 497 424 531
rect 368 463 424 497
rect 368 429 379 463
rect 413 429 424 463
rect 368 367 424 429
rect 454 595 510 619
rect 454 561 465 595
rect 499 561 510 595
rect 454 511 510 561
rect 454 477 465 511
rect 499 477 510 511
rect 454 425 510 477
rect 454 391 465 425
rect 499 391 510 425
rect 454 367 510 391
rect 540 599 596 619
rect 540 565 551 599
rect 585 565 596 599
rect 540 531 596 565
rect 540 497 551 531
rect 585 497 596 531
rect 540 463 596 497
rect 540 429 551 463
rect 585 429 596 463
rect 540 367 596 429
rect 626 595 682 619
rect 626 561 637 595
rect 671 561 682 595
rect 626 511 682 561
rect 626 477 637 511
rect 671 477 682 511
rect 626 425 682 477
rect 626 391 637 425
rect 671 391 682 425
rect 626 367 682 391
rect 712 599 768 619
rect 712 565 723 599
rect 757 565 768 599
rect 712 531 768 565
rect 712 497 723 531
rect 757 497 768 531
rect 712 463 768 497
rect 712 429 723 463
rect 757 429 768 463
rect 712 367 768 429
rect 798 595 854 619
rect 798 561 809 595
rect 843 561 854 595
rect 798 511 854 561
rect 798 477 809 511
rect 843 477 854 511
rect 798 425 854 477
rect 798 391 809 425
rect 843 391 854 425
rect 798 367 854 391
rect 884 599 937 619
rect 884 565 895 599
rect 929 565 937 599
rect 884 531 937 565
rect 884 497 895 531
rect 929 497 937 531
rect 884 463 937 497
rect 884 429 895 463
rect 929 429 937 463
rect 884 367 937 429
<< ndiffc >>
rect 35 72 69 106
rect 121 72 155 106
rect 207 72 241 106
rect 293 72 327 106
rect 379 63 413 97
rect 465 72 499 106
rect 551 63 585 97
rect 637 72 671 106
rect 723 63 757 97
rect 809 72 843 106
rect 896 63 930 97
<< pdiffc >>
rect 35 561 69 595
rect 35 477 69 511
rect 35 391 69 425
rect 121 561 155 595
rect 121 477 155 511
rect 121 391 155 425
rect 207 561 241 595
rect 207 477 241 511
rect 207 391 241 425
rect 293 561 327 595
rect 293 477 327 511
rect 293 391 327 425
rect 379 565 413 599
rect 379 497 413 531
rect 379 429 413 463
rect 465 561 499 595
rect 465 477 499 511
rect 465 391 499 425
rect 551 565 585 599
rect 551 497 585 531
rect 551 429 585 463
rect 637 561 671 595
rect 637 477 671 511
rect 637 391 671 425
rect 723 565 757 599
rect 723 497 757 531
rect 723 429 757 463
rect 809 561 843 595
rect 809 477 843 511
rect 809 391 843 425
rect 895 565 929 599
rect 895 497 929 531
rect 895 429 929 463
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 252 619 282 645
rect 338 619 368 645
rect 424 619 454 645
rect 510 619 540 645
rect 596 619 626 645
rect 682 619 712 645
rect 768 619 798 645
rect 854 619 884 645
rect 80 314 110 367
rect 166 314 196 367
rect 21 298 196 314
rect 21 264 37 298
rect 71 264 196 298
rect 21 230 196 264
rect 21 196 37 230
rect 71 196 196 230
rect 21 180 196 196
rect 80 131 110 180
rect 166 131 196 180
rect 252 297 282 367
rect 338 297 368 367
rect 424 297 454 367
rect 510 297 540 367
rect 596 297 626 367
rect 682 297 712 367
rect 768 297 798 367
rect 854 297 884 367
rect 252 281 884 297
rect 252 247 292 281
rect 326 247 360 281
rect 394 247 428 281
rect 462 247 496 281
rect 530 247 564 281
rect 598 247 632 281
rect 666 247 884 281
rect 252 231 884 247
rect 252 131 282 231
rect 338 131 368 231
rect 424 131 454 231
rect 510 131 540 231
rect 596 131 626 231
rect 682 131 712 231
rect 768 131 798 231
rect 854 131 884 231
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 424 21 454 47
rect 510 21 540 47
rect 596 21 626 47
rect 682 21 712 47
rect 768 21 798 47
rect 854 21 884 47
<< polycont >>
rect 37 264 71 298
rect 37 196 71 230
rect 292 247 326 281
rect 360 247 394 281
rect 428 247 462 281
rect 496 247 530 281
rect 564 247 598 281
rect 632 247 666 281
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 19 595 78 611
rect 19 579 35 595
rect 19 545 33 579
rect 69 561 78 595
rect 67 545 78 561
rect 19 511 78 545
rect 19 477 35 511
rect 69 477 78 511
rect 19 425 78 477
rect 19 391 35 425
rect 69 391 78 425
rect 19 375 78 391
rect 114 595 164 615
rect 114 561 121 595
rect 155 561 164 595
rect 114 511 164 561
rect 114 477 121 511
rect 155 477 164 511
rect 114 425 164 477
rect 114 391 121 425
rect 155 391 164 425
rect 17 298 80 314
rect 17 264 37 298
rect 71 264 80 298
rect 17 230 80 264
rect 17 196 37 230
rect 71 196 80 230
rect 17 156 80 196
rect 114 297 164 391
rect 198 595 250 611
rect 198 561 207 595
rect 241 579 250 595
rect 198 545 208 561
rect 242 545 250 579
rect 198 511 250 545
rect 198 477 207 511
rect 241 477 250 511
rect 198 425 250 477
rect 198 391 207 425
rect 241 391 250 425
rect 198 375 250 391
rect 284 595 336 615
rect 284 561 293 595
rect 327 561 336 595
rect 284 511 336 561
rect 284 477 293 511
rect 327 477 336 511
rect 284 425 336 477
rect 284 391 293 425
rect 327 391 336 425
rect 370 599 422 615
rect 370 579 379 599
rect 370 545 378 579
rect 413 565 422 599
rect 412 545 422 565
rect 370 531 422 545
rect 370 497 379 531
rect 413 497 422 531
rect 370 463 422 497
rect 370 429 379 463
rect 413 429 422 463
rect 370 413 422 429
rect 456 595 508 615
rect 456 561 465 595
rect 499 561 508 595
rect 456 511 508 561
rect 456 477 465 511
rect 499 477 508 511
rect 456 425 508 477
rect 284 379 336 391
rect 456 391 465 425
rect 499 391 508 425
rect 542 599 594 615
rect 542 579 551 599
rect 542 545 550 579
rect 585 565 594 599
rect 584 545 594 565
rect 542 531 594 545
rect 542 497 551 531
rect 585 497 594 531
rect 542 463 594 497
rect 542 429 551 463
rect 585 429 594 463
rect 542 413 594 429
rect 628 595 680 615
rect 628 561 637 595
rect 671 561 680 595
rect 628 511 680 561
rect 628 477 637 511
rect 671 477 680 511
rect 628 425 680 477
rect 456 379 508 391
rect 628 391 637 425
rect 671 391 680 425
rect 714 599 766 615
rect 714 579 723 599
rect 714 545 721 579
rect 757 565 766 599
rect 755 545 766 565
rect 714 531 766 545
rect 714 497 723 531
rect 757 497 766 531
rect 714 463 766 497
rect 714 429 723 463
rect 757 429 766 463
rect 714 413 766 429
rect 800 595 852 615
rect 800 561 809 595
rect 843 561 852 595
rect 800 511 852 561
rect 800 477 809 511
rect 843 477 852 511
rect 800 425 852 477
rect 628 379 680 391
rect 800 391 809 425
rect 843 391 852 425
rect 886 599 945 615
rect 886 565 895 599
rect 929 579 945 599
rect 886 545 898 565
rect 932 545 945 579
rect 886 531 945 545
rect 886 497 895 531
rect 929 497 945 531
rect 886 463 945 497
rect 886 429 895 463
rect 929 429 945 463
rect 886 413 945 429
rect 800 379 852 391
rect 284 331 946 379
rect 114 281 718 297
rect 114 247 292 281
rect 326 247 360 281
rect 394 247 428 281
rect 462 247 496 281
rect 530 247 564 281
rect 598 247 632 281
rect 666 247 718 281
rect 114 231 718 247
rect 29 106 78 122
rect 29 72 35 106
rect 69 72 78 106
rect 29 17 78 72
rect 114 106 164 231
rect 752 195 946 331
rect 284 147 946 195
rect 114 72 121 106
rect 155 72 164 106
rect 114 53 164 72
rect 198 106 250 122
rect 198 72 207 106
rect 241 72 250 106
rect 198 17 250 72
rect 284 106 336 147
rect 284 72 293 106
rect 327 72 336 106
rect 284 56 336 72
rect 370 97 422 113
rect 370 63 379 97
rect 413 63 422 97
rect 370 17 422 63
rect 456 106 508 147
rect 456 72 465 106
rect 499 72 508 106
rect 456 56 508 72
rect 542 97 594 113
rect 542 63 551 97
rect 585 63 594 97
rect 542 17 594 63
rect 628 106 680 147
rect 628 72 637 106
rect 671 72 680 106
rect 628 56 680 72
rect 714 97 766 113
rect 714 63 723 97
rect 757 63 766 97
rect 714 17 766 63
rect 800 106 852 147
rect 800 72 809 106
rect 843 72 852 106
rect 800 56 852 72
rect 886 97 946 113
rect 886 63 896 97
rect 930 63 946 97
rect 886 17 946 63
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 33 561 35 579
rect 35 561 67 579
rect 33 545 67 561
rect 208 561 241 579
rect 241 561 242 579
rect 208 545 242 561
rect 378 565 379 579
rect 379 565 412 579
rect 378 545 412 565
rect 550 565 551 579
rect 551 565 584 579
rect 550 545 584 565
rect 721 565 723 579
rect 723 565 755 579
rect 721 545 755 565
rect 898 565 929 579
rect 929 565 932 579
rect 898 545 932 565
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 14 579 1042 589
rect 14 545 33 579
rect 67 545 208 579
rect 242 545 378 579
rect 412 545 550 579
rect 584 545 721 579
rect 755 545 898 579
rect 932 545 1042 579
rect 14 538 1042 545
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 bufkapwr_8
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 14 538 1042 589 0 FreeSans 200 0 0 0 KAPWR
port 2 nsew power bidirectional
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y
string GDS_END 2549290
string GDS_START 2539800
<< end >>
