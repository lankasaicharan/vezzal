magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 25 49 767 167
rect 0 0 768 49
<< scnmos >>
rect 108 57 138 141
rect 180 57 210 141
rect 266 57 296 141
rect 338 57 368 141
rect 424 57 454 141
rect 496 57 526 141
rect 582 57 612 141
rect 654 57 684 141
<< scpmoshvt >>
rect 164 409 214 609
rect 393 409 443 609
rect 491 409 541 609
rect 605 409 655 609
<< ndiff >>
rect 51 116 108 141
rect 51 82 63 116
rect 97 82 108 116
rect 51 57 108 82
rect 138 57 180 141
rect 210 112 266 141
rect 210 78 221 112
rect 255 78 266 112
rect 210 57 266 78
rect 296 57 338 141
rect 368 116 424 141
rect 368 82 379 116
rect 413 82 424 116
rect 368 57 424 82
rect 454 57 496 141
rect 526 112 582 141
rect 526 78 537 112
rect 571 78 582 112
rect 526 57 582 78
rect 612 57 654 141
rect 684 116 741 141
rect 684 82 695 116
rect 729 82 741 116
rect 684 57 741 82
<< pdiff >>
rect 107 597 164 609
rect 107 563 119 597
rect 153 563 164 597
rect 107 526 164 563
rect 107 492 119 526
rect 153 492 164 526
rect 107 455 164 492
rect 107 421 119 455
rect 153 421 164 455
rect 107 409 164 421
rect 214 597 393 609
rect 214 563 225 597
rect 259 563 393 597
rect 214 526 393 563
rect 214 492 225 526
rect 259 492 393 526
rect 214 455 393 492
rect 214 421 225 455
rect 259 421 393 455
rect 214 409 393 421
rect 443 409 491 609
rect 541 409 605 609
rect 655 597 712 609
rect 655 563 666 597
rect 700 563 712 597
rect 655 463 712 563
rect 655 429 666 463
rect 700 429 712 463
rect 655 409 712 429
<< ndiffc >>
rect 63 82 97 116
rect 221 78 255 112
rect 379 82 413 116
rect 537 78 571 112
rect 695 82 729 116
<< pdiffc >>
rect 119 563 153 597
rect 119 492 153 526
rect 119 421 153 455
rect 225 563 259 597
rect 225 492 259 526
rect 225 421 259 455
rect 666 563 700 597
rect 666 429 700 463
<< poly >>
rect 164 609 214 635
rect 393 609 443 635
rect 491 609 541 635
rect 605 609 655 635
rect 164 368 214 409
rect 393 377 443 409
rect 491 377 541 409
rect 605 377 655 409
rect 180 352 271 368
rect 180 318 221 352
rect 255 318 271 352
rect 180 284 271 318
rect 180 264 221 284
rect 108 250 221 264
rect 255 250 271 284
rect 108 234 271 250
rect 338 361 423 377
rect 338 327 354 361
rect 388 327 423 361
rect 338 293 423 327
rect 338 259 354 293
rect 388 259 423 293
rect 338 243 423 259
rect 491 361 557 377
rect 491 327 507 361
rect 541 327 557 361
rect 491 293 557 327
rect 491 259 507 293
rect 541 259 557 293
rect 491 243 557 259
rect 605 361 671 377
rect 605 327 621 361
rect 655 327 671 361
rect 605 293 671 327
rect 605 259 621 293
rect 655 259 671 293
rect 605 243 671 259
rect 108 141 138 234
rect 180 141 210 234
rect 338 186 368 243
rect 491 186 521 243
rect 605 186 635 243
rect 266 156 368 186
rect 266 141 296 156
rect 338 141 368 156
rect 424 156 526 186
rect 424 141 454 156
rect 496 141 526 156
rect 582 156 684 186
rect 582 141 612 156
rect 654 141 684 156
rect 108 31 138 57
rect 180 31 210 57
rect 266 31 296 57
rect 338 31 368 57
rect 424 31 454 57
rect 496 31 526 57
rect 582 31 612 57
rect 654 31 684 57
<< polycont >>
rect 221 318 255 352
rect 221 250 255 284
rect 354 327 388 361
rect 354 259 388 293
rect 507 327 541 361
rect 507 259 541 293
rect 621 327 655 361
rect 621 259 655 293
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 25 597 169 613
rect 25 563 119 597
rect 153 563 169 597
rect 25 526 169 563
rect 25 492 119 526
rect 153 492 169 526
rect 25 455 169 492
rect 25 421 119 455
rect 153 421 169 455
rect 25 116 169 421
rect 209 597 275 649
rect 209 563 225 597
rect 259 563 275 597
rect 650 597 745 613
rect 209 526 275 563
rect 209 492 225 526
rect 259 492 275 526
rect 209 455 275 492
rect 209 421 225 455
rect 259 421 275 455
rect 209 405 275 421
rect 205 352 271 368
rect 205 318 221 352
rect 255 318 271 352
rect 205 284 271 318
rect 205 250 221 284
rect 255 250 271 284
rect 205 207 271 250
rect 313 361 455 578
rect 313 327 354 361
rect 388 327 455 361
rect 313 293 455 327
rect 313 259 354 293
rect 388 259 455 293
rect 313 243 455 259
rect 491 361 557 578
rect 650 563 666 597
rect 700 563 745 597
rect 650 463 745 563
rect 650 429 666 463
rect 700 429 745 463
rect 650 413 745 429
rect 491 327 507 361
rect 541 327 557 361
rect 491 293 557 327
rect 491 259 507 293
rect 541 259 557 293
rect 491 243 557 259
rect 601 361 671 377
rect 601 327 621 361
rect 655 327 671 361
rect 601 293 671 327
rect 601 259 621 293
rect 655 259 671 293
rect 601 243 671 259
rect 711 207 745 413
rect 205 173 745 207
rect 25 82 63 116
rect 97 88 169 116
rect 205 112 271 137
rect 97 82 113 88
rect 25 53 113 82
rect 205 78 221 112
rect 255 78 271 112
rect 205 17 271 78
rect 363 116 429 173
rect 363 82 379 116
rect 413 82 429 116
rect 363 53 429 82
rect 521 112 587 137
rect 521 78 537 112
rect 571 78 587 112
rect 521 17 587 78
rect 679 116 745 173
rect 679 82 695 116
rect 729 82 745 116
rect 679 53 745 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or3_lp
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3175784
string GDS_START 3167202
<< end >>
