magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4946 1975
<< nwell >>
rect -38 331 3686 704
rect 512 271 718 331
<< pwell >>
rect 1749 273 1851 281
rect 1749 247 2768 273
rect 1163 241 3261 247
rect 11 205 677 229
rect 11 177 923 205
rect 1163 177 3647 241
rect 11 49 3647 177
rect 0 0 3648 49
<< scnmos >>
rect 94 119 124 203
rect 172 119 202 203
rect 293 119 323 203
rect 407 119 437 203
rect 564 119 594 203
rect 810 95 840 179
rect 1047 67 1077 151
rect 1243 137 1273 221
rect 1329 137 1359 221
rect 1452 137 1482 221
rect 1640 93 1670 221
rect 1730 93 1760 221
rect 1840 93 1870 221
rect 2086 119 2116 247
rect 2188 119 2218 247
rect 2337 163 2367 247
rect 2415 163 2445 247
rect 2544 119 2574 247
rect 2662 119 2692 247
rect 2757 71 2787 199
rect 2955 137 2985 221
rect 3057 53 3087 221
rect 3143 53 3173 221
rect 3346 47 3376 131
rect 3448 47 3478 215
rect 3534 47 3564 215
<< scpmoshvt >>
rect 113 481 143 609
rect 215 481 245 609
rect 293 481 323 609
rect 407 481 437 609
rect 598 307 628 435
rect 810 411 840 539
rect 1047 469 1077 597
rect 1243 463 1273 547
rect 1345 463 1375 547
rect 1423 463 1453 547
rect 1652 379 1682 547
rect 1766 379 1796 547
rect 1844 379 1874 547
rect 2086 379 2116 547
rect 2181 428 2211 596
rect 2283 506 2313 590
rect 2452 506 2482 590
rect 2598 451 2628 619
rect 2684 451 2714 619
rect 2762 451 2792 619
rect 2954 367 2984 495
rect 3056 367 3086 619
rect 3142 367 3172 619
rect 3346 396 3376 524
rect 3448 367 3478 619
rect 3534 367 3564 619
<< ndiff >>
rect 37 178 94 203
rect 37 144 49 178
rect 83 144 94 178
rect 37 119 94 144
rect 124 119 172 203
rect 202 178 293 203
rect 202 144 213 178
rect 247 144 293 178
rect 202 119 293 144
rect 323 119 407 203
rect 437 175 564 203
rect 437 141 481 175
rect 515 141 564 175
rect 437 119 564 141
rect 594 178 651 203
rect 1775 243 1825 255
rect 1775 221 1783 243
rect 594 144 605 178
rect 639 144 651 178
rect 594 119 651 144
rect 737 154 810 179
rect 737 120 749 154
rect 783 120 810 154
rect 737 95 810 120
rect 840 154 897 179
rect 840 120 851 154
rect 885 120 897 154
rect 1189 196 1243 221
rect 1189 162 1198 196
rect 1232 162 1243 196
rect 840 95 897 120
rect 978 126 1047 151
rect 978 92 990 126
rect 1024 92 1047 126
rect 978 67 1047 92
rect 1077 126 1135 151
rect 1189 137 1243 162
rect 1273 196 1329 221
rect 1273 162 1284 196
rect 1318 162 1329 196
rect 1273 137 1329 162
rect 1359 137 1452 221
rect 1482 137 1640 221
rect 1077 92 1092 126
rect 1126 92 1135 126
rect 1077 67 1135 92
rect 1497 114 1640 137
rect 1497 80 1509 114
rect 1543 93 1640 114
rect 1670 178 1730 221
rect 1670 144 1681 178
rect 1715 144 1730 178
rect 1670 93 1730 144
rect 1760 209 1783 221
rect 1817 221 1825 243
rect 1817 209 1840 221
rect 1760 93 1840 209
rect 1870 174 1931 221
rect 1870 140 1885 174
rect 1919 140 1931 174
rect 1870 93 1931 140
rect 2029 166 2086 247
rect 2029 132 2041 166
rect 2075 132 2086 166
rect 2029 119 2086 132
rect 2116 119 2188 247
rect 2218 235 2337 247
rect 2218 201 2276 235
rect 2310 201 2337 235
rect 2218 165 2337 201
rect 2218 131 2276 165
rect 2310 163 2337 165
rect 2367 163 2415 247
rect 2445 163 2544 247
rect 2310 131 2322 163
rect 2218 119 2322 131
rect 2471 119 2544 163
rect 2574 119 2662 247
rect 2692 199 2742 247
rect 2692 180 2757 199
rect 2692 146 2712 180
rect 2746 146 2757 180
rect 2692 119 2757 146
rect 2471 114 2529 119
rect 1543 80 1555 93
rect 1497 68 1555 80
rect 2471 80 2483 114
rect 2517 80 2529 114
rect 2589 114 2647 119
rect 2471 68 2529 80
rect 2589 80 2601 114
rect 2635 80 2647 114
rect 2589 68 2647 80
rect 2707 71 2757 119
rect 2787 132 2844 199
rect 2898 196 2955 221
rect 2898 162 2910 196
rect 2944 162 2955 196
rect 2898 137 2955 162
rect 2985 209 3057 221
rect 2985 175 3012 209
rect 3046 175 3057 209
rect 2985 137 3057 175
rect 2787 98 2798 132
rect 2832 98 2844 132
rect 2787 71 2844 98
rect 3000 99 3057 137
rect 3000 65 3012 99
rect 3046 65 3057 99
rect 3000 53 3057 65
rect 3087 209 3143 221
rect 3087 175 3098 209
rect 3132 175 3143 209
rect 3087 103 3143 175
rect 3087 69 3098 103
rect 3132 69 3143 103
rect 3087 53 3143 69
rect 3173 209 3235 221
rect 3173 175 3189 209
rect 3223 175 3235 209
rect 3173 99 3235 175
rect 3391 185 3448 215
rect 3391 151 3403 185
rect 3437 151 3448 185
rect 3391 131 3448 151
rect 3173 65 3189 99
rect 3223 65 3235 99
rect 3173 53 3235 65
rect 3289 106 3346 131
rect 3289 72 3301 106
rect 3335 72 3346 106
rect 3289 47 3346 72
rect 3376 93 3448 131
rect 3376 59 3403 93
rect 3437 59 3448 93
rect 3376 47 3448 59
rect 3478 203 3534 215
rect 3478 169 3489 203
rect 3523 169 3534 203
rect 3478 103 3534 169
rect 3478 69 3489 103
rect 3523 69 3534 103
rect 3478 47 3534 69
rect 3564 203 3621 215
rect 3564 169 3575 203
rect 3609 169 3621 203
rect 3564 93 3621 169
rect 3564 59 3575 93
rect 3609 59 3621 93
rect 3564 47 3621 59
<< pdiff >>
rect 56 597 113 609
rect 56 563 68 597
rect 102 563 113 597
rect 56 527 113 563
rect 56 493 68 527
rect 102 493 113 527
rect 56 481 113 493
rect 143 565 215 609
rect 143 531 170 565
rect 204 531 215 565
rect 143 481 215 531
rect 245 481 293 609
rect 323 535 407 609
rect 323 501 346 535
rect 380 501 407 535
rect 323 481 407 501
rect 437 597 494 609
rect 437 563 448 597
rect 482 563 494 597
rect 437 527 494 563
rect 437 493 448 527
rect 482 493 494 527
rect 437 481 494 493
rect 548 535 606 547
rect 548 501 560 535
rect 594 501 606 535
rect 548 489 606 501
rect 736 527 810 539
rect 736 493 745 527
rect 779 493 810 527
rect 548 435 578 489
rect 548 307 598 435
rect 628 354 682 435
rect 736 411 810 493
rect 840 527 927 539
rect 840 493 885 527
rect 919 493 927 527
rect 840 457 927 493
rect 840 423 885 457
rect 919 423 927 457
rect 840 411 927 423
rect 981 469 1047 597
rect 1077 585 1131 597
rect 1077 551 1088 585
rect 1122 551 1131 585
rect 1077 469 1131 551
rect 2131 547 2181 596
rect 1189 522 1243 547
rect 1189 488 1198 522
rect 1232 488 1243 522
rect 981 413 1032 469
rect 981 379 990 413
rect 1024 379 1032 413
rect 981 367 1032 379
rect 628 320 639 354
rect 673 320 682 354
rect 628 307 682 320
rect 1189 463 1243 488
rect 1273 522 1345 547
rect 1273 488 1300 522
rect 1334 488 1345 522
rect 1273 463 1345 488
rect 1375 463 1423 547
rect 1453 535 1652 547
rect 1453 501 1607 535
rect 1641 501 1652 535
rect 1453 463 1652 501
rect 1595 379 1652 463
rect 1682 535 1766 547
rect 1682 501 1721 535
rect 1755 501 1766 535
rect 1682 465 1766 501
rect 1682 431 1721 465
rect 1755 431 1766 465
rect 1682 379 1766 431
rect 1796 379 1844 547
rect 1874 535 2086 547
rect 1874 501 1918 535
rect 1952 501 2086 535
rect 1874 425 2086 501
rect 1874 391 1918 425
rect 1952 391 2086 425
rect 1874 379 2086 391
rect 2116 428 2181 547
rect 2211 590 2268 596
rect 2544 590 2598 619
rect 2211 506 2283 590
rect 2313 506 2452 590
rect 2482 575 2598 590
rect 2482 541 2553 575
rect 2587 541 2598 575
rect 2482 506 2598 541
rect 2211 500 2268 506
rect 2211 466 2222 500
rect 2256 466 2268 500
rect 2211 428 2268 466
rect 2116 379 2166 428
rect 2544 451 2598 506
rect 2628 597 2684 619
rect 2628 563 2639 597
rect 2673 563 2684 597
rect 2628 497 2684 563
rect 2628 463 2639 497
rect 2673 463 2684 497
rect 2628 451 2684 463
rect 2714 451 2762 619
rect 2792 602 2846 619
rect 2792 568 2803 602
rect 2837 568 2846 602
rect 2792 451 2846 568
rect 2999 602 3056 619
rect 2999 568 3011 602
rect 3045 568 3056 602
rect 2999 495 3056 568
rect 2900 442 2954 495
rect 2900 408 2909 442
rect 2943 408 2954 442
rect 2900 367 2954 408
rect 2984 367 3056 495
rect 3086 597 3142 619
rect 3086 563 3097 597
rect 3131 563 3142 597
rect 3086 505 3142 563
rect 3086 471 3097 505
rect 3131 471 3142 505
rect 3086 413 3142 471
rect 3086 379 3097 413
rect 3131 379 3142 413
rect 3086 367 3142 379
rect 3172 607 3232 619
rect 3172 573 3189 607
rect 3223 573 3232 607
rect 3172 510 3232 573
rect 3391 607 3448 619
rect 3391 573 3403 607
rect 3437 573 3448 607
rect 3391 524 3448 573
rect 3172 476 3189 510
rect 3223 476 3232 510
rect 3172 413 3232 476
rect 3172 379 3189 413
rect 3223 379 3232 413
rect 3292 512 3346 524
rect 3292 478 3301 512
rect 3335 478 3346 512
rect 3292 442 3346 478
rect 3292 408 3301 442
rect 3335 408 3346 442
rect 3292 396 3346 408
rect 3376 510 3448 524
rect 3376 476 3403 510
rect 3437 476 3448 510
rect 3376 413 3448 476
rect 3376 396 3403 413
rect 3172 367 3232 379
rect 3391 379 3403 396
rect 3437 379 3448 413
rect 3391 367 3448 379
rect 3478 597 3534 619
rect 3478 563 3489 597
rect 3523 563 3534 597
rect 3478 505 3534 563
rect 3478 471 3489 505
rect 3523 471 3534 505
rect 3478 413 3534 471
rect 3478 379 3489 413
rect 3523 379 3534 413
rect 3478 367 3534 379
rect 3564 607 3621 619
rect 3564 573 3575 607
rect 3609 573 3621 607
rect 3564 510 3621 573
rect 3564 476 3575 510
rect 3609 476 3621 510
rect 3564 413 3621 476
rect 3564 379 3575 413
rect 3609 379 3621 413
rect 3564 367 3621 379
<< ndiffc >>
rect 49 144 83 178
rect 213 144 247 178
rect 481 141 515 175
rect 605 144 639 178
rect 749 120 783 154
rect 851 120 885 154
rect 1198 162 1232 196
rect 990 92 1024 126
rect 1284 162 1318 196
rect 1092 92 1126 126
rect 1509 80 1543 114
rect 1681 144 1715 178
rect 1783 209 1817 243
rect 1885 140 1919 174
rect 2041 132 2075 166
rect 2276 201 2310 235
rect 2276 131 2310 165
rect 2712 146 2746 180
rect 2483 80 2517 114
rect 2601 80 2635 114
rect 2910 162 2944 196
rect 3012 175 3046 209
rect 2798 98 2832 132
rect 3012 65 3046 99
rect 3098 175 3132 209
rect 3098 69 3132 103
rect 3189 175 3223 209
rect 3403 151 3437 185
rect 3189 65 3223 99
rect 3301 72 3335 106
rect 3403 59 3437 93
rect 3489 169 3523 203
rect 3489 69 3523 103
rect 3575 169 3609 203
rect 3575 59 3609 93
<< pdiffc >>
rect 68 563 102 597
rect 68 493 102 527
rect 170 531 204 565
rect 346 501 380 535
rect 448 563 482 597
rect 448 493 482 527
rect 560 501 594 535
rect 745 493 779 527
rect 885 493 919 527
rect 885 423 919 457
rect 1088 551 1122 585
rect 1198 488 1232 522
rect 990 379 1024 413
rect 639 320 673 354
rect 1300 488 1334 522
rect 1607 501 1641 535
rect 1721 501 1755 535
rect 1721 431 1755 465
rect 1918 501 1952 535
rect 1918 391 1952 425
rect 2553 541 2587 575
rect 2222 466 2256 500
rect 2639 563 2673 597
rect 2639 463 2673 497
rect 2803 568 2837 602
rect 3011 568 3045 602
rect 2909 408 2943 442
rect 3097 563 3131 597
rect 3097 471 3131 505
rect 3097 379 3131 413
rect 3189 573 3223 607
rect 3403 573 3437 607
rect 3189 476 3223 510
rect 3189 379 3223 413
rect 3301 478 3335 512
rect 3301 408 3335 442
rect 3403 476 3437 510
rect 3403 379 3437 413
rect 3489 563 3523 597
rect 3489 471 3523 505
rect 3489 379 3523 413
rect 3575 573 3609 607
rect 3575 476 3609 510
rect 3575 379 3609 413
<< poly >>
rect 113 609 143 635
rect 215 609 245 635
rect 293 609 323 635
rect 407 609 437 635
rect 1047 612 1273 642
rect 1047 597 1077 612
rect 810 539 840 565
rect 113 455 143 481
rect 94 425 143 455
rect 94 377 124 425
rect 215 377 245 481
rect 44 361 124 377
rect 44 327 60 361
rect 94 327 124 361
rect 44 293 124 327
rect 44 259 60 293
rect 94 259 124 293
rect 44 243 124 259
rect 94 203 124 243
rect 172 361 245 377
rect 172 327 195 361
rect 229 327 245 361
rect 172 293 245 327
rect 172 259 195 293
rect 229 259 245 293
rect 172 243 245 259
rect 293 359 323 481
rect 407 401 437 481
rect 598 435 628 461
rect 407 371 480 401
rect 293 343 359 359
rect 293 309 309 343
rect 343 309 359 343
rect 293 275 359 309
rect 172 203 202 243
rect 293 241 309 275
rect 343 241 359 275
rect 450 355 516 371
rect 450 321 466 355
rect 500 321 516 355
rect 450 287 516 321
rect 1243 547 1273 612
rect 1345 615 2211 645
rect 2598 619 2628 645
rect 2684 619 2714 645
rect 2762 619 2792 645
rect 3056 619 3086 645
rect 3142 619 3172 645
rect 3448 619 3478 645
rect 3534 619 3564 645
rect 1345 547 1375 615
rect 2181 596 2211 615
rect 1423 547 1453 573
rect 1652 547 1682 573
rect 1766 547 1796 573
rect 1844 547 1874 573
rect 2086 547 2116 573
rect 810 356 840 411
rect 774 340 840 356
rect 450 267 466 287
rect 293 225 359 241
rect 407 253 466 267
rect 500 253 516 287
rect 407 237 516 253
rect 598 248 628 307
rect 293 203 323 225
rect 407 203 437 237
rect 564 218 628 248
rect 774 306 790 340
rect 824 306 840 340
rect 1047 335 1077 469
rect 1243 437 1273 463
rect 774 272 840 306
rect 774 238 790 272
rect 824 238 840 272
rect 774 222 840 238
rect 564 203 594 218
rect 810 179 840 222
rect 888 319 1077 335
rect 888 285 904 319
rect 938 285 1077 319
rect 888 251 1077 285
rect 1123 389 1189 397
rect 1345 389 1375 463
rect 1423 431 1453 463
rect 1423 415 1546 431
rect 1423 401 1496 415
rect 1123 381 1375 389
rect 1123 347 1139 381
rect 1173 359 1375 381
rect 1452 381 1496 401
rect 1530 381 1546 415
rect 1452 365 1546 381
rect 2283 590 2313 616
rect 2452 590 2482 616
rect 2283 491 2313 506
rect 2283 461 2404 491
rect 2338 458 2404 461
rect 2452 458 2482 506
rect 2181 413 2211 428
rect 2338 424 2354 458
rect 2388 424 2404 458
rect 2181 383 2296 413
rect 1173 347 1189 359
rect 1123 313 1189 347
rect 1123 279 1139 313
rect 1173 279 1189 313
rect 1123 263 1189 279
rect 888 217 904 251
rect 938 217 1077 251
rect 1243 221 1273 359
rect 1329 293 1404 309
rect 1329 259 1354 293
rect 1388 259 1404 293
rect 1329 243 1404 259
rect 1329 221 1359 243
rect 1452 221 1482 365
rect 1652 309 1682 379
rect 1766 347 1796 379
rect 1730 331 1796 347
rect 1622 293 1688 309
rect 1622 259 1638 293
rect 1672 259 1688 293
rect 1622 243 1688 259
rect 1730 297 1746 331
rect 1780 297 1796 331
rect 1730 281 1796 297
rect 1640 221 1670 243
rect 1730 221 1760 281
rect 1844 266 1874 379
rect 2086 347 2116 379
rect 2034 331 2116 347
rect 2034 297 2050 331
rect 2084 297 2116 331
rect 2034 281 2116 297
rect 888 201 1077 217
rect 94 93 124 119
rect 172 51 202 119
rect 293 93 323 119
rect 407 93 437 119
rect 564 51 594 119
rect 1047 151 1077 201
rect 810 69 840 95
rect 1243 111 1273 137
rect 172 21 594 51
rect 1047 52 1077 67
rect 1329 52 1359 137
rect 1452 111 1482 137
rect 1840 236 1874 266
rect 2086 247 2116 281
rect 2158 319 2224 335
rect 2158 285 2174 319
rect 2208 285 2224 319
rect 2158 269 2224 285
rect 2266 292 2296 383
rect 2338 390 2404 424
rect 2338 356 2354 390
rect 2388 356 2404 390
rect 2338 340 2404 356
rect 2446 442 2512 458
rect 2954 495 2984 521
rect 2446 408 2462 442
rect 2496 408 2512 442
rect 2598 436 2628 451
rect 2446 392 2512 408
rect 2560 406 2628 436
rect 2446 292 2476 392
rect 2560 335 2590 406
rect 2684 358 2714 451
rect 2188 247 2218 269
rect 2266 262 2367 292
rect 2337 247 2367 262
rect 2415 262 2476 292
rect 2524 319 2590 335
rect 2524 285 2540 319
rect 2574 285 2590 319
rect 2632 342 2714 358
rect 2632 308 2648 342
rect 2682 308 2714 342
rect 2632 292 2714 308
rect 2762 409 2792 451
rect 2762 393 2868 409
rect 2762 359 2818 393
rect 2852 359 2868 393
rect 3346 524 3376 550
rect 3346 381 3376 396
rect 2762 325 2868 359
rect 2954 335 2984 367
rect 2524 269 2590 285
rect 2415 247 2445 262
rect 2544 247 2574 269
rect 2662 247 2692 292
rect 2762 291 2818 325
rect 2852 291 2868 325
rect 2762 275 2868 291
rect 2918 319 2984 335
rect 3056 327 3086 367
rect 2918 285 2934 319
rect 2968 299 2984 319
rect 3033 311 3099 327
rect 2968 285 2985 299
rect 1840 221 1870 236
rect 2337 137 2367 163
rect 2415 137 2445 163
rect 2762 244 2792 275
rect 2918 269 2985 285
rect 2757 214 2792 244
rect 2955 221 2985 269
rect 3033 277 3049 311
rect 3083 291 3099 311
rect 3142 291 3172 367
rect 3250 351 3376 381
rect 3250 291 3280 351
rect 3448 303 3478 367
rect 3083 277 3280 291
rect 3033 261 3280 277
rect 3057 221 3087 261
rect 3143 221 3173 261
rect 2757 199 2787 214
rect 2086 93 2116 119
rect 2188 93 2218 119
rect 1640 67 1670 93
rect 1730 67 1760 93
rect 1047 22 1359 52
rect 1840 51 1870 93
rect 2544 93 2574 119
rect 2662 93 2692 119
rect 2955 111 2985 137
rect 2757 51 2787 71
rect 3250 189 3280 261
rect 3387 287 3478 303
rect 3387 253 3403 287
rect 3437 267 3478 287
rect 3534 267 3564 367
rect 3437 253 3564 267
rect 3387 237 3564 253
rect 3448 215 3478 237
rect 3534 215 3564 237
rect 3250 159 3376 189
rect 3346 131 3376 159
rect 1840 21 2787 51
rect 3057 27 3087 53
rect 3143 27 3173 53
rect 3346 21 3376 47
rect 3448 21 3478 47
rect 3534 21 3564 47
<< polycont >>
rect 60 327 94 361
rect 60 259 94 293
rect 195 327 229 361
rect 195 259 229 293
rect 309 309 343 343
rect 309 241 343 275
rect 466 321 500 355
rect 466 253 500 287
rect 790 306 824 340
rect 790 238 824 272
rect 904 285 938 319
rect 1139 347 1173 381
rect 1496 381 1530 415
rect 2354 424 2388 458
rect 1139 279 1173 313
rect 904 217 938 251
rect 1354 259 1388 293
rect 1638 259 1672 293
rect 1746 297 1780 331
rect 2050 297 2084 331
rect 2174 285 2208 319
rect 2354 356 2388 390
rect 2462 408 2496 442
rect 2540 285 2574 319
rect 2648 308 2682 342
rect 2818 359 2852 393
rect 2818 291 2852 325
rect 2934 285 2968 319
rect 3049 277 3083 311
rect 3403 253 3437 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3648 683
rect 52 597 118 613
rect 52 563 68 597
rect 102 563 118 597
rect 52 527 118 563
rect 52 493 68 527
rect 102 493 118 527
rect 52 447 118 493
rect 154 565 220 649
rect 154 531 170 565
rect 204 531 220 565
rect 154 483 220 531
rect 260 597 498 613
rect 260 579 448 597
rect 260 447 294 579
rect 432 563 448 579
rect 482 563 498 597
rect 52 413 294 447
rect 330 535 396 543
rect 330 501 346 535
rect 380 501 396 535
rect 330 441 396 501
rect 432 527 498 563
rect 432 493 448 527
rect 482 493 498 527
rect 432 477 498 493
rect 544 535 610 649
rect 544 501 560 535
rect 594 501 610 535
rect 544 485 610 501
rect 729 527 779 649
rect 729 493 745 527
rect 729 477 779 493
rect 815 579 1036 613
rect 815 441 849 579
rect 330 407 849 441
rect 885 527 954 543
rect 919 493 954 527
rect 885 457 954 493
rect 1002 499 1036 579
rect 1072 585 1138 649
rect 1072 551 1088 585
rect 1122 551 1138 585
rect 1072 535 1138 551
rect 1182 522 1248 551
rect 1182 499 1198 522
rect 1002 488 1198 499
rect 1232 488 1248 522
rect 1002 465 1248 488
rect 1182 459 1248 465
rect 919 423 954 457
rect 25 361 110 377
rect 25 327 60 361
rect 94 327 110 361
rect 25 293 110 327
rect 25 259 60 293
rect 94 259 110 293
rect 25 243 110 259
rect 179 361 263 377
rect 179 327 195 361
rect 229 327 263 361
rect 179 293 263 327
rect 179 259 195 293
rect 229 259 263 293
rect 179 243 263 259
rect 299 343 359 359
rect 299 309 309 343
rect 343 309 359 343
rect 299 275 359 309
rect 299 241 309 275
rect 343 241 359 275
rect 33 178 99 207
rect 33 144 49 178
rect 83 144 99 178
rect 33 17 99 144
rect 197 178 263 207
rect 197 144 213 178
rect 247 144 263 178
rect 299 162 359 241
rect 197 126 263 144
rect 395 126 429 407
rect 465 355 689 371
rect 465 321 466 355
rect 500 354 689 355
rect 500 321 639 354
rect 465 320 639 321
rect 673 320 689 354
rect 465 303 689 320
rect 465 287 516 303
rect 465 253 466 287
rect 500 253 516 287
rect 465 237 516 253
rect 197 92 429 126
rect 465 175 531 201
rect 465 141 481 175
rect 515 141 531 175
rect 465 17 531 141
rect 589 178 689 303
rect 774 340 840 356
rect 774 306 790 340
rect 824 306 840 340
rect 774 272 840 306
rect 774 238 790 272
rect 824 238 840 272
rect 774 222 840 238
rect 885 319 954 423
rect 885 285 904 319
rect 938 285 954 319
rect 885 251 954 285
rect 885 217 904 251
rect 938 217 954 251
rect 885 201 954 217
rect 990 413 1040 429
rect 1024 397 1040 413
rect 1024 381 1178 397
rect 1024 379 1139 381
rect 990 363 1139 379
rect 885 183 919 201
rect 589 144 605 178
rect 639 144 689 178
rect 589 115 689 144
rect 733 154 799 183
rect 733 120 749 154
rect 783 120 799 154
rect 733 17 799 120
rect 835 154 919 183
rect 990 155 1040 363
rect 1123 347 1139 363
rect 1173 347 1178 381
rect 1123 313 1178 347
rect 1123 279 1139 313
rect 1173 279 1178 313
rect 1123 263 1178 279
rect 1214 225 1248 459
rect 1182 196 1248 225
rect 1182 162 1198 196
rect 1232 162 1248 196
rect 835 120 851 154
rect 885 120 919 154
rect 835 91 919 120
rect 974 126 1040 155
rect 974 92 990 126
rect 1024 92 1040 126
rect 974 63 1040 92
rect 1076 126 1142 155
rect 1182 133 1248 162
rect 1284 522 1350 551
rect 1284 488 1300 522
rect 1334 488 1350 522
rect 1284 449 1350 488
rect 1591 535 1657 649
rect 1591 501 1607 535
rect 1641 501 1657 535
rect 1591 485 1657 501
rect 1705 535 1866 551
rect 1705 501 1721 535
rect 1755 501 1866 535
rect 1705 465 1866 501
rect 1705 449 1721 465
rect 1284 415 1459 449
rect 1284 196 1318 415
rect 1425 329 1459 415
rect 1495 431 1721 449
rect 1755 431 1866 465
rect 1495 415 1866 431
rect 1495 381 1496 415
rect 1530 381 1531 415
rect 1495 365 1531 381
rect 1567 345 1796 379
rect 1567 329 1601 345
rect 1354 293 1389 309
rect 1425 295 1601 329
rect 1741 331 1796 345
rect 1388 259 1389 293
rect 1354 200 1389 259
rect 1637 293 1703 309
rect 1637 259 1638 293
rect 1672 276 1703 293
rect 1741 297 1746 331
rect 1780 297 1796 331
rect 1741 281 1796 297
rect 1832 323 1866 415
rect 1902 535 1968 649
rect 1902 501 1918 535
rect 1952 501 1968 535
rect 1902 425 1968 501
rect 1902 391 1918 425
rect 1952 391 1968 425
rect 1902 375 1968 391
rect 2136 579 2404 613
rect 2034 331 2100 341
rect 2034 323 2050 331
rect 1832 297 2050 323
rect 2084 297 2100 331
rect 1832 289 2100 297
rect 2136 335 2170 579
rect 2206 500 2294 543
rect 2206 466 2222 500
rect 2256 466 2294 500
rect 2206 424 2294 466
rect 2136 319 2224 335
rect 1637 242 1663 259
rect 1697 242 1703 276
rect 1832 245 1866 289
rect 2136 285 2174 319
rect 2208 285 2224 319
rect 2136 253 2224 285
rect 1637 236 1703 242
rect 1767 243 1866 245
rect 1767 209 1783 243
rect 1817 211 1866 243
rect 1971 219 2224 253
rect 2260 251 2294 424
rect 2338 458 2404 579
rect 2537 575 2587 649
rect 2537 541 2553 575
rect 2537 494 2587 541
rect 2623 597 2689 613
rect 2623 563 2639 597
rect 2673 563 2689 597
rect 2623 512 2689 563
rect 2787 602 2853 649
rect 2787 568 2803 602
rect 2837 568 2853 602
rect 2787 548 2853 568
rect 2995 602 3061 649
rect 2995 568 3011 602
rect 3045 568 3061 602
rect 2995 548 3061 568
rect 3097 597 3153 613
rect 3131 563 3153 597
rect 2623 497 3061 512
rect 2623 463 2639 497
rect 2673 478 3061 497
rect 2673 463 2689 478
rect 2623 458 2689 463
rect 2338 424 2354 458
rect 2388 424 2404 458
rect 2338 390 2404 424
rect 2446 442 2689 458
rect 2446 408 2462 442
rect 2496 424 2689 442
rect 2496 408 2512 424
rect 2446 392 2512 408
rect 2338 356 2354 390
rect 2388 356 2404 390
rect 2338 340 2404 356
rect 2521 319 2590 356
rect 2521 285 2540 319
rect 2574 285 2590 319
rect 2521 276 2590 285
rect 2260 235 2326 251
rect 2521 242 2527 276
rect 2561 242 2590 276
rect 2521 236 2590 242
rect 2626 342 2697 358
rect 2626 308 2648 342
rect 2682 308 2697 342
rect 2626 292 2697 308
rect 1817 209 1833 211
rect 1354 166 1629 200
rect 1284 133 1318 162
rect 1076 92 1092 126
rect 1126 92 1142 126
rect 1076 17 1142 92
rect 1493 114 1559 130
rect 1493 80 1509 114
rect 1543 80 1559 114
rect 1493 17 1559 80
rect 1595 87 1629 166
rect 1665 178 1731 200
rect 1767 193 1833 209
rect 1665 144 1681 178
rect 1715 157 1731 178
rect 1869 174 1935 175
rect 1869 157 1885 174
rect 1715 144 1885 157
rect 1665 140 1885 144
rect 1919 140 1935 174
rect 1665 123 1935 140
rect 1971 87 2005 219
rect 2260 201 2276 235
rect 2310 201 2326 235
rect 2260 200 2326 201
rect 2626 200 2660 292
rect 2733 233 2767 478
rect 1595 53 2005 87
rect 2041 166 2091 183
rect 2075 132 2091 166
rect 2041 17 2091 132
rect 2260 166 2660 200
rect 2696 199 2767 233
rect 2803 408 2909 442
rect 2943 408 2959 442
rect 2803 393 2959 408
rect 2803 359 2818 393
rect 2852 392 2959 393
rect 2852 359 2868 392
rect 2803 325 2868 359
rect 2803 291 2818 325
rect 2852 291 2868 325
rect 2803 233 2868 291
rect 2905 319 2984 356
rect 2905 285 2934 319
rect 2968 285 2984 319
rect 2905 269 2984 285
rect 3027 327 3061 478
rect 3097 505 3153 563
rect 3131 471 3153 505
rect 3097 413 3153 471
rect 3131 379 3153 413
rect 3097 363 3153 379
rect 3189 607 3239 649
rect 3223 573 3239 607
rect 3189 510 3239 573
rect 3387 607 3437 649
rect 3387 573 3403 607
rect 3223 476 3239 510
rect 3189 413 3239 476
rect 3223 379 3239 413
rect 3189 363 3239 379
rect 3285 512 3351 528
rect 3285 478 3301 512
rect 3335 478 3351 512
rect 3285 442 3351 478
rect 3285 408 3301 442
rect 3335 408 3351 442
rect 3027 311 3083 327
rect 3027 277 3049 311
rect 3027 261 3083 277
rect 2803 199 2960 233
rect 3119 225 3153 363
rect 3285 303 3351 408
rect 3387 510 3437 573
rect 3387 476 3403 510
rect 3387 413 3437 476
rect 3387 379 3403 413
rect 3387 363 3437 379
rect 3473 597 3539 613
rect 3473 563 3489 597
rect 3523 563 3539 597
rect 3473 505 3539 563
rect 3473 471 3489 505
rect 3523 471 3539 505
rect 3473 413 3539 471
rect 3473 379 3489 413
rect 3523 379 3539 413
rect 3285 287 3437 303
rect 3285 253 3403 287
rect 3285 237 3437 253
rect 2696 180 2762 199
rect 2260 165 2326 166
rect 2260 131 2276 165
rect 2310 131 2326 165
rect 2260 115 2326 131
rect 2696 146 2712 180
rect 2746 146 2762 180
rect 2894 196 2960 199
rect 2467 114 2533 130
rect 2467 80 2483 114
rect 2517 80 2533 114
rect 2467 17 2533 80
rect 2585 114 2651 130
rect 2696 123 2762 146
rect 2798 132 2848 163
rect 2894 162 2910 196
rect 2944 162 2960 196
rect 2894 133 2960 162
rect 2996 209 3046 225
rect 2996 175 3012 209
rect 2585 80 2601 114
rect 2635 87 2651 114
rect 2832 98 2848 132
rect 2798 87 2848 98
rect 2635 80 2848 87
rect 2585 53 2848 80
rect 2996 99 3046 175
rect 2996 65 3012 99
rect 2996 17 3046 65
rect 3082 209 3153 225
rect 3082 175 3098 209
rect 3132 175 3153 209
rect 3082 103 3153 175
rect 3082 69 3098 103
rect 3132 69 3153 103
rect 3082 53 3153 69
rect 3189 209 3239 225
rect 3223 175 3239 209
rect 3189 99 3239 175
rect 3223 65 3239 99
rect 3189 17 3239 65
rect 3285 106 3351 237
rect 3473 203 3539 379
rect 3575 607 3625 649
rect 3609 573 3625 607
rect 3575 510 3625 573
rect 3609 476 3625 510
rect 3575 413 3625 476
rect 3609 379 3625 413
rect 3575 363 3625 379
rect 3285 72 3301 106
rect 3335 72 3351 106
rect 3285 59 3351 72
rect 3387 185 3437 201
rect 3387 151 3403 185
rect 3387 93 3437 151
rect 3387 59 3403 93
rect 3387 17 3437 59
rect 3473 169 3489 203
rect 3523 169 3539 203
rect 3473 103 3539 169
rect 3473 69 3489 103
rect 3523 69 3539 103
rect 3473 53 3539 69
rect 3575 203 3625 219
rect 3609 169 3625 203
rect 3575 93 3625 169
rect 3609 59 3625 93
rect 3575 17 3625 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3648 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 3583 649 3617 683
rect 1663 259 1672 276
rect 1672 259 1697 276
rect 1663 242 1697 259
rect 2527 242 2561 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
<< metal1 >>
rect 0 683 3648 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3648 683
rect 0 617 3648 649
rect 1651 276 1709 282
rect 1651 242 1663 276
rect 1697 273 1709 276
rect 2515 276 2573 282
rect 2515 273 2527 276
rect 1697 245 2527 273
rect 1697 242 1709 245
rect 1651 236 1709 242
rect 2515 242 2527 245
rect 2561 242 2573 276
rect 2515 236 2573 242
rect 0 17 3648 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3648 17
rect 0 -49 3648 -17
<< labels >>
flabel pwell s 0 0 3648 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 3648 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfbbn_2
flabel comment s 1055 266 1055 266 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 3648 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 3648 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 2911 316 2945 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 2527 316 2561 350 0 FreeSans 340 0 0 0 SET_B
port 6 nsew signal input
flabel locali s 3487 94 3521 128 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 3487 168 3521 202 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 3487 242 3521 276 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 3487 316 3521 350 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 3487 390 3521 424 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 3487 464 3521 498 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 3487 538 3521 572 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 3103 390 3137 424 0 FreeSans 340 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 3103 464 3137 498 0 FreeSans 340 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 3103 538 3137 572 0 FreeSans 340 0 0 0 Q_N
port 12 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3648 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2967930
string GDS_START 2943182
<< end >>
