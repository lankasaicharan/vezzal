magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 103 228 292 248
rect 103 210 959 228
rect 1 49 959 210
rect 0 0 960 49
<< scpmos >>
rect 83 368 119 536
rect 190 368 226 592
rect 419 424 455 592
rect 519 424 555 592
rect 629 424 665 592
rect 719 424 755 592
rect 833 424 869 592
<< nmoslvt >>
rect 84 74 114 184
rect 179 74 209 222
rect 425 74 455 202
rect 503 74 533 202
rect 617 74 647 202
rect 719 74 749 202
rect 846 92 876 202
<< ndiff >>
rect 129 184 179 222
rect 27 146 84 184
rect 27 112 39 146
rect 73 112 84 146
rect 27 74 84 112
rect 114 142 179 184
rect 114 108 125 142
rect 159 108 179 142
rect 114 74 179 108
rect 209 210 266 222
rect 209 176 220 210
rect 254 176 266 210
rect 209 120 266 176
rect 209 86 220 120
rect 254 86 266 120
rect 209 74 266 86
rect 368 190 425 202
rect 368 156 380 190
rect 414 156 425 190
rect 368 120 425 156
rect 368 86 380 120
rect 414 86 425 120
rect 368 74 425 86
rect 455 74 503 202
rect 533 74 617 202
rect 647 74 719 202
rect 749 120 846 202
rect 749 86 772 120
rect 806 92 846 120
rect 876 164 933 202
rect 876 130 887 164
rect 921 130 933 164
rect 876 92 933 130
rect 806 86 831 92
rect 749 74 831 86
<< pdiff >>
rect 134 573 190 592
rect 134 539 146 573
rect 180 539 190 573
rect 134 536 190 539
rect 27 524 83 536
rect 27 490 39 524
rect 73 490 83 524
rect 27 440 83 490
rect 27 406 39 440
rect 73 406 83 440
rect 27 368 83 406
rect 119 368 190 536
rect 226 414 309 592
rect 363 573 419 592
rect 363 539 375 573
rect 409 539 419 573
rect 363 424 419 539
rect 455 580 519 592
rect 455 546 475 580
rect 509 546 519 580
rect 455 470 519 546
rect 455 436 475 470
rect 509 436 519 470
rect 455 424 519 436
rect 555 584 629 592
rect 555 550 575 584
rect 609 550 629 584
rect 555 508 629 550
rect 555 474 575 508
rect 609 474 629 508
rect 555 424 629 474
rect 665 580 719 592
rect 665 546 675 580
rect 709 546 719 580
rect 665 470 719 546
rect 665 436 675 470
rect 709 436 719 470
rect 665 424 719 436
rect 755 580 833 592
rect 755 546 779 580
rect 813 546 833 580
rect 755 495 833 546
rect 755 461 779 495
rect 813 461 833 495
rect 755 424 833 461
rect 869 580 925 592
rect 869 546 879 580
rect 913 546 925 580
rect 869 470 925 546
rect 869 436 879 470
rect 913 436 925 470
rect 869 424 925 436
rect 226 380 249 414
rect 283 380 309 414
rect 226 368 309 380
<< ndiffc >>
rect 39 112 73 146
rect 125 108 159 142
rect 220 176 254 210
rect 220 86 254 120
rect 380 156 414 190
rect 380 86 414 120
rect 772 86 806 120
rect 887 130 921 164
<< pdiffc >>
rect 146 539 180 573
rect 39 490 73 524
rect 39 406 73 440
rect 375 539 409 573
rect 475 546 509 580
rect 475 436 509 470
rect 575 550 609 584
rect 575 474 609 508
rect 675 546 709 580
rect 675 436 709 470
rect 779 546 813 580
rect 779 461 813 495
rect 879 546 913 580
rect 879 436 913 470
rect 249 380 283 414
<< poly >>
rect 190 592 226 618
rect 419 592 455 618
rect 519 592 555 618
rect 629 592 665 618
rect 719 592 755 618
rect 833 592 869 618
rect 83 536 119 562
rect 419 392 455 424
rect 351 376 455 392
rect 83 326 119 368
rect 21 310 119 326
rect 21 276 37 310
rect 71 276 119 310
rect 190 326 226 368
rect 351 342 367 376
rect 401 342 455 376
rect 519 358 555 424
rect 629 372 665 424
rect 719 372 755 424
rect 190 310 309 326
rect 190 290 259 310
rect 21 260 119 276
rect 179 276 259 290
rect 293 276 309 310
rect 179 260 309 276
rect 351 308 455 342
rect 351 274 367 308
rect 401 274 455 308
rect 84 184 114 260
rect 179 222 209 260
rect 351 258 455 274
rect 425 202 455 258
rect 503 342 569 358
rect 503 308 519 342
rect 553 308 569 342
rect 503 274 569 308
rect 503 240 519 274
rect 553 240 569 274
rect 503 224 569 240
rect 611 356 677 372
rect 611 322 627 356
rect 661 322 677 356
rect 611 288 677 322
rect 611 254 627 288
rect 661 254 677 288
rect 611 238 677 254
rect 719 356 785 372
rect 719 322 735 356
rect 769 322 785 356
rect 719 288 785 322
rect 719 254 735 288
rect 769 254 785 288
rect 833 326 869 424
rect 833 310 939 326
rect 833 276 889 310
rect 923 276 939 310
rect 833 260 939 276
rect 719 238 785 254
rect 503 202 533 224
rect 617 202 647 238
rect 719 202 749 238
rect 846 202 876 260
rect 84 48 114 74
rect 179 48 209 74
rect 425 48 455 74
rect 503 48 533 74
rect 617 48 647 74
rect 719 48 749 74
rect 846 66 876 92
<< polycont >>
rect 37 276 71 310
rect 367 342 401 376
rect 259 276 293 310
rect 367 274 401 308
rect 519 308 553 342
rect 519 240 553 274
rect 627 322 661 356
rect 627 254 661 288
rect 735 322 769 356
rect 735 254 769 288
rect 889 276 923 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 130 573 196 649
rect 23 524 89 540
rect 130 539 146 573
rect 180 539 196 573
rect 130 532 196 539
rect 359 573 425 649
rect 359 539 375 573
rect 409 539 425 573
rect 359 532 425 539
rect 459 580 525 596
rect 459 546 475 580
rect 509 546 525 580
rect 23 490 39 524
rect 73 498 89 524
rect 73 490 409 498
rect 23 464 409 490
rect 23 440 148 464
rect 23 406 39 440
rect 73 406 148 440
rect 23 390 148 406
rect 21 310 80 356
rect 21 276 37 310
rect 71 276 80 310
rect 21 260 80 276
rect 114 226 148 390
rect 23 192 148 226
rect 182 414 313 430
rect 182 380 249 414
rect 283 380 313 414
rect 182 364 313 380
rect 356 376 409 464
rect 459 470 525 546
rect 559 584 625 649
rect 559 550 575 584
rect 609 550 625 584
rect 559 508 625 550
rect 559 474 575 508
rect 609 474 625 508
rect 659 580 725 596
rect 659 546 675 580
rect 709 546 725 580
rect 459 440 475 470
rect 182 226 216 364
rect 356 342 367 376
rect 401 342 409 376
rect 250 310 322 326
rect 250 276 259 310
rect 293 276 322 310
rect 250 260 322 276
rect 182 210 254 226
rect 182 192 220 210
rect 23 146 73 192
rect 216 176 220 192
rect 23 112 39 146
rect 23 70 73 112
rect 109 142 175 158
rect 109 108 125 142
rect 159 108 175 142
rect 109 17 175 108
rect 216 120 254 176
rect 288 206 322 260
rect 356 308 409 342
rect 356 274 367 308
rect 401 274 409 308
rect 356 258 409 274
rect 443 436 475 440
rect 509 440 525 470
rect 659 470 725 546
rect 659 440 675 470
rect 509 436 675 440
rect 709 436 725 470
rect 763 580 829 649
rect 763 546 779 580
rect 813 546 829 580
rect 763 495 829 546
rect 763 461 779 495
rect 813 461 829 495
rect 763 458 829 461
rect 863 580 929 596
rect 863 546 879 580
rect 913 546 929 580
rect 863 470 929 546
rect 443 406 725 436
rect 863 436 879 470
rect 913 436 929 470
rect 863 424 929 436
rect 443 206 477 406
rect 812 390 929 424
rect 288 190 477 206
rect 288 172 380 190
rect 216 86 220 120
rect 216 70 254 86
rect 364 156 380 172
rect 414 156 477 190
rect 511 342 569 358
rect 511 308 519 342
rect 553 308 569 342
rect 511 274 569 308
rect 511 240 519 274
rect 553 240 569 274
rect 511 204 569 240
rect 603 356 669 372
rect 603 322 627 356
rect 661 322 669 356
rect 603 288 669 322
rect 603 254 627 288
rect 661 254 669 288
rect 603 238 669 254
rect 703 356 778 372
rect 703 322 735 356
rect 769 322 778 356
rect 703 288 778 322
rect 703 254 735 288
rect 769 254 778 288
rect 703 238 778 254
rect 812 206 846 390
rect 880 310 939 356
rect 880 276 889 310
rect 923 276 939 310
rect 880 260 939 276
rect 812 204 937 206
rect 511 170 937 204
rect 364 120 477 156
rect 871 164 937 170
rect 364 86 380 120
rect 414 86 477 120
rect 364 70 477 86
rect 744 120 822 136
rect 744 86 772 120
rect 806 86 822 120
rect 871 130 887 164
rect 921 130 937 164
rect 871 88 937 130
rect 744 17 822 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4bb_1
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 3088518
string GDS_START 3080798
<< end >>
