magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 7 49 1500 241
rect 0 0 1536 49
<< scnmos >>
rect 86 47 116 215
rect 172 47 202 215
rect 258 47 288 215
rect 344 47 374 215
rect 430 47 460 215
rect 516 47 546 215
rect 602 47 632 215
rect 688 47 718 215
rect 785 47 815 215
rect 871 47 901 215
rect 957 47 987 215
rect 1043 47 1073 215
rect 1129 47 1159 215
rect 1215 47 1245 215
rect 1301 47 1331 215
rect 1387 47 1417 215
<< scpmoshvt >>
rect 89 367 119 619
rect 175 367 205 619
rect 261 367 291 619
rect 347 367 377 619
rect 433 367 463 619
rect 519 367 549 619
rect 605 367 635 619
rect 691 367 721 619
rect 791 367 821 619
rect 877 367 907 619
rect 963 367 993 619
rect 1049 367 1079 619
rect 1135 367 1165 619
rect 1221 367 1251 619
rect 1307 367 1337 619
rect 1393 367 1423 619
<< ndiff >>
rect 33 203 86 215
rect 33 169 41 203
rect 75 169 86 203
rect 33 101 86 169
rect 33 67 41 101
rect 75 67 86 101
rect 33 47 86 67
rect 116 165 172 215
rect 116 131 127 165
rect 161 131 172 165
rect 116 93 172 131
rect 116 59 127 93
rect 161 59 172 93
rect 116 47 172 59
rect 202 203 258 215
rect 202 169 213 203
rect 247 169 258 203
rect 202 101 258 169
rect 202 67 213 101
rect 247 67 258 101
rect 202 47 258 67
rect 288 165 344 215
rect 288 131 299 165
rect 333 131 344 165
rect 288 93 344 131
rect 288 59 299 93
rect 333 59 344 93
rect 288 47 344 59
rect 374 203 430 215
rect 374 169 385 203
rect 419 169 430 203
rect 374 101 430 169
rect 374 67 385 101
rect 419 67 430 101
rect 374 47 430 67
rect 460 165 516 215
rect 460 131 471 165
rect 505 131 516 165
rect 460 93 516 131
rect 460 59 471 93
rect 505 59 516 93
rect 460 47 516 59
rect 546 203 602 215
rect 546 169 557 203
rect 591 169 602 203
rect 546 101 602 169
rect 546 67 557 101
rect 591 67 602 101
rect 546 47 602 67
rect 632 165 688 215
rect 632 131 643 165
rect 677 131 688 165
rect 632 93 688 131
rect 632 59 643 93
rect 677 59 688 93
rect 632 47 688 59
rect 718 203 785 215
rect 718 169 729 203
rect 763 169 785 203
rect 718 101 785 169
rect 718 67 729 101
rect 763 67 785 101
rect 718 47 785 67
rect 815 169 871 215
rect 815 135 826 169
rect 860 135 871 169
rect 815 47 871 135
rect 901 91 957 215
rect 901 57 912 91
rect 946 57 957 91
rect 901 47 957 57
rect 987 165 1043 215
rect 987 131 998 165
rect 1032 131 1043 165
rect 987 47 1043 131
rect 1073 91 1129 215
rect 1073 57 1084 91
rect 1118 57 1129 91
rect 1073 47 1129 57
rect 1159 165 1215 215
rect 1159 131 1170 165
rect 1204 131 1215 165
rect 1159 47 1215 131
rect 1245 91 1301 215
rect 1245 57 1256 91
rect 1290 57 1301 91
rect 1245 47 1301 57
rect 1331 165 1387 215
rect 1331 131 1342 165
rect 1376 131 1387 165
rect 1331 47 1387 131
rect 1417 91 1474 215
rect 1417 57 1428 91
rect 1462 57 1474 91
rect 1417 47 1474 57
<< pdiff >>
rect 36 607 89 619
rect 36 573 44 607
rect 78 573 89 607
rect 36 506 89 573
rect 36 472 44 506
rect 78 472 89 506
rect 36 413 89 472
rect 36 379 44 413
rect 78 379 89 413
rect 36 367 89 379
rect 119 599 175 619
rect 119 565 130 599
rect 164 565 175 599
rect 119 505 175 565
rect 119 471 130 505
rect 164 471 175 505
rect 119 413 175 471
rect 119 379 130 413
rect 164 379 175 413
rect 119 367 175 379
rect 205 576 261 619
rect 205 542 216 576
rect 250 542 261 576
rect 205 367 261 542
rect 291 599 347 619
rect 291 565 302 599
rect 336 565 347 599
rect 291 508 347 565
rect 291 474 302 508
rect 336 474 347 508
rect 291 367 347 474
rect 377 508 433 619
rect 377 474 388 508
rect 422 474 433 508
rect 377 367 433 474
rect 463 600 519 619
rect 463 566 474 600
rect 508 566 519 600
rect 463 367 519 566
rect 549 508 605 619
rect 549 474 560 508
rect 594 474 605 508
rect 549 367 605 474
rect 635 600 691 619
rect 635 566 646 600
rect 680 566 691 600
rect 635 367 691 566
rect 721 578 791 619
rect 721 544 741 578
rect 775 544 791 578
rect 721 367 791 544
rect 821 599 877 619
rect 821 565 832 599
rect 866 565 877 599
rect 821 529 877 565
rect 821 495 832 529
rect 866 495 877 529
rect 821 459 877 495
rect 821 425 832 459
rect 866 425 877 459
rect 821 367 877 425
rect 907 607 963 619
rect 907 573 918 607
rect 952 573 963 607
rect 907 520 963 573
rect 907 486 918 520
rect 952 486 963 520
rect 907 367 963 486
rect 993 597 1049 619
rect 993 563 1004 597
rect 1038 563 1049 597
rect 993 529 1049 563
rect 993 495 1004 529
rect 1038 495 1049 529
rect 993 459 1049 495
rect 993 425 1004 459
rect 1038 425 1049 459
rect 993 367 1049 425
rect 1079 540 1135 619
rect 1079 506 1090 540
rect 1124 506 1135 540
rect 1079 413 1135 506
rect 1079 379 1090 413
rect 1124 379 1135 413
rect 1079 367 1135 379
rect 1165 599 1221 619
rect 1165 565 1176 599
rect 1210 565 1221 599
rect 1165 504 1221 565
rect 1165 470 1176 504
rect 1210 470 1221 504
rect 1165 367 1221 470
rect 1251 540 1307 619
rect 1251 506 1262 540
rect 1296 506 1307 540
rect 1251 413 1307 506
rect 1251 379 1262 413
rect 1296 379 1307 413
rect 1251 367 1307 379
rect 1337 599 1393 619
rect 1337 565 1348 599
rect 1382 565 1393 599
rect 1337 529 1393 565
rect 1337 495 1348 529
rect 1382 495 1393 529
rect 1337 459 1393 495
rect 1337 425 1348 459
rect 1382 425 1393 459
rect 1337 367 1393 425
rect 1423 607 1476 619
rect 1423 573 1434 607
rect 1468 573 1476 607
rect 1423 529 1476 573
rect 1423 495 1434 529
rect 1468 495 1476 529
rect 1423 455 1476 495
rect 1423 421 1434 455
rect 1468 421 1476 455
rect 1423 367 1476 421
<< ndiffc >>
rect 41 169 75 203
rect 41 67 75 101
rect 127 131 161 165
rect 127 59 161 93
rect 213 169 247 203
rect 213 67 247 101
rect 299 131 333 165
rect 299 59 333 93
rect 385 169 419 203
rect 385 67 419 101
rect 471 131 505 165
rect 471 59 505 93
rect 557 169 591 203
rect 557 67 591 101
rect 643 131 677 165
rect 643 59 677 93
rect 729 169 763 203
rect 729 67 763 101
rect 826 135 860 169
rect 912 57 946 91
rect 998 131 1032 165
rect 1084 57 1118 91
rect 1170 131 1204 165
rect 1256 57 1290 91
rect 1342 131 1376 165
rect 1428 57 1462 91
<< pdiffc >>
rect 44 573 78 607
rect 44 472 78 506
rect 44 379 78 413
rect 130 565 164 599
rect 130 471 164 505
rect 130 379 164 413
rect 216 542 250 576
rect 302 565 336 599
rect 302 474 336 508
rect 388 474 422 508
rect 474 566 508 600
rect 560 474 594 508
rect 646 566 680 600
rect 741 544 775 578
rect 832 565 866 599
rect 832 495 866 529
rect 832 425 866 459
rect 918 573 952 607
rect 918 486 952 520
rect 1004 563 1038 597
rect 1004 495 1038 529
rect 1004 425 1038 459
rect 1090 506 1124 540
rect 1090 379 1124 413
rect 1176 565 1210 599
rect 1176 470 1210 504
rect 1262 506 1296 540
rect 1262 379 1296 413
rect 1348 565 1382 599
rect 1348 495 1382 529
rect 1348 425 1382 459
rect 1434 573 1468 607
rect 1434 495 1468 529
rect 1434 421 1468 455
<< poly >>
rect 89 619 119 645
rect 175 619 205 645
rect 261 619 291 645
rect 347 619 377 645
rect 433 619 463 645
rect 519 619 549 645
rect 605 619 635 645
rect 691 619 721 645
rect 791 619 821 645
rect 877 619 907 645
rect 963 619 993 645
rect 1049 619 1079 645
rect 1135 619 1165 645
rect 1221 619 1251 645
rect 1307 619 1337 645
rect 1393 619 1423 645
rect 89 325 119 367
rect 175 325 205 367
rect 261 325 291 367
rect 347 335 377 367
rect 433 335 463 367
rect 519 335 549 367
rect 605 335 635 367
rect 21 309 291 325
rect 21 275 37 309
rect 71 275 105 309
rect 139 275 173 309
rect 207 275 241 309
rect 275 275 291 309
rect 21 259 291 275
rect 344 319 635 335
rect 691 321 721 367
rect 791 321 821 367
rect 877 321 907 367
rect 963 321 993 367
rect 1049 321 1079 367
rect 1135 321 1165 367
rect 1221 321 1251 367
rect 1307 321 1337 367
rect 344 285 378 319
rect 412 285 446 319
rect 480 285 514 319
rect 548 285 582 319
rect 616 305 635 319
rect 677 305 743 321
rect 616 285 632 305
rect 344 269 632 285
rect 86 215 116 259
rect 172 215 202 259
rect 258 215 288 259
rect 344 215 374 269
rect 430 215 460 269
rect 516 215 546 269
rect 602 215 632 269
rect 677 271 693 305
rect 727 271 743 305
rect 791 305 993 321
rect 791 285 807 305
rect 677 255 743 271
rect 785 271 807 285
rect 841 271 875 305
rect 909 271 943 305
rect 977 271 993 305
rect 785 255 993 271
rect 1043 305 1337 321
rect 1043 271 1077 305
rect 1111 271 1145 305
rect 1179 271 1213 305
rect 1247 271 1281 305
rect 1315 271 1337 305
rect 1393 303 1423 367
rect 1043 255 1337 271
rect 1387 287 1453 303
rect 688 215 718 255
rect 785 215 815 255
rect 871 215 901 255
rect 957 215 987 255
rect 1043 215 1073 255
rect 1129 215 1159 255
rect 1215 215 1245 255
rect 1301 215 1331 255
rect 1387 253 1403 287
rect 1437 253 1453 287
rect 1387 237 1453 253
rect 1387 215 1417 237
rect 86 21 116 47
rect 172 21 202 47
rect 258 21 288 47
rect 344 21 374 47
rect 430 21 460 47
rect 516 21 546 47
rect 602 21 632 47
rect 688 21 718 47
rect 785 21 815 47
rect 871 21 901 47
rect 957 21 987 47
rect 1043 21 1073 47
rect 1129 21 1159 47
rect 1215 21 1245 47
rect 1301 21 1331 47
rect 1387 21 1417 47
<< polycont >>
rect 37 275 71 309
rect 105 275 139 309
rect 173 275 207 309
rect 241 275 275 309
rect 378 285 412 319
rect 446 285 480 319
rect 514 285 548 319
rect 582 285 616 319
rect 693 271 727 305
rect 807 271 841 305
rect 875 271 909 305
rect 943 271 977 305
rect 1077 271 1111 305
rect 1145 271 1179 305
rect 1213 271 1247 305
rect 1281 271 1315 305
rect 1403 253 1437 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 28 607 86 649
rect 28 573 44 607
rect 78 573 86 607
rect 28 506 86 573
rect 28 472 44 506
rect 78 472 86 506
rect 28 413 86 472
rect 28 379 44 413
rect 78 379 86 413
rect 28 363 86 379
rect 120 599 166 615
rect 120 565 130 599
rect 164 565 166 599
rect 120 505 166 565
rect 200 576 266 649
rect 200 542 216 576
rect 250 542 266 576
rect 200 526 266 542
rect 300 600 696 615
rect 300 599 474 600
rect 300 565 302 599
rect 336 566 474 599
rect 508 566 646 600
rect 680 566 696 600
rect 336 565 696 566
rect 300 558 696 565
rect 730 578 792 649
rect 120 471 130 505
rect 164 492 166 505
rect 300 508 340 558
rect 730 544 741 578
rect 775 544 792 578
rect 730 528 792 544
rect 826 599 868 615
rect 826 565 832 599
rect 866 565 868 599
rect 826 529 868 565
rect 300 492 302 508
rect 164 474 302 492
rect 336 474 340 508
rect 164 471 340 474
rect 120 458 340 471
rect 384 508 610 524
rect 384 474 388 508
rect 422 474 560 508
rect 594 494 610 508
rect 826 495 832 529
rect 866 495 868 529
rect 594 474 792 494
rect 384 458 792 474
rect 120 413 171 458
rect 120 379 130 413
rect 164 379 171 413
rect 120 363 171 379
rect 205 390 711 424
rect 205 326 291 390
rect 21 309 291 326
rect 21 275 37 309
rect 71 275 105 309
rect 139 275 173 309
rect 207 275 241 309
rect 275 275 291 309
rect 21 269 291 275
rect 362 319 641 350
rect 362 285 378 319
rect 412 285 446 319
rect 480 285 514 319
rect 548 285 582 319
rect 616 285 641 319
rect 362 269 641 285
rect 677 305 711 390
rect 758 375 792 458
rect 826 459 868 495
rect 902 607 968 649
rect 902 573 918 607
rect 952 573 968 607
rect 902 520 968 573
rect 902 486 918 520
rect 952 486 968 520
rect 902 479 968 486
rect 1002 599 1384 615
rect 1002 597 1176 599
rect 1002 563 1004 597
rect 1038 581 1176 597
rect 1038 563 1040 581
rect 1002 529 1040 563
rect 1174 565 1176 581
rect 1210 581 1348 599
rect 1210 565 1212 581
rect 1002 495 1004 529
rect 1038 495 1040 529
rect 826 425 832 459
rect 866 445 868 459
rect 1002 459 1040 495
rect 1002 445 1004 459
rect 866 425 1004 445
rect 1038 425 1040 459
rect 826 409 1040 425
rect 1074 540 1140 547
rect 1074 506 1090 540
rect 1124 506 1140 540
rect 1074 420 1140 506
rect 1174 504 1212 565
rect 1346 565 1348 581
rect 1382 565 1384 599
rect 1174 470 1176 504
rect 1210 470 1212 504
rect 1174 454 1212 470
rect 1246 540 1312 547
rect 1246 506 1262 540
rect 1296 506 1312 540
rect 1246 420 1312 506
rect 1074 413 1312 420
rect 1074 379 1090 413
rect 1124 386 1262 413
rect 1124 379 1128 386
rect 1074 375 1128 379
rect 758 341 1128 375
rect 1258 379 1262 386
rect 1296 379 1312 413
rect 1346 529 1384 565
rect 1346 495 1348 529
rect 1382 495 1384 529
rect 1346 459 1384 495
rect 1346 425 1348 459
rect 1382 425 1384 459
rect 1346 409 1384 425
rect 1418 607 1484 649
rect 1418 573 1434 607
rect 1468 573 1484 607
rect 1418 529 1484 573
rect 1418 495 1434 529
rect 1468 495 1484 529
rect 1418 455 1484 495
rect 1418 421 1434 455
rect 1468 421 1484 455
rect 1258 375 1312 379
rect 1162 307 1224 352
rect 1258 341 1507 375
rect 791 305 1025 307
rect 677 271 693 305
rect 727 271 743 305
rect 791 271 807 305
rect 841 271 875 305
rect 909 271 943 305
rect 977 271 1025 305
rect 677 269 743 271
rect 799 242 1025 271
rect 1061 305 1331 307
rect 1061 271 1077 305
rect 1111 271 1145 305
rect 1179 271 1213 305
rect 1247 271 1281 305
rect 1315 271 1331 305
rect 1061 269 1331 271
rect 1386 287 1439 303
rect 977 235 1025 242
rect 1386 253 1403 287
rect 1437 253 1439 287
rect 1386 235 1439 253
rect 25 203 763 235
rect 25 169 41 203
rect 75 201 213 203
rect 75 169 77 201
rect 25 101 77 169
rect 211 169 213 201
rect 247 201 385 203
rect 247 169 249 201
rect 25 67 41 101
rect 75 67 77 101
rect 25 51 77 67
rect 111 131 127 165
rect 161 131 177 165
rect 111 93 177 131
rect 111 59 127 93
rect 161 59 177 93
rect 111 17 177 59
rect 211 101 249 169
rect 383 169 385 201
rect 419 201 557 203
rect 419 169 421 201
rect 211 67 213 101
rect 247 67 249 101
rect 211 51 249 67
rect 283 131 299 165
rect 333 131 349 165
rect 283 93 349 131
rect 283 59 299 93
rect 333 59 349 93
rect 283 17 349 59
rect 383 101 421 169
rect 555 169 557 201
rect 591 201 729 203
rect 591 169 593 201
rect 383 67 385 101
rect 419 67 421 101
rect 383 51 421 67
rect 455 131 471 165
rect 505 131 521 165
rect 455 93 521 131
rect 455 59 471 93
rect 505 59 521 93
rect 455 17 521 59
rect 555 101 593 169
rect 727 169 729 201
rect 555 67 557 101
rect 591 67 593 101
rect 555 51 593 67
rect 627 131 643 165
rect 677 131 693 165
rect 627 93 693 131
rect 627 59 643 93
rect 677 59 693 93
rect 627 17 693 59
rect 727 101 763 169
rect 797 169 943 208
rect 977 201 1439 235
rect 797 135 826 169
rect 860 167 943 169
rect 1473 167 1507 341
rect 860 165 1507 167
rect 860 135 998 165
rect 797 131 998 135
rect 1032 131 1170 165
rect 1204 131 1342 165
rect 1376 131 1507 165
rect 797 129 1507 131
rect 727 67 729 101
rect 763 91 1478 95
rect 763 67 912 91
rect 727 57 912 67
rect 946 57 1084 91
rect 1118 57 1256 91
rect 1290 57 1428 91
rect 1462 57 1478 91
rect 727 51 1478 57
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o22ai_4
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1205024
string GDS_START 1192062
<< end >>
