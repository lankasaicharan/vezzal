magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
rect 1606 285 1814 331
<< pwell >>
rect 291 184 742 229
rect 15 157 742 184
rect 983 157 1616 201
rect 15 49 1616 157
rect 1806 49 2096 241
rect 0 0 2112 49
<< scnmos >>
rect 94 74 124 158
rect 180 74 210 158
rect 370 119 400 203
rect 456 119 486 203
rect 542 119 572 203
rect 614 119 644 203
rect 823 47 853 131
rect 895 47 925 131
rect 1080 47 1110 175
rect 1152 47 1182 175
rect 1257 91 1287 175
rect 1329 91 1359 175
rect 1401 91 1431 175
rect 1503 91 1533 175
rect 1885 131 1915 215
rect 1987 47 2017 215
<< scpmoshvt >>
rect 86 463 116 591
rect 172 463 202 591
rect 380 463 410 547
rect 466 463 496 547
rect 552 463 582 547
rect 624 463 654 547
rect 732 463 762 547
rect 818 463 848 547
rect 955 379 985 547
rect 1145 417 1175 501
rect 1250 417 1280 585
rect 1465 463 1495 547
rect 1551 463 1581 547
rect 1695 321 1725 405
rect 1885 367 1915 495
rect 2002 367 2032 619
<< ndiff >>
rect 317 178 370 203
rect 41 128 94 158
rect 41 94 49 128
rect 83 94 94 128
rect 41 74 94 94
rect 124 118 180 158
rect 124 84 135 118
rect 169 84 180 118
rect 124 74 180 84
rect 210 132 263 158
rect 210 98 221 132
rect 255 98 263 132
rect 317 144 325 178
rect 359 144 370 178
rect 317 119 370 144
rect 400 178 456 203
rect 400 144 411 178
rect 445 144 456 178
rect 400 119 456 144
rect 486 179 542 203
rect 486 145 497 179
rect 531 145 542 179
rect 486 119 542 145
rect 572 119 614 203
rect 644 151 716 203
rect 644 119 674 151
rect 210 74 263 98
rect 666 117 674 119
rect 708 117 716 151
rect 1009 161 1080 175
rect 1009 131 1035 161
rect 666 105 716 117
rect 770 106 823 131
rect 770 72 778 106
rect 812 72 823 106
rect 770 47 823 72
rect 853 47 895 131
rect 925 127 1035 131
rect 1069 127 1080 161
rect 925 106 1080 127
rect 925 72 936 106
rect 970 93 1080 106
rect 970 72 1035 93
rect 925 59 1035 72
rect 1069 59 1080 93
rect 925 47 1080 59
rect 1110 47 1152 175
rect 1182 163 1257 175
rect 1182 129 1204 163
rect 1238 129 1257 163
rect 1182 95 1257 129
rect 1182 61 1193 95
rect 1227 91 1257 95
rect 1287 91 1329 175
rect 1359 91 1401 175
rect 1431 142 1503 175
rect 1431 108 1442 142
rect 1476 108 1503 142
rect 1431 91 1503 108
rect 1533 143 1590 175
rect 1533 109 1548 143
rect 1582 109 1590 143
rect 1533 91 1590 109
rect 1227 61 1235 91
rect 1832 190 1885 215
rect 1832 156 1840 190
rect 1874 156 1885 190
rect 1832 131 1885 156
rect 1915 203 1987 215
rect 1915 169 1930 203
rect 1964 169 1987 203
rect 1915 131 1987 169
rect 1182 47 1235 61
rect 1934 94 1987 131
rect 1934 60 1942 94
rect 1976 60 1987 94
rect 1934 47 1987 60
rect 2017 203 2070 215
rect 2017 169 2028 203
rect 2062 169 2070 203
rect 2017 101 2070 169
rect 2017 67 2028 101
rect 2062 67 2070 101
rect 2017 47 2070 67
<< pdiff >>
rect 33 577 86 591
rect 33 543 41 577
rect 75 543 86 577
rect 33 509 86 543
rect 33 475 41 509
rect 75 475 86 509
rect 33 463 86 475
rect 116 579 172 591
rect 116 545 127 579
rect 161 545 172 579
rect 116 511 172 545
rect 116 477 127 511
rect 161 477 172 511
rect 116 463 172 477
rect 202 577 255 591
rect 202 543 213 577
rect 247 543 255 577
rect 1302 603 1352 615
rect 1302 585 1310 603
rect 202 509 255 543
rect 202 475 213 509
rect 247 475 255 509
rect 202 463 255 475
rect 327 522 380 547
rect 327 488 335 522
rect 369 488 380 522
rect 327 463 380 488
rect 410 522 466 547
rect 410 488 421 522
rect 455 488 466 522
rect 410 463 466 488
rect 496 521 552 547
rect 496 487 507 521
rect 541 487 552 521
rect 496 463 552 487
rect 582 463 624 547
rect 654 522 732 547
rect 654 488 675 522
rect 709 488 732 522
rect 654 463 732 488
rect 762 522 818 547
rect 762 488 773 522
rect 807 488 818 522
rect 762 463 818 488
rect 848 535 955 547
rect 848 501 859 535
rect 893 501 955 535
rect 848 471 955 501
rect 848 463 910 471
rect 902 437 910 463
rect 944 437 955 471
rect 902 379 955 437
rect 985 535 1038 547
rect 985 501 996 535
rect 1030 501 1038 535
rect 1197 501 1250 585
rect 985 461 1038 501
rect 985 427 996 461
rect 1030 427 1038 461
rect 985 379 1038 427
rect 1092 475 1145 501
rect 1092 441 1100 475
rect 1134 441 1145 475
rect 1092 417 1145 441
rect 1175 463 1250 501
rect 1175 429 1200 463
rect 1234 429 1250 463
rect 1175 417 1250 429
rect 1280 569 1310 585
rect 1344 569 1352 603
rect 1280 417 1352 569
rect 1412 529 1465 547
rect 1412 495 1420 529
rect 1454 495 1465 529
rect 1412 463 1465 495
rect 1495 537 1551 547
rect 1495 503 1506 537
rect 1540 503 1551 537
rect 1495 463 1551 503
rect 1581 522 1634 547
rect 1581 488 1592 522
rect 1626 488 1634 522
rect 1581 463 1634 488
rect 1949 607 2002 619
rect 1949 573 1957 607
rect 1991 573 2002 607
rect 1949 514 2002 573
rect 1949 495 1957 514
rect 1832 481 1885 495
rect 1832 447 1840 481
rect 1874 447 1885 481
rect 1832 413 1885 447
rect 1642 369 1695 405
rect 1642 335 1650 369
rect 1684 335 1695 369
rect 1642 321 1695 335
rect 1725 367 1778 405
rect 1832 379 1840 413
rect 1874 379 1885 413
rect 1832 367 1885 379
rect 1915 480 1957 495
rect 1991 480 2002 514
rect 1915 421 2002 480
rect 1915 387 1938 421
rect 1972 387 2002 421
rect 1915 367 2002 387
rect 2032 599 2085 619
rect 2032 565 2043 599
rect 2077 565 2085 599
rect 2032 502 2085 565
rect 2032 468 2043 502
rect 2077 468 2085 502
rect 2032 420 2085 468
rect 2032 386 2043 420
rect 2077 386 2085 420
rect 2032 367 2085 386
rect 1725 333 1736 367
rect 1770 333 1778 367
rect 1725 321 1778 333
<< ndiffc >>
rect 49 94 83 128
rect 135 84 169 118
rect 221 98 255 132
rect 325 144 359 178
rect 411 144 445 178
rect 497 145 531 179
rect 674 117 708 151
rect 778 72 812 106
rect 1035 127 1069 161
rect 936 72 970 106
rect 1035 59 1069 93
rect 1204 129 1238 163
rect 1193 61 1227 95
rect 1442 108 1476 142
rect 1548 109 1582 143
rect 1840 156 1874 190
rect 1930 169 1964 203
rect 1942 60 1976 94
rect 2028 169 2062 203
rect 2028 67 2062 101
<< pdiffc >>
rect 41 543 75 577
rect 41 475 75 509
rect 127 545 161 579
rect 127 477 161 511
rect 213 543 247 577
rect 213 475 247 509
rect 335 488 369 522
rect 421 488 455 522
rect 507 487 541 521
rect 675 488 709 522
rect 773 488 807 522
rect 859 501 893 535
rect 910 437 944 471
rect 996 501 1030 535
rect 996 427 1030 461
rect 1100 441 1134 475
rect 1200 429 1234 463
rect 1310 569 1344 603
rect 1420 495 1454 529
rect 1506 503 1540 537
rect 1592 488 1626 522
rect 1957 573 1991 607
rect 1840 447 1874 481
rect 1650 335 1684 369
rect 1840 379 1874 413
rect 1957 480 1991 514
rect 1938 387 1972 421
rect 2043 565 2077 599
rect 2043 468 2077 502
rect 2043 386 2077 420
rect 1736 333 1770 367
<< poly >>
rect 86 591 116 617
rect 172 615 1280 645
rect 1367 615 1782 645
rect 2002 619 2032 645
rect 172 591 202 615
rect 380 547 410 573
rect 466 547 496 573
rect 552 547 582 615
rect 1250 585 1280 615
rect 624 547 654 573
rect 732 547 762 573
rect 818 547 848 573
rect 955 547 985 573
rect 86 440 116 463
rect 29 410 116 440
rect 29 248 59 410
rect 172 362 202 463
rect 380 441 410 463
rect 107 346 202 362
rect 107 312 123 346
rect 157 326 202 346
rect 287 415 410 441
rect 287 381 303 415
rect 337 411 410 415
rect 337 381 353 411
rect 157 312 210 326
rect 107 296 210 312
rect 29 232 138 248
rect 29 198 88 232
rect 122 198 138 232
rect 29 182 138 198
rect 94 158 124 182
rect 180 158 210 296
rect 287 255 353 381
rect 466 369 496 463
rect 552 437 582 463
rect 395 353 496 369
rect 395 319 411 353
rect 445 333 496 353
rect 624 431 654 463
rect 624 415 690 431
rect 624 381 640 415
rect 674 381 690 415
rect 624 365 690 381
rect 445 319 572 333
rect 395 303 572 319
rect 287 225 400 255
rect 370 203 400 225
rect 456 203 486 229
rect 542 203 572 303
rect 624 291 654 365
rect 732 323 762 463
rect 818 431 848 463
rect 804 415 870 431
rect 804 381 820 415
rect 854 381 870 415
rect 804 365 870 381
rect 1145 501 1175 527
rect 732 307 798 323
rect 614 275 687 291
rect 614 241 637 275
rect 671 241 687 275
rect 732 273 748 307
rect 782 297 798 307
rect 955 297 985 379
rect 1145 335 1175 417
rect 1250 395 1280 417
rect 1367 402 1397 615
rect 1465 547 1495 615
rect 1716 597 1782 615
rect 1551 547 1581 573
rect 1716 563 1732 597
rect 1766 563 1782 597
rect 1716 529 1782 563
rect 1716 495 1732 529
rect 1766 495 1782 529
rect 1885 495 1915 521
rect 1716 479 1782 495
rect 1465 437 1495 463
rect 1250 365 1287 395
rect 1075 319 1175 335
rect 782 273 1033 297
rect 732 267 1033 273
rect 1075 285 1091 319
rect 1125 299 1175 319
rect 1125 285 1182 299
rect 1075 269 1182 285
rect 732 257 853 267
rect 614 225 687 241
rect 614 203 644 225
rect 370 93 400 119
rect 94 48 124 74
rect 180 51 210 74
rect 456 51 486 119
rect 542 93 572 119
rect 614 93 644 119
rect 823 131 853 257
rect 1003 227 1033 267
rect 895 203 961 219
rect 895 169 911 203
rect 945 169 961 203
rect 1003 197 1110 227
rect 1080 175 1110 197
rect 1152 175 1182 269
rect 1257 175 1287 365
rect 1329 372 1397 402
rect 1551 383 1581 463
rect 1695 405 1725 431
rect 1329 175 1359 372
rect 1455 367 1581 383
rect 1455 333 1471 367
rect 1505 333 1581 367
rect 1455 299 1581 333
rect 1455 279 1471 299
rect 1401 265 1471 279
rect 1505 265 1581 299
rect 1695 267 1725 321
rect 1885 267 1915 367
rect 2002 329 2032 367
rect 1401 249 1581 265
rect 1629 251 1915 267
rect 1957 313 2032 329
rect 1957 279 1973 313
rect 2007 279 2032 313
rect 1957 263 2032 279
rect 1401 175 1431 249
rect 1629 217 1645 251
rect 1679 237 1915 251
rect 1679 217 1695 237
rect 1503 175 1533 201
rect 1629 183 1695 217
rect 1885 215 1915 237
rect 1987 215 2017 263
rect 895 153 961 169
rect 895 131 925 153
rect 180 21 486 51
rect 1629 149 1645 183
rect 1679 149 1695 183
rect 1257 65 1287 91
rect 1329 65 1359 91
rect 1401 65 1431 91
rect 1503 69 1533 91
rect 1629 69 1695 149
rect 1885 105 1915 131
rect 823 21 853 47
rect 895 21 925 47
rect 1080 21 1110 47
rect 1152 21 1182 47
rect 1503 39 1695 69
rect 1987 21 2017 47
<< polycont >>
rect 123 312 157 346
rect 303 381 337 415
rect 88 198 122 232
rect 411 319 445 353
rect 640 381 674 415
rect 820 381 854 415
rect 637 241 671 275
rect 748 273 782 307
rect 1732 563 1766 597
rect 1732 495 1766 529
rect 1091 285 1125 319
rect 911 169 945 203
rect 1471 333 1505 367
rect 1471 265 1505 299
rect 1973 279 2007 313
rect 1645 217 1679 251
rect 1645 149 1679 183
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 18 577 79 593
rect 18 543 41 577
rect 75 543 79 577
rect 18 509 79 543
rect 18 475 41 509
rect 75 475 79 509
rect 18 362 79 475
rect 113 579 175 649
rect 113 545 127 579
rect 161 545 175 579
rect 113 511 175 545
rect 113 477 127 511
rect 161 477 175 511
rect 113 461 175 477
rect 209 577 251 593
rect 209 543 213 577
rect 247 543 251 577
rect 209 509 251 543
rect 209 475 213 509
rect 247 475 251 509
rect 18 346 173 362
rect 18 312 123 346
rect 157 312 173 346
rect 209 337 251 475
rect 319 522 379 649
rect 319 488 335 522
rect 369 488 379 522
rect 319 472 379 488
rect 413 522 457 538
rect 413 488 421 522
rect 455 488 457 522
rect 287 415 367 438
rect 287 381 303 415
rect 337 381 367 415
rect 413 437 457 488
rect 491 521 585 537
rect 491 487 507 521
rect 541 487 585 521
rect 491 471 585 487
rect 659 522 716 649
rect 659 488 675 522
rect 709 488 716 522
rect 659 472 716 488
rect 750 522 823 538
rect 750 488 773 522
rect 807 488 823 522
rect 750 472 823 488
rect 857 535 946 649
rect 857 501 859 535
rect 893 501 946 535
rect 413 403 515 437
rect 287 371 367 381
rect 401 353 447 369
rect 401 337 411 353
rect 209 319 411 337
rect 445 319 447 353
rect 18 134 52 312
rect 209 303 447 319
rect 88 232 175 278
rect 122 198 175 232
rect 88 168 175 198
rect 209 276 271 303
rect 209 242 223 276
rect 257 242 271 276
rect 481 269 515 403
rect 18 128 99 134
rect 18 94 49 128
rect 83 94 99 128
rect 18 78 99 94
rect 133 118 173 134
rect 133 84 135 118
rect 169 84 173 118
rect 133 17 173 84
rect 209 132 271 242
rect 403 235 515 269
rect 551 345 585 471
rect 750 431 784 472
rect 857 471 946 501
rect 894 437 910 471
rect 944 437 946 471
rect 624 415 784 431
rect 624 381 640 415
rect 674 381 784 415
rect 624 379 784 381
rect 818 415 860 431
rect 894 421 946 437
rect 980 603 1360 615
rect 980 569 1310 603
rect 1344 569 1360 603
rect 980 567 1360 569
rect 980 535 1046 567
rect 980 501 996 535
rect 1030 501 1046 535
rect 1506 537 1540 649
rect 980 461 1046 501
rect 980 427 996 461
rect 1030 427 1046 461
rect 980 421 1046 427
rect 1084 529 1470 533
rect 1084 499 1420 529
rect 1084 475 1150 499
rect 1404 495 1420 499
rect 1454 495 1470 529
rect 1404 487 1470 495
rect 1506 487 1540 503
rect 1576 522 1628 538
rect 1576 488 1592 522
rect 1626 488 1628 522
rect 1084 441 1100 475
rect 1134 441 1150 475
rect 1084 425 1150 441
rect 1184 463 1281 465
rect 1184 429 1200 463
rect 1234 453 1281 463
rect 1576 453 1628 488
rect 1234 429 1628 453
rect 1184 421 1628 429
rect 1247 419 1628 421
rect 818 381 820 415
rect 854 387 860 415
rect 854 383 1211 387
rect 854 381 1521 383
rect 818 367 1521 381
rect 818 353 1471 367
rect 551 311 784 345
rect 209 98 221 132
rect 255 98 271 132
rect 209 82 271 98
rect 309 178 369 194
rect 309 144 325 178
rect 359 144 369 178
rect 309 17 369 144
rect 403 178 447 235
rect 551 195 585 311
rect 732 307 784 311
rect 403 144 411 178
rect 445 144 447 178
rect 403 128 447 144
rect 481 179 585 195
rect 621 275 687 277
rect 621 241 637 275
rect 671 241 687 275
rect 732 273 748 307
rect 782 273 784 307
rect 732 257 784 273
rect 621 221 687 241
rect 621 187 816 221
rect 481 145 497 179
rect 531 145 585 179
rect 481 129 585 145
rect 658 151 724 153
rect 658 117 674 151
rect 708 117 724 151
rect 658 17 724 117
rect 762 106 816 187
rect 854 219 888 353
rect 1177 333 1471 353
rect 1505 333 1521 367
rect 1075 285 1091 319
rect 1125 285 1141 319
rect 1075 276 1141 285
rect 1121 242 1141 276
rect 1177 299 1521 333
rect 1177 265 1471 299
rect 1505 265 1521 299
rect 1177 249 1521 265
rect 1555 267 1610 419
rect 1662 385 1696 649
rect 1646 369 1696 385
rect 1646 335 1650 369
rect 1684 335 1696 369
rect 1646 317 1696 335
rect 1730 597 1786 613
rect 1730 563 1732 597
rect 1766 563 1786 597
rect 1730 529 1786 563
rect 1730 495 1732 529
rect 1766 495 1786 529
rect 1912 607 2007 649
rect 1912 573 1957 607
rect 1991 573 2007 607
rect 1912 514 2007 573
rect 1730 367 1786 495
rect 1730 333 1736 367
rect 1770 333 1786 367
rect 1555 251 1695 267
rect 854 203 961 219
rect 1555 217 1645 251
rect 1679 217 1695 251
rect 1555 215 1695 217
rect 854 169 911 203
rect 945 169 961 203
rect 1177 183 1695 215
rect 1177 181 1645 183
rect 1013 161 1085 177
rect 1013 127 1035 161
rect 1069 127 1085 161
rect 1013 122 1085 127
rect 762 72 778 106
rect 812 72 816 106
rect 762 56 816 72
rect 920 106 1085 122
rect 920 72 936 106
rect 970 93 1085 106
rect 970 72 1035 93
rect 920 59 1035 72
rect 1069 59 1085 93
rect 920 17 1085 59
rect 1177 163 1261 181
rect 1177 129 1204 163
rect 1238 129 1261 163
rect 1632 149 1645 181
rect 1679 149 1695 183
rect 1177 95 1261 129
rect 1177 61 1193 95
rect 1227 61 1261 95
rect 1177 57 1261 61
rect 1426 142 1492 147
rect 1426 108 1442 142
rect 1476 108 1492 142
rect 1426 17 1492 108
rect 1532 143 1598 147
rect 1532 109 1548 143
rect 1582 109 1598 143
rect 1632 133 1695 149
rect 1532 97 1598 109
rect 1730 97 1786 333
rect 1824 481 1878 497
rect 1824 447 1840 481
rect 1874 447 1878 481
rect 1824 413 1878 447
rect 1824 379 1840 413
rect 1874 379 1878 413
rect 1824 329 1878 379
rect 1912 480 1957 514
rect 1991 480 2007 514
rect 1912 421 2007 480
rect 1912 387 1938 421
rect 1972 387 2007 421
rect 1912 365 2007 387
rect 2041 599 2095 615
rect 2041 565 2043 599
rect 2077 565 2095 599
rect 2041 502 2095 565
rect 2041 468 2043 502
rect 2077 468 2095 502
rect 2041 420 2095 468
rect 2041 386 2043 420
rect 2077 386 2095 420
rect 1824 313 2007 329
rect 1824 279 1973 313
rect 1824 263 2007 279
rect 1824 190 1878 263
rect 2041 219 2095 386
rect 1824 156 1840 190
rect 1874 156 1878 190
rect 1824 140 1878 156
rect 1914 203 1985 219
rect 1914 169 1930 203
rect 1964 169 1985 203
rect 1532 63 1786 97
rect 1914 94 1985 169
rect 1914 60 1942 94
rect 1976 60 1985 94
rect 1914 17 1985 60
rect 2019 203 2095 219
rect 2019 169 2028 203
rect 2062 169 2095 203
rect 2019 101 2095 169
rect 2019 67 2028 101
rect 2062 67 2095 101
rect 2019 51 2095 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 223 242 257 276
rect 1087 242 1121 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 211 276 269 282
rect 211 242 223 276
rect 257 273 269 276
rect 1075 276 1133 282
rect 1075 273 1087 276
rect 257 245 1087 273
rect 257 242 269 245
rect 211 236 269 242
rect 1075 242 1087 245
rect 1121 242 1133 276
rect 1075 236 1133 242
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfstp_1
flabel comment s 636 331 636 331 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 464 2081 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 538 2081 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 89728
string GDS_START 73662
<< end >>
