magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 60 49 1628 241
rect 0 0 1632 49
<< scnmos >>
rect 139 47 169 215
rect 225 47 255 215
rect 311 47 341 215
rect 397 47 427 215
rect 573 47 603 215
rect 659 47 689 215
rect 745 47 775 215
rect 831 47 861 215
rect 917 47 947 215
rect 1003 47 1033 215
rect 1089 47 1119 215
rect 1175 47 1205 215
rect 1261 47 1291 215
rect 1347 47 1377 215
rect 1433 47 1463 215
rect 1519 47 1549 215
<< scpmoshvt >>
rect 125 367 155 619
rect 211 367 241 619
rect 297 367 327 619
rect 383 367 413 619
rect 469 367 499 619
rect 555 367 585 619
rect 641 367 671 619
rect 727 367 757 619
rect 917 367 947 619
rect 1003 367 1033 619
rect 1089 367 1119 619
rect 1175 367 1205 619
rect 1261 367 1291 619
rect 1347 367 1377 619
rect 1433 367 1463 619
rect 1519 367 1549 619
<< ndiff >>
rect 86 203 139 215
rect 86 169 94 203
rect 128 169 139 203
rect 86 93 139 169
rect 86 59 94 93
rect 128 59 139 93
rect 86 47 139 59
rect 169 203 225 215
rect 169 169 180 203
rect 214 169 225 203
rect 169 101 225 169
rect 169 67 180 101
rect 214 67 225 101
rect 169 47 225 67
rect 255 164 311 215
rect 255 130 266 164
rect 300 130 311 164
rect 255 93 311 130
rect 255 59 266 93
rect 300 59 311 93
rect 255 47 311 59
rect 341 203 397 215
rect 341 169 352 203
rect 386 169 397 203
rect 341 101 397 169
rect 341 67 352 101
rect 386 67 397 101
rect 341 47 397 67
rect 427 124 573 215
rect 427 90 438 124
rect 472 90 528 124
rect 562 90 573 124
rect 427 47 573 90
rect 603 171 659 215
rect 603 137 614 171
rect 648 137 659 171
rect 603 103 659 137
rect 603 69 614 103
rect 648 69 659 103
rect 603 47 659 69
rect 689 124 745 215
rect 689 90 700 124
rect 734 90 745 124
rect 689 47 745 90
rect 775 171 831 215
rect 775 137 786 171
rect 820 137 831 171
rect 775 103 831 137
rect 775 69 786 103
rect 820 69 831 103
rect 775 47 831 69
rect 861 124 917 215
rect 861 90 872 124
rect 906 90 917 124
rect 861 47 917 90
rect 947 171 1003 215
rect 947 137 958 171
rect 992 137 1003 171
rect 947 103 1003 137
rect 947 69 958 103
rect 992 69 1003 103
rect 947 47 1003 69
rect 1033 124 1089 215
rect 1033 90 1044 124
rect 1078 90 1089 124
rect 1033 47 1089 90
rect 1119 171 1175 215
rect 1119 137 1130 171
rect 1164 137 1175 171
rect 1119 103 1175 137
rect 1119 69 1130 103
rect 1164 69 1175 103
rect 1119 47 1175 69
rect 1205 124 1261 215
rect 1205 90 1216 124
rect 1250 90 1261 124
rect 1205 47 1261 90
rect 1291 183 1347 215
rect 1291 149 1302 183
rect 1336 149 1347 183
rect 1291 103 1347 149
rect 1291 69 1302 103
rect 1336 69 1347 103
rect 1291 47 1347 69
rect 1377 124 1433 215
rect 1377 90 1388 124
rect 1422 90 1433 124
rect 1377 47 1433 90
rect 1463 203 1519 215
rect 1463 169 1474 203
rect 1508 169 1519 203
rect 1463 101 1519 169
rect 1463 67 1474 101
rect 1508 67 1519 101
rect 1463 47 1519 67
rect 1549 167 1602 215
rect 1549 133 1560 167
rect 1594 133 1602 167
rect 1549 93 1602 133
rect 1549 59 1560 93
rect 1594 59 1602 93
rect 1549 47 1602 59
<< pdiff >>
rect 72 597 125 619
rect 72 563 80 597
rect 114 563 125 597
rect 72 515 125 563
rect 72 481 80 515
rect 114 481 125 515
rect 72 434 125 481
rect 72 400 80 434
rect 114 400 125 434
rect 72 367 125 400
rect 155 607 211 619
rect 155 573 166 607
rect 200 573 211 607
rect 155 502 211 573
rect 155 468 166 502
rect 200 468 211 502
rect 155 367 211 468
rect 241 597 297 619
rect 241 563 252 597
rect 286 563 297 597
rect 241 515 297 563
rect 241 481 252 515
rect 286 481 297 515
rect 241 434 297 481
rect 241 400 252 434
rect 286 400 297 434
rect 241 367 297 400
rect 327 607 383 619
rect 327 573 338 607
rect 372 573 383 607
rect 327 493 383 573
rect 327 459 338 493
rect 372 459 383 493
rect 327 367 383 459
rect 413 597 469 619
rect 413 563 424 597
rect 458 563 469 597
rect 413 515 469 563
rect 413 481 424 515
rect 458 481 469 515
rect 413 434 469 481
rect 413 400 424 434
rect 458 400 469 434
rect 413 367 469 400
rect 499 529 555 619
rect 499 495 510 529
rect 544 495 555 529
rect 499 413 555 495
rect 499 379 510 413
rect 544 379 555 413
rect 499 367 555 379
rect 585 597 641 619
rect 585 563 596 597
rect 630 563 641 597
rect 585 529 641 563
rect 585 495 596 529
rect 630 495 641 529
rect 585 461 641 495
rect 585 427 596 461
rect 630 427 641 461
rect 585 367 641 427
rect 671 529 727 619
rect 671 495 682 529
rect 716 495 727 529
rect 671 413 727 495
rect 671 379 682 413
rect 716 379 727 413
rect 671 367 727 379
rect 757 597 810 619
rect 757 563 768 597
rect 802 563 810 597
rect 757 529 810 563
rect 757 495 768 529
rect 802 495 810 529
rect 757 461 810 495
rect 757 427 768 461
rect 802 427 810 461
rect 757 367 810 427
rect 864 599 917 619
rect 864 565 872 599
rect 906 565 917 599
rect 864 520 917 565
rect 864 486 872 520
rect 906 486 917 520
rect 864 445 917 486
rect 864 411 872 445
rect 906 411 917 445
rect 864 367 917 411
rect 947 531 1003 619
rect 947 497 958 531
rect 992 497 1003 531
rect 947 413 1003 497
rect 947 379 958 413
rect 992 379 1003 413
rect 947 367 1003 379
rect 1033 599 1089 619
rect 1033 565 1044 599
rect 1078 565 1089 599
rect 1033 520 1089 565
rect 1033 486 1044 520
rect 1078 486 1089 520
rect 1033 445 1089 486
rect 1033 411 1044 445
rect 1078 411 1089 445
rect 1033 367 1089 411
rect 1119 531 1175 619
rect 1119 497 1130 531
rect 1164 497 1175 531
rect 1119 413 1175 497
rect 1119 379 1130 413
rect 1164 379 1175 413
rect 1119 367 1175 379
rect 1205 599 1261 619
rect 1205 565 1216 599
rect 1250 565 1261 599
rect 1205 520 1261 565
rect 1205 486 1216 520
rect 1250 486 1261 520
rect 1205 445 1261 486
rect 1205 411 1216 445
rect 1250 411 1261 445
rect 1205 367 1261 411
rect 1291 531 1347 619
rect 1291 497 1302 531
rect 1336 497 1347 531
rect 1291 413 1347 497
rect 1291 379 1302 413
rect 1336 379 1347 413
rect 1291 367 1347 379
rect 1377 599 1433 619
rect 1377 565 1388 599
rect 1422 565 1433 599
rect 1377 520 1433 565
rect 1377 486 1388 520
rect 1422 486 1433 520
rect 1377 445 1433 486
rect 1377 411 1388 445
rect 1422 411 1433 445
rect 1377 367 1433 411
rect 1463 531 1519 619
rect 1463 497 1474 531
rect 1508 497 1519 531
rect 1463 413 1519 497
rect 1463 379 1474 413
rect 1508 379 1519 413
rect 1463 367 1519 379
rect 1549 599 1602 619
rect 1549 565 1560 599
rect 1594 565 1602 599
rect 1549 520 1602 565
rect 1549 486 1560 520
rect 1594 486 1602 520
rect 1549 445 1602 486
rect 1549 411 1560 445
rect 1594 411 1602 445
rect 1549 367 1602 411
<< ndiffc >>
rect 94 169 128 203
rect 94 59 128 93
rect 180 169 214 203
rect 180 67 214 101
rect 266 130 300 164
rect 266 59 300 93
rect 352 169 386 203
rect 352 67 386 101
rect 438 90 472 124
rect 528 90 562 124
rect 614 137 648 171
rect 614 69 648 103
rect 700 90 734 124
rect 786 137 820 171
rect 786 69 820 103
rect 872 90 906 124
rect 958 137 992 171
rect 958 69 992 103
rect 1044 90 1078 124
rect 1130 137 1164 171
rect 1130 69 1164 103
rect 1216 90 1250 124
rect 1302 149 1336 183
rect 1302 69 1336 103
rect 1388 90 1422 124
rect 1474 169 1508 203
rect 1474 67 1508 101
rect 1560 133 1594 167
rect 1560 59 1594 93
<< pdiffc >>
rect 80 563 114 597
rect 80 481 114 515
rect 80 400 114 434
rect 166 573 200 607
rect 166 468 200 502
rect 252 563 286 597
rect 252 481 286 515
rect 252 400 286 434
rect 338 573 372 607
rect 338 459 372 493
rect 424 563 458 597
rect 424 481 458 515
rect 424 400 458 434
rect 510 495 544 529
rect 510 379 544 413
rect 596 563 630 597
rect 596 495 630 529
rect 596 427 630 461
rect 682 495 716 529
rect 682 379 716 413
rect 768 563 802 597
rect 768 495 802 529
rect 768 427 802 461
rect 872 565 906 599
rect 872 486 906 520
rect 872 411 906 445
rect 958 497 992 531
rect 958 379 992 413
rect 1044 565 1078 599
rect 1044 486 1078 520
rect 1044 411 1078 445
rect 1130 497 1164 531
rect 1130 379 1164 413
rect 1216 565 1250 599
rect 1216 486 1250 520
rect 1216 411 1250 445
rect 1302 497 1336 531
rect 1302 379 1336 413
rect 1388 565 1422 599
rect 1388 486 1422 520
rect 1388 411 1422 445
rect 1474 497 1508 531
rect 1474 379 1508 413
rect 1560 565 1594 599
rect 1560 486 1594 520
rect 1560 411 1594 445
<< poly >>
rect 125 619 155 645
rect 211 619 241 645
rect 297 619 327 645
rect 383 619 413 645
rect 469 619 499 645
rect 555 619 585 645
rect 641 619 671 645
rect 727 619 757 645
rect 917 619 947 645
rect 1003 619 1033 645
rect 1089 619 1119 645
rect 1175 619 1205 645
rect 1261 619 1291 645
rect 1347 619 1377 645
rect 1433 619 1463 645
rect 1519 619 1549 645
rect 125 325 155 367
rect 211 325 241 367
rect 297 325 327 367
rect 383 325 413 367
rect 469 345 499 367
rect 555 345 585 367
rect 641 345 671 367
rect 727 345 757 367
rect 21 309 427 325
rect 21 275 37 309
rect 71 275 105 309
rect 139 275 173 309
rect 207 275 241 309
rect 275 275 309 309
rect 343 275 377 309
rect 411 275 427 309
rect 21 237 427 275
rect 469 315 757 345
rect 469 287 875 315
rect 469 253 485 287
rect 519 253 553 287
rect 587 253 621 287
rect 655 253 689 287
rect 723 253 757 287
rect 791 253 825 287
rect 859 253 875 287
rect 469 237 875 253
rect 917 303 947 367
rect 1003 303 1033 367
rect 1089 303 1119 367
rect 1175 303 1205 367
rect 917 287 1205 303
rect 917 253 951 287
rect 985 253 1019 287
rect 1053 253 1087 287
rect 1121 253 1155 287
rect 1189 253 1205 287
rect 917 237 1205 253
rect 139 215 169 237
rect 225 215 255 237
rect 311 215 341 237
rect 397 215 427 237
rect 573 215 603 237
rect 659 215 689 237
rect 745 215 775 237
rect 831 215 861 237
rect 917 215 947 237
rect 1003 215 1033 237
rect 1089 215 1119 237
rect 1175 215 1205 237
rect 1261 321 1291 367
rect 1347 321 1377 367
rect 1433 321 1463 367
rect 1519 321 1549 367
rect 1261 305 1549 321
rect 1261 271 1277 305
rect 1311 271 1345 305
rect 1379 271 1413 305
rect 1447 271 1481 305
rect 1515 271 1549 305
rect 1261 255 1549 271
rect 1261 215 1291 255
rect 1347 215 1377 255
rect 1433 215 1463 255
rect 1519 215 1549 255
rect 139 21 169 47
rect 225 21 255 47
rect 311 21 341 47
rect 397 21 427 47
rect 573 21 603 47
rect 659 21 689 47
rect 745 21 775 47
rect 831 21 861 47
rect 917 21 947 47
rect 1003 21 1033 47
rect 1089 21 1119 47
rect 1175 21 1205 47
rect 1261 21 1291 47
rect 1347 21 1377 47
rect 1433 21 1463 47
rect 1519 21 1549 47
<< polycont >>
rect 37 275 71 309
rect 105 275 139 309
rect 173 275 207 309
rect 241 275 275 309
rect 309 275 343 309
rect 377 275 411 309
rect 485 253 519 287
rect 553 253 587 287
rect 621 253 655 287
rect 689 253 723 287
rect 757 253 791 287
rect 825 253 859 287
rect 951 253 985 287
rect 1019 253 1053 287
rect 1087 253 1121 287
rect 1155 253 1189 287
rect 1277 271 1311 305
rect 1345 271 1379 305
rect 1413 271 1447 305
rect 1481 271 1515 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 64 597 116 613
rect 64 563 80 597
rect 114 563 116 597
rect 64 515 116 563
rect 64 481 80 515
rect 114 481 116 515
rect 64 434 116 481
rect 150 607 216 649
rect 150 573 166 607
rect 200 573 216 607
rect 150 502 216 573
rect 150 468 166 502
rect 200 468 216 502
rect 150 452 216 468
rect 250 597 288 613
rect 250 563 252 597
rect 286 563 288 597
rect 250 515 288 563
rect 250 481 252 515
rect 286 481 288 515
rect 64 400 80 434
rect 114 418 116 434
rect 250 434 288 481
rect 322 607 388 649
rect 322 573 338 607
rect 372 573 388 607
rect 322 493 388 573
rect 322 459 338 493
rect 372 459 388 493
rect 322 452 388 459
rect 422 597 818 613
rect 422 563 424 597
rect 458 579 596 597
rect 458 563 469 579
rect 422 515 469 563
rect 580 563 596 579
rect 630 579 768 597
rect 630 563 646 579
rect 422 481 424 515
rect 458 481 469 515
rect 250 418 252 434
rect 114 400 252 418
rect 286 418 288 434
rect 422 434 469 481
rect 422 418 424 434
rect 286 400 424 418
rect 458 400 469 434
rect 64 384 469 400
rect 503 529 546 545
rect 503 495 510 529
rect 544 495 546 529
rect 503 413 546 495
rect 503 379 510 413
rect 544 379 546 413
rect 580 529 646 563
rect 757 563 768 579
rect 802 563 818 597
rect 580 495 596 529
rect 630 495 646 529
rect 580 461 646 495
rect 580 427 596 461
rect 630 427 646 461
rect 580 411 646 427
rect 680 529 723 545
rect 680 495 682 529
rect 716 495 723 529
rect 680 413 723 495
rect 503 375 546 379
rect 680 379 682 413
rect 716 379 723 413
rect 757 529 818 563
rect 757 495 768 529
rect 802 495 818 529
rect 757 461 818 495
rect 757 427 768 461
rect 802 427 818 461
rect 757 411 818 427
rect 856 599 1610 615
rect 856 565 872 599
rect 906 581 1044 599
rect 906 565 922 581
rect 856 520 922 565
rect 1028 565 1044 581
rect 1078 581 1216 599
rect 1078 565 1094 581
rect 856 486 872 520
rect 906 486 922 520
rect 856 445 922 486
rect 856 411 872 445
rect 906 411 922 445
rect 956 531 994 547
rect 956 497 958 531
rect 992 497 994 531
rect 956 413 994 497
rect 680 375 723 379
rect 956 379 958 413
rect 992 379 994 413
rect 1028 520 1094 565
rect 1200 565 1216 581
rect 1250 581 1388 599
rect 1250 565 1266 581
rect 1028 486 1044 520
rect 1078 486 1094 520
rect 1028 445 1094 486
rect 1028 411 1044 445
rect 1078 411 1094 445
rect 1128 531 1164 547
rect 1128 497 1130 531
rect 1128 413 1164 497
rect 956 375 994 379
rect 1128 379 1130 413
rect 1200 520 1266 565
rect 1372 565 1388 581
rect 1422 581 1560 599
rect 1422 565 1438 581
rect 1200 486 1216 520
rect 1250 486 1266 520
rect 1200 445 1266 486
rect 1200 411 1216 445
rect 1250 411 1266 445
rect 1300 531 1338 547
rect 1300 497 1302 531
rect 1336 497 1338 531
rect 1300 413 1338 497
rect 1128 375 1164 379
rect 21 309 427 350
rect 503 341 1164 375
rect 1300 379 1302 413
rect 1336 379 1338 413
rect 1372 520 1438 565
rect 1544 565 1560 581
rect 1594 565 1610 599
rect 1372 486 1388 520
rect 1422 486 1438 520
rect 1372 445 1438 486
rect 1372 411 1388 445
rect 1422 411 1438 445
rect 1472 531 1510 547
rect 1472 497 1474 531
rect 1508 497 1510 531
rect 1472 413 1510 497
rect 1300 375 1338 379
rect 1472 379 1474 413
rect 1508 379 1510 413
rect 1544 520 1610 565
rect 1544 486 1560 520
rect 1594 486 1610 520
rect 1544 445 1610 486
rect 1544 411 1560 445
rect 1594 411 1610 445
rect 1472 375 1510 379
rect 1300 339 1614 375
rect 21 275 37 309
rect 71 275 105 309
rect 139 275 173 309
rect 207 275 241 309
rect 275 275 309 309
rect 343 275 377 309
rect 411 275 427 309
rect 21 269 427 275
rect 469 287 875 307
rect 469 253 485 287
rect 519 253 553 287
rect 587 253 621 287
rect 655 253 689 287
rect 723 253 757 287
rect 791 253 825 287
rect 859 253 875 287
rect 469 242 875 253
rect 935 287 1217 307
rect 935 253 951 287
rect 985 253 1019 287
rect 1053 253 1087 287
rect 1121 253 1155 287
rect 1189 253 1217 287
rect 935 242 1217 253
rect 1261 271 1277 305
rect 1311 271 1345 305
rect 1379 271 1413 305
rect 1447 271 1481 305
rect 1515 271 1531 305
rect 1261 242 1429 271
rect 1565 237 1614 339
rect 78 203 139 219
rect 78 169 94 203
rect 128 169 139 203
rect 78 93 139 169
rect 78 59 94 93
rect 128 59 139 93
rect 78 17 139 59
rect 173 208 386 235
rect 1463 208 1614 237
rect 173 203 1614 208
rect 173 169 180 203
rect 214 201 352 203
rect 214 169 216 201
rect 173 101 216 169
rect 350 169 352 201
rect 386 183 1474 203
rect 386 174 1302 183
rect 386 169 388 174
rect 173 67 180 101
rect 214 67 216 101
rect 173 51 216 67
rect 250 164 316 167
rect 250 130 266 164
rect 300 130 316 164
rect 250 93 316 130
rect 250 59 266 93
rect 300 59 316 93
rect 250 17 316 59
rect 350 101 388 169
rect 611 171 650 174
rect 350 67 352 101
rect 386 67 388 101
rect 350 51 388 67
rect 422 124 577 140
rect 422 90 438 124
rect 472 90 528 124
rect 562 90 577 124
rect 422 17 577 90
rect 611 137 614 171
rect 648 137 650 171
rect 784 171 822 174
rect 611 103 650 137
rect 611 69 614 103
rect 648 69 650 103
rect 611 53 650 69
rect 684 124 750 140
rect 684 90 700 124
rect 734 90 750 124
rect 684 17 750 90
rect 784 137 786 171
rect 820 137 822 171
rect 956 171 994 174
rect 784 103 822 137
rect 784 69 786 103
rect 820 69 822 103
rect 784 53 822 69
rect 856 124 922 140
rect 856 90 872 124
rect 906 90 922 124
rect 856 17 922 90
rect 956 137 958 171
rect 992 137 994 171
rect 1128 171 1166 174
rect 956 103 994 137
rect 956 69 958 103
rect 992 69 994 103
rect 956 53 994 69
rect 1028 124 1094 140
rect 1028 90 1044 124
rect 1078 90 1094 124
rect 1028 17 1094 90
rect 1128 137 1130 171
rect 1164 137 1166 171
rect 1300 149 1302 174
rect 1336 174 1474 183
rect 1336 149 1338 174
rect 1128 103 1166 137
rect 1128 69 1130 103
rect 1164 69 1166 103
rect 1128 53 1166 69
rect 1200 124 1266 140
rect 1200 90 1216 124
rect 1250 90 1266 124
rect 1200 17 1266 90
rect 1300 103 1338 149
rect 1472 169 1474 174
rect 1508 201 1614 203
rect 1508 169 1510 201
rect 1300 69 1302 103
rect 1336 69 1338 103
rect 1300 53 1338 69
rect 1372 124 1438 140
rect 1372 90 1388 124
rect 1422 90 1438 124
rect 1372 17 1438 90
rect 1472 101 1510 169
rect 1472 67 1474 101
rect 1508 67 1510 101
rect 1472 51 1510 67
rect 1544 133 1560 167
rect 1594 133 1610 167
rect 1544 93 1610 133
rect 1544 59 1560 93
rect 1594 59 1610 93
rect 1544 17 1610 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4173264
string GDS_START 4159276
<< end >>
