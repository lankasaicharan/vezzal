magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2034 1852
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 684 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 173 47 203 177
rect 284 47 314 177
rect 378 47 408 177
rect 472 47 502 177
rect 576 47 606 177
<< scpmoshvt >>
rect 93 297 129 497
rect 175 297 211 497
rect 286 297 322 497
rect 380 297 416 497
rect 474 297 510 497
rect 568 297 604 497
<< ndiff >>
rect 27 99 89 177
rect 27 65 35 99
rect 69 65 89 99
rect 27 47 89 65
rect 119 165 173 177
rect 119 131 129 165
rect 163 131 173 165
rect 119 97 173 131
rect 119 63 129 97
rect 163 63 173 97
rect 119 47 173 63
rect 203 132 284 177
rect 203 98 232 132
rect 266 98 284 132
rect 203 47 284 98
rect 314 165 378 177
rect 314 131 334 165
rect 368 131 378 165
rect 314 97 378 131
rect 314 63 334 97
rect 368 63 378 97
rect 314 47 378 63
rect 408 97 472 177
rect 408 63 428 97
rect 462 63 472 97
rect 408 47 472 63
rect 502 165 576 177
rect 502 131 522 165
rect 556 131 576 165
rect 502 97 576 131
rect 502 63 522 97
rect 556 63 576 97
rect 502 47 576 63
rect 606 97 658 177
rect 606 63 616 97
rect 650 63 658 97
rect 606 47 658 63
<< pdiff >>
rect 35 477 93 497
rect 35 443 47 477
rect 81 443 93 477
rect 35 409 93 443
rect 35 375 47 409
rect 81 375 93 409
rect 35 341 93 375
rect 35 307 47 341
rect 81 307 93 341
rect 35 297 93 307
rect 129 297 175 497
rect 211 487 286 497
rect 211 453 232 487
rect 266 453 286 487
rect 211 419 286 453
rect 211 385 232 419
rect 266 385 286 419
rect 211 297 286 385
rect 322 485 380 497
rect 322 451 334 485
rect 368 451 380 485
rect 322 417 380 451
rect 322 383 334 417
rect 368 383 380 417
rect 322 297 380 383
rect 416 485 474 497
rect 416 451 428 485
rect 462 451 474 485
rect 416 297 474 451
rect 510 485 568 497
rect 510 451 522 485
rect 556 451 568 485
rect 510 417 568 451
rect 510 383 522 417
rect 556 383 568 417
rect 510 349 568 383
rect 510 315 522 349
rect 556 315 568 349
rect 510 297 568 315
rect 604 485 662 497
rect 604 451 616 485
rect 650 451 662 485
rect 604 417 662 451
rect 604 383 616 417
rect 650 383 662 417
rect 604 297 662 383
<< ndiffc >>
rect 35 65 69 99
rect 129 131 163 165
rect 129 63 163 97
rect 232 98 266 132
rect 334 131 368 165
rect 334 63 368 97
rect 428 63 462 97
rect 522 131 556 165
rect 522 63 556 97
rect 616 63 650 97
<< pdiffc >>
rect 47 443 81 477
rect 47 375 81 409
rect 47 307 81 341
rect 232 453 266 487
rect 232 385 266 419
rect 334 451 368 485
rect 334 383 368 417
rect 428 451 462 485
rect 522 451 556 485
rect 522 383 556 417
rect 522 315 556 349
rect 616 451 650 485
rect 616 383 650 417
<< poly >>
rect 93 497 129 523
rect 175 497 211 523
rect 286 497 322 523
rect 380 497 416 523
rect 474 497 510 523
rect 568 497 604 523
rect 93 282 129 297
rect 175 282 211 297
rect 286 282 322 297
rect 380 282 416 297
rect 474 282 510 297
rect 568 282 604 297
rect 91 265 131 282
rect 25 249 131 265
rect 25 215 35 249
rect 69 215 131 249
rect 25 199 131 215
rect 173 265 213 282
rect 284 265 324 282
rect 378 265 418 282
rect 472 265 512 282
rect 566 265 606 282
rect 173 249 237 265
rect 173 215 183 249
rect 217 215 237 249
rect 173 199 237 215
rect 284 249 606 265
rect 284 215 328 249
rect 362 215 396 249
rect 430 215 474 249
rect 508 215 606 249
rect 284 199 606 215
rect 89 177 119 199
rect 173 177 203 199
rect 284 177 314 199
rect 378 177 408 199
rect 472 177 502 199
rect 576 177 606 199
rect 89 21 119 47
rect 173 21 203 47
rect 284 21 314 47
rect 378 21 408 47
rect 472 21 502 47
rect 576 21 606 47
<< polycont >>
rect 35 215 69 249
rect 183 215 217 249
rect 328 215 362 249
rect 396 215 430 249
rect 474 215 508 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 31 477 103 493
rect 31 443 47 477
rect 81 443 103 477
rect 31 409 103 443
rect 31 375 47 409
rect 81 375 103 409
rect 31 341 103 375
rect 232 487 266 527
rect 232 419 266 453
rect 232 367 266 385
rect 318 485 394 493
rect 318 451 334 485
rect 368 451 394 485
rect 318 417 394 451
rect 428 485 462 527
rect 428 435 462 451
rect 506 485 582 493
rect 506 451 522 485
rect 556 451 582 485
rect 318 383 334 417
rect 368 401 394 417
rect 506 417 582 451
rect 506 401 522 417
rect 368 383 522 401
rect 556 383 582 417
rect 318 367 582 383
rect 616 485 650 527
rect 616 417 650 451
rect 616 367 650 383
rect 31 307 47 341
rect 81 333 103 341
rect 506 349 582 367
rect 81 307 353 333
rect 31 299 353 307
rect 506 315 522 349
rect 556 333 582 349
rect 556 315 634 333
rect 506 299 634 315
rect 18 249 69 265
rect 18 215 35 249
rect 18 153 69 215
rect 103 165 149 299
rect 183 249 268 265
rect 217 215 268 249
rect 302 249 353 299
rect 302 215 328 249
rect 362 215 396 249
rect 430 215 474 249
rect 508 215 524 249
rect 183 199 268 215
rect 565 181 634 299
rect 318 165 634 181
rect 103 131 129 165
rect 163 131 179 165
rect 21 99 69 119
rect 21 65 35 99
rect 21 17 69 65
rect 103 97 179 131
rect 103 63 129 97
rect 163 63 179 97
rect 103 58 179 63
rect 232 132 266 165
rect 232 17 266 98
rect 318 131 334 165
rect 368 147 522 165
rect 368 131 394 147
rect 318 97 394 131
rect 506 131 522 147
rect 556 147 634 165
rect 556 131 582 147
rect 318 63 334 97
rect 368 63 394 97
rect 318 53 394 63
rect 428 97 462 113
rect 428 17 462 63
rect 506 97 582 131
rect 506 63 522 97
rect 556 63 582 97
rect 506 53 582 63
rect 616 97 650 113
rect 616 17 650 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 581 289 615 323 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or2_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2605972
string GDS_START 2599918
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
