magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 7 49 1151 251
rect 0 0 1152 49
<< scnmos >>
rect 86 57 116 225
rect 172 57 202 225
rect 258 57 288 225
rect 344 57 374 225
rect 430 57 460 225
rect 516 57 546 225
rect 606 57 636 225
rect 698 57 728 225
rect 784 57 814 225
rect 870 57 900 225
rect 956 57 986 225
rect 1042 57 1072 225
<< scpmoshvt >>
rect 90 367 120 619
rect 176 367 206 619
rect 262 367 292 619
rect 348 367 378 619
rect 434 367 464 619
rect 520 367 550 619
rect 606 367 636 619
rect 692 367 722 619
rect 784 367 814 619
rect 870 367 900 619
rect 956 367 986 619
rect 1042 367 1072 619
<< ndiff >>
rect 33 213 86 225
rect 33 179 41 213
rect 75 179 86 213
rect 33 103 86 179
rect 33 69 41 103
rect 75 69 86 103
rect 33 57 86 69
rect 116 169 172 225
rect 116 135 127 169
rect 161 135 172 169
rect 116 57 172 135
rect 202 177 258 225
rect 202 143 213 177
rect 247 143 258 177
rect 202 103 258 143
rect 202 69 213 103
rect 247 69 258 103
rect 202 57 258 69
rect 288 169 344 225
rect 288 135 299 169
rect 333 135 344 169
rect 288 57 344 135
rect 374 213 430 225
rect 374 179 385 213
rect 419 179 430 213
rect 374 103 430 179
rect 374 69 385 103
rect 419 69 430 103
rect 374 57 430 69
rect 460 183 516 225
rect 460 149 471 183
rect 505 149 516 183
rect 460 103 516 149
rect 460 69 471 103
rect 505 69 516 103
rect 460 57 516 69
rect 546 179 606 225
rect 546 145 561 179
rect 595 145 606 179
rect 546 57 606 145
rect 636 183 698 225
rect 636 149 651 183
rect 685 149 698 183
rect 636 101 698 149
rect 636 67 651 101
rect 685 67 698 101
rect 636 57 698 67
rect 728 99 784 225
rect 728 65 739 99
rect 773 65 784 99
rect 728 57 784 65
rect 814 183 870 225
rect 814 149 825 183
rect 859 149 870 183
rect 814 57 870 149
rect 900 111 956 225
rect 900 77 911 111
rect 945 77 956 111
rect 900 57 956 77
rect 986 183 1042 225
rect 986 149 997 183
rect 1031 149 1042 183
rect 986 57 1042 149
rect 1072 213 1125 225
rect 1072 179 1083 213
rect 1117 179 1125 213
rect 1072 103 1125 179
rect 1072 69 1083 103
rect 1117 69 1125 103
rect 1072 57 1125 69
<< pdiff >>
rect 37 607 90 619
rect 37 573 45 607
rect 79 573 90 607
rect 37 514 90 573
rect 37 480 45 514
rect 79 480 90 514
rect 37 418 90 480
rect 37 384 45 418
rect 79 384 90 418
rect 37 367 90 384
rect 120 599 176 619
rect 120 565 131 599
rect 165 565 176 599
rect 120 519 176 565
rect 120 485 131 519
rect 165 485 176 519
rect 120 434 176 485
rect 120 400 131 434
rect 165 400 176 434
rect 120 367 176 400
rect 206 607 262 619
rect 206 573 217 607
rect 251 573 262 607
rect 206 488 262 573
rect 206 454 217 488
rect 251 454 262 488
rect 206 367 262 454
rect 292 599 348 619
rect 292 565 303 599
rect 337 565 348 599
rect 292 519 348 565
rect 292 485 303 519
rect 337 485 348 519
rect 292 434 348 485
rect 292 400 303 434
rect 337 400 348 434
rect 292 367 348 400
rect 378 611 434 619
rect 378 577 389 611
rect 423 577 434 611
rect 378 534 434 577
rect 378 500 389 534
rect 423 500 434 534
rect 378 457 434 500
rect 378 423 389 457
rect 423 423 434 457
rect 378 367 434 423
rect 464 599 520 619
rect 464 565 475 599
rect 509 565 520 599
rect 464 508 520 565
rect 464 474 475 508
rect 509 474 520 508
rect 464 413 520 474
rect 464 379 475 413
rect 509 379 520 413
rect 464 367 520 379
rect 550 568 606 619
rect 550 534 561 568
rect 595 534 606 568
rect 550 367 606 534
rect 636 599 692 619
rect 636 565 647 599
rect 681 565 692 599
rect 636 508 692 565
rect 636 474 647 508
rect 681 474 692 508
rect 636 367 692 474
rect 722 568 784 619
rect 722 534 733 568
rect 767 534 784 568
rect 722 367 784 534
rect 814 599 870 619
rect 814 565 825 599
rect 859 565 870 599
rect 814 508 870 565
rect 814 474 825 508
rect 859 474 870 508
rect 814 367 870 474
rect 900 568 956 619
rect 900 534 911 568
rect 945 534 956 568
rect 900 367 956 534
rect 986 599 1042 619
rect 986 565 997 599
rect 1031 565 1042 599
rect 986 508 1042 565
rect 986 474 997 508
rect 1031 474 1042 508
rect 986 367 1042 474
rect 1072 607 1125 619
rect 1072 573 1083 607
rect 1117 573 1125 607
rect 1072 492 1125 573
rect 1072 458 1083 492
rect 1117 458 1125 492
rect 1072 367 1125 458
<< ndiffc >>
rect 41 179 75 213
rect 41 69 75 103
rect 127 135 161 169
rect 213 143 247 177
rect 213 69 247 103
rect 299 135 333 169
rect 385 179 419 213
rect 385 69 419 103
rect 471 149 505 183
rect 471 69 505 103
rect 561 145 595 179
rect 651 149 685 183
rect 651 67 685 101
rect 739 65 773 99
rect 825 149 859 183
rect 911 77 945 111
rect 997 149 1031 183
rect 1083 179 1117 213
rect 1083 69 1117 103
<< pdiffc >>
rect 45 573 79 607
rect 45 480 79 514
rect 45 384 79 418
rect 131 565 165 599
rect 131 485 165 519
rect 131 400 165 434
rect 217 573 251 607
rect 217 454 251 488
rect 303 565 337 599
rect 303 485 337 519
rect 303 400 337 434
rect 389 577 423 611
rect 389 500 423 534
rect 389 423 423 457
rect 475 565 509 599
rect 475 474 509 508
rect 475 379 509 413
rect 561 534 595 568
rect 647 565 681 599
rect 647 474 681 508
rect 733 534 767 568
rect 825 565 859 599
rect 825 474 859 508
rect 911 534 945 568
rect 997 565 1031 599
rect 997 474 1031 508
rect 1083 573 1117 607
rect 1083 458 1117 492
<< poly >>
rect 90 619 120 645
rect 176 619 206 645
rect 262 619 292 645
rect 348 619 378 645
rect 434 619 464 645
rect 520 619 550 645
rect 606 619 636 645
rect 692 619 722 645
rect 784 619 814 645
rect 870 619 900 645
rect 956 619 986 645
rect 1042 619 1072 645
rect 90 335 120 367
rect 176 335 206 367
rect 262 335 292 367
rect 348 335 378 367
rect 434 335 464 367
rect 520 335 550 367
rect 606 335 636 367
rect 692 335 722 367
rect 784 335 814 367
rect 870 335 900 367
rect 956 335 986 367
rect 60 319 378 335
rect 60 285 76 319
rect 110 285 144 319
rect 178 285 212 319
rect 246 305 378 319
rect 430 319 636 335
rect 246 285 374 305
rect 60 269 374 285
rect 86 225 116 269
rect 172 225 202 269
rect 258 225 288 269
rect 344 225 374 269
rect 430 285 450 319
rect 484 285 518 319
rect 552 285 586 319
rect 620 285 636 319
rect 430 269 636 285
rect 678 319 986 335
rect 678 285 694 319
rect 728 285 762 319
rect 796 285 830 319
rect 864 285 898 319
rect 932 285 986 319
rect 678 269 986 285
rect 430 225 460 269
rect 516 225 546 269
rect 606 225 636 269
rect 698 225 728 269
rect 784 225 814 269
rect 870 225 900 269
rect 956 225 986 269
rect 1042 335 1072 367
rect 1042 319 1108 335
rect 1042 285 1058 319
rect 1092 285 1108 319
rect 1042 269 1108 285
rect 1042 225 1072 269
rect 86 31 116 57
rect 172 31 202 57
rect 258 31 288 57
rect 344 31 374 57
rect 430 31 460 57
rect 516 31 546 57
rect 606 31 636 57
rect 698 31 728 57
rect 784 31 814 57
rect 870 31 900 57
rect 956 31 986 57
rect 1042 31 1072 57
<< polycont >>
rect 76 285 110 319
rect 144 285 178 319
rect 212 285 246 319
rect 450 285 484 319
rect 518 285 552 319
rect 586 285 620 319
rect 694 285 728 319
rect 762 285 796 319
rect 830 285 864 319
rect 898 285 932 319
rect 1058 285 1092 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 29 607 95 649
rect 29 573 45 607
rect 79 573 95 607
rect 29 514 95 573
rect 29 480 45 514
rect 79 480 95 514
rect 29 418 95 480
rect 29 384 45 418
rect 79 384 95 418
rect 129 599 167 615
rect 129 565 131 599
rect 165 565 167 599
rect 129 519 167 565
rect 129 485 131 519
rect 165 485 167 519
rect 129 434 167 485
rect 201 607 267 649
rect 201 573 217 607
rect 251 573 267 607
rect 201 488 267 573
rect 201 454 217 488
rect 251 454 267 488
rect 301 599 339 615
rect 301 565 303 599
rect 337 565 339 599
rect 301 519 339 565
rect 301 485 303 519
rect 337 485 339 519
rect 129 400 131 434
rect 165 420 167 434
rect 301 434 339 485
rect 301 420 303 434
rect 165 400 303 420
rect 337 400 339 434
rect 373 611 439 649
rect 373 577 389 611
rect 423 577 439 611
rect 373 534 439 577
rect 373 500 389 534
rect 423 500 439 534
rect 373 457 439 500
rect 373 423 389 457
rect 423 423 439 457
rect 473 599 509 615
rect 473 565 475 599
rect 473 508 509 565
rect 545 568 611 649
rect 545 534 561 568
rect 595 534 611 568
rect 545 526 611 534
rect 645 599 683 615
rect 645 565 647 599
rect 681 565 683 599
rect 473 474 475 508
rect 645 508 683 565
rect 717 568 783 649
rect 717 534 733 568
rect 767 534 783 568
rect 717 526 783 534
rect 821 599 861 615
rect 821 565 825 599
rect 859 565 861 599
rect 645 492 647 508
rect 509 474 647 492
rect 681 492 683 508
rect 821 508 861 565
rect 895 568 961 649
rect 895 534 911 568
rect 945 534 961 568
rect 895 526 961 534
rect 995 599 1033 615
rect 995 565 997 599
rect 1031 565 1033 599
rect 821 492 825 508
rect 681 474 825 492
rect 859 492 861 508
rect 995 508 1033 565
rect 995 492 997 508
rect 859 474 997 492
rect 1031 474 1033 508
rect 473 458 1033 474
rect 1067 607 1133 649
rect 1067 573 1083 607
rect 1117 573 1133 607
rect 1067 492 1133 573
rect 1067 458 1083 492
rect 1117 458 1133 492
rect 129 389 339 400
rect 473 413 525 458
rect 473 389 475 413
rect 129 384 475 389
rect 299 379 475 384
rect 509 379 525 413
rect 299 355 525 379
rect 559 384 1086 424
rect 17 319 262 350
rect 17 285 76 319
rect 110 285 144 319
rect 178 285 212 319
rect 246 285 262 319
rect 17 279 262 285
rect 299 285 400 355
rect 559 321 636 384
rect 434 319 636 321
rect 434 285 450 319
rect 484 285 518 319
rect 552 285 586 319
rect 620 285 636 319
rect 678 319 986 350
rect 678 285 694 319
rect 728 285 762 319
rect 796 285 830 319
rect 864 285 898 319
rect 932 285 986 319
rect 1040 341 1086 384
rect 1040 319 1108 341
rect 1040 285 1058 319
rect 1092 285 1108 319
rect 299 245 342 285
rect 25 213 85 229
rect 25 179 41 213
rect 75 179 85 213
rect 25 103 85 179
rect 119 211 342 245
rect 119 169 163 211
rect 119 135 127 169
rect 161 135 163 169
rect 119 119 163 135
rect 197 143 213 177
rect 247 143 263 177
rect 25 69 41 103
rect 75 85 85 103
rect 197 103 263 143
rect 297 169 342 211
rect 297 135 299 169
rect 333 135 342 169
rect 297 119 342 135
rect 376 217 1133 251
rect 376 213 421 217
rect 376 179 385 213
rect 419 179 421 213
rect 197 85 213 103
rect 75 69 213 85
rect 247 85 263 103
rect 376 103 421 179
rect 376 85 385 103
rect 247 69 385 85
rect 419 69 421 103
rect 25 51 421 69
rect 455 149 471 183
rect 505 149 521 183
rect 455 103 521 149
rect 555 179 601 217
rect 1081 213 1133 217
rect 555 145 561 179
rect 595 145 601 179
rect 555 129 601 145
rect 635 149 651 183
rect 685 149 825 183
rect 859 149 997 183
rect 1031 149 1047 183
rect 455 69 471 103
rect 505 85 521 103
rect 635 101 701 149
rect 813 140 871 149
rect 986 140 1047 149
rect 1081 179 1083 213
rect 1117 179 1133 213
rect 635 85 651 101
rect 505 69 651 85
rect 455 67 651 69
rect 685 67 701 101
rect 455 51 701 67
rect 735 99 789 115
rect 735 65 739 99
rect 773 65 789 99
rect 735 17 789 65
rect 895 111 961 115
rect 895 77 911 111
rect 945 77 961 111
rect 895 17 961 77
rect 1081 103 1133 179
rect 1081 69 1083 103
rect 1117 69 1133 103
rect 1081 53 1133 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand3_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 411942
string GDS_START 401742
<< end >>
