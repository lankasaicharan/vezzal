magic
tech sky130A
magscale 1 2
timestamp 1627202617
<< checkpaint >>
rect -1298 -1308 2494 1852
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 98 157 940 203
rect 1 21 1195 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 174 47 204 177
rect 258 47 288 177
rect 342 47 372 177
rect 426 47 456 177
rect 526 47 556 177
rect 622 47 652 177
rect 736 47 766 177
rect 832 47 862 177
rect 1087 47 1117 131
<< scpmoshvt >>
rect 79 413 109 497
rect 174 297 204 497
rect 258 297 288 497
rect 342 297 372 497
rect 426 297 456 497
rect 526 297 556 497
rect 622 297 652 497
rect 736 297 766 497
rect 832 297 862 497
rect 1087 413 1117 497
<< ndiff >>
rect 124 131 174 177
rect 27 101 79 131
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 93 174 131
rect 109 59 130 93
rect 164 59 174 93
rect 109 47 174 59
rect 204 101 258 177
rect 204 67 214 101
rect 248 67 258 101
rect 204 47 258 67
rect 288 94 342 177
rect 288 60 298 94
rect 332 60 342 94
rect 288 47 342 60
rect 372 101 426 177
rect 372 67 382 101
rect 416 67 426 101
rect 372 47 426 67
rect 456 89 526 177
rect 456 55 470 89
rect 504 55 526 89
rect 456 47 526 55
rect 556 47 622 177
rect 652 47 736 177
rect 766 47 832 177
rect 862 162 914 177
rect 862 128 872 162
rect 906 128 914 162
rect 862 94 914 128
rect 862 60 872 94
rect 906 60 914 94
rect 862 47 914 60
rect 1003 93 1087 131
rect 1003 59 1011 93
rect 1045 59 1087 93
rect 1003 47 1087 59
rect 1117 101 1169 131
rect 1117 67 1127 101
rect 1161 67 1169 101
rect 1117 47 1169 67
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 413 79 443
rect 109 485 174 497
rect 109 451 119 485
rect 153 451 174 485
rect 109 413 174 451
rect 124 297 174 413
rect 204 343 258 497
rect 204 309 214 343
rect 248 309 258 343
rect 204 297 258 309
rect 288 485 342 497
rect 288 451 298 485
rect 332 451 342 485
rect 288 297 342 451
rect 372 343 426 497
rect 372 309 382 343
rect 416 309 426 343
rect 372 297 426 309
rect 456 485 526 497
rect 456 451 466 485
rect 500 451 526 485
rect 456 297 526 451
rect 556 343 622 497
rect 556 309 578 343
rect 612 309 622 343
rect 556 297 622 309
rect 652 485 736 497
rect 652 451 682 485
rect 716 451 736 485
rect 652 297 736 451
rect 766 343 832 497
rect 766 309 780 343
rect 814 309 832 343
rect 766 297 832 309
rect 862 485 1087 497
rect 862 451 888 485
rect 922 451 956 485
rect 990 451 1024 485
rect 1058 451 1087 485
rect 862 413 1087 451
rect 1117 477 1169 497
rect 1117 443 1127 477
rect 1161 443 1169 477
rect 1117 413 1169 443
rect 862 297 914 413
<< ndiffc >>
rect 35 67 69 101
rect 130 59 164 93
rect 214 67 248 101
rect 298 60 332 94
rect 382 67 416 101
rect 470 55 504 89
rect 872 128 906 162
rect 872 60 906 94
rect 1011 59 1045 93
rect 1127 67 1161 101
<< pdiffc >>
rect 35 443 69 477
rect 119 451 153 485
rect 214 309 248 343
rect 298 451 332 485
rect 382 309 416 343
rect 466 451 500 485
rect 578 309 612 343
rect 682 451 716 485
rect 780 309 814 343
rect 888 451 922 485
rect 956 451 990 485
rect 1024 451 1058 485
rect 1127 443 1161 477
<< poly >>
rect 79 497 109 523
rect 174 497 204 523
rect 258 497 288 523
rect 342 497 372 523
rect 426 497 456 523
rect 526 497 556 523
rect 622 497 652 523
rect 736 497 766 523
rect 832 497 862 523
rect 1087 497 1117 523
rect 79 265 109 413
rect 174 275 204 297
rect 258 275 288 297
rect 342 275 372 297
rect 426 275 456 297
rect 76 249 130 265
rect 76 215 86 249
rect 120 215 130 249
rect 76 199 130 215
rect 174 259 456 275
rect 526 265 556 297
rect 622 265 652 297
rect 736 265 766 297
rect 832 265 862 297
rect 1087 265 1117 413
rect 174 249 484 259
rect 174 215 298 249
rect 332 215 366 249
rect 400 215 434 249
rect 468 215 484 249
rect 174 205 484 215
rect 526 249 580 265
rect 526 215 536 249
rect 570 215 580 249
rect 79 131 109 199
rect 174 177 204 205
rect 258 177 288 205
rect 342 177 372 205
rect 426 177 456 205
rect 526 199 580 215
rect 622 249 694 265
rect 622 215 650 249
rect 684 215 694 249
rect 622 199 694 215
rect 736 249 790 265
rect 736 215 746 249
rect 780 215 790 249
rect 736 199 790 215
rect 832 249 1044 265
rect 832 215 990 249
rect 1024 215 1044 249
rect 832 199 1044 215
rect 1087 249 1141 265
rect 1087 215 1097 249
rect 1131 215 1141 249
rect 1087 199 1141 215
rect 526 177 556 199
rect 622 177 652 199
rect 736 177 766 199
rect 832 177 862 199
rect 1087 131 1117 199
rect 79 21 109 47
rect 174 21 204 47
rect 258 21 288 47
rect 342 21 372 47
rect 426 21 456 47
rect 526 21 556 47
rect 622 21 652 47
rect 736 21 766 47
rect 832 21 862 47
rect 1087 21 1117 47
<< polycont >>
rect 86 215 120 249
rect 298 215 332 249
rect 366 215 400 249
rect 434 215 468 249
rect 536 215 570 249
rect 650 215 684 249
rect 746 215 780 249
rect 990 215 1024 249
rect 1097 215 1131 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 477 69 493
rect 17 443 35 477
rect 103 485 169 527
rect 103 451 119 485
rect 153 451 169 485
rect 282 485 348 527
rect 282 451 298 485
rect 332 451 348 485
rect 450 485 516 527
rect 450 451 466 485
rect 500 451 516 485
rect 666 485 732 527
rect 666 451 682 485
rect 716 451 732 485
rect 872 485 1074 527
rect 872 451 888 485
rect 922 451 956 485
rect 990 451 1024 485
rect 1058 451 1074 485
rect 1127 477 1161 493
rect 17 417 69 443
rect 1127 417 1161 443
rect 17 383 898 417
rect 17 117 52 383
rect 86 249 156 327
rect 120 215 156 249
rect 86 153 156 215
rect 192 309 214 343
rect 248 309 382 343
rect 416 309 432 343
rect 466 309 578 343
rect 612 309 780 343
rect 814 309 830 343
rect 192 164 248 309
rect 466 249 500 309
rect 864 265 898 383
rect 282 215 298 249
rect 332 215 366 249
rect 400 215 434 249
rect 468 215 500 249
rect 192 130 416 164
rect 17 101 69 117
rect 17 67 35 101
rect 214 101 248 130
rect 17 51 69 67
rect 114 93 180 94
rect 114 59 130 93
rect 164 59 180 93
rect 114 17 180 59
rect 382 101 416 130
rect 466 157 500 215
rect 536 249 616 265
rect 570 215 616 249
rect 536 199 616 215
rect 650 249 709 265
rect 684 215 709 249
rect 466 123 588 157
rect 650 151 709 215
rect 746 249 898 265
rect 780 231 898 249
rect 990 383 1161 417
rect 990 249 1024 383
rect 746 199 780 215
rect 990 165 1024 215
rect 1097 249 1169 324
rect 1131 215 1169 249
rect 1097 199 1169 215
rect 214 51 248 67
rect 282 60 298 94
rect 332 60 348 94
rect 282 17 348 60
rect 554 94 588 123
rect 851 128 872 162
rect 906 128 922 162
rect 990 131 1161 165
rect 851 94 922 128
rect 382 51 416 67
rect 454 55 470 89
rect 504 55 520 89
rect 554 60 872 94
rect 906 60 922 94
rect 1127 101 1161 131
rect 454 17 520 55
rect 995 59 1011 93
rect 1045 59 1061 93
rect 995 17 1061 59
rect 1127 51 1161 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 674 221 708 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 674 153 708 187 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 1132 289 1166 323 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 1132 221 1166 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 214 289 248 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 122 153 156 187 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel locali s 122 289 156 323 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel locali s 214 153 248 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 and4bb_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 3093466
string GDS_START 3084808
string path 0.000 0.000 29.900 0.000 
<< end >>
