magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 1004 241 1631 263
rect 31 49 1631 241
rect 0 0 1632 49
<< scnmos >>
rect 110 47 140 215
rect 196 47 226 215
rect 282 47 312 215
rect 368 47 398 215
rect 454 47 484 215
rect 540 47 570 215
rect 626 47 656 215
rect 714 47 744 215
rect 806 47 836 215
rect 892 47 922 215
rect 978 47 1008 215
rect 1110 69 1140 237
rect 1196 69 1226 237
rect 1314 69 1344 237
rect 1400 69 1430 237
rect 1518 69 1548 237
<< scpmoshvt >>
rect 110 367 140 619
rect 196 367 226 619
rect 282 367 312 619
rect 368 367 398 619
rect 454 367 484 619
rect 540 367 570 619
rect 626 367 656 619
rect 712 367 742 619
rect 806 367 836 619
rect 892 367 922 619
rect 978 367 1008 619
rect 1064 367 1094 619
rect 1150 367 1180 619
rect 1236 367 1266 619
rect 1390 367 1420 619
rect 1476 367 1506 619
<< ndiff >>
rect 1030 215 1110 237
rect 57 203 110 215
rect 57 169 65 203
rect 99 169 110 203
rect 57 101 110 169
rect 57 67 65 101
rect 99 67 110 101
rect 57 47 110 67
rect 140 161 196 215
rect 140 127 151 161
rect 185 127 196 161
rect 140 89 196 127
rect 140 55 151 89
rect 185 55 196 89
rect 140 47 196 55
rect 226 203 282 215
rect 226 169 237 203
rect 271 169 282 203
rect 226 101 282 169
rect 226 67 237 101
rect 271 67 282 101
rect 226 47 282 67
rect 312 157 368 215
rect 312 123 323 157
rect 357 123 368 157
rect 312 89 368 123
rect 312 55 323 89
rect 357 55 368 89
rect 312 47 368 55
rect 398 203 454 215
rect 398 169 409 203
rect 443 169 454 203
rect 398 101 454 169
rect 398 67 409 101
rect 443 67 454 101
rect 398 47 454 67
rect 484 161 540 215
rect 484 127 495 161
rect 529 127 540 161
rect 484 89 540 127
rect 484 55 495 89
rect 529 55 540 89
rect 484 47 540 55
rect 570 203 626 215
rect 570 169 581 203
rect 615 169 626 203
rect 570 101 626 169
rect 570 67 581 101
rect 615 67 626 101
rect 570 47 626 67
rect 656 160 714 215
rect 656 126 667 160
rect 701 126 714 160
rect 656 89 714 126
rect 656 55 667 89
rect 701 55 714 89
rect 656 47 714 55
rect 744 203 806 215
rect 744 169 757 203
rect 791 169 806 203
rect 744 101 806 169
rect 744 67 757 101
rect 791 67 806 101
rect 744 47 806 67
rect 836 159 892 215
rect 836 125 847 159
rect 881 125 892 159
rect 836 91 892 125
rect 836 57 847 91
rect 881 57 892 91
rect 836 47 892 57
rect 922 175 978 215
rect 922 141 933 175
rect 967 141 978 175
rect 922 47 978 141
rect 1008 89 1110 215
rect 1008 55 1042 89
rect 1076 69 1110 89
rect 1140 229 1196 237
rect 1140 195 1151 229
rect 1185 195 1196 229
rect 1140 69 1196 195
rect 1226 89 1314 237
rect 1226 69 1253 89
rect 1076 55 1088 69
rect 1008 47 1088 55
rect 1241 55 1253 69
rect 1287 69 1314 89
rect 1344 229 1400 237
rect 1344 195 1355 229
rect 1389 195 1400 229
rect 1344 69 1400 195
rect 1430 89 1518 237
rect 1430 69 1457 89
rect 1287 55 1299 69
rect 1241 47 1299 55
rect 1445 55 1457 69
rect 1491 69 1518 89
rect 1548 179 1605 237
rect 1548 145 1559 179
rect 1593 145 1605 179
rect 1548 111 1605 145
rect 1548 77 1559 111
rect 1593 77 1605 111
rect 1548 69 1605 77
rect 1491 55 1503 69
rect 1445 47 1503 55
<< pdiff >>
rect 57 607 110 619
rect 57 573 65 607
rect 99 573 110 607
rect 57 505 110 573
rect 57 471 65 505
rect 99 471 110 505
rect 57 413 110 471
rect 57 379 65 413
rect 99 379 110 413
rect 57 367 110 379
rect 140 599 196 619
rect 140 565 151 599
rect 185 565 196 599
rect 140 505 196 565
rect 140 471 151 505
rect 185 471 196 505
rect 140 413 196 471
rect 140 379 151 413
rect 185 379 196 413
rect 140 367 196 379
rect 226 580 282 619
rect 226 546 237 580
rect 271 546 282 580
rect 226 367 282 546
rect 312 599 368 619
rect 312 565 323 599
rect 357 565 368 599
rect 312 508 368 565
rect 312 474 323 508
rect 357 474 368 508
rect 312 367 368 474
rect 398 510 454 619
rect 398 476 409 510
rect 443 476 454 510
rect 398 367 454 476
rect 484 600 540 619
rect 484 566 495 600
rect 529 566 540 600
rect 484 367 540 566
rect 570 498 626 619
rect 570 464 581 498
rect 615 464 626 498
rect 570 367 626 464
rect 656 586 712 619
rect 656 552 667 586
rect 701 552 712 586
rect 656 367 712 552
rect 742 578 806 619
rect 742 544 757 578
rect 791 544 806 578
rect 742 367 806 544
rect 836 599 892 619
rect 836 565 847 599
rect 881 565 892 599
rect 836 518 892 565
rect 836 484 847 518
rect 881 484 892 518
rect 836 436 892 484
rect 836 402 847 436
rect 881 402 892 436
rect 836 367 892 402
rect 922 566 978 619
rect 922 532 933 566
rect 967 532 978 566
rect 922 367 978 532
rect 1008 599 1064 619
rect 1008 565 1019 599
rect 1053 565 1064 599
rect 1008 489 1064 565
rect 1008 455 1019 489
rect 1053 455 1064 489
rect 1008 367 1064 455
rect 1094 572 1150 619
rect 1094 538 1105 572
rect 1139 538 1150 572
rect 1094 367 1150 538
rect 1180 599 1236 619
rect 1180 565 1191 599
rect 1225 565 1236 599
rect 1180 488 1236 565
rect 1180 454 1191 488
rect 1225 454 1236 488
rect 1180 367 1236 454
rect 1266 578 1390 619
rect 1266 544 1277 578
rect 1311 544 1345 578
rect 1379 544 1390 578
rect 1266 367 1390 544
rect 1420 599 1476 619
rect 1420 565 1431 599
rect 1465 565 1476 599
rect 1420 492 1476 565
rect 1420 458 1431 492
rect 1465 458 1476 492
rect 1420 367 1476 458
rect 1506 582 1559 619
rect 1506 548 1517 582
rect 1551 548 1559 582
rect 1506 367 1559 548
<< ndiffc >>
rect 65 169 99 203
rect 65 67 99 101
rect 151 127 185 161
rect 151 55 185 89
rect 237 169 271 203
rect 237 67 271 101
rect 323 123 357 157
rect 323 55 357 89
rect 409 169 443 203
rect 409 67 443 101
rect 495 127 529 161
rect 495 55 529 89
rect 581 169 615 203
rect 581 67 615 101
rect 667 126 701 160
rect 667 55 701 89
rect 757 169 791 203
rect 757 67 791 101
rect 847 125 881 159
rect 847 57 881 91
rect 933 141 967 175
rect 1042 55 1076 89
rect 1151 195 1185 229
rect 1253 55 1287 89
rect 1355 195 1389 229
rect 1457 55 1491 89
rect 1559 145 1593 179
rect 1559 77 1593 111
<< pdiffc >>
rect 65 573 99 607
rect 65 471 99 505
rect 65 379 99 413
rect 151 565 185 599
rect 151 471 185 505
rect 151 379 185 413
rect 237 546 271 580
rect 323 565 357 599
rect 323 474 357 508
rect 409 476 443 510
rect 495 566 529 600
rect 581 464 615 498
rect 667 552 701 586
rect 757 544 791 578
rect 847 565 881 599
rect 847 484 881 518
rect 847 402 881 436
rect 933 532 967 566
rect 1019 565 1053 599
rect 1019 455 1053 489
rect 1105 538 1139 572
rect 1191 565 1225 599
rect 1191 454 1225 488
rect 1277 544 1311 578
rect 1345 544 1379 578
rect 1431 565 1465 599
rect 1431 458 1465 492
rect 1517 548 1551 582
<< poly >>
rect 110 619 140 645
rect 196 619 226 645
rect 282 619 312 645
rect 368 619 398 645
rect 454 619 484 645
rect 540 619 570 645
rect 626 619 656 645
rect 712 619 742 645
rect 806 619 836 645
rect 892 619 922 645
rect 978 619 1008 645
rect 1064 619 1094 645
rect 1150 619 1180 645
rect 1236 619 1266 645
rect 1390 619 1420 645
rect 1476 619 1506 645
rect 110 325 140 367
rect 196 325 226 367
rect 282 325 312 367
rect 42 309 312 325
rect 42 275 58 309
rect 92 275 126 309
rect 160 275 194 309
rect 228 275 262 309
rect 296 275 312 309
rect 42 259 312 275
rect 110 215 140 259
rect 196 215 226 259
rect 282 215 312 259
rect 368 345 398 367
rect 454 345 484 367
rect 540 345 570 367
rect 626 345 656 367
rect 368 319 656 345
rect 712 335 742 367
rect 806 335 836 367
rect 892 335 922 367
rect 978 335 1008 367
rect 368 285 387 319
rect 421 285 455 319
rect 489 285 523 319
rect 557 285 591 319
rect 625 285 656 319
rect 368 269 656 285
rect 698 319 764 335
rect 698 285 714 319
rect 748 285 764 319
rect 698 269 764 285
rect 806 319 1008 335
rect 806 285 822 319
rect 856 285 890 319
rect 924 285 958 319
rect 992 285 1008 319
rect 806 269 1008 285
rect 1064 335 1094 367
rect 1150 335 1180 367
rect 1236 335 1266 367
rect 1390 335 1420 367
rect 1064 319 1420 335
rect 1064 285 1087 319
rect 1121 285 1155 319
rect 1189 285 1223 319
rect 1257 285 1291 319
rect 1325 285 1359 319
rect 1393 299 1420 319
rect 1476 335 1506 367
rect 1476 319 1548 335
rect 1476 305 1494 319
rect 1393 285 1430 299
rect 1064 269 1430 285
rect 1478 285 1494 305
rect 1528 285 1548 319
rect 1478 269 1548 285
rect 368 215 398 269
rect 454 215 484 269
rect 540 215 570 269
rect 626 215 656 269
rect 714 215 744 269
rect 806 215 836 269
rect 892 215 922 269
rect 978 215 1008 269
rect 1110 237 1140 269
rect 1196 237 1226 269
rect 1314 237 1344 269
rect 1400 237 1430 269
rect 1518 237 1548 269
rect 110 21 140 47
rect 196 21 226 47
rect 282 21 312 47
rect 368 21 398 47
rect 454 21 484 47
rect 540 21 570 47
rect 626 21 656 47
rect 714 21 744 47
rect 806 21 836 47
rect 892 21 922 47
rect 978 21 1008 47
rect 1110 43 1140 69
rect 1196 43 1226 69
rect 1314 43 1344 69
rect 1400 43 1430 69
rect 1518 43 1548 69
<< polycont >>
rect 58 275 92 309
rect 126 275 160 309
rect 194 275 228 309
rect 262 275 296 309
rect 387 285 421 319
rect 455 285 489 319
rect 523 285 557 319
rect 591 285 625 319
rect 714 285 748 319
rect 822 285 856 319
rect 890 285 924 319
rect 958 285 992 319
rect 1087 285 1121 319
rect 1155 285 1189 319
rect 1223 285 1257 319
rect 1291 285 1325 319
rect 1359 285 1393 319
rect 1494 285 1528 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 49 607 107 649
rect 49 573 65 607
rect 99 573 107 607
rect 49 505 107 573
rect 49 471 65 505
rect 99 471 107 505
rect 49 413 107 471
rect 49 379 65 413
rect 99 379 107 413
rect 49 363 107 379
rect 141 599 185 615
rect 141 565 151 599
rect 141 505 185 565
rect 221 580 287 649
rect 221 546 237 580
rect 271 546 287 580
rect 221 538 287 546
rect 321 600 705 615
rect 321 599 495 600
rect 321 565 323 599
rect 357 566 495 599
rect 529 586 705 600
rect 529 566 667 586
rect 357 565 667 566
rect 321 562 667 565
rect 141 471 151 505
rect 321 508 361 562
rect 663 552 667 562
rect 701 552 705 586
rect 663 536 705 552
rect 741 578 807 649
rect 741 544 757 578
rect 791 544 807 578
rect 741 536 807 544
rect 841 599 883 615
rect 841 565 847 599
rect 881 565 883 599
rect 321 504 323 508
rect 185 474 323 504
rect 357 474 361 508
rect 185 471 361 474
rect 141 458 361 471
rect 405 510 447 526
rect 405 476 409 510
rect 443 502 447 510
rect 841 518 883 565
rect 917 566 983 649
rect 917 532 933 566
rect 967 532 983 566
rect 917 522 983 532
rect 1017 599 1062 615
rect 1017 565 1019 599
rect 1053 565 1062 599
rect 841 502 847 518
rect 443 498 847 502
rect 443 476 581 498
rect 405 464 581 476
rect 615 484 847 498
rect 881 488 883 518
rect 1017 489 1062 565
rect 1096 572 1146 649
rect 1096 538 1105 572
rect 1139 538 1146 572
rect 1096 522 1146 538
rect 1180 599 1227 615
rect 1180 565 1191 599
rect 1225 565 1227 599
rect 1017 488 1019 489
rect 881 484 1019 488
rect 615 464 1019 484
rect 405 458 1019 464
rect 141 413 185 458
rect 843 455 1019 458
rect 1053 488 1062 489
rect 1180 501 1227 565
rect 1261 578 1395 649
rect 1261 544 1277 578
rect 1311 544 1345 578
rect 1379 544 1395 578
rect 1261 535 1395 544
rect 1429 599 1467 615
rect 1429 565 1431 599
rect 1465 565 1467 599
rect 1429 501 1467 565
rect 1501 582 1567 649
rect 1501 548 1517 582
rect 1551 548 1567 582
rect 1501 535 1567 548
rect 1180 492 1614 501
rect 1180 488 1431 492
rect 1053 455 1191 488
rect 843 454 1191 455
rect 1225 458 1431 488
rect 1465 458 1614 492
rect 1225 454 1614 458
rect 843 436 885 454
rect 141 379 151 413
rect 141 363 185 379
rect 223 385 756 424
rect 843 402 847 436
rect 881 402 885 436
rect 843 386 885 402
rect 991 386 1544 420
rect 223 326 312 385
rect 42 309 312 326
rect 42 275 58 309
rect 92 275 126 309
rect 160 275 194 309
rect 228 275 262 309
rect 296 275 312 309
rect 371 319 666 350
rect 371 285 387 319
rect 421 285 455 319
rect 489 285 523 319
rect 557 285 591 319
rect 625 285 666 319
rect 700 319 756 385
rect 991 352 1025 386
rect 700 285 714 319
rect 748 285 756 319
rect 42 269 312 275
rect 700 269 756 285
rect 790 319 1025 352
rect 790 285 822 319
rect 856 285 890 319
rect 924 285 958 319
rect 992 285 1025 319
rect 1071 319 1409 352
rect 1071 285 1087 319
rect 1121 285 1155 319
rect 1189 285 1223 319
rect 1257 285 1291 319
rect 1325 285 1359 319
rect 1393 285 1409 319
rect 1478 319 1544 386
rect 1478 285 1494 319
rect 1528 285 1544 319
rect 790 269 1025 285
rect 1578 251 1614 454
rect 61 203 983 235
rect 61 169 65 203
rect 99 199 237 203
rect 99 169 101 199
rect 61 101 101 169
rect 235 169 237 199
rect 271 199 409 203
rect 271 169 273 199
rect 61 67 65 101
rect 99 67 101 101
rect 61 51 101 67
rect 135 161 201 165
rect 135 127 151 161
rect 185 127 201 161
rect 135 89 201 127
rect 135 55 151 89
rect 185 55 201 89
rect 135 17 201 55
rect 235 101 273 169
rect 407 169 409 199
rect 443 199 581 203
rect 443 169 445 199
rect 235 67 237 101
rect 271 67 273 101
rect 235 51 273 67
rect 307 157 373 161
rect 307 123 323 157
rect 357 123 373 157
rect 307 89 373 123
rect 307 55 323 89
rect 357 55 373 89
rect 307 17 373 55
rect 407 101 445 169
rect 579 169 581 199
rect 615 199 757 203
rect 615 169 617 199
rect 407 67 409 101
rect 443 67 445 101
rect 407 51 445 67
rect 479 161 545 165
rect 479 127 495 161
rect 529 127 545 161
rect 479 89 545 127
rect 479 55 495 89
rect 529 55 545 89
rect 479 17 545 55
rect 579 101 617 169
rect 751 169 757 199
rect 791 199 983 203
rect 791 169 797 199
rect 579 67 581 101
rect 615 67 617 101
rect 579 51 617 67
rect 651 160 717 165
rect 651 126 667 160
rect 701 126 717 160
rect 651 89 717 126
rect 651 55 667 89
rect 701 55 717 89
rect 651 17 717 55
rect 751 101 797 169
rect 931 175 983 199
rect 1135 229 1614 251
rect 1135 195 1151 229
rect 1185 195 1355 229
rect 1389 215 1614 229
rect 1389 195 1405 215
rect 1135 193 1405 195
rect 751 67 757 101
rect 791 67 797 101
rect 751 51 797 67
rect 831 159 897 165
rect 831 125 847 159
rect 881 125 897 159
rect 931 141 933 175
rect 967 159 983 175
rect 1543 179 1609 181
rect 1543 159 1559 179
rect 967 145 1559 159
rect 1593 145 1609 179
rect 967 141 1609 145
rect 931 125 1609 141
rect 831 91 897 125
rect 1543 111 1609 125
rect 831 57 847 91
rect 881 89 1507 91
rect 881 57 1042 89
rect 831 55 1042 57
rect 1076 55 1253 89
rect 1287 55 1457 89
rect 1491 55 1507 89
rect 1543 77 1559 111
rect 1593 77 1609 111
rect 1543 73 1609 77
rect 831 53 1507 55
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o211ai_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 464 1217 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1279 464 1313 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1375 464 1409 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1471 464 1505 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6780132
string GDS_START 6766446
<< end >>
