magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 1 49 491 241
rect 0 0 576 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 296 47 326 215
rect 382 47 412 215
<< scpmoshvt >>
rect 80 367 110 619
rect 176 367 206 619
rect 274 367 304 619
rect 382 367 412 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 93 80 169
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 203 166 215
rect 110 169 121 203
rect 155 169 166 203
rect 110 101 166 169
rect 110 67 121 101
rect 155 67 166 101
rect 110 47 166 67
rect 196 174 296 215
rect 196 140 229 174
rect 263 140 296 174
rect 196 93 296 140
rect 196 59 229 93
rect 263 59 296 93
rect 196 47 296 59
rect 326 203 382 215
rect 326 169 337 203
rect 371 169 382 203
rect 326 101 382 169
rect 326 67 337 101
rect 371 67 382 101
rect 326 47 382 67
rect 412 174 465 215
rect 412 140 423 174
rect 457 140 465 174
rect 412 93 465 140
rect 412 59 423 93
rect 457 59 465 93
rect 412 47 465 59
<< pdiff >>
rect 27 607 80 619
rect 27 573 35 607
rect 69 573 80 607
rect 27 512 80 573
rect 27 478 35 512
rect 69 478 80 512
rect 27 418 80 478
rect 27 384 35 418
rect 69 384 80 418
rect 27 367 80 384
rect 110 367 176 619
rect 206 367 274 619
rect 304 367 382 619
rect 412 607 465 619
rect 412 573 423 607
rect 457 573 465 607
rect 412 513 465 573
rect 412 479 423 513
rect 457 479 465 513
rect 412 420 465 479
rect 412 386 423 420
rect 457 386 465 420
rect 412 367 465 386
<< ndiffc >>
rect 35 169 69 203
rect 35 59 69 93
rect 121 169 155 203
rect 121 67 155 101
rect 229 140 263 174
rect 229 59 263 93
rect 337 169 371 203
rect 337 67 371 101
rect 423 140 457 174
rect 423 59 457 93
<< pdiffc >>
rect 35 573 69 607
rect 35 478 69 512
rect 35 384 69 418
rect 423 573 457 607
rect 423 479 457 513
rect 423 386 457 420
<< poly >>
rect 80 619 110 645
rect 176 619 206 645
rect 274 619 304 645
rect 382 619 412 645
rect 80 335 110 367
rect 176 335 206 367
rect 274 335 304 367
rect 42 319 110 335
rect 42 285 59 319
rect 93 285 110 319
rect 42 269 110 285
rect 152 319 218 335
rect 152 285 168 319
rect 202 285 218 319
rect 152 269 218 285
rect 260 319 326 335
rect 260 285 276 319
rect 310 285 326 319
rect 260 269 326 285
rect 80 215 110 269
rect 166 215 196 269
rect 296 215 326 269
rect 382 308 412 367
rect 382 292 506 308
rect 382 258 456 292
rect 490 258 506 292
rect 382 242 506 258
rect 382 215 412 242
rect 80 21 110 47
rect 166 21 196 47
rect 296 21 326 47
rect 382 21 412 47
<< polycont >>
rect 59 285 93 319
rect 168 285 202 319
rect 276 285 310 319
rect 456 258 490 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 19 607 85 649
rect 19 573 35 607
rect 69 573 85 607
rect 388 607 473 615
rect 19 512 85 573
rect 19 478 35 512
rect 69 478 85 512
rect 19 418 85 478
rect 19 384 35 418
rect 69 384 85 418
rect 119 384 184 582
rect 127 380 184 384
rect 17 319 93 350
rect 17 285 59 319
rect 127 319 218 380
rect 282 342 354 582
rect 127 285 168 319
rect 202 285 218 319
rect 260 319 354 342
rect 260 285 276 319
rect 310 285 354 319
rect 388 573 423 607
rect 457 573 473 607
rect 388 513 473 573
rect 388 479 423 513
rect 457 479 473 513
rect 388 420 473 479
rect 388 386 423 420
rect 457 386 473 420
rect 17 269 93 285
rect 388 247 422 386
rect 19 203 85 219
rect 19 169 35 203
rect 69 169 85 203
rect 19 93 85 169
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 119 213 422 247
rect 456 292 545 352
rect 490 258 545 292
rect 456 213 545 258
rect 119 203 171 213
rect 119 169 121 203
rect 155 169 171 203
rect 321 203 373 213
rect 119 101 171 169
rect 119 67 121 101
rect 155 67 171 101
rect 119 51 171 67
rect 213 174 279 179
rect 213 140 229 174
rect 263 140 279 174
rect 213 93 279 140
rect 213 59 229 93
rect 263 59 279 93
rect 213 17 279 59
rect 321 169 337 203
rect 371 169 373 203
rect 321 101 373 169
rect 321 67 337 101
rect 371 67 373 101
rect 321 51 373 67
rect 407 174 473 179
rect 407 140 423 174
rect 457 140 473 174
rect 407 93 473 140
rect 407 59 423 93
rect 457 59 473 93
rect 407 17 473 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4_1
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4159220
string GDS_START 4152948
<< end >>
