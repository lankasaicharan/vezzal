magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
rect 952 313 1160 331
<< pwell >>
rect 1155 241 1343 255
rect 33 157 307 239
rect 940 157 1343 241
rect 33 49 1343 157
rect 0 0 1344 49
<< scnmos >>
rect 112 129 142 213
rect 198 129 228 213
rect 540 47 570 131
rect 626 47 656 131
rect 698 47 728 131
rect 806 47 836 131
rect 914 47 944 131
rect 1019 47 1049 215
rect 1234 61 1264 229
<< scpmoshvt >>
rect 112 481 142 609
rect 198 481 228 609
rect 395 481 425 609
rect 554 481 584 609
rect 626 481 656 609
rect 734 481 764 565
rect 842 481 872 565
rect 1041 349 1071 601
rect 1234 367 1264 619
<< ndiff >>
rect 59 185 112 213
rect 59 151 67 185
rect 101 151 112 185
rect 59 129 112 151
rect 142 185 198 213
rect 142 151 153 185
rect 187 151 198 185
rect 142 129 198 151
rect 228 199 281 213
rect 228 165 239 199
rect 273 165 281 199
rect 228 129 281 165
rect 966 201 1019 215
rect 966 167 974 201
rect 1008 167 1019 201
rect 966 131 1019 167
rect 487 109 540 131
rect 487 75 495 109
rect 529 75 540 109
rect 487 47 540 75
rect 570 94 626 131
rect 570 60 581 94
rect 615 60 626 94
rect 570 47 626 60
rect 656 47 698 131
rect 728 89 806 131
rect 728 55 761 89
rect 795 55 806 89
rect 728 47 806 55
rect 836 47 914 131
rect 944 93 1019 131
rect 944 59 968 93
rect 1002 59 1019 93
rect 944 47 1019 59
rect 1049 199 1102 215
rect 1049 165 1060 199
rect 1094 165 1102 199
rect 1049 101 1102 165
rect 1049 67 1060 101
rect 1094 67 1102 101
rect 1049 47 1102 67
rect 1181 201 1234 229
rect 1181 167 1189 201
rect 1223 167 1234 201
rect 1181 107 1234 167
rect 1181 73 1189 107
rect 1223 73 1234 107
rect 1181 61 1234 73
rect 1264 212 1317 229
rect 1264 178 1275 212
rect 1309 178 1317 212
rect 1264 107 1317 178
rect 1264 73 1275 107
rect 1309 73 1317 107
rect 1264 61 1317 73
<< pdiff >>
rect 59 597 112 609
rect 59 563 67 597
rect 101 563 112 597
rect 59 527 112 563
rect 59 493 67 527
rect 101 493 112 527
rect 59 481 112 493
rect 142 597 198 609
rect 142 563 153 597
rect 187 563 198 597
rect 142 527 198 563
rect 142 493 153 527
rect 187 493 198 527
rect 142 481 198 493
rect 228 597 281 609
rect 228 563 239 597
rect 273 563 281 597
rect 228 527 281 563
rect 228 493 239 527
rect 273 493 281 527
rect 228 481 281 493
rect 342 531 395 609
rect 342 497 350 531
rect 384 497 395 531
rect 342 481 395 497
rect 425 593 554 609
rect 425 559 490 593
rect 524 559 554 593
rect 425 481 554 559
rect 584 481 626 609
rect 656 593 709 609
rect 1181 607 1234 619
rect 656 559 667 593
rect 701 565 709 593
rect 988 589 1041 601
rect 988 565 996 589
rect 701 559 734 565
rect 656 481 734 559
rect 764 481 842 565
rect 872 555 996 565
rect 1030 555 1041 589
rect 872 540 1041 555
rect 872 506 890 540
rect 924 521 1041 540
rect 924 506 996 521
rect 872 487 996 506
rect 1030 487 1041 521
rect 872 481 1041 487
rect 988 349 1041 481
rect 1071 589 1124 601
rect 1071 555 1082 589
rect 1116 555 1124 589
rect 1071 493 1124 555
rect 1071 459 1082 493
rect 1116 459 1124 493
rect 1071 395 1124 459
rect 1071 361 1082 395
rect 1116 361 1124 395
rect 1181 573 1189 607
rect 1223 573 1234 607
rect 1181 508 1234 573
rect 1181 474 1189 508
rect 1223 474 1234 508
rect 1181 413 1234 474
rect 1181 379 1189 413
rect 1223 379 1234 413
rect 1181 367 1234 379
rect 1264 599 1317 619
rect 1264 565 1275 599
rect 1309 565 1317 599
rect 1264 506 1317 565
rect 1264 472 1275 506
rect 1309 472 1317 506
rect 1264 413 1317 472
rect 1264 379 1275 413
rect 1309 379 1317 413
rect 1264 367 1317 379
rect 1071 349 1124 361
<< ndiffc >>
rect 67 151 101 185
rect 153 151 187 185
rect 239 165 273 199
rect 974 167 1008 201
rect 495 75 529 109
rect 581 60 615 94
rect 761 55 795 89
rect 968 59 1002 93
rect 1060 165 1094 199
rect 1060 67 1094 101
rect 1189 167 1223 201
rect 1189 73 1223 107
rect 1275 178 1309 212
rect 1275 73 1309 107
<< pdiffc >>
rect 67 563 101 597
rect 67 493 101 527
rect 153 563 187 597
rect 153 493 187 527
rect 239 563 273 597
rect 239 493 273 527
rect 350 497 384 531
rect 490 559 524 593
rect 667 559 701 593
rect 996 555 1030 589
rect 890 506 924 540
rect 996 487 1030 521
rect 1082 555 1116 589
rect 1082 459 1116 493
rect 1082 361 1116 395
rect 1189 573 1223 607
rect 1189 474 1223 508
rect 1189 379 1223 413
rect 1275 565 1309 599
rect 1275 472 1309 506
rect 1275 379 1309 413
<< poly >>
rect 112 609 142 635
rect 198 609 228 635
rect 395 609 425 635
rect 554 609 584 635
rect 626 609 656 635
rect 1041 601 1071 627
rect 1234 619 1264 645
rect 734 565 764 591
rect 842 565 872 591
rect 112 301 142 481
rect 84 285 150 301
rect 84 251 100 285
rect 134 251 150 285
rect 84 235 150 251
rect 198 265 228 481
rect 395 317 425 481
rect 554 387 584 481
rect 512 371 584 387
rect 512 337 528 371
rect 562 337 584 371
rect 389 301 455 317
rect 389 267 405 301
rect 439 267 455 301
rect 198 235 333 265
rect 112 213 142 235
rect 198 213 228 235
rect 112 103 142 129
rect 198 103 228 129
rect 303 109 333 235
rect 389 233 455 267
rect 389 199 405 233
rect 439 199 455 233
rect 512 303 584 337
rect 626 441 656 481
rect 734 445 764 481
rect 626 425 692 441
rect 626 391 642 425
rect 676 391 692 425
rect 626 357 692 391
rect 734 429 800 445
rect 734 395 750 429
rect 784 395 800 429
rect 842 443 872 481
rect 842 427 956 443
rect 842 413 906 427
rect 734 379 800 395
rect 890 393 906 413
rect 940 393 956 427
rect 890 377 956 393
rect 626 323 642 357
rect 676 337 692 357
rect 676 323 836 337
rect 626 307 836 323
rect 512 269 528 303
rect 562 269 584 303
rect 512 259 584 269
rect 806 287 836 307
rect 806 271 872 287
rect 512 229 656 259
rect 389 187 455 199
rect 389 157 570 187
rect 540 131 570 157
rect 626 131 656 229
rect 698 233 764 249
rect 698 199 714 233
rect 748 199 764 233
rect 698 183 764 199
rect 806 237 822 271
rect 856 237 872 271
rect 806 203 872 237
rect 698 131 728 183
rect 806 169 822 203
rect 856 169 872 203
rect 806 153 872 169
rect 806 131 836 153
rect 914 131 944 377
rect 1041 317 1071 349
rect 1234 317 1264 367
rect 992 301 1071 317
rect 992 267 1008 301
rect 1042 267 1071 301
rect 992 251 1071 267
rect 1185 301 1264 317
rect 1185 267 1201 301
rect 1235 267 1264 301
rect 1185 251 1264 267
rect 1019 215 1049 251
rect 1234 229 1264 251
rect 303 93 369 109
rect 303 59 319 93
rect 353 59 369 93
rect 303 43 369 59
rect 540 21 570 47
rect 626 21 656 47
rect 698 21 728 47
rect 806 21 836 47
rect 914 21 944 47
rect 1019 21 1049 47
rect 1234 35 1264 61
<< polycont >>
rect 100 251 134 285
rect 528 337 562 371
rect 405 267 439 301
rect 405 199 439 233
rect 642 391 676 425
rect 750 395 784 429
rect 906 393 940 427
rect 642 323 676 357
rect 528 269 562 303
rect 714 199 748 233
rect 822 237 856 271
rect 822 169 856 203
rect 1008 267 1042 301
rect 1201 267 1235 301
rect 319 59 353 93
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 30 597 110 613
rect 30 563 67 597
rect 101 563 110 597
rect 30 527 110 563
rect 30 493 67 527
rect 101 493 110 527
rect 30 373 110 493
rect 144 597 196 649
rect 144 563 153 597
rect 187 563 196 597
rect 144 527 196 563
rect 144 493 153 527
rect 187 493 196 527
rect 144 477 196 493
rect 230 597 454 615
rect 230 563 239 597
rect 273 581 454 597
rect 273 563 289 581
rect 230 527 289 563
rect 230 493 239 527
rect 273 493 289 527
rect 230 477 289 493
rect 346 531 386 547
rect 346 497 350 531
rect 384 497 386 531
rect 346 441 386 497
rect 420 509 454 581
rect 488 593 540 649
rect 488 559 490 593
rect 524 559 540 593
rect 488 543 540 559
rect 651 593 856 613
rect 651 559 667 593
rect 701 559 856 593
rect 651 543 856 559
rect 420 475 784 509
rect 346 425 692 441
rect 346 407 642 425
rect 626 391 642 407
rect 676 391 692 425
rect 30 371 578 373
rect 30 337 528 371
rect 562 337 578 371
rect 30 335 578 337
rect 30 201 66 335
rect 512 303 578 335
rect 626 357 692 391
rect 626 323 642 357
rect 676 323 692 357
rect 626 307 692 323
rect 734 429 784 475
rect 734 395 750 429
rect 100 285 355 301
rect 134 251 355 285
rect 100 235 355 251
rect 389 267 405 301
rect 439 267 455 301
rect 512 269 528 303
rect 562 269 578 303
rect 512 267 578 269
rect 389 233 455 267
rect 734 249 784 395
rect 818 357 856 543
rect 890 589 1038 649
rect 1173 607 1235 649
rect 890 555 996 589
rect 1030 555 1038 589
rect 890 540 1038 555
rect 924 521 1038 540
rect 924 506 996 521
rect 890 490 996 506
rect 990 487 996 490
rect 1030 487 1038 521
rect 990 461 1038 487
rect 1072 589 1132 605
rect 1072 555 1082 589
rect 1116 555 1132 589
rect 1072 493 1132 555
rect 1072 459 1082 493
rect 1116 459 1132 493
rect 890 427 956 443
rect 1072 427 1132 459
rect 890 393 906 427
rect 940 395 1132 427
rect 940 393 1082 395
rect 890 391 956 393
rect 1078 361 1082 393
rect 1116 361 1132 395
rect 1173 573 1189 607
rect 1223 573 1235 607
rect 1173 508 1235 573
rect 1173 474 1189 508
rect 1223 474 1235 508
rect 1173 413 1235 474
rect 1173 379 1189 413
rect 1223 379 1235 413
rect 1173 363 1235 379
rect 1269 599 1327 615
rect 1269 565 1275 599
rect 1309 565 1327 599
rect 1269 506 1327 565
rect 1269 472 1275 506
rect 1309 472 1327 506
rect 1269 413 1327 472
rect 1269 379 1275 413
rect 1309 379 1327 413
rect 818 323 1042 357
rect 892 301 1042 323
rect 698 233 784 249
rect 389 201 405 233
rect 30 185 110 201
rect 30 151 67 185
rect 101 151 110 185
rect 30 135 110 151
rect 144 185 189 201
rect 144 151 153 185
rect 187 151 189 185
rect 223 199 405 201
rect 439 199 714 233
rect 748 199 784 233
rect 818 271 858 287
rect 818 237 822 271
rect 856 237 858 271
rect 818 203 858 237
rect 223 165 239 199
rect 273 165 455 199
rect 818 169 822 203
rect 856 169 858 203
rect 818 165 858 169
rect 223 162 455 165
rect 144 17 189 151
rect 491 131 858 165
rect 892 267 1008 301
rect 892 251 1042 267
rect 1078 317 1132 361
rect 1078 301 1235 317
rect 1078 267 1201 301
rect 1078 251 1235 267
rect 223 93 457 128
rect 223 59 319 93
rect 353 59 457 93
rect 491 109 529 131
rect 491 75 495 109
rect 491 59 529 75
rect 565 94 631 97
rect 565 60 581 94
rect 615 60 631 94
rect 892 93 926 251
rect 565 17 631 60
rect 745 89 926 93
rect 745 55 761 89
rect 795 55 926 89
rect 960 201 1022 217
rect 1078 215 1112 251
rect 960 167 974 201
rect 1008 167 1022 201
rect 960 93 1022 167
rect 960 59 968 93
rect 1002 59 1022 93
rect 960 17 1022 59
rect 1056 199 1112 215
rect 1056 165 1060 199
rect 1094 165 1112 199
rect 1056 101 1112 165
rect 1056 67 1060 101
rect 1094 67 1112 101
rect 1056 51 1112 67
rect 1173 201 1235 217
rect 1173 167 1189 201
rect 1223 167 1235 201
rect 1173 107 1235 167
rect 1173 73 1189 107
rect 1223 73 1235 107
rect 1173 17 1235 73
rect 1269 212 1327 379
rect 1269 178 1275 212
rect 1309 178 1327 212
rect 1269 107 1327 178
rect 1269 73 1275 107
rect 1309 73 1327 107
rect 1269 57 1327 73
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlxtn_1
flabel comment s 763 327 763 327 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1279 94 1313 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 168 1313 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 464 1313 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 538 1313 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 626102
string GDS_START 614650
<< end >>
