magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
rect 427 319 901 331
<< pwell >>
rect 19 241 379 274
rect 19 49 1323 241
rect 0 0 1344 49
<< scnmos >>
rect 98 164 128 248
rect 270 164 300 248
rect 516 47 546 215
rect 602 47 632 215
rect 688 47 718 215
rect 774 47 804 215
rect 956 47 986 215
rect 1042 47 1072 215
rect 1128 47 1158 215
rect 1214 47 1244 215
<< scpmoshvt >>
rect 102 512 132 596
rect 256 512 286 596
rect 516 355 546 607
rect 602 355 632 607
rect 688 355 718 607
rect 782 355 812 607
rect 972 367 1002 619
rect 1058 367 1088 619
rect 1144 367 1174 619
rect 1230 367 1260 619
<< ndiff >>
rect 45 223 98 248
rect 45 189 53 223
rect 87 189 98 223
rect 45 164 98 189
rect 128 209 270 248
rect 128 175 141 209
rect 175 175 270 209
rect 128 164 270 175
rect 300 236 353 248
rect 300 202 311 236
rect 345 202 353 236
rect 300 164 353 202
rect 463 93 516 215
rect 463 59 471 93
rect 505 59 516 93
rect 463 47 516 59
rect 546 207 602 215
rect 546 173 557 207
rect 591 173 602 207
rect 546 101 602 173
rect 546 67 557 101
rect 591 67 602 101
rect 546 47 602 67
rect 632 165 688 215
rect 632 131 643 165
rect 677 131 688 165
rect 632 89 688 131
rect 632 55 643 89
rect 677 55 688 89
rect 632 47 688 55
rect 718 203 774 215
rect 718 169 729 203
rect 763 169 774 203
rect 718 101 774 169
rect 718 67 729 101
rect 763 67 774 101
rect 718 47 774 67
rect 804 126 956 215
rect 804 92 815 126
rect 849 92 911 126
rect 945 92 956 126
rect 804 47 956 92
rect 986 203 1042 215
rect 986 169 997 203
rect 1031 169 1042 203
rect 986 101 1042 169
rect 986 67 997 101
rect 1031 67 1042 101
rect 986 47 1042 67
rect 1072 177 1128 215
rect 1072 143 1083 177
rect 1117 143 1128 177
rect 1072 93 1128 143
rect 1072 59 1083 93
rect 1117 59 1128 93
rect 1072 47 1128 59
rect 1158 203 1214 215
rect 1158 169 1169 203
rect 1203 169 1214 203
rect 1158 101 1214 169
rect 1158 67 1169 101
rect 1203 67 1214 101
rect 1158 47 1214 67
rect 1244 203 1297 215
rect 1244 169 1255 203
rect 1289 169 1297 203
rect 1244 93 1297 169
rect 1244 59 1255 93
rect 1289 59 1297 93
rect 1244 47 1297 59
<< pdiff >>
rect 49 571 102 596
rect 49 537 57 571
rect 91 537 102 571
rect 49 512 102 537
rect 132 574 256 596
rect 132 540 143 574
rect 177 540 211 574
rect 245 540 256 574
rect 132 512 256 540
rect 286 584 355 596
rect 286 550 297 584
rect 331 550 355 584
rect 286 512 355 550
rect 463 595 516 607
rect 463 561 471 595
rect 505 561 516 595
rect 463 503 516 561
rect 463 469 471 503
rect 505 469 516 503
rect 463 401 516 469
rect 463 367 471 401
rect 505 367 516 401
rect 463 355 516 367
rect 546 547 602 607
rect 546 513 557 547
rect 591 513 602 547
rect 546 477 602 513
rect 546 443 557 477
rect 591 443 602 477
rect 546 401 602 443
rect 546 367 557 401
rect 591 367 602 401
rect 546 355 602 367
rect 632 593 688 607
rect 632 559 643 593
rect 677 559 688 593
rect 632 525 688 559
rect 632 491 643 525
rect 677 491 688 525
rect 632 453 688 491
rect 632 419 643 453
rect 677 419 688 453
rect 632 355 688 419
rect 718 595 782 607
rect 718 561 733 595
rect 767 561 782 595
rect 718 509 782 561
rect 718 475 733 509
rect 767 475 782 509
rect 718 355 782 475
rect 812 531 865 607
rect 812 497 823 531
rect 857 497 865 531
rect 812 453 865 497
rect 812 419 823 453
rect 857 419 865 453
rect 812 355 865 419
rect 919 531 972 619
rect 919 497 927 531
rect 961 497 972 531
rect 919 413 972 497
rect 919 379 927 413
rect 961 379 972 413
rect 919 367 972 379
rect 1002 599 1058 619
rect 1002 565 1013 599
rect 1047 565 1058 599
rect 1002 522 1058 565
rect 1002 488 1013 522
rect 1047 488 1058 522
rect 1002 439 1058 488
rect 1002 405 1013 439
rect 1047 405 1058 439
rect 1002 367 1058 405
rect 1088 599 1144 619
rect 1088 565 1099 599
rect 1133 565 1144 599
rect 1088 504 1144 565
rect 1088 470 1099 504
rect 1133 470 1144 504
rect 1088 413 1144 470
rect 1088 379 1099 413
rect 1133 379 1144 413
rect 1088 367 1144 379
rect 1174 607 1230 619
rect 1174 573 1185 607
rect 1219 573 1230 607
rect 1174 523 1230 573
rect 1174 489 1185 523
rect 1219 489 1230 523
rect 1174 439 1230 489
rect 1174 405 1185 439
rect 1219 405 1230 439
rect 1174 367 1230 405
rect 1260 599 1313 619
rect 1260 565 1271 599
rect 1305 565 1313 599
rect 1260 504 1313 565
rect 1260 470 1271 504
rect 1305 470 1313 504
rect 1260 413 1313 470
rect 1260 379 1271 413
rect 1305 379 1313 413
rect 1260 367 1313 379
<< ndiffc >>
rect 53 189 87 223
rect 141 175 175 209
rect 311 202 345 236
rect 471 59 505 93
rect 557 173 591 207
rect 557 67 591 101
rect 643 131 677 165
rect 643 55 677 89
rect 729 169 763 203
rect 729 67 763 101
rect 815 92 849 126
rect 911 92 945 126
rect 997 169 1031 203
rect 997 67 1031 101
rect 1083 143 1117 177
rect 1083 59 1117 93
rect 1169 169 1203 203
rect 1169 67 1203 101
rect 1255 169 1289 203
rect 1255 59 1289 93
<< pdiffc >>
rect 57 537 91 571
rect 143 540 177 574
rect 211 540 245 574
rect 297 550 331 584
rect 471 561 505 595
rect 471 469 505 503
rect 471 367 505 401
rect 557 513 591 547
rect 557 443 591 477
rect 557 367 591 401
rect 643 559 677 593
rect 643 491 677 525
rect 643 419 677 453
rect 733 561 767 595
rect 733 475 767 509
rect 823 497 857 531
rect 823 419 857 453
rect 927 497 961 531
rect 927 379 961 413
rect 1013 565 1047 599
rect 1013 488 1047 522
rect 1013 405 1047 439
rect 1099 565 1133 599
rect 1099 470 1133 504
rect 1099 379 1133 413
rect 1185 573 1219 607
rect 1185 489 1219 523
rect 1185 405 1219 439
rect 1271 565 1305 599
rect 1271 470 1305 504
rect 1271 379 1305 413
<< poly >>
rect 102 596 132 622
rect 256 596 286 622
rect 516 607 546 633
rect 602 607 632 633
rect 688 607 718 633
rect 782 607 812 633
rect 972 619 1002 645
rect 1058 619 1088 645
rect 1144 619 1174 645
rect 1230 619 1260 645
rect 102 450 132 512
rect 256 450 286 512
rect 98 434 177 450
rect 98 400 127 434
rect 161 400 177 434
rect 98 366 177 400
rect 98 332 127 366
rect 161 332 177 366
rect 98 316 177 332
rect 234 434 300 450
rect 234 400 250 434
rect 284 400 300 434
rect 234 366 300 400
rect 234 332 250 366
rect 284 332 300 366
rect 234 316 300 332
rect 98 248 128 316
rect 270 248 300 316
rect 375 304 441 320
rect 375 270 391 304
rect 425 270 441 304
rect 375 267 441 270
rect 516 267 546 355
rect 602 267 632 355
rect 688 317 718 355
rect 782 317 812 355
rect 972 345 1002 367
rect 1058 345 1088 367
rect 375 237 632 267
rect 674 301 812 317
rect 940 315 1002 345
rect 1050 315 1088 345
rect 940 303 1086 315
rect 674 267 715 301
rect 749 267 812 301
rect 674 251 812 267
rect 891 287 1086 303
rect 891 253 907 287
rect 941 253 1086 287
rect 1144 303 1174 367
rect 1230 303 1260 367
rect 1144 287 1296 303
rect 1144 267 1246 287
rect 375 236 441 237
rect 375 202 391 236
rect 425 202 441 236
rect 516 215 546 237
rect 602 215 632 237
rect 688 215 718 251
rect 774 215 804 251
rect 891 237 1086 253
rect 1128 253 1246 267
rect 1280 253 1296 287
rect 1128 237 1296 253
rect 956 215 986 237
rect 1042 215 1072 237
rect 1128 215 1158 237
rect 1214 215 1244 237
rect 375 186 441 202
rect 98 138 128 164
rect 270 138 300 164
rect 516 21 546 47
rect 602 21 632 47
rect 688 21 718 47
rect 774 21 804 47
rect 956 21 986 47
rect 1042 21 1072 47
rect 1128 21 1158 47
rect 1214 21 1244 47
<< polycont >>
rect 127 400 161 434
rect 127 332 161 366
rect 250 400 284 434
rect 250 332 284 366
rect 391 270 425 304
rect 715 267 749 301
rect 907 253 941 287
rect 391 202 425 236
rect 1246 253 1280 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 37 571 93 587
rect 37 537 57 571
rect 91 537 93 571
rect 37 521 93 537
rect 127 574 261 649
rect 127 540 143 574
rect 177 540 211 574
rect 245 540 261 574
rect 127 534 261 540
rect 295 584 395 600
rect 295 550 297 584
rect 331 550 395 584
rect 295 534 395 550
rect 37 282 87 521
rect 121 434 177 450
rect 121 400 127 434
rect 161 400 177 434
rect 121 366 177 400
rect 121 332 127 366
rect 161 332 177 366
rect 121 316 177 332
rect 211 434 284 500
rect 211 400 250 434
rect 211 366 284 400
rect 211 332 250 366
rect 211 316 284 332
rect 361 320 395 534
rect 455 595 683 615
rect 455 561 471 595
rect 505 593 683 595
rect 505 581 643 593
rect 505 561 507 581
rect 455 503 507 561
rect 641 559 643 581
rect 677 559 683 593
rect 455 469 471 503
rect 505 469 507 503
rect 455 401 507 469
rect 455 367 471 401
rect 505 367 507 401
rect 455 351 507 367
rect 541 513 557 547
rect 591 513 607 547
rect 541 477 607 513
rect 541 443 557 477
rect 591 443 607 477
rect 541 401 607 443
rect 641 525 683 559
rect 641 491 643 525
rect 677 491 683 525
rect 641 453 683 491
rect 717 599 1063 615
rect 717 595 1013 599
rect 717 561 733 595
rect 767 581 1013 595
rect 767 561 783 581
rect 717 509 783 561
rect 997 565 1013 581
rect 1047 565 1063 599
rect 717 475 733 509
rect 767 475 783 509
rect 717 471 783 475
rect 817 531 873 547
rect 817 497 823 531
rect 857 497 873 531
rect 641 419 643 453
rect 677 437 683 453
rect 817 453 873 497
rect 817 437 823 453
rect 677 419 823 437
rect 857 419 873 453
rect 641 403 873 419
rect 911 531 963 547
rect 911 497 927 531
rect 961 497 963 531
rect 911 413 963 497
rect 541 367 557 401
rect 591 369 607 401
rect 911 379 927 413
rect 961 379 963 413
rect 997 522 1063 565
rect 997 488 1013 522
rect 1047 488 1063 522
rect 997 439 1063 488
rect 997 405 1013 439
rect 1047 405 1063 439
rect 1097 599 1135 615
rect 1097 565 1099 599
rect 1133 565 1135 599
rect 1097 504 1135 565
rect 1097 470 1099 504
rect 1133 470 1135 504
rect 1097 413 1135 470
rect 911 371 963 379
rect 1097 379 1099 413
rect 1133 379 1135 413
rect 1169 607 1235 649
rect 1169 573 1185 607
rect 1219 573 1235 607
rect 1169 523 1235 573
rect 1169 489 1185 523
rect 1219 489 1235 523
rect 1169 439 1235 489
rect 1169 405 1185 439
rect 1219 405 1235 439
rect 1269 599 1321 615
rect 1269 565 1271 599
rect 1305 565 1321 599
rect 1269 504 1321 565
rect 1269 470 1271 504
rect 1305 470 1321 504
rect 1269 413 1321 470
rect 1097 371 1135 379
rect 1269 379 1271 413
rect 1305 379 1321 413
rect 1269 371 1321 379
rect 591 367 846 369
rect 541 335 846 367
rect 911 337 1321 371
rect 361 304 441 320
rect 37 248 259 282
rect 361 270 391 304
rect 425 270 441 304
rect 361 252 441 270
rect 37 223 87 248
rect 37 189 53 223
rect 37 173 87 189
rect 123 209 191 214
rect 123 175 141 209
rect 175 175 191 209
rect 123 17 191 175
rect 225 166 259 248
rect 295 236 441 252
rect 295 202 311 236
rect 345 202 391 236
rect 425 202 441 236
rect 295 200 441 202
rect 477 267 715 301
rect 749 267 765 301
rect 477 166 511 267
rect 799 233 846 335
rect 880 287 943 303
rect 880 253 907 287
rect 941 253 943 287
rect 880 237 943 253
rect 1239 287 1327 303
rect 1239 253 1246 287
rect 1280 253 1327 287
rect 225 132 511 166
rect 555 207 846 233
rect 555 173 557 207
rect 591 203 846 207
rect 977 213 1205 247
rect 1239 237 1327 253
rect 977 203 1033 213
rect 591 199 729 203
rect 591 173 593 199
rect 555 101 593 173
rect 727 169 729 199
rect 763 169 997 203
rect 1031 169 1033 203
rect 1167 203 1205 213
rect 727 168 1033 169
rect 455 93 521 98
rect 455 59 471 93
rect 505 59 521 93
rect 455 17 521 59
rect 555 67 557 101
rect 591 67 593 101
rect 555 51 593 67
rect 627 131 643 165
rect 677 131 693 165
rect 627 89 693 131
rect 627 55 643 89
rect 677 55 693 89
rect 627 17 693 55
rect 727 101 765 168
rect 727 67 729 101
rect 763 67 765 101
rect 727 51 765 67
rect 799 126 961 134
rect 799 92 815 126
rect 849 92 911 126
rect 945 92 961 126
rect 799 17 961 92
rect 995 101 1033 168
rect 995 67 997 101
rect 1031 67 1033 101
rect 995 51 1033 67
rect 1067 143 1083 177
rect 1117 143 1133 177
rect 1067 93 1133 143
rect 1067 59 1083 93
rect 1117 59 1133 93
rect 1067 17 1133 59
rect 1167 169 1169 203
rect 1203 169 1205 203
rect 1167 101 1205 169
rect 1167 67 1169 101
rect 1203 67 1205 101
rect 1167 51 1205 67
rect 1239 169 1255 203
rect 1289 169 1305 203
rect 1239 93 1305 169
rect 1239 59 1255 93
rect 1289 59 1305 93
rect 1239 17 1305 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4bb_2
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3396978
string GDS_START 3385662
<< end >>
