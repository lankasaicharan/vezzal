magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 768 210 957 248
rect 6 49 957 210
rect 0 0 960 49
<< scnmos >>
rect 89 74 119 184
rect 203 74 233 184
rect 413 74 443 184
rect 510 74 540 184
rect 623 74 653 184
rect 723 74 753 184
rect 844 74 874 222
<< scpmoshvt >>
rect 86 424 116 592
rect 186 424 216 592
rect 416 378 446 578
rect 500 378 530 578
rect 596 378 626 578
rect 704 378 734 578
rect 821 368 851 592
<< ndiff >>
rect 794 184 844 222
rect 32 146 89 184
rect 32 112 44 146
rect 78 112 89 146
rect 32 74 89 112
rect 119 131 203 184
rect 119 97 144 131
rect 178 97 203 131
rect 119 74 203 97
rect 233 140 290 184
rect 233 106 244 140
rect 278 106 290 140
rect 233 74 290 106
rect 353 120 413 184
rect 353 86 365 120
rect 399 86 413 120
rect 353 74 413 86
rect 443 146 510 184
rect 443 112 465 146
rect 499 112 510 146
rect 443 74 510 112
rect 540 120 623 184
rect 540 86 571 120
rect 605 86 623 120
rect 540 74 623 86
rect 653 146 723 184
rect 653 112 678 146
rect 712 112 723 146
rect 653 74 723 112
rect 753 136 844 184
rect 753 102 778 136
rect 812 102 844 136
rect 753 74 844 102
rect 874 210 931 222
rect 874 176 885 210
rect 919 176 931 210
rect 874 120 931 176
rect 874 86 885 120
rect 919 86 931 120
rect 874 74 931 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 470 86 546
rect 27 436 39 470
rect 73 436 86 470
rect 27 424 86 436
rect 116 580 186 592
rect 116 546 139 580
rect 173 546 186 580
rect 116 424 186 546
rect 216 428 303 592
rect 752 580 821 592
rect 752 578 764 580
rect 216 424 251 428
rect 234 394 251 424
rect 285 394 303 428
rect 234 382 303 394
rect 357 531 416 578
rect 357 497 369 531
rect 403 497 416 531
rect 357 424 416 497
rect 357 390 369 424
rect 403 390 416 424
rect 357 378 416 390
rect 446 378 500 578
rect 530 378 596 578
rect 626 378 704 578
rect 734 546 764 578
rect 798 546 821 580
rect 734 510 821 546
rect 734 476 764 510
rect 798 476 821 510
rect 734 440 821 476
rect 734 406 764 440
rect 798 406 821 440
rect 734 378 821 406
rect 768 368 821 378
rect 851 580 910 592
rect 851 546 864 580
rect 898 546 910 580
rect 851 497 910 546
rect 851 463 864 497
rect 898 463 910 497
rect 851 414 910 463
rect 851 380 864 414
rect 898 380 910 414
rect 851 368 910 380
<< ndiffc >>
rect 44 112 78 146
rect 144 97 178 131
rect 244 106 278 140
rect 365 86 399 120
rect 465 112 499 146
rect 571 86 605 120
rect 678 112 712 146
rect 778 102 812 136
rect 885 176 919 210
rect 885 86 919 120
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 139 546 173 580
rect 251 394 285 428
rect 369 497 403 531
rect 369 390 403 424
rect 764 546 798 580
rect 764 476 798 510
rect 764 406 798 440
rect 864 546 898 580
rect 864 463 898 497
rect 864 380 898 414
<< poly >>
rect 86 592 116 618
rect 186 592 216 618
rect 416 578 446 604
rect 500 578 530 604
rect 596 578 626 604
rect 704 578 734 604
rect 821 592 851 618
rect 86 409 116 424
rect 186 409 216 424
rect 83 326 119 409
rect 25 310 119 326
rect 25 276 41 310
rect 75 276 119 310
rect 25 260 119 276
rect 89 184 119 260
rect 183 344 219 409
rect 416 363 446 378
rect 500 363 530 378
rect 596 363 626 378
rect 704 363 734 378
rect 183 328 259 344
rect 413 340 449 363
rect 183 294 209 328
rect 243 294 259 328
rect 183 260 259 294
rect 183 226 209 260
rect 243 226 259 260
rect 183 210 259 226
rect 315 332 449 340
rect 315 324 443 332
rect 315 290 331 324
rect 365 290 443 324
rect 497 304 533 363
rect 593 336 629 363
rect 701 336 737 363
rect 821 353 851 368
rect 593 320 659 336
rect 315 256 443 290
rect 315 222 331 256
rect 365 222 443 256
rect 485 288 551 304
rect 485 254 501 288
rect 535 254 551 288
rect 593 286 609 320
rect 643 286 659 320
rect 593 270 659 286
rect 701 320 767 336
rect 818 326 854 353
rect 701 286 717 320
rect 751 286 767 320
rect 701 270 767 286
rect 809 310 875 326
rect 809 276 825 310
rect 859 276 875 310
rect 485 238 551 254
rect 203 184 233 210
rect 315 206 443 222
rect 413 184 443 206
rect 510 184 540 238
rect 623 184 653 270
rect 723 184 753 270
rect 809 260 875 276
rect 844 222 874 260
rect 89 48 119 74
rect 203 48 233 74
rect 413 48 443 74
rect 510 48 540 74
rect 623 48 653 74
rect 723 48 753 74
rect 844 48 874 74
<< polycont >>
rect 41 276 75 310
rect 209 294 243 328
rect 209 226 243 260
rect 331 290 365 324
rect 331 222 365 256
rect 501 254 535 288
rect 609 286 643 320
rect 717 286 751 320
rect 825 276 859 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 496 89 546
rect 123 580 189 649
rect 123 546 139 580
rect 173 546 189 580
rect 123 530 189 546
rect 223 581 551 615
rect 223 496 257 581
rect 23 470 257 496
rect 23 436 39 470
rect 73 462 257 470
rect 369 531 449 547
rect 403 497 449 531
rect 73 436 159 462
rect 23 420 159 436
rect 25 310 91 356
rect 25 276 41 310
rect 75 276 91 310
rect 25 260 91 276
rect 125 226 159 420
rect 230 394 251 428
rect 285 394 331 428
rect 230 378 331 394
rect 28 192 159 226
rect 193 328 263 344
rect 193 294 209 328
rect 243 294 263 328
rect 193 260 263 294
rect 193 226 209 260
rect 243 226 263 260
rect 193 210 263 226
rect 297 340 331 378
rect 369 424 449 497
rect 403 390 449 424
rect 369 374 449 390
rect 297 324 381 340
rect 297 290 331 324
rect 365 290 381 324
rect 297 256 381 290
rect 297 222 331 256
rect 365 222 381 256
rect 297 206 381 222
rect 28 146 94 192
rect 297 176 331 206
rect 28 112 44 146
rect 78 112 94 146
rect 28 70 94 112
rect 128 131 194 158
rect 128 97 144 131
rect 178 97 194 131
rect 128 17 194 97
rect 228 140 331 176
rect 415 204 449 374
rect 485 288 551 581
rect 748 580 814 649
rect 485 254 501 288
rect 535 254 551 288
rect 593 320 659 578
rect 748 546 764 580
rect 798 546 814 580
rect 748 510 814 546
rect 748 476 764 510
rect 798 476 814 510
rect 748 440 814 476
rect 748 406 764 440
rect 798 406 814 440
rect 748 390 814 406
rect 848 580 943 596
rect 848 546 864 580
rect 898 546 943 580
rect 848 497 943 546
rect 848 463 864 497
rect 898 463 943 497
rect 848 414 943 463
rect 848 380 864 414
rect 898 380 943 414
rect 848 364 943 380
rect 593 286 609 320
rect 643 286 659 320
rect 593 270 659 286
rect 697 320 767 356
rect 697 286 717 320
rect 751 286 767 320
rect 697 270 767 286
rect 801 310 875 326
rect 801 276 825 310
rect 859 276 875 310
rect 485 238 551 254
rect 801 260 875 276
rect 801 236 835 260
rect 662 204 835 236
rect 909 226 943 364
rect 415 202 835 204
rect 869 210 943 226
rect 415 170 728 202
rect 228 106 244 140
rect 278 106 331 140
rect 449 146 515 170
rect 228 70 331 106
rect 365 120 415 136
rect 399 86 415 120
rect 365 17 415 86
rect 449 112 465 146
rect 499 112 515 146
rect 662 146 728 170
rect 869 176 885 210
rect 919 176 943 210
rect 449 70 515 112
rect 549 120 628 136
rect 549 86 571 120
rect 605 86 628 120
rect 549 17 628 86
rect 662 112 678 146
rect 712 112 728 146
rect 662 70 728 112
rect 762 136 828 168
rect 762 102 778 136
rect 812 102 828 136
rect 762 17 828 102
rect 869 120 943 176
rect 869 86 885 120
rect 919 86 943 120
rect 869 70 943 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or4bb_1
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 94 929 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 3861602
string GDS_START 3853266
<< end >>
