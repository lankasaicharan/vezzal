magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 191 245 1009 259
rect 1 49 1009 245
rect 0 0 1056 49
<< scnmos >>
rect 80 51 110 219
rect 270 65 300 233
rect 356 65 386 233
rect 456 65 486 233
rect 556 65 586 233
rect 642 65 672 233
rect 728 65 758 233
rect 814 65 844 233
rect 900 65 930 233
<< scpmoshvt >>
rect 80 367 110 619
rect 254 367 284 619
rect 340 367 370 619
rect 442 367 472 619
rect 528 367 558 619
rect 642 367 672 619
rect 740 367 770 619
rect 826 367 856 619
rect 912 367 942 619
<< ndiff >>
rect 217 221 270 233
rect 27 207 80 219
rect 27 173 35 207
rect 69 173 80 207
rect 27 101 80 173
rect 27 67 35 101
rect 69 67 80 101
rect 27 51 80 67
rect 110 171 163 219
rect 110 137 121 171
rect 155 137 163 171
rect 110 97 163 137
rect 110 63 121 97
rect 155 63 163 97
rect 217 187 225 221
rect 259 187 270 221
rect 217 111 270 187
rect 217 77 225 111
rect 259 77 270 111
rect 217 65 270 77
rect 300 225 356 233
rect 300 191 311 225
rect 345 191 356 225
rect 300 155 356 191
rect 300 121 311 155
rect 345 121 356 155
rect 300 65 356 121
rect 386 183 456 233
rect 386 149 411 183
rect 445 149 456 183
rect 386 107 456 149
rect 386 73 411 107
rect 445 73 456 107
rect 386 65 456 73
rect 486 225 556 233
rect 486 191 511 225
rect 545 191 556 225
rect 486 155 556 191
rect 486 121 511 155
rect 545 121 556 155
rect 486 65 556 121
rect 586 225 642 233
rect 586 191 597 225
rect 631 191 642 225
rect 586 107 642 191
rect 586 73 597 107
rect 631 73 642 107
rect 586 65 642 73
rect 672 183 728 233
rect 672 149 683 183
rect 717 149 728 183
rect 672 107 728 149
rect 672 73 683 107
rect 717 73 728 107
rect 672 65 728 73
rect 758 221 814 233
rect 758 187 769 221
rect 803 187 814 221
rect 758 107 814 187
rect 758 73 769 107
rect 803 73 814 107
rect 758 65 814 73
rect 844 181 900 233
rect 844 147 855 181
rect 889 147 900 181
rect 844 107 900 147
rect 844 73 855 107
rect 889 73 900 107
rect 844 65 900 73
rect 930 221 983 233
rect 930 187 941 221
rect 975 187 983 221
rect 930 111 983 187
rect 930 77 941 111
rect 975 77 983 111
rect 930 65 983 77
rect 110 51 163 63
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 519 80 565
rect 27 485 35 519
rect 69 485 80 519
rect 27 436 80 485
rect 27 402 35 436
rect 69 402 80 436
rect 27 367 80 402
rect 110 607 254 619
rect 110 573 121 607
rect 155 573 209 607
rect 243 573 254 607
rect 110 506 254 573
rect 110 488 209 506
rect 110 454 121 488
rect 155 472 209 488
rect 243 472 254 506
rect 155 454 254 472
rect 110 410 254 454
rect 110 376 209 410
rect 243 376 254 410
rect 110 367 254 376
rect 284 599 340 619
rect 284 565 295 599
rect 329 565 340 599
rect 284 506 340 565
rect 284 472 295 506
rect 329 472 340 506
rect 284 410 340 472
rect 284 376 295 410
rect 329 376 340 410
rect 284 367 340 376
rect 370 611 442 619
rect 370 577 389 611
rect 423 577 442 611
rect 370 533 442 577
rect 370 499 389 533
rect 423 499 442 533
rect 370 455 442 499
rect 370 421 389 455
rect 423 421 442 455
rect 370 367 442 421
rect 472 599 528 619
rect 472 565 483 599
rect 517 565 528 599
rect 472 506 528 565
rect 472 472 483 506
rect 517 472 528 506
rect 472 410 528 472
rect 472 376 483 410
rect 517 376 528 410
rect 472 367 528 376
rect 558 611 642 619
rect 558 577 583 611
rect 617 577 642 611
rect 558 492 642 577
rect 558 458 583 492
rect 617 458 642 492
rect 558 367 642 458
rect 672 599 740 619
rect 672 565 688 599
rect 722 565 740 599
rect 672 513 740 565
rect 672 479 688 513
rect 722 479 740 513
rect 672 436 740 479
rect 672 402 688 436
rect 722 402 740 436
rect 672 367 740 402
rect 770 607 826 619
rect 770 573 781 607
rect 815 573 826 607
rect 770 504 826 573
rect 770 470 781 504
rect 815 470 826 504
rect 770 367 826 470
rect 856 599 912 619
rect 856 565 867 599
rect 901 565 912 599
rect 856 517 912 565
rect 856 483 867 517
rect 901 483 912 517
rect 856 436 912 483
rect 856 402 867 436
rect 901 402 912 436
rect 856 367 912 402
rect 942 607 995 619
rect 942 573 953 607
rect 987 573 995 607
rect 942 515 995 573
rect 942 481 953 515
rect 987 481 995 515
rect 942 420 995 481
rect 942 386 953 420
rect 987 386 995 420
rect 942 367 995 386
<< ndiffc >>
rect 35 173 69 207
rect 35 67 69 101
rect 121 137 155 171
rect 121 63 155 97
rect 225 187 259 221
rect 225 77 259 111
rect 311 191 345 225
rect 311 121 345 155
rect 411 149 445 183
rect 411 73 445 107
rect 511 191 545 225
rect 511 121 545 155
rect 597 191 631 225
rect 597 73 631 107
rect 683 149 717 183
rect 683 73 717 107
rect 769 187 803 221
rect 769 73 803 107
rect 855 147 889 181
rect 855 73 889 107
rect 941 187 975 221
rect 941 77 975 111
<< pdiffc >>
rect 35 565 69 599
rect 35 485 69 519
rect 35 402 69 436
rect 121 573 155 607
rect 209 573 243 607
rect 121 454 155 488
rect 209 472 243 506
rect 209 376 243 410
rect 295 565 329 599
rect 295 472 329 506
rect 295 376 329 410
rect 389 577 423 611
rect 389 499 423 533
rect 389 421 423 455
rect 483 565 517 599
rect 483 472 517 506
rect 483 376 517 410
rect 583 577 617 611
rect 583 458 617 492
rect 688 565 722 599
rect 688 479 722 513
rect 688 402 722 436
rect 781 573 815 607
rect 781 470 815 504
rect 867 565 901 599
rect 867 483 901 517
rect 867 402 901 436
rect 953 573 987 607
rect 953 481 987 515
rect 953 386 987 420
<< poly >>
rect 80 619 110 645
rect 254 619 284 645
rect 340 619 370 645
rect 442 619 472 645
rect 528 619 558 645
rect 642 619 672 645
rect 740 619 770 645
rect 826 619 856 645
rect 912 619 942 645
rect 80 325 110 367
rect 254 335 284 367
rect 340 335 370 367
rect 442 335 472 367
rect 528 335 558 367
rect 642 335 672 367
rect 740 335 770 367
rect 826 335 856 367
rect 912 335 942 367
rect 33 309 110 325
rect 33 275 49 309
rect 83 275 110 309
rect 33 259 110 275
rect 152 319 586 335
rect 152 285 168 319
rect 202 285 236 319
rect 270 285 304 319
rect 338 285 372 319
rect 406 285 440 319
rect 474 285 586 319
rect 152 269 586 285
rect 80 219 110 259
rect 270 233 300 269
rect 356 233 386 269
rect 456 233 486 269
rect 556 233 586 269
rect 642 319 988 335
rect 642 285 666 319
rect 700 285 734 319
rect 768 285 802 319
rect 836 285 870 319
rect 904 285 938 319
rect 972 285 988 319
rect 642 269 988 285
rect 642 233 672 269
rect 728 233 758 269
rect 814 233 844 269
rect 900 233 930 269
rect 80 25 110 51
rect 270 39 300 65
rect 356 39 386 65
rect 456 39 486 65
rect 556 39 586 65
rect 642 39 672 65
rect 728 39 758 65
rect 814 39 844 65
rect 900 39 930 65
<< polycont >>
rect 49 275 83 309
rect 168 285 202 319
rect 236 285 270 319
rect 304 285 338 319
rect 372 285 406 319
rect 440 285 474 319
rect 666 285 700 319
rect 734 285 768 319
rect 802 285 836 319
rect 870 285 904 319
rect 938 285 972 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 19 599 71 615
rect 19 565 35 599
rect 69 565 71 599
rect 19 519 71 565
rect 19 485 35 519
rect 69 485 71 519
rect 19 436 71 485
rect 105 607 253 649
rect 105 573 121 607
rect 155 573 209 607
rect 243 573 253 607
rect 105 506 253 573
rect 105 488 209 506
rect 105 454 121 488
rect 155 472 209 488
rect 243 472 253 506
rect 155 454 253 472
rect 19 402 35 436
rect 69 420 71 436
rect 69 402 167 420
rect 19 386 167 402
rect 31 309 99 352
rect 31 275 49 309
rect 83 275 99 309
rect 31 273 99 275
rect 133 319 167 386
rect 201 410 253 454
rect 201 376 209 410
rect 243 376 253 410
rect 201 360 253 376
rect 287 599 339 615
rect 287 565 295 599
rect 329 565 339 599
rect 287 506 339 565
rect 287 472 295 506
rect 329 472 339 506
rect 287 410 339 472
rect 373 611 439 649
rect 373 577 389 611
rect 423 577 439 611
rect 373 533 439 577
rect 373 499 389 533
rect 423 499 439 533
rect 373 455 439 499
rect 373 421 389 455
rect 423 421 439 455
rect 473 599 533 615
rect 473 565 483 599
rect 517 565 533 599
rect 473 506 533 565
rect 473 472 483 506
rect 517 472 533 506
rect 473 424 533 472
rect 567 611 633 649
rect 567 577 583 611
rect 617 577 633 611
rect 567 492 633 577
rect 567 458 583 492
rect 617 458 633 492
rect 672 599 738 615
rect 672 565 688 599
rect 722 565 738 599
rect 672 513 738 565
rect 672 479 688 513
rect 722 479 738 513
rect 672 436 738 479
rect 772 607 825 649
rect 772 573 781 607
rect 815 573 825 607
rect 772 504 825 573
rect 772 470 781 504
rect 815 470 825 504
rect 772 454 825 470
rect 859 599 903 615
rect 859 565 867 599
rect 901 565 903 599
rect 859 517 903 565
rect 859 483 867 517
rect 901 483 903 517
rect 672 424 688 436
rect 287 376 295 410
rect 329 387 339 410
rect 473 410 688 424
rect 473 387 483 410
rect 329 376 483 387
rect 517 402 688 410
rect 722 420 738 436
rect 859 436 903 483
rect 859 420 867 436
rect 722 402 867 420
rect 901 402 903 436
rect 517 386 903 402
rect 937 607 1003 649
rect 937 573 953 607
rect 987 573 1003 607
rect 937 515 1003 573
rect 937 481 953 515
rect 987 481 1003 515
rect 937 420 1003 481
rect 937 386 953 420
rect 987 386 1003 420
rect 517 376 616 386
rect 287 353 616 376
rect 133 285 168 319
rect 202 285 236 319
rect 270 285 304 319
rect 338 285 372 319
rect 406 285 440 319
rect 474 285 490 319
rect 524 288 616 353
rect 650 319 1036 352
rect 133 239 167 285
rect 524 251 561 288
rect 650 285 666 319
rect 700 285 734 319
rect 768 285 802 319
rect 836 285 870 319
rect 904 285 938 319
rect 972 285 1036 319
rect 19 207 167 239
rect 19 173 35 207
rect 69 205 167 207
rect 209 221 261 237
rect 19 101 69 173
rect 209 187 225 221
rect 259 187 261 221
rect 19 67 35 101
rect 19 51 69 67
rect 105 137 121 171
rect 155 137 171 171
rect 105 97 171 137
rect 105 63 121 97
rect 155 63 171 97
rect 105 17 171 63
rect 209 111 261 187
rect 295 225 561 251
rect 295 191 311 225
rect 345 217 511 225
rect 345 191 361 217
rect 295 155 361 191
rect 495 191 511 217
rect 545 191 561 225
rect 295 121 311 155
rect 345 121 361 155
rect 395 149 411 183
rect 445 149 461 183
rect 209 77 225 111
rect 259 85 261 111
rect 395 107 461 149
rect 495 155 561 191
rect 495 121 511 155
rect 545 121 561 155
rect 595 225 991 251
rect 595 191 597 225
rect 631 221 991 225
rect 631 217 769 221
rect 631 191 633 217
rect 395 85 411 107
rect 259 77 411 85
rect 209 73 411 77
rect 445 85 461 107
rect 595 107 633 191
rect 767 187 769 217
rect 803 215 941 221
rect 803 187 805 215
rect 595 85 597 107
rect 445 73 597 85
rect 631 73 633 107
rect 209 51 633 73
rect 667 149 683 183
rect 717 149 733 183
rect 667 107 733 149
rect 667 73 683 107
rect 717 73 733 107
rect 667 17 733 73
rect 767 107 805 187
rect 939 187 941 215
rect 975 187 991 221
rect 767 73 769 107
rect 803 73 805 107
rect 767 57 805 73
rect 839 147 855 181
rect 889 147 905 181
rect 839 107 905 147
rect 839 73 855 107
rect 889 73 905 107
rect 839 17 905 73
rect 939 111 991 187
rect 939 77 941 111
rect 975 77 991 111
rect 939 61 991 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2b_4
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4440312
string GDS_START 4430774
<< end >>
