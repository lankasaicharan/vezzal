magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 2 49 849 157
rect 0 0 864 49
<< scnmos >>
rect 85 47 115 131
rect 157 47 187 131
rect 264 47 294 131
rect 342 47 372 131
rect 420 47 450 131
rect 506 47 536 131
rect 578 47 608 131
rect 664 47 694 131
rect 736 47 766 131
<< scpmoshvt >>
rect 101 414 151 614
rect 207 414 257 614
rect 313 414 363 614
rect 440 414 490 614
rect 546 414 596 614
rect 701 414 751 614
<< ndiff >>
rect 28 110 85 131
rect 28 76 40 110
rect 74 76 85 110
rect 28 47 85 76
rect 115 47 157 131
rect 187 105 264 131
rect 187 71 219 105
rect 253 71 264 105
rect 187 47 264 71
rect 294 47 342 131
rect 372 47 420 131
rect 450 111 506 131
rect 450 77 461 111
rect 495 77 506 111
rect 450 47 506 77
rect 536 47 578 131
rect 608 105 664 131
rect 608 71 619 105
rect 653 71 664 105
rect 608 47 664 71
rect 694 47 736 131
rect 766 111 823 131
rect 766 77 777 111
rect 811 77 823 111
rect 766 47 823 77
<< pdiff >>
rect 44 597 101 614
rect 44 563 56 597
rect 90 563 101 597
rect 44 528 101 563
rect 44 494 56 528
rect 90 494 101 528
rect 44 460 101 494
rect 44 426 56 460
rect 90 426 101 460
rect 44 414 101 426
rect 151 602 207 614
rect 151 568 162 602
rect 196 568 207 602
rect 151 531 207 568
rect 151 497 162 531
rect 196 497 207 531
rect 151 460 207 497
rect 151 426 162 460
rect 196 426 207 460
rect 151 414 207 426
rect 257 597 313 614
rect 257 563 268 597
rect 302 563 313 597
rect 257 528 313 563
rect 257 494 268 528
rect 302 494 313 528
rect 257 460 313 494
rect 257 426 268 460
rect 302 426 313 460
rect 257 414 313 426
rect 363 602 440 614
rect 363 568 374 602
rect 408 568 440 602
rect 363 530 440 568
rect 363 496 374 530
rect 408 496 440 530
rect 363 414 440 496
rect 490 597 546 614
rect 490 563 501 597
rect 535 563 546 597
rect 490 528 546 563
rect 490 494 501 528
rect 535 494 546 528
rect 490 460 546 494
rect 490 426 501 460
rect 535 426 546 460
rect 490 414 546 426
rect 596 414 701 614
rect 751 597 808 614
rect 751 563 762 597
rect 796 563 808 597
rect 751 528 808 563
rect 751 494 762 528
rect 796 494 808 528
rect 751 460 808 494
rect 751 426 762 460
rect 796 426 808 460
rect 751 414 808 426
<< ndiffc >>
rect 40 76 74 110
rect 219 71 253 105
rect 461 77 495 111
rect 619 71 653 105
rect 777 77 811 111
<< pdiffc >>
rect 56 563 90 597
rect 56 494 90 528
rect 56 426 90 460
rect 162 568 196 602
rect 162 497 196 531
rect 162 426 196 460
rect 268 563 302 597
rect 268 494 302 528
rect 268 426 302 460
rect 374 568 408 602
rect 374 496 408 530
rect 501 563 535 597
rect 501 494 535 528
rect 501 426 535 460
rect 762 563 796 597
rect 762 494 796 528
rect 762 426 796 460
<< poly >>
rect 101 614 151 640
rect 207 614 257 640
rect 313 614 363 640
rect 440 614 490 640
rect 546 614 596 640
rect 701 614 751 640
rect 101 352 151 414
rect 207 374 257 414
rect 313 374 363 414
rect 440 374 490 414
rect 199 358 265 374
rect 101 304 131 352
rect 199 324 215 358
rect 249 324 265 358
rect 85 288 157 304
rect 85 254 107 288
rect 141 254 157 288
rect 85 220 157 254
rect 199 290 265 324
rect 199 256 215 290
rect 249 256 265 290
rect 199 240 265 256
rect 307 358 373 374
rect 307 324 323 358
rect 357 324 373 358
rect 307 290 373 324
rect 307 256 323 290
rect 357 256 373 290
rect 307 240 373 256
rect 421 358 490 374
rect 421 324 437 358
rect 471 324 490 358
rect 421 290 490 324
rect 421 256 437 290
rect 471 256 490 290
rect 421 240 490 256
rect 546 382 596 414
rect 546 366 653 382
rect 546 332 603 366
rect 637 332 653 366
rect 546 298 653 332
rect 546 264 603 298
rect 637 264 653 298
rect 546 248 653 264
rect 701 374 751 414
rect 701 358 767 374
rect 701 324 717 358
rect 751 324 767 358
rect 701 290 767 324
rect 701 256 717 290
rect 751 256 767 290
rect 85 186 107 220
rect 141 192 157 220
rect 141 186 187 192
rect 85 162 187 186
rect 85 131 115 162
rect 157 131 187 162
rect 235 176 265 240
rect 235 146 294 176
rect 264 131 294 146
rect 342 131 372 240
rect 421 176 451 240
rect 546 176 576 248
rect 701 240 767 256
rect 701 176 731 240
rect 420 146 451 176
rect 506 146 608 176
rect 420 131 450 146
rect 506 131 536 146
rect 578 131 608 146
rect 664 146 766 176
rect 664 131 694 146
rect 736 131 766 146
rect 85 21 115 47
rect 157 21 187 47
rect 264 21 294 47
rect 342 21 372 47
rect 420 21 450 47
rect 506 21 536 47
rect 578 21 608 47
rect 664 21 694 47
rect 736 21 766 47
<< polycont >>
rect 215 324 249 358
rect 107 254 141 288
rect 215 256 249 290
rect 323 324 357 358
rect 323 256 357 290
rect 437 324 471 358
rect 437 256 471 290
rect 603 332 637 366
rect 603 264 637 298
rect 717 324 751 358
rect 717 256 751 290
rect 107 186 141 220
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 21 597 106 613
rect 21 563 56 597
rect 90 563 106 597
rect 21 528 106 563
rect 21 494 56 528
rect 90 494 106 528
rect 21 460 106 494
rect 21 426 56 460
rect 90 426 106 460
rect 21 410 106 426
rect 146 602 212 649
rect 146 568 162 602
rect 196 568 212 602
rect 146 531 212 568
rect 146 497 162 531
rect 196 497 212 531
rect 146 460 212 497
rect 146 426 162 460
rect 196 426 212 460
rect 146 410 212 426
rect 252 597 318 613
rect 252 563 268 597
rect 302 563 318 597
rect 252 528 318 563
rect 252 494 268 528
rect 302 494 318 528
rect 252 460 318 494
rect 358 602 424 649
rect 358 568 374 602
rect 408 568 424 602
rect 358 530 424 568
rect 358 496 374 530
rect 408 496 424 530
rect 358 480 424 496
rect 485 597 551 613
rect 485 563 501 597
rect 535 563 551 597
rect 746 597 837 613
rect 485 528 551 563
rect 485 494 501 528
rect 535 494 551 528
rect 252 426 268 460
rect 302 444 318 460
rect 485 460 551 494
rect 485 444 501 460
rect 302 426 501 444
rect 535 426 551 460
rect 252 410 551 426
rect 21 134 55 410
rect 199 358 265 374
rect 199 324 215 358
rect 249 324 265 358
rect 91 288 157 304
rect 91 254 107 288
rect 141 254 157 288
rect 91 220 157 254
rect 199 290 265 324
rect 199 256 215 290
rect 249 256 265 290
rect 199 240 265 256
rect 307 358 373 374
rect 307 324 323 358
rect 357 324 373 358
rect 307 290 373 324
rect 307 256 323 290
rect 357 256 373 290
rect 307 240 373 256
rect 409 358 551 374
rect 409 324 437 358
rect 471 324 551 358
rect 409 290 551 324
rect 409 256 437 290
rect 471 256 551 290
rect 409 240 551 256
rect 587 366 653 578
rect 746 563 762 597
rect 796 563 837 597
rect 746 528 837 563
rect 746 494 762 528
rect 796 494 837 528
rect 746 460 837 494
rect 746 426 762 460
rect 796 426 837 460
rect 746 410 837 426
rect 587 332 603 366
rect 637 332 653 366
rect 587 298 653 332
rect 587 264 603 298
rect 637 264 653 298
rect 587 248 653 264
rect 697 358 767 374
rect 697 324 717 358
rect 751 324 767 358
rect 697 290 767 324
rect 697 256 717 290
rect 751 256 767 290
rect 697 240 767 256
rect 91 186 107 220
rect 141 204 157 220
rect 803 204 837 410
rect 141 186 837 204
rect 91 170 837 186
rect 21 110 167 134
rect 21 76 40 110
rect 74 76 167 110
rect 21 53 167 76
rect 203 105 269 134
rect 203 71 219 105
rect 253 71 269 105
rect 203 17 269 71
rect 445 111 511 170
rect 445 77 461 111
rect 495 77 511 111
rect 445 53 511 77
rect 603 105 669 134
rect 603 71 619 105
rect 653 71 669 105
rect 603 17 669 71
rect 761 111 827 170
rect 761 77 777 111
rect 811 77 827 111
rect 761 53 827 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a311o_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3935262
string GDS_START 3927174
<< end >>
