magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1778 1975
<< nwell >>
rect -38 331 518 704
<< pwell >>
rect 14 49 472 157
rect 0 0 480 49
<< scnmos >>
rect 93 47 123 131
rect 171 47 201 131
rect 249 47 279 131
rect 363 47 393 131
<< scpmoshvt >>
rect 80 473 110 601
rect 166 473 196 601
rect 252 473 282 601
rect 338 473 368 601
<< ndiff >>
rect 40 103 93 131
rect 40 69 48 103
rect 82 69 93 103
rect 40 47 93 69
rect 123 47 171 131
rect 201 47 249 131
rect 279 106 363 131
rect 279 72 305 106
rect 339 72 363 106
rect 279 47 363 72
rect 393 106 446 131
rect 393 72 404 106
rect 438 72 446 106
rect 393 47 446 72
<< pdiff >>
rect 27 587 80 601
rect 27 553 35 587
rect 69 553 80 587
rect 27 519 80 553
rect 27 485 35 519
rect 69 485 80 519
rect 27 473 80 485
rect 110 589 166 601
rect 110 555 121 589
rect 155 555 166 589
rect 110 519 166 555
rect 110 485 121 519
rect 155 485 166 519
rect 110 473 166 485
rect 196 531 252 601
rect 196 497 207 531
rect 241 497 252 531
rect 196 473 252 497
rect 282 589 338 601
rect 282 555 293 589
rect 327 555 338 589
rect 282 519 338 555
rect 282 485 293 519
rect 327 485 338 519
rect 282 473 338 485
rect 368 589 421 601
rect 368 555 379 589
rect 413 555 421 589
rect 368 519 421 555
rect 368 485 379 519
rect 413 485 421 519
rect 368 473 421 485
<< ndiffc >>
rect 48 69 82 103
rect 305 72 339 106
rect 404 72 438 106
<< pdiffc >>
rect 35 553 69 587
rect 35 485 69 519
rect 121 555 155 589
rect 121 485 155 519
rect 207 497 241 531
rect 293 555 327 589
rect 293 485 327 519
rect 379 555 413 589
rect 379 485 413 519
<< poly >>
rect 80 601 110 627
rect 166 601 196 627
rect 252 601 282 627
rect 338 601 368 627
rect 80 443 110 473
rect 57 413 110 443
rect 57 325 87 413
rect 166 365 196 473
rect 21 309 87 325
rect 21 275 37 309
rect 71 275 87 309
rect 21 241 87 275
rect 21 207 37 241
rect 71 207 87 241
rect 135 349 201 365
rect 135 315 151 349
rect 185 315 201 349
rect 135 281 201 315
rect 252 302 282 473
rect 338 380 368 473
rect 338 350 393 380
rect 363 325 393 350
rect 363 309 455 325
rect 135 247 151 281
rect 185 247 201 281
rect 135 231 201 247
rect 21 191 87 207
rect 57 183 87 191
rect 57 153 123 183
rect 93 131 123 153
rect 171 131 201 231
rect 249 286 315 302
rect 249 252 265 286
rect 299 252 315 286
rect 249 218 315 252
rect 249 184 265 218
rect 299 184 315 218
rect 249 168 315 184
rect 363 275 405 309
rect 439 275 455 309
rect 363 241 455 275
rect 363 207 405 241
rect 439 207 455 241
rect 363 191 455 207
rect 249 131 279 168
rect 363 131 393 191
rect 93 21 123 47
rect 171 21 201 47
rect 249 21 279 47
rect 363 21 393 47
<< polycont >>
rect 37 275 71 309
rect 37 207 71 241
rect 151 315 185 349
rect 151 247 185 281
rect 265 252 299 286
rect 265 184 299 218
rect 405 275 439 309
rect 405 207 439 241
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 19 587 78 649
rect 19 553 35 587
rect 69 553 78 587
rect 19 519 78 553
rect 19 485 35 519
rect 69 485 78 519
rect 19 433 78 485
rect 112 589 335 615
rect 112 555 121 589
rect 155 581 293 589
rect 155 555 164 581
rect 112 519 164 555
rect 284 555 293 581
rect 327 555 335 589
rect 112 485 121 519
rect 155 485 164 519
rect 112 469 164 485
rect 198 531 250 547
rect 198 497 207 531
rect 241 497 250 531
rect 198 433 250 497
rect 284 519 335 555
rect 284 485 293 519
rect 327 485 335 519
rect 284 469 335 485
rect 369 589 463 605
rect 369 555 379 589
rect 413 555 463 589
rect 369 519 463 555
rect 369 485 379 519
rect 413 485 463 519
rect 369 435 463 485
rect 19 399 250 433
rect 335 390 463 435
rect 17 309 91 364
rect 17 275 37 309
rect 71 275 91 309
rect 17 241 91 275
rect 17 207 37 241
rect 71 207 91 241
rect 17 153 91 207
rect 125 349 185 365
rect 125 315 151 349
rect 125 281 185 315
rect 125 247 151 281
rect 25 103 91 119
rect 25 69 48 103
rect 82 69 91 103
rect 125 78 185 247
rect 219 286 301 365
rect 219 252 265 286
rect 299 252 301 286
rect 219 218 301 252
rect 219 184 265 218
rect 299 184 301 218
rect 219 157 301 184
rect 335 123 369 390
rect 403 309 463 356
rect 403 275 405 309
rect 439 275 463 309
rect 403 241 463 275
rect 403 207 405 241
rect 439 207 463 241
rect 403 168 463 207
rect 275 106 369 123
rect 25 17 91 69
rect 275 72 305 106
rect 339 72 369 106
rect 275 56 369 72
rect 403 106 459 122
rect 403 72 404 106
rect 438 72 459 106
rect 403 17 459 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a31oi_0
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3455646
string GDS_START 3449088
<< end >>
