magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 1 49 958 248
rect 0 0 960 49
<< scpmos >>
rect 84 368 120 592
rect 174 368 210 592
rect 264 368 300 592
rect 354 368 390 592
rect 561 368 597 592
rect 651 368 687 592
rect 751 368 787 592
rect 841 368 877 592
<< nmoslvt >>
rect 84 74 114 222
rect 198 74 228 222
rect 284 74 314 222
rect 398 74 428 222
rect 484 74 514 222
rect 659 74 689 222
rect 745 74 775 222
rect 841 74 871 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 149 198 222
rect 114 115 139 149
rect 173 115 198 149
rect 114 74 198 115
rect 228 210 284 222
rect 228 176 239 210
rect 273 176 284 210
rect 228 120 284 176
rect 228 86 239 120
rect 273 86 284 120
rect 228 74 284 86
rect 314 149 398 222
rect 314 115 339 149
rect 373 115 398 149
rect 314 74 398 115
rect 428 210 484 222
rect 428 176 439 210
rect 473 176 484 210
rect 428 120 484 176
rect 428 86 439 120
rect 473 86 484 120
rect 428 74 484 86
rect 514 84 659 222
rect 514 74 569 84
rect 529 50 569 74
rect 603 74 659 84
rect 689 136 745 222
rect 689 102 700 136
rect 734 102 745 136
rect 689 74 745 102
rect 775 172 841 222
rect 775 138 786 172
rect 820 138 841 172
rect 775 74 841 138
rect 871 202 932 222
rect 871 168 886 202
rect 920 168 932 202
rect 871 120 932 168
rect 871 86 886 120
rect 920 86 932 120
rect 871 74 932 86
rect 603 50 644 74
rect 529 38 644 50
<< pdiff >>
rect 28 580 84 592
rect 28 546 40 580
rect 74 546 84 580
rect 28 510 84 546
rect 28 476 40 510
rect 74 476 84 510
rect 28 440 84 476
rect 28 406 40 440
rect 74 406 84 440
rect 28 368 84 406
rect 120 580 174 592
rect 120 546 130 580
rect 164 546 174 580
rect 120 508 174 546
rect 120 474 130 508
rect 164 474 174 508
rect 120 368 174 474
rect 210 580 264 592
rect 210 546 220 580
rect 254 546 264 580
rect 210 510 264 546
rect 210 476 220 510
rect 254 476 264 510
rect 210 440 264 476
rect 210 406 220 440
rect 254 406 264 440
rect 210 368 264 406
rect 300 580 354 592
rect 300 546 310 580
rect 344 546 354 580
rect 300 508 354 546
rect 300 474 310 508
rect 344 474 354 508
rect 300 368 354 474
rect 390 531 446 592
rect 390 497 400 531
rect 434 497 446 531
rect 390 440 446 497
rect 390 406 400 440
rect 434 406 446 440
rect 390 368 446 406
rect 505 531 561 592
rect 505 497 517 531
rect 551 497 561 531
rect 505 414 561 497
rect 505 380 517 414
rect 551 380 561 414
rect 505 368 561 380
rect 597 580 651 592
rect 597 546 607 580
rect 641 546 651 580
rect 597 508 651 546
rect 597 474 607 508
rect 641 474 651 508
rect 597 368 651 474
rect 687 580 751 592
rect 687 546 707 580
rect 741 546 751 580
rect 687 510 751 546
rect 687 476 707 510
rect 741 476 751 510
rect 687 440 751 476
rect 687 406 707 440
rect 741 406 751 440
rect 687 368 751 406
rect 787 580 841 592
rect 787 546 797 580
rect 831 546 841 580
rect 787 488 841 546
rect 787 454 797 488
rect 831 454 841 488
rect 787 368 841 454
rect 877 580 933 592
rect 877 546 887 580
rect 921 546 933 580
rect 877 500 933 546
rect 877 466 887 500
rect 921 466 933 500
rect 877 420 933 466
rect 877 386 887 420
rect 921 386 933 420
rect 877 368 933 386
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 115 173 149
rect 239 176 273 210
rect 239 86 273 120
rect 339 115 373 149
rect 439 176 473 210
rect 439 86 473 120
rect 569 50 603 84
rect 700 102 734 136
rect 786 138 820 172
rect 886 168 920 202
rect 886 86 920 120
<< pdiffc >>
rect 40 546 74 580
rect 40 476 74 510
rect 40 406 74 440
rect 130 546 164 580
rect 130 474 164 508
rect 220 546 254 580
rect 220 476 254 510
rect 220 406 254 440
rect 310 546 344 580
rect 310 474 344 508
rect 400 497 434 531
rect 400 406 434 440
rect 517 497 551 531
rect 517 380 551 414
rect 607 546 641 580
rect 607 474 641 508
rect 707 546 741 580
rect 707 476 741 510
rect 707 406 741 440
rect 797 546 831 580
rect 797 454 831 488
rect 887 546 921 580
rect 887 466 921 500
rect 887 386 921 420
<< poly >>
rect 84 592 120 618
rect 174 592 210 618
rect 264 592 300 618
rect 354 592 390 618
rect 561 592 597 618
rect 651 592 687 618
rect 751 592 787 618
rect 841 592 877 618
rect 84 336 120 368
rect 174 336 210 368
rect 84 320 210 336
rect 84 286 100 320
rect 134 286 210 320
rect 264 345 300 368
rect 354 345 390 368
rect 264 320 390 345
rect 264 315 329 320
rect 84 270 210 286
rect 84 222 114 270
rect 180 267 210 270
rect 284 286 329 315
rect 363 300 390 320
rect 561 336 597 368
rect 651 336 687 368
rect 751 336 787 368
rect 841 336 877 368
rect 561 320 689 336
rect 561 300 639 320
rect 363 286 428 300
rect 284 270 428 286
rect 180 237 228 267
rect 198 222 228 237
rect 284 222 314 270
rect 398 222 428 270
rect 484 286 639 300
rect 673 286 689 320
rect 484 270 689 286
rect 484 222 514 270
rect 659 222 689 270
rect 737 326 877 336
rect 737 320 939 326
rect 737 286 753 320
rect 787 286 821 320
rect 855 310 939 320
rect 855 286 889 310
rect 737 276 889 286
rect 923 276 939 310
rect 737 260 939 276
rect 745 222 775 260
rect 841 222 871 260
rect 84 48 114 74
rect 198 48 228 74
rect 284 48 314 74
rect 398 48 428 74
rect 484 48 514 74
rect 659 48 689 74
rect 745 48 775 74
rect 841 48 871 74
<< polycont >>
rect 100 286 134 320
rect 329 286 363 320
rect 639 286 673 320
rect 753 286 787 320
rect 821 286 855 320
rect 889 276 923 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 24 580 74 596
rect 24 546 40 580
rect 24 510 74 546
rect 24 476 40 510
rect 24 440 74 476
rect 114 580 164 649
rect 114 546 130 580
rect 114 508 164 546
rect 114 474 130 508
rect 114 458 164 474
rect 204 580 270 596
rect 204 546 220 580
rect 254 546 270 580
rect 204 510 270 546
rect 204 476 220 510
rect 254 476 270 510
rect 24 406 40 440
rect 204 440 270 476
rect 310 581 657 615
rect 310 580 344 581
rect 591 580 657 581
rect 310 508 344 546
rect 310 458 344 474
rect 384 531 450 547
rect 384 497 400 531
rect 434 497 450 531
rect 204 424 220 440
rect 74 406 220 424
rect 254 424 270 440
rect 384 440 450 497
rect 384 424 400 440
rect 254 406 400 424
rect 434 406 450 440
rect 24 390 450 406
rect 501 531 551 547
rect 501 497 517 531
rect 501 424 551 497
rect 591 546 607 580
rect 641 546 657 580
rect 591 508 657 546
rect 591 474 607 508
rect 641 474 657 508
rect 591 458 657 474
rect 691 580 757 596
rect 691 546 707 580
rect 741 546 757 580
rect 691 510 757 546
rect 691 476 707 510
rect 741 476 757 510
rect 691 440 757 476
rect 691 424 707 440
rect 501 414 707 424
rect 501 380 517 414
rect 551 406 707 414
rect 741 406 757 440
rect 797 580 831 649
rect 797 488 831 546
rect 797 438 831 454
rect 871 580 937 596
rect 871 546 887 580
rect 921 546 937 580
rect 871 500 937 546
rect 871 466 887 500
rect 921 466 937 500
rect 551 404 757 406
rect 871 420 937 466
rect 871 404 887 420
rect 551 390 887 404
rect 551 380 567 390
rect 501 364 567 380
rect 723 386 887 390
rect 921 386 937 420
rect 723 370 937 386
rect 25 320 263 356
rect 25 286 100 320
rect 134 286 263 320
rect 25 270 263 286
rect 313 320 455 356
rect 313 286 329 320
rect 363 286 455 320
rect 313 270 455 286
rect 533 236 567 364
rect 601 320 689 356
rect 601 286 639 320
rect 673 286 689 320
rect 601 270 689 286
rect 737 320 939 336
rect 737 286 753 320
rect 787 286 821 320
rect 855 310 939 320
rect 855 286 889 310
rect 737 276 889 286
rect 923 276 939 310
rect 737 270 939 276
rect 873 236 939 270
rect 23 210 489 236
rect 23 176 39 210
rect 73 202 239 210
rect 73 176 89 202
rect 23 120 89 176
rect 223 176 239 202
rect 273 202 439 210
rect 273 176 289 202
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 149 189 165
rect 123 115 139 149
rect 173 115 189 149
rect 123 17 189 115
rect 223 120 289 176
rect 423 176 439 202
rect 473 176 489 210
rect 533 202 836 236
rect 423 168 489 176
rect 770 172 836 202
rect 223 86 239 120
rect 273 86 289 120
rect 223 70 289 86
rect 323 149 389 165
rect 323 115 339 149
rect 373 115 389 149
rect 323 17 389 115
rect 423 136 734 168
rect 423 134 700 136
rect 423 120 489 134
rect 423 86 439 120
rect 473 86 489 120
rect 684 102 700 134
rect 770 138 786 172
rect 820 138 836 172
rect 770 122 836 138
rect 870 168 886 202
rect 920 168 936 202
rect 423 70 489 86
rect 525 84 648 100
rect 525 50 569 84
rect 603 50 648 84
rect 684 85 734 102
rect 870 120 936 168
rect 870 86 886 120
rect 920 86 936 120
rect 870 85 936 86
rect 684 51 936 85
rect 525 17 648 50
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o31ai_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 308896
string GDS_START 300372
<< end >>
