magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 16 49 1494 241
rect 0 0 1536 49
<< scnmos >>
rect 95 47 125 215
rect 181 47 211 215
rect 267 47 297 215
rect 353 47 383 215
rect 439 47 469 215
rect 525 47 555 215
rect 611 47 641 215
rect 697 47 727 215
rect 783 47 813 215
rect 869 47 899 215
rect 955 47 985 215
rect 1041 47 1071 215
rect 1127 47 1157 215
rect 1213 47 1243 215
rect 1299 47 1329 215
rect 1385 47 1415 215
<< scpmoshvt >>
rect 95 367 125 619
rect 181 367 211 619
rect 267 367 297 619
rect 353 367 383 619
rect 439 367 469 619
rect 525 367 555 619
rect 611 367 641 619
rect 697 367 727 619
rect 783 367 813 619
rect 869 367 899 619
rect 955 367 985 619
rect 1041 367 1071 619
rect 1127 367 1157 619
rect 1213 367 1243 619
rect 1299 367 1329 619
rect 1385 367 1415 619
<< ndiff >>
rect 42 185 95 215
rect 42 151 50 185
rect 84 151 95 185
rect 42 111 95 151
rect 42 77 50 111
rect 84 77 95 111
rect 42 47 95 77
rect 125 185 181 215
rect 125 151 136 185
rect 170 151 181 185
rect 125 111 181 151
rect 125 77 136 111
rect 170 77 181 111
rect 125 47 181 77
rect 211 185 267 215
rect 211 151 222 185
rect 256 151 267 185
rect 211 111 267 151
rect 211 77 222 111
rect 256 77 267 111
rect 211 47 267 77
rect 297 185 353 215
rect 297 151 308 185
rect 342 151 353 185
rect 297 111 353 151
rect 297 77 308 111
rect 342 77 353 111
rect 297 47 353 77
rect 383 185 439 215
rect 383 151 394 185
rect 428 151 439 185
rect 383 111 439 151
rect 383 77 394 111
rect 428 77 439 111
rect 383 47 439 77
rect 469 185 525 215
rect 469 151 480 185
rect 514 151 525 185
rect 469 111 525 151
rect 469 77 480 111
rect 514 77 525 111
rect 469 47 525 77
rect 555 185 611 215
rect 555 151 566 185
rect 600 151 611 185
rect 555 111 611 151
rect 555 77 566 111
rect 600 77 611 111
rect 555 47 611 77
rect 641 185 697 215
rect 641 151 652 185
rect 686 151 697 185
rect 641 111 697 151
rect 641 77 652 111
rect 686 77 697 111
rect 641 47 697 77
rect 727 185 783 215
rect 727 151 738 185
rect 772 151 783 185
rect 727 111 783 151
rect 727 77 738 111
rect 772 77 783 111
rect 727 47 783 77
rect 813 185 869 215
rect 813 151 824 185
rect 858 151 869 185
rect 813 111 869 151
rect 813 77 824 111
rect 858 77 869 111
rect 813 47 869 77
rect 899 185 955 215
rect 899 151 910 185
rect 944 151 955 185
rect 899 111 955 151
rect 899 77 910 111
rect 944 77 955 111
rect 899 47 955 77
rect 985 185 1041 215
rect 985 151 996 185
rect 1030 151 1041 185
rect 985 111 1041 151
rect 985 77 996 111
rect 1030 77 1041 111
rect 985 47 1041 77
rect 1071 185 1127 215
rect 1071 151 1082 185
rect 1116 151 1127 185
rect 1071 111 1127 151
rect 1071 77 1082 111
rect 1116 77 1127 111
rect 1071 47 1127 77
rect 1157 185 1213 215
rect 1157 151 1168 185
rect 1202 151 1213 185
rect 1157 111 1213 151
rect 1157 77 1168 111
rect 1202 77 1213 111
rect 1157 47 1213 77
rect 1243 185 1299 215
rect 1243 151 1254 185
rect 1288 151 1299 185
rect 1243 111 1299 151
rect 1243 77 1254 111
rect 1288 77 1299 111
rect 1243 47 1299 77
rect 1329 185 1385 215
rect 1329 151 1340 185
rect 1374 151 1385 185
rect 1329 111 1385 151
rect 1329 77 1340 111
rect 1374 77 1385 111
rect 1329 47 1385 77
rect 1415 185 1468 215
rect 1415 151 1426 185
rect 1460 151 1468 185
rect 1415 111 1468 151
rect 1415 77 1426 111
rect 1460 77 1468 111
rect 1415 47 1468 77
<< pdiff >>
rect 42 596 95 619
rect 42 562 50 596
rect 84 562 95 596
rect 42 512 95 562
rect 42 478 50 512
rect 84 478 95 512
rect 42 434 95 478
rect 42 400 50 434
rect 84 400 95 434
rect 42 367 95 400
rect 125 594 181 619
rect 125 560 136 594
rect 170 560 181 594
rect 125 510 181 560
rect 125 476 136 510
rect 170 476 181 510
rect 125 426 181 476
rect 125 392 136 426
rect 170 392 181 426
rect 125 367 181 392
rect 211 596 267 619
rect 211 562 222 596
rect 256 562 267 596
rect 211 512 267 562
rect 211 478 222 512
rect 256 478 267 512
rect 211 434 267 478
rect 211 400 222 434
rect 256 400 267 434
rect 211 367 267 400
rect 297 594 353 619
rect 297 560 308 594
rect 342 560 353 594
rect 297 510 353 560
rect 297 476 308 510
rect 342 476 353 510
rect 297 426 353 476
rect 297 392 308 426
rect 342 392 353 426
rect 297 367 353 392
rect 383 596 439 619
rect 383 562 394 596
rect 428 562 439 596
rect 383 512 439 562
rect 383 478 394 512
rect 428 478 439 512
rect 383 434 439 478
rect 383 400 394 434
rect 428 400 439 434
rect 383 367 439 400
rect 469 594 525 619
rect 469 560 480 594
rect 514 560 525 594
rect 469 510 525 560
rect 469 476 480 510
rect 514 476 525 510
rect 469 426 525 476
rect 469 392 480 426
rect 514 392 525 426
rect 469 367 525 392
rect 555 596 611 619
rect 555 562 566 596
rect 600 562 611 596
rect 555 512 611 562
rect 555 478 566 512
rect 600 478 611 512
rect 555 434 611 478
rect 555 400 566 434
rect 600 400 611 434
rect 555 367 611 400
rect 641 594 697 619
rect 641 560 652 594
rect 686 560 697 594
rect 641 510 697 560
rect 641 476 652 510
rect 686 476 697 510
rect 641 426 697 476
rect 641 392 652 426
rect 686 392 697 426
rect 641 367 697 392
rect 727 596 783 619
rect 727 562 738 596
rect 772 562 783 596
rect 727 512 783 562
rect 727 478 738 512
rect 772 478 783 512
rect 727 434 783 478
rect 727 400 738 434
rect 772 400 783 434
rect 727 367 783 400
rect 813 594 869 619
rect 813 560 824 594
rect 858 560 869 594
rect 813 510 869 560
rect 813 476 824 510
rect 858 476 869 510
rect 813 426 869 476
rect 813 392 824 426
rect 858 392 869 426
rect 813 367 869 392
rect 899 596 955 619
rect 899 562 910 596
rect 944 562 955 596
rect 899 512 955 562
rect 899 478 910 512
rect 944 478 955 512
rect 899 434 955 478
rect 899 400 910 434
rect 944 400 955 434
rect 899 367 955 400
rect 985 594 1041 619
rect 985 560 996 594
rect 1030 560 1041 594
rect 985 510 1041 560
rect 985 476 996 510
rect 1030 476 1041 510
rect 985 426 1041 476
rect 985 392 996 426
rect 1030 392 1041 426
rect 985 367 1041 392
rect 1071 596 1127 619
rect 1071 562 1082 596
rect 1116 562 1127 596
rect 1071 512 1127 562
rect 1071 478 1082 512
rect 1116 478 1127 512
rect 1071 434 1127 478
rect 1071 400 1082 434
rect 1116 400 1127 434
rect 1071 367 1127 400
rect 1157 594 1213 619
rect 1157 560 1168 594
rect 1202 560 1213 594
rect 1157 510 1213 560
rect 1157 476 1168 510
rect 1202 476 1213 510
rect 1157 426 1213 476
rect 1157 392 1168 426
rect 1202 392 1213 426
rect 1157 367 1213 392
rect 1243 596 1299 619
rect 1243 562 1254 596
rect 1288 562 1299 596
rect 1243 512 1299 562
rect 1243 478 1254 512
rect 1288 478 1299 512
rect 1243 434 1299 478
rect 1243 400 1254 434
rect 1288 400 1299 434
rect 1243 367 1299 400
rect 1329 594 1385 619
rect 1329 560 1340 594
rect 1374 560 1385 594
rect 1329 510 1385 560
rect 1329 476 1340 510
rect 1374 476 1385 510
rect 1329 426 1385 476
rect 1329 392 1340 426
rect 1374 392 1385 426
rect 1329 367 1385 392
rect 1415 596 1472 619
rect 1415 562 1426 596
rect 1460 562 1472 596
rect 1415 512 1472 562
rect 1415 478 1426 512
rect 1460 478 1472 512
rect 1415 434 1472 478
rect 1415 400 1426 434
rect 1460 400 1472 434
rect 1415 367 1472 400
<< ndiffc >>
rect 50 151 84 185
rect 50 77 84 111
rect 136 151 170 185
rect 136 77 170 111
rect 222 151 256 185
rect 222 77 256 111
rect 308 151 342 185
rect 308 77 342 111
rect 394 151 428 185
rect 394 77 428 111
rect 480 151 514 185
rect 480 77 514 111
rect 566 151 600 185
rect 566 77 600 111
rect 652 151 686 185
rect 652 77 686 111
rect 738 151 772 185
rect 738 77 772 111
rect 824 151 858 185
rect 824 77 858 111
rect 910 151 944 185
rect 910 77 944 111
rect 996 151 1030 185
rect 996 77 1030 111
rect 1082 151 1116 185
rect 1082 77 1116 111
rect 1168 151 1202 185
rect 1168 77 1202 111
rect 1254 151 1288 185
rect 1254 77 1288 111
rect 1340 151 1374 185
rect 1340 77 1374 111
rect 1426 151 1460 185
rect 1426 77 1460 111
<< pdiffc >>
rect 50 562 84 596
rect 50 478 84 512
rect 50 400 84 434
rect 136 560 170 594
rect 136 476 170 510
rect 136 392 170 426
rect 222 562 256 596
rect 222 478 256 512
rect 222 400 256 434
rect 308 560 342 594
rect 308 476 342 510
rect 308 392 342 426
rect 394 562 428 596
rect 394 478 428 512
rect 394 400 428 434
rect 480 560 514 594
rect 480 476 514 510
rect 480 392 514 426
rect 566 562 600 596
rect 566 478 600 512
rect 566 400 600 434
rect 652 560 686 594
rect 652 476 686 510
rect 652 392 686 426
rect 738 562 772 596
rect 738 478 772 512
rect 738 400 772 434
rect 824 560 858 594
rect 824 476 858 510
rect 824 392 858 426
rect 910 562 944 596
rect 910 478 944 512
rect 910 400 944 434
rect 996 560 1030 594
rect 996 476 1030 510
rect 996 392 1030 426
rect 1082 562 1116 596
rect 1082 478 1116 512
rect 1082 400 1116 434
rect 1168 560 1202 594
rect 1168 476 1202 510
rect 1168 392 1202 426
rect 1254 562 1288 596
rect 1254 478 1288 512
rect 1254 400 1288 434
rect 1340 560 1374 594
rect 1340 476 1374 510
rect 1340 392 1374 426
rect 1426 562 1460 596
rect 1426 478 1460 512
rect 1426 400 1460 434
<< poly >>
rect 95 619 125 645
rect 181 619 211 645
rect 267 619 297 645
rect 353 619 383 645
rect 439 619 469 645
rect 525 619 555 645
rect 611 619 641 645
rect 697 619 727 645
rect 783 619 813 645
rect 869 619 899 645
rect 955 619 985 645
rect 1041 619 1071 645
rect 1127 619 1157 645
rect 1213 619 1243 645
rect 1299 619 1329 645
rect 1385 619 1415 645
rect 95 345 125 367
rect 181 345 211 367
rect 267 345 297 367
rect 353 345 383 367
rect 439 345 469 367
rect 525 345 555 367
rect 611 345 641 367
rect 697 345 727 367
rect 783 345 813 367
rect 869 345 899 367
rect 955 345 985 367
rect 1041 345 1071 367
rect 1127 345 1157 367
rect 1213 345 1243 367
rect 1299 345 1329 367
rect 1385 345 1415 367
rect 95 317 1415 345
rect 95 283 222 317
rect 256 283 394 317
rect 428 283 566 317
rect 600 283 738 317
rect 772 283 910 317
rect 944 283 1082 317
rect 1116 283 1254 317
rect 1288 283 1415 317
rect 95 267 1415 283
rect 95 215 125 267
rect 181 215 211 267
rect 267 215 297 267
rect 353 215 383 267
rect 439 215 469 267
rect 525 215 555 267
rect 611 215 641 267
rect 697 215 727 267
rect 783 215 813 267
rect 869 215 899 267
rect 955 215 985 267
rect 1041 215 1071 267
rect 1127 215 1157 267
rect 1213 215 1243 267
rect 1299 215 1329 267
rect 1385 215 1415 267
rect 95 21 125 47
rect 181 21 211 47
rect 267 21 297 47
rect 353 21 383 47
rect 439 21 469 47
rect 525 21 555 47
rect 611 21 641 47
rect 697 21 727 47
rect 783 21 813 47
rect 869 21 899 47
rect 955 21 985 47
rect 1041 21 1071 47
rect 1127 21 1157 47
rect 1213 21 1243 47
rect 1299 21 1329 47
rect 1385 21 1415 47
<< polycont >>
rect 222 283 256 317
rect 394 283 428 317
rect 566 283 600 317
rect 738 283 772 317
rect 910 283 944 317
rect 1082 283 1116 317
rect 1254 283 1288 317
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 34 596 93 649
rect 34 562 50 596
rect 84 562 93 596
rect 34 512 93 562
rect 34 478 50 512
rect 84 478 93 512
rect 34 434 93 478
rect 34 400 50 434
rect 84 400 93 434
rect 34 384 93 400
rect 127 594 179 610
rect 127 560 136 594
rect 170 560 179 594
rect 127 510 179 560
rect 127 476 136 510
rect 170 476 179 510
rect 127 426 179 476
rect 127 390 136 426
rect 170 390 179 426
rect 34 185 93 201
rect 34 151 50 185
rect 84 151 93 185
rect 34 111 93 151
rect 34 77 50 111
rect 84 77 93 111
rect 34 17 93 77
rect 127 185 179 390
rect 213 596 265 649
rect 213 562 222 596
rect 256 562 265 596
rect 213 512 265 562
rect 213 478 222 512
rect 256 478 265 512
rect 213 434 265 478
rect 213 400 222 434
rect 256 400 265 434
rect 213 384 265 400
rect 299 594 351 610
rect 299 560 308 594
rect 342 560 351 594
rect 299 510 351 560
rect 299 476 308 510
rect 342 476 351 510
rect 299 426 351 476
rect 299 390 308 426
rect 342 390 351 426
rect 213 283 222 350
rect 256 283 265 350
rect 213 267 265 283
rect 127 151 136 185
rect 170 151 179 185
rect 127 111 179 151
rect 127 77 136 111
rect 170 77 179 111
rect 127 61 179 77
rect 213 185 265 201
rect 213 151 222 185
rect 256 151 265 185
rect 213 111 265 151
rect 213 77 222 111
rect 256 77 265 111
rect 213 17 265 77
rect 299 185 351 390
rect 385 596 437 649
rect 385 562 394 596
rect 428 562 437 596
rect 385 512 437 562
rect 385 478 394 512
rect 428 478 437 512
rect 385 434 437 478
rect 385 400 394 434
rect 428 400 437 434
rect 385 384 437 400
rect 471 594 523 610
rect 471 560 480 594
rect 514 560 523 594
rect 471 510 523 560
rect 471 476 480 510
rect 514 476 523 510
rect 471 426 523 476
rect 471 390 480 426
rect 514 390 523 426
rect 385 283 394 350
rect 428 283 437 350
rect 385 267 437 283
rect 299 151 308 185
rect 342 151 351 185
rect 299 111 351 151
rect 299 77 308 111
rect 342 77 351 111
rect 299 61 351 77
rect 385 185 437 201
rect 385 151 394 185
rect 428 151 437 185
rect 385 111 437 151
rect 385 77 394 111
rect 428 77 437 111
rect 385 17 437 77
rect 471 185 523 390
rect 557 596 609 649
rect 557 562 566 596
rect 600 562 609 596
rect 557 512 609 562
rect 557 478 566 512
rect 600 478 609 512
rect 557 434 609 478
rect 557 400 566 434
rect 600 400 609 434
rect 557 384 609 400
rect 643 594 695 610
rect 643 560 652 594
rect 686 560 695 594
rect 643 510 695 560
rect 643 476 652 510
rect 686 476 695 510
rect 643 426 695 476
rect 643 390 652 426
rect 686 390 695 426
rect 557 283 566 350
rect 600 283 609 350
rect 557 267 609 283
rect 471 151 480 185
rect 514 151 523 185
rect 471 111 523 151
rect 471 77 480 111
rect 514 77 523 111
rect 471 61 523 77
rect 557 185 609 201
rect 557 151 566 185
rect 600 151 609 185
rect 557 111 609 151
rect 557 77 566 111
rect 600 77 609 111
rect 557 17 609 77
rect 643 185 695 390
rect 729 596 781 649
rect 729 562 738 596
rect 772 562 781 596
rect 729 512 781 562
rect 729 478 738 512
rect 772 478 781 512
rect 729 434 781 478
rect 729 400 738 434
rect 772 400 781 434
rect 729 384 781 400
rect 815 594 867 610
rect 815 560 824 594
rect 858 560 867 594
rect 815 510 867 560
rect 815 476 824 510
rect 858 476 867 510
rect 815 426 867 476
rect 815 390 824 426
rect 858 390 867 426
rect 729 283 738 350
rect 772 283 781 350
rect 729 267 781 283
rect 643 151 652 185
rect 686 151 695 185
rect 643 111 695 151
rect 643 77 652 111
rect 686 77 695 111
rect 643 61 695 77
rect 729 185 781 201
rect 729 151 738 185
rect 772 151 781 185
rect 729 111 781 151
rect 729 77 738 111
rect 772 77 781 111
rect 729 17 781 77
rect 815 185 867 390
rect 901 596 953 649
rect 901 562 910 596
rect 944 562 953 596
rect 901 512 953 562
rect 901 478 910 512
rect 944 478 953 512
rect 901 434 953 478
rect 901 400 910 434
rect 944 400 953 434
rect 901 384 953 400
rect 987 594 1039 610
rect 987 560 996 594
rect 1030 560 1039 594
rect 987 510 1039 560
rect 987 476 996 510
rect 1030 476 1039 510
rect 987 426 1039 476
rect 987 390 996 426
rect 1030 390 1039 426
rect 901 283 910 350
rect 944 283 953 350
rect 901 267 953 283
rect 815 151 824 185
rect 858 151 867 185
rect 815 111 867 151
rect 815 77 824 111
rect 858 77 867 111
rect 815 61 867 77
rect 901 185 953 201
rect 901 151 910 185
rect 944 151 953 185
rect 901 111 953 151
rect 901 77 910 111
rect 944 77 953 111
rect 901 17 953 77
rect 987 185 1039 390
rect 1073 596 1125 649
rect 1073 562 1082 596
rect 1116 562 1125 596
rect 1073 512 1125 562
rect 1073 478 1082 512
rect 1116 478 1125 512
rect 1073 434 1125 478
rect 1073 400 1082 434
rect 1116 400 1125 434
rect 1073 384 1125 400
rect 1159 594 1211 610
rect 1159 560 1168 594
rect 1202 560 1211 594
rect 1159 510 1211 560
rect 1159 476 1168 510
rect 1202 476 1211 510
rect 1159 426 1211 476
rect 1159 390 1168 426
rect 1202 390 1211 426
rect 1073 283 1082 350
rect 1116 283 1125 350
rect 1073 267 1125 283
rect 987 151 996 185
rect 1030 151 1039 185
rect 987 111 1039 151
rect 987 77 996 111
rect 1030 77 1039 111
rect 987 61 1039 77
rect 1073 185 1125 201
rect 1073 151 1082 185
rect 1116 151 1125 185
rect 1073 111 1125 151
rect 1073 77 1082 111
rect 1116 77 1125 111
rect 1073 17 1125 77
rect 1159 185 1211 390
rect 1245 596 1297 649
rect 1245 562 1254 596
rect 1288 562 1297 596
rect 1245 512 1297 562
rect 1245 478 1254 512
rect 1288 478 1297 512
rect 1245 434 1297 478
rect 1245 400 1254 434
rect 1288 400 1297 434
rect 1245 384 1297 400
rect 1331 594 1383 610
rect 1331 560 1340 594
rect 1374 560 1383 594
rect 1331 510 1383 560
rect 1331 476 1340 510
rect 1374 476 1383 510
rect 1331 426 1383 476
rect 1331 390 1340 426
rect 1374 390 1383 426
rect 1245 283 1254 350
rect 1288 283 1297 350
rect 1245 267 1297 283
rect 1159 151 1168 185
rect 1202 151 1211 185
rect 1159 111 1211 151
rect 1159 77 1168 111
rect 1202 77 1211 111
rect 1159 61 1211 77
rect 1245 185 1297 201
rect 1245 151 1254 185
rect 1288 151 1297 185
rect 1245 111 1297 151
rect 1245 77 1254 111
rect 1288 77 1297 111
rect 1245 17 1297 77
rect 1331 185 1383 390
rect 1417 596 1476 649
rect 1417 562 1426 596
rect 1460 562 1476 596
rect 1417 512 1476 562
rect 1417 478 1426 512
rect 1460 478 1476 512
rect 1417 434 1476 478
rect 1417 400 1426 434
rect 1460 400 1476 434
rect 1417 384 1476 400
rect 1331 151 1340 185
rect 1374 151 1383 185
rect 1331 111 1383 151
rect 1331 77 1340 111
rect 1374 77 1383 111
rect 1331 61 1383 77
rect 1417 185 1476 201
rect 1417 151 1426 185
rect 1460 151 1476 185
rect 1417 111 1476 151
rect 1417 77 1426 111
rect 1460 77 1476 111
rect 1417 17 1476 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 136 392 170 424
rect 136 390 170 392
rect 308 392 342 424
rect 308 390 342 392
rect 222 317 256 350
rect 222 316 256 317
rect 480 392 514 424
rect 480 390 514 392
rect 394 317 428 350
rect 394 316 428 317
rect 652 392 686 424
rect 652 390 686 392
rect 566 317 600 350
rect 566 316 600 317
rect 824 392 858 424
rect 824 390 858 392
rect 738 317 772 350
rect 738 316 772 317
rect 996 392 1030 424
rect 996 390 1030 392
rect 910 317 944 350
rect 910 316 944 317
rect 1168 392 1202 424
rect 1168 390 1202 392
rect 1082 317 1116 350
rect 1082 316 1116 317
rect 1340 392 1374 424
rect 1340 390 1374 392
rect 1254 317 1288 350
rect 1254 316 1288 317
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 560 100 617
rect 124 424 1386 430
rect 124 390 136 424
rect 170 390 308 424
rect 342 390 480 424
rect 514 390 652 424
rect 686 390 824 424
rect 858 390 996 424
rect 1030 390 1168 424
rect 1202 390 1340 424
rect 1374 390 1386 424
rect 124 384 1386 390
rect 210 350 1300 356
rect 210 316 222 350
rect 256 316 394 350
rect 428 316 566 350
rect 600 316 738 350
rect 772 316 910 350
rect 944 316 1082 350
rect 1116 316 1254 350
rect 1288 316 1300 350
rect 210 310 1300 316
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 inv_16
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 124 384 1386 430 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel metal1 s 210 310 1300 356 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
rlabel metal1 s 0 617 1536 715 1 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 560 100 617 1 VPB
port 4 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5455290
string GDS_START 5442082
<< end >>
