magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 11 243 285 273
rect 11 49 928 243
rect 0 0 960 49
<< scnmos >>
rect 90 79 120 247
rect 176 79 206 247
rect 423 49 453 217
rect 531 49 561 217
rect 603 49 633 217
rect 711 49 741 217
rect 819 49 849 217
<< scpmoshvt >>
rect 90 367 120 619
rect 176 367 206 619
rect 423 367 453 619
rect 509 367 539 619
rect 603 367 633 619
rect 733 367 763 619
rect 819 367 849 619
<< ndiff >>
rect 37 235 90 247
rect 37 201 45 235
rect 79 201 90 235
rect 37 125 90 201
rect 37 91 45 125
rect 79 91 90 125
rect 37 79 90 91
rect 120 212 176 247
rect 120 178 131 212
rect 165 178 176 212
rect 120 144 176 178
rect 120 110 131 144
rect 165 110 176 144
rect 120 79 176 110
rect 206 235 259 247
rect 206 201 217 235
rect 251 201 259 235
rect 206 125 259 201
rect 206 91 217 125
rect 251 91 259 125
rect 206 79 259 91
rect 370 205 423 217
rect 370 171 378 205
rect 412 171 423 205
rect 370 101 423 171
rect 370 67 378 101
rect 412 67 423 101
rect 370 49 423 67
rect 453 165 531 217
rect 453 131 475 165
rect 509 131 531 165
rect 453 91 531 131
rect 453 57 475 91
rect 509 57 531 91
rect 453 49 531 57
rect 561 49 603 217
rect 633 49 711 217
rect 741 49 819 217
rect 849 205 902 217
rect 849 171 860 205
rect 894 171 902 205
rect 849 101 902 171
rect 849 67 860 101
rect 894 67 902 101
rect 849 49 902 67
<< pdiff >>
rect 37 607 90 619
rect 37 573 45 607
rect 79 573 90 607
rect 37 506 90 573
rect 37 472 45 506
rect 79 472 90 506
rect 37 413 90 472
rect 37 379 45 413
rect 79 379 90 413
rect 37 367 90 379
rect 120 549 176 619
rect 120 515 131 549
rect 165 515 176 549
rect 120 481 176 515
rect 120 447 131 481
rect 165 447 176 481
rect 120 413 176 447
rect 120 379 131 413
rect 165 379 176 413
rect 120 367 176 379
rect 206 607 259 619
rect 206 573 217 607
rect 251 573 259 607
rect 206 509 259 573
rect 206 475 217 509
rect 251 475 259 509
rect 206 419 259 475
rect 206 385 217 419
rect 251 385 259 419
rect 206 367 259 385
rect 370 599 423 619
rect 370 565 378 599
rect 412 565 423 599
rect 370 516 423 565
rect 370 482 378 516
rect 412 482 423 516
rect 370 434 423 482
rect 370 400 378 434
rect 412 400 423 434
rect 370 367 423 400
rect 453 599 509 619
rect 453 565 464 599
rect 498 565 509 599
rect 453 515 509 565
rect 453 481 464 515
rect 498 481 509 515
rect 453 436 509 481
rect 453 402 464 436
rect 498 402 509 436
rect 453 367 509 402
rect 539 607 603 619
rect 539 573 554 607
rect 588 573 603 607
rect 539 494 603 573
rect 539 460 554 494
rect 588 460 603 494
rect 539 367 603 460
rect 633 599 733 619
rect 633 565 668 599
rect 702 565 733 599
rect 633 511 733 565
rect 633 477 668 511
rect 702 477 733 511
rect 633 420 733 477
rect 633 386 668 420
rect 702 386 733 420
rect 633 367 733 386
rect 763 607 819 619
rect 763 573 774 607
rect 808 573 819 607
rect 763 494 819 573
rect 763 460 774 494
rect 808 460 819 494
rect 763 367 819 460
rect 849 599 902 619
rect 849 565 860 599
rect 894 565 902 599
rect 849 518 902 565
rect 849 484 860 518
rect 894 484 902 518
rect 849 436 902 484
rect 849 402 860 436
rect 894 402 902 436
rect 849 367 902 402
<< ndiffc >>
rect 45 201 79 235
rect 45 91 79 125
rect 131 178 165 212
rect 131 110 165 144
rect 217 201 251 235
rect 217 91 251 125
rect 378 171 412 205
rect 378 67 412 101
rect 475 131 509 165
rect 475 57 509 91
rect 860 171 894 205
rect 860 67 894 101
<< pdiffc >>
rect 45 573 79 607
rect 45 472 79 506
rect 45 379 79 413
rect 131 515 165 549
rect 131 447 165 481
rect 131 379 165 413
rect 217 573 251 607
rect 217 475 251 509
rect 217 385 251 419
rect 378 565 412 599
rect 378 482 412 516
rect 378 400 412 434
rect 464 565 498 599
rect 464 481 498 515
rect 464 402 498 436
rect 554 573 588 607
rect 554 460 588 494
rect 668 565 702 599
rect 668 477 702 511
rect 668 386 702 420
rect 774 573 808 607
rect 774 460 808 494
rect 860 565 894 599
rect 860 484 894 518
rect 860 402 894 436
<< poly >>
rect 90 619 120 645
rect 176 619 206 645
rect 423 619 453 645
rect 509 619 539 645
rect 603 619 633 645
rect 733 619 763 645
rect 819 619 849 645
rect 90 299 120 367
rect 176 335 206 367
rect 423 335 453 367
rect 509 335 539 367
rect 603 335 633 367
rect 733 335 763 367
rect 176 319 255 335
rect 176 299 205 319
rect 90 285 205 299
rect 239 285 255 319
rect 90 269 255 285
rect 387 319 453 335
rect 387 285 403 319
rect 437 285 453 319
rect 387 269 453 285
rect 495 319 561 335
rect 495 285 511 319
rect 545 285 561 319
rect 495 269 561 285
rect 90 247 120 269
rect 176 247 206 269
rect 423 217 453 269
rect 531 217 561 269
rect 603 319 669 335
rect 603 285 619 319
rect 653 285 669 319
rect 603 269 669 285
rect 711 319 777 335
rect 711 285 727 319
rect 761 285 777 319
rect 711 269 777 285
rect 819 325 849 367
rect 819 309 935 325
rect 819 275 885 309
rect 919 275 935 309
rect 603 217 633 269
rect 711 217 741 269
rect 819 259 935 275
rect 819 217 849 259
rect 90 53 120 79
rect 176 53 206 79
rect 423 23 453 49
rect 531 23 561 49
rect 603 23 633 49
rect 711 23 741 49
rect 819 23 849 49
<< polycont >>
rect 205 285 239 319
rect 403 285 437 319
rect 511 285 545 319
rect 619 285 653 319
rect 727 285 761 319
rect 885 275 919 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 29 607 86 649
rect 29 573 45 607
rect 79 573 86 607
rect 201 607 267 649
rect 29 506 86 573
rect 29 472 45 506
rect 79 472 86 506
rect 29 413 86 472
rect 29 379 45 413
rect 79 379 86 413
rect 29 363 86 379
rect 120 549 167 595
rect 120 515 131 549
rect 165 515 167 549
rect 120 481 167 515
rect 120 447 131 481
rect 165 447 167 481
rect 120 413 167 447
rect 120 379 131 413
rect 165 379 167 413
rect 29 235 86 251
rect 29 201 45 235
rect 79 201 86 235
rect 29 125 86 201
rect 29 91 45 125
rect 79 91 86 125
rect 29 17 86 91
rect 120 212 167 379
rect 201 573 217 607
rect 251 573 267 607
rect 201 509 267 573
rect 201 475 217 509
rect 251 475 267 509
rect 201 419 267 475
rect 362 599 416 615
rect 362 565 378 599
rect 412 565 416 599
rect 362 516 416 565
rect 362 482 378 516
rect 412 482 416 516
rect 362 434 416 482
rect 362 420 378 434
rect 201 385 217 419
rect 251 385 267 419
rect 201 369 267 385
rect 333 400 378 420
rect 412 400 416 434
rect 333 384 416 400
rect 460 599 504 615
rect 460 565 464 599
rect 498 565 504 599
rect 460 515 504 565
rect 460 481 464 515
rect 498 481 504 515
rect 460 436 504 481
rect 538 607 604 649
rect 538 573 554 607
rect 588 573 604 607
rect 538 494 604 573
rect 538 460 554 494
rect 588 460 604 494
rect 538 454 604 460
rect 652 599 718 615
rect 652 565 668 599
rect 702 565 718 599
rect 652 511 718 565
rect 652 477 668 511
rect 702 477 718 511
rect 460 402 464 436
rect 498 420 504 436
rect 652 420 718 477
rect 758 607 824 649
rect 758 573 774 607
rect 808 573 824 607
rect 758 494 824 573
rect 758 460 774 494
rect 808 460 824 494
rect 758 454 824 460
rect 858 599 910 615
rect 858 565 860 599
rect 894 565 910 599
rect 858 518 910 565
rect 858 484 860 518
rect 894 484 910 518
rect 858 436 910 484
rect 858 420 860 436
rect 498 402 668 420
rect 460 386 668 402
rect 702 402 860 420
rect 894 402 910 436
rect 702 386 910 402
rect 460 384 910 386
rect 333 335 367 384
rect 205 319 367 335
rect 239 285 367 319
rect 205 269 367 285
rect 401 319 461 350
rect 401 285 403 319
rect 437 285 461 319
rect 401 269 461 285
rect 495 319 561 350
rect 495 285 511 319
rect 545 285 561 319
rect 495 269 561 285
rect 595 319 661 350
rect 595 285 619 319
rect 653 285 661 319
rect 595 269 661 285
rect 695 319 835 350
rect 695 285 727 319
rect 761 285 835 319
rect 695 269 835 285
rect 869 309 942 350
rect 869 275 885 309
rect 919 275 942 309
rect 869 269 942 275
rect 120 178 131 212
rect 165 178 167 212
rect 120 144 167 178
rect 120 110 131 144
rect 165 110 167 144
rect 120 72 167 110
rect 201 201 217 235
rect 251 201 267 235
rect 201 125 267 201
rect 201 91 217 125
rect 251 91 267 125
rect 201 17 267 91
rect 301 233 367 269
rect 301 205 910 233
rect 301 171 378 205
rect 412 199 860 205
rect 412 171 416 199
rect 301 101 416 171
rect 844 171 860 199
rect 894 171 910 205
rect 301 67 378 101
rect 412 67 416 101
rect 301 51 416 67
rect 459 131 475 165
rect 509 131 525 165
rect 459 91 525 131
rect 459 57 475 91
rect 509 57 525 91
rect 459 17 525 57
rect 844 101 910 171
rect 844 67 860 101
rect 894 67 910 101
rect 844 51 910 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a41o_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5486522
string GDS_START 5477640
<< end >>
