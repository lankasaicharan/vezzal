magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
rect 804 329 1012 331
<< pwell >>
rect 485 184 973 243
rect 1351 184 1627 249
rect 485 180 1627 184
rect 1 49 1627 180
rect 0 0 1632 49
<< scnmos >>
rect 80 70 110 154
rect 166 70 196 154
rect 252 70 282 154
rect 584 133 614 217
rect 670 133 700 217
rect 742 133 772 217
rect 860 49 890 217
rect 1058 74 1088 158
rect 1144 74 1174 158
rect 1216 74 1246 158
rect 1432 55 1462 223
rect 1518 55 1548 223
<< scpmoshvt >>
rect 80 468 110 596
rect 152 468 182 596
rect 381 417 411 545
rect 630 457 660 541
rect 716 457 746 541
rect 788 457 818 541
rect 893 365 923 617
rect 1087 429 1117 557
rect 1205 429 1235 557
rect 1291 429 1321 557
rect 1432 367 1462 619
rect 1518 367 1548 619
<< ndiff >>
rect 27 126 80 154
rect 27 92 35 126
rect 69 92 80 126
rect 27 70 80 92
rect 110 129 166 154
rect 110 95 121 129
rect 155 95 166 129
rect 110 70 166 95
rect 196 129 252 154
rect 196 95 207 129
rect 241 95 252 129
rect 196 70 252 95
rect 282 129 335 154
rect 282 95 293 129
rect 327 95 335 129
rect 282 70 335 95
rect 511 207 584 217
rect 511 173 523 207
rect 557 173 584 207
rect 511 133 584 173
rect 614 207 670 217
rect 614 173 625 207
rect 659 173 670 207
rect 614 133 670 173
rect 700 133 742 217
rect 772 133 860 217
rect 787 71 860 133
rect 787 37 799 71
rect 833 49 860 71
rect 890 207 947 217
rect 890 173 901 207
rect 935 173 947 207
rect 890 49 947 173
rect 1377 175 1432 223
rect 1005 123 1058 158
rect 1005 89 1013 123
rect 1047 89 1058 123
rect 1005 74 1058 89
rect 1088 126 1144 158
rect 1088 92 1099 126
rect 1133 92 1144 126
rect 1088 74 1144 92
rect 1174 74 1216 158
rect 1246 128 1299 158
rect 1246 94 1257 128
rect 1291 94 1299 128
rect 1246 74 1299 94
rect 1377 141 1385 175
rect 1419 141 1432 175
rect 1377 101 1432 141
rect 833 37 845 49
rect 787 27 845 37
rect 1377 67 1385 101
rect 1419 67 1432 101
rect 1377 55 1432 67
rect 1462 212 1518 223
rect 1462 178 1473 212
rect 1507 178 1518 212
rect 1462 101 1518 178
rect 1462 67 1473 101
rect 1507 67 1518 101
rect 1462 55 1518 67
rect 1548 209 1601 223
rect 1548 175 1559 209
rect 1593 175 1601 209
rect 1548 101 1601 175
rect 1548 67 1559 101
rect 1593 67 1601 101
rect 1548 55 1601 67
<< pdiff >>
rect 27 584 80 596
rect 27 550 35 584
rect 69 550 80 584
rect 27 516 80 550
rect 27 482 35 516
rect 69 482 80 516
rect 27 468 80 482
rect 110 468 152 596
rect 182 582 235 596
rect 182 548 193 582
rect 227 548 235 582
rect 182 514 235 548
rect 182 480 193 514
rect 227 480 235 514
rect 182 468 235 480
rect 295 537 381 545
rect 295 503 309 537
rect 343 503 381 537
rect 295 488 381 503
rect 331 417 381 488
rect 411 529 509 545
rect 840 605 893 617
rect 840 571 848 605
rect 882 571 893 605
rect 840 541 893 571
rect 411 495 461 529
rect 495 495 509 529
rect 411 459 509 495
rect 411 425 461 459
rect 495 425 509 459
rect 577 515 630 541
rect 577 481 585 515
rect 619 481 630 515
rect 577 457 630 481
rect 660 515 716 541
rect 660 481 671 515
rect 705 481 716 515
rect 660 457 716 481
rect 746 457 788 541
rect 818 529 893 541
rect 818 495 829 529
rect 863 495 893 529
rect 818 457 893 495
rect 411 417 509 425
rect 840 451 893 457
rect 840 417 848 451
rect 882 417 893 451
rect 840 365 893 417
rect 923 599 976 617
rect 923 565 934 599
rect 968 565 976 599
rect 1132 609 1190 619
rect 923 500 976 565
rect 1132 575 1144 609
rect 1178 575 1190 609
rect 1375 607 1432 619
rect 1132 557 1190 575
rect 1375 573 1387 607
rect 1421 573 1432 607
rect 1375 557 1432 573
rect 923 466 934 500
rect 968 466 976 500
rect 923 411 976 466
rect 1030 473 1087 557
rect 1030 439 1042 473
rect 1076 439 1087 473
rect 1030 429 1087 439
rect 1117 429 1205 557
rect 1235 549 1291 557
rect 1235 515 1246 549
rect 1280 515 1291 549
rect 1235 481 1291 515
rect 1235 447 1246 481
rect 1280 447 1291 481
rect 1235 429 1291 447
rect 1321 545 1432 557
rect 1321 511 1332 545
rect 1366 511 1432 545
rect 1321 429 1432 511
rect 923 377 934 411
rect 968 377 976 411
rect 923 365 976 377
rect 1375 367 1432 429
rect 1462 409 1518 619
rect 1462 375 1473 409
rect 1507 375 1518 409
rect 1462 367 1518 375
rect 1548 561 1601 619
rect 1548 527 1559 561
rect 1593 527 1601 561
rect 1548 367 1601 527
<< ndiffc >>
rect 35 92 69 126
rect 121 95 155 129
rect 207 95 241 129
rect 293 95 327 129
rect 523 173 557 207
rect 625 173 659 207
rect 799 37 833 71
rect 901 173 935 207
rect 1013 89 1047 123
rect 1099 92 1133 126
rect 1257 94 1291 128
rect 1385 141 1419 175
rect 1385 67 1419 101
rect 1473 178 1507 212
rect 1473 67 1507 101
rect 1559 175 1593 209
rect 1559 67 1593 101
<< pdiffc >>
rect 35 550 69 584
rect 35 482 69 516
rect 193 548 227 582
rect 193 480 227 514
rect 309 503 343 537
rect 848 571 882 605
rect 461 495 495 529
rect 461 425 495 459
rect 585 481 619 515
rect 671 481 705 515
rect 829 495 863 529
rect 848 417 882 451
rect 934 565 968 599
rect 1144 575 1178 609
rect 1387 573 1421 607
rect 934 466 968 500
rect 1042 439 1076 473
rect 1246 515 1280 549
rect 1246 447 1280 481
rect 1332 511 1366 545
rect 934 377 968 411
rect 1473 375 1507 409
rect 1559 527 1593 561
<< poly >>
rect 80 596 110 622
rect 152 596 182 622
rect 250 615 746 645
rect 893 617 923 643
rect 1432 619 1462 645
rect 1518 619 1548 645
rect 250 473 280 615
rect 381 545 411 571
rect 80 310 110 468
rect 152 395 182 468
rect 250 443 316 473
rect 152 379 237 395
rect 152 365 187 379
rect 31 294 110 310
rect 31 260 47 294
rect 81 260 110 294
rect 31 226 110 260
rect 31 192 47 226
rect 81 192 110 226
rect 31 176 110 192
rect 80 154 110 176
rect 166 345 187 365
rect 221 345 237 379
rect 166 311 237 345
rect 166 277 187 311
rect 221 277 237 311
rect 166 261 237 277
rect 286 269 316 443
rect 630 541 660 567
rect 716 541 746 615
rect 788 541 818 567
rect 630 425 660 457
rect 716 431 746 457
rect 381 269 411 417
rect 524 395 660 425
rect 524 383 554 395
rect 788 383 818 457
rect 453 367 554 383
rect 453 333 469 367
rect 503 347 554 367
rect 742 367 818 383
rect 503 333 700 347
rect 453 317 700 333
rect 166 154 196 261
rect 286 239 614 269
rect 286 206 447 239
rect 584 217 614 239
rect 670 217 700 317
rect 742 333 758 367
rect 792 333 818 367
rect 1087 557 1117 583
rect 1205 557 1235 583
rect 1291 557 1321 583
rect 1087 371 1117 429
rect 1205 371 1235 429
rect 1291 397 1321 429
rect 742 317 818 333
rect 742 217 772 317
rect 893 311 923 365
rect 1087 341 1235 371
rect 1277 381 1343 397
rect 1277 347 1293 381
rect 1327 347 1343 381
rect 1087 314 1174 341
rect 860 295 926 311
rect 860 261 876 295
rect 910 261 926 295
rect 860 245 926 261
rect 1058 298 1174 314
rect 1058 264 1087 298
rect 1121 264 1174 298
rect 1277 313 1343 347
rect 1277 293 1293 313
rect 860 217 890 245
rect 1058 230 1174 264
rect 252 176 447 206
rect 252 154 282 176
rect 381 155 447 176
rect 381 121 397 155
rect 431 121 447 155
rect 381 87 447 121
rect 584 107 614 133
rect 670 107 700 133
rect 742 107 772 133
rect 80 44 110 70
rect 166 44 196 70
rect 252 44 282 70
rect 381 53 397 87
rect 431 53 447 87
rect 381 37 447 53
rect 1058 196 1087 230
rect 1121 196 1174 230
rect 1058 180 1174 196
rect 1058 158 1088 180
rect 1144 158 1174 180
rect 1216 279 1293 293
rect 1327 279 1343 313
rect 1216 263 1343 279
rect 1432 289 1462 367
rect 1518 325 1548 367
rect 1518 309 1609 325
rect 1518 289 1559 309
rect 1432 275 1559 289
rect 1593 275 1609 309
rect 1216 158 1246 263
rect 1432 259 1609 275
rect 1432 223 1462 259
rect 1518 223 1548 259
rect 860 23 890 49
rect 1058 48 1088 74
rect 1144 48 1174 74
rect 1216 48 1246 74
rect 1432 29 1462 55
rect 1518 29 1548 55
<< polycont >>
rect 47 260 81 294
rect 47 192 81 226
rect 187 345 221 379
rect 187 277 221 311
rect 469 333 503 367
rect 758 333 792 367
rect 1293 347 1327 381
rect 876 261 910 295
rect 1087 264 1121 298
rect 397 121 431 155
rect 397 53 431 87
rect 1087 196 1121 230
rect 1293 279 1327 313
rect 1559 275 1593 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 19 584 83 649
rect 19 550 35 584
rect 69 550 83 584
rect 19 516 83 550
rect 19 482 35 516
rect 69 482 83 516
rect 19 466 83 482
rect 117 582 243 598
rect 117 548 193 582
rect 227 548 243 582
rect 117 514 243 548
rect 117 480 193 514
rect 227 480 243 514
rect 293 537 359 649
rect 293 503 309 537
rect 343 503 359 537
rect 293 501 359 503
rect 393 579 627 613
rect 117 467 243 480
rect 393 467 427 579
rect 117 433 427 467
rect 461 529 505 545
rect 495 495 505 529
rect 461 459 505 495
rect 17 294 83 432
rect 17 260 47 294
rect 81 260 83 294
rect 17 226 83 260
rect 17 192 47 226
rect 81 192 83 226
rect 17 168 83 192
rect 117 186 151 433
rect 495 425 505 459
rect 185 379 263 395
rect 461 383 505 425
rect 185 345 187 379
rect 221 345 263 379
rect 185 311 263 345
rect 185 277 187 311
rect 221 277 263 311
rect 185 261 263 277
rect 297 367 505 383
rect 297 333 469 367
rect 503 333 505 367
rect 297 317 505 333
rect 539 515 627 579
rect 809 605 898 649
rect 809 571 848 605
rect 882 571 898 605
rect 539 481 585 515
rect 619 481 627 515
rect 539 465 627 481
rect 661 515 709 531
rect 661 481 671 515
rect 705 481 709 515
rect 297 225 343 317
rect 539 225 573 465
rect 661 279 709 481
rect 809 529 898 571
rect 809 495 829 529
rect 863 495 898 529
rect 809 451 898 495
rect 809 417 848 451
rect 882 417 898 451
rect 932 599 984 615
rect 932 565 934 599
rect 968 565 984 599
rect 1128 609 1194 649
rect 1128 575 1144 609
rect 1178 575 1194 609
rect 1316 607 1437 649
rect 1316 573 1387 607
rect 1421 573 1437 607
rect 932 541 984 565
rect 1230 549 1282 565
rect 932 507 1191 541
rect 932 500 980 507
rect 932 466 934 500
rect 968 466 980 500
rect 932 411 980 466
rect 932 383 934 411
rect 743 377 934 383
rect 968 377 980 411
rect 743 367 980 377
rect 743 333 758 367
rect 792 349 980 367
rect 792 333 808 349
rect 743 317 808 333
rect 860 295 912 311
rect 860 279 876 295
rect 117 148 164 186
rect 19 126 85 134
rect 19 92 35 126
rect 69 92 85 126
rect 19 17 85 92
rect 119 129 164 148
rect 119 95 121 129
rect 155 95 164 129
rect 119 79 164 95
rect 198 129 250 145
rect 198 95 207 129
rect 241 95 250 129
rect 198 17 250 95
rect 284 129 343 225
rect 507 207 573 225
rect 507 173 523 207
rect 557 173 573 207
rect 609 261 876 279
rect 910 261 912 295
rect 609 245 912 261
rect 609 207 709 245
rect 946 211 980 349
rect 609 173 625 207
rect 659 173 709 207
rect 885 207 980 211
rect 885 173 901 207
rect 935 173 980 207
rect 1014 439 1042 473
rect 1076 439 1092 473
rect 1014 423 1092 439
rect 284 95 293 129
rect 327 95 343 129
rect 284 79 343 95
rect 381 155 447 171
rect 381 121 397 155
rect 431 139 447 155
rect 1014 139 1049 423
rect 1157 381 1191 507
rect 1230 515 1246 549
rect 1280 515 1282 549
rect 1230 481 1282 515
rect 1316 545 1437 573
rect 1316 511 1332 545
rect 1366 511 1437 545
rect 1543 561 1609 649
rect 1543 527 1559 561
rect 1593 527 1609 561
rect 1543 511 1609 527
rect 1230 447 1246 481
rect 1280 477 1282 481
rect 1280 447 1609 477
rect 1230 443 1609 447
rect 1230 415 1423 443
rect 1083 313 1123 366
rect 1157 347 1293 381
rect 1327 347 1343 381
rect 1277 313 1343 347
rect 1083 298 1158 313
rect 1083 264 1087 298
rect 1121 264 1158 298
rect 1277 279 1293 313
rect 1327 279 1343 313
rect 1277 277 1343 279
rect 1083 230 1158 264
rect 1379 243 1423 415
rect 1457 375 1473 409
rect 1507 375 1523 409
rect 1457 371 1523 375
rect 1083 196 1087 230
rect 1121 196 1158 230
rect 1083 168 1158 196
rect 1241 209 1423 243
rect 1469 212 1523 371
rect 1557 309 1609 443
rect 1557 275 1559 309
rect 1593 275 1609 309
rect 1557 259 1609 275
rect 431 123 1049 139
rect 431 121 1013 123
rect 381 105 1013 121
rect 381 87 447 105
rect 381 53 397 87
rect 431 53 447 87
rect 997 89 1013 105
rect 1047 89 1049 123
rect 997 73 1049 89
rect 1083 126 1149 134
rect 1083 92 1099 126
rect 1133 92 1149 126
rect 381 51 447 53
rect 783 37 799 71
rect 833 37 849 71
rect 783 17 849 37
rect 1083 17 1149 92
rect 1241 128 1307 209
rect 1469 178 1473 212
rect 1507 178 1523 212
rect 1241 94 1257 128
rect 1291 94 1307 128
rect 1241 90 1307 94
rect 1369 141 1385 175
rect 1419 141 1435 175
rect 1369 101 1435 141
rect 1369 67 1385 101
rect 1419 67 1435 101
rect 1369 17 1435 67
rect 1469 101 1523 178
rect 1469 67 1473 101
rect 1507 67 1523 101
rect 1469 51 1523 67
rect 1557 209 1609 225
rect 1557 175 1559 209
rect 1593 175 1609 209
rect 1557 101 1609 175
rect 1557 67 1559 101
rect 1593 67 1609 101
rect 1557 17 1609 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdlclkp_2
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 1471 94 1505 128 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1471 168 1505 202 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1477732
string GDS_START 1465172
<< end >>
