magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2494 1852
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 2 21 1164 203
rect 29 -17 63 21
<< scnmos >>
rect 90 47 120 177
rect 184 47 214 177
rect 382 47 412 177
rect 466 47 496 177
rect 570 47 600 177
rect 664 47 694 177
rect 774 47 804 177
rect 858 47 888 177
rect 962 47 992 177
rect 1056 47 1086 177
<< scpmoshvt >>
rect 82 297 118 497
rect 176 297 212 497
rect 374 297 410 497
rect 468 297 504 497
rect 562 297 598 497
rect 656 297 692 497
rect 766 297 802 497
rect 860 297 896 497
rect 954 297 990 497
rect 1048 297 1084 497
<< ndiff >>
rect 28 163 90 177
rect 28 129 36 163
rect 70 129 90 163
rect 28 95 90 129
rect 28 61 36 95
rect 70 61 90 95
rect 28 47 90 61
rect 120 163 184 177
rect 120 129 130 163
rect 164 129 184 163
rect 120 47 184 129
rect 214 163 266 177
rect 214 129 224 163
rect 258 129 266 163
rect 214 95 266 129
rect 214 61 224 95
rect 258 61 266 95
rect 214 47 266 61
rect 320 95 382 177
rect 320 61 328 95
rect 362 61 382 95
rect 320 47 382 61
rect 412 163 466 177
rect 412 129 422 163
rect 456 129 466 163
rect 412 47 466 129
rect 496 95 570 177
rect 496 61 516 95
rect 550 61 570 95
rect 496 47 570 61
rect 600 163 664 177
rect 600 129 610 163
rect 644 129 664 163
rect 600 47 664 129
rect 694 163 774 177
rect 694 129 713 163
rect 747 129 774 163
rect 694 95 774 129
rect 694 61 713 95
rect 747 61 774 95
rect 694 47 774 61
rect 804 95 858 177
rect 804 61 814 95
rect 848 61 858 95
rect 804 47 858 61
rect 888 163 962 177
rect 888 129 908 163
rect 942 129 962 163
rect 888 95 962 129
rect 888 61 908 95
rect 942 61 962 95
rect 888 47 962 61
rect 992 95 1056 177
rect 992 61 1002 95
rect 1036 61 1056 95
rect 992 47 1056 61
rect 1086 163 1138 177
rect 1086 129 1096 163
rect 1130 129 1138 163
rect 1086 95 1138 129
rect 1086 61 1096 95
rect 1130 61 1138 95
rect 1086 47 1138 61
<< pdiff >>
rect 28 483 82 497
rect 28 449 36 483
rect 70 449 82 483
rect 28 415 82 449
rect 28 381 36 415
rect 70 381 82 415
rect 28 347 82 381
rect 28 313 36 347
rect 70 313 82 347
rect 28 297 82 313
rect 118 477 176 497
rect 118 443 130 477
rect 164 443 176 477
rect 118 409 176 443
rect 118 375 130 409
rect 164 375 176 409
rect 118 341 176 375
rect 118 307 130 341
rect 164 307 176 341
rect 118 297 176 307
rect 212 477 374 497
rect 212 443 224 477
rect 258 443 328 477
rect 362 443 374 477
rect 212 297 374 443
rect 410 477 468 497
rect 410 443 422 477
rect 456 443 468 477
rect 410 297 468 443
rect 504 409 562 497
rect 504 375 516 409
rect 550 375 562 409
rect 504 297 562 375
rect 598 477 656 497
rect 598 443 610 477
rect 644 443 656 477
rect 598 297 656 443
rect 692 477 766 497
rect 692 443 704 477
rect 738 443 766 477
rect 692 297 766 443
rect 802 477 860 497
rect 802 443 814 477
rect 848 443 860 477
rect 802 297 860 443
rect 896 409 954 497
rect 896 375 908 409
rect 942 375 954 409
rect 896 297 954 375
rect 990 477 1048 497
rect 990 443 1002 477
rect 1036 443 1048 477
rect 990 409 1048 443
rect 990 375 1002 409
rect 1036 375 1048 409
rect 990 297 1048 375
rect 1084 477 1143 497
rect 1084 443 1097 477
rect 1131 443 1143 477
rect 1084 409 1143 443
rect 1084 375 1097 409
rect 1131 375 1143 409
rect 1084 341 1143 375
rect 1084 307 1097 341
rect 1131 307 1143 341
rect 1084 297 1143 307
<< ndiffc >>
rect 36 129 70 163
rect 36 61 70 95
rect 130 129 164 163
rect 224 129 258 163
rect 224 61 258 95
rect 328 61 362 95
rect 422 129 456 163
rect 516 61 550 95
rect 610 129 644 163
rect 713 129 747 163
rect 713 61 747 95
rect 814 61 848 95
rect 908 129 942 163
rect 908 61 942 95
rect 1002 61 1036 95
rect 1096 129 1130 163
rect 1096 61 1130 95
<< pdiffc >>
rect 36 449 70 483
rect 36 381 70 415
rect 36 313 70 347
rect 130 443 164 477
rect 130 375 164 409
rect 130 307 164 341
rect 224 443 258 477
rect 328 443 362 477
rect 422 443 456 477
rect 516 375 550 409
rect 610 443 644 477
rect 704 443 738 477
rect 814 443 848 477
rect 908 375 942 409
rect 1002 443 1036 477
rect 1002 375 1036 409
rect 1097 443 1131 477
rect 1097 375 1131 409
rect 1097 307 1131 341
<< poly >>
rect 82 497 118 523
rect 176 497 212 523
rect 374 497 410 523
rect 468 497 504 523
rect 562 497 598 523
rect 656 497 692 523
rect 766 497 802 523
rect 860 497 896 523
rect 954 497 990 523
rect 1048 497 1084 523
rect 82 282 118 297
rect 176 282 212 297
rect 374 282 410 297
rect 468 282 504 297
rect 562 282 598 297
rect 656 282 692 297
rect 766 282 802 297
rect 860 282 896 297
rect 954 282 990 297
rect 1048 282 1084 297
rect 80 265 120 282
rect 174 265 214 282
rect 372 265 412 282
rect 466 265 506 282
rect 560 265 600 282
rect 654 265 694 282
rect 764 265 804 282
rect 858 265 898 282
rect 952 265 992 282
rect 1046 265 1086 282
rect 21 249 214 265
rect 21 215 37 249
rect 71 215 214 249
rect 21 199 214 215
rect 360 249 424 265
rect 360 215 370 249
rect 404 215 424 249
rect 360 199 424 215
rect 466 249 600 265
rect 466 215 516 249
rect 550 215 600 249
rect 466 199 600 215
rect 642 249 706 265
rect 642 215 652 249
rect 686 215 706 249
rect 642 199 706 215
rect 752 249 816 265
rect 752 215 762 249
rect 796 215 816 249
rect 752 199 816 215
rect 858 249 992 265
rect 858 215 908 249
rect 942 215 992 249
rect 858 199 992 215
rect 1034 249 1098 265
rect 1034 215 1044 249
rect 1078 215 1098 249
rect 1034 199 1098 215
rect 90 177 120 199
rect 184 177 214 199
rect 382 177 412 199
rect 466 177 496 199
rect 570 177 600 199
rect 664 177 694 199
rect 774 177 804 199
rect 858 177 888 199
rect 962 177 992 199
rect 1056 177 1086 199
rect 90 21 120 47
rect 184 21 214 47
rect 382 21 412 47
rect 466 21 496 47
rect 570 21 600 47
rect 664 21 694 47
rect 774 21 804 47
rect 858 21 888 47
rect 962 21 992 47
rect 1056 21 1086 47
<< polycont >>
rect 37 215 71 249
rect 370 215 404 249
rect 516 215 550 249
rect 652 215 686 249
rect 762 215 796 249
rect 908 215 942 249
rect 1044 215 1078 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 28 483 78 527
rect 28 449 36 483
rect 70 449 78 483
rect 28 415 78 449
rect 28 381 36 415
rect 70 381 78 415
rect 28 347 78 381
rect 28 313 36 347
rect 70 313 78 347
rect 28 291 78 313
rect 122 477 172 493
rect 122 443 130 477
rect 164 443 172 477
rect 122 409 172 443
rect 216 477 370 527
rect 216 443 224 477
rect 258 443 328 477
rect 362 443 370 477
rect 216 425 370 443
rect 414 477 652 493
rect 414 443 422 477
rect 456 459 610 477
rect 456 443 464 459
rect 414 425 464 443
rect 602 443 610 459
rect 644 443 652 477
rect 602 425 652 443
rect 696 477 762 527
rect 696 443 704 477
rect 738 443 762 477
rect 696 425 762 443
rect 806 477 1044 493
rect 806 443 814 477
rect 848 459 1002 477
rect 848 443 856 459
rect 806 425 856 443
rect 994 443 1002 459
rect 1036 443 1044 477
rect 122 375 130 409
rect 164 391 172 409
rect 508 409 558 425
rect 508 391 516 409
rect 164 375 516 391
rect 550 391 558 409
rect 900 409 950 425
rect 900 391 908 409
rect 550 375 908 391
rect 942 375 950 409
rect 122 357 950 375
rect 994 409 1044 443
rect 994 375 1002 409
rect 1036 375 1044 409
rect 994 357 1044 375
rect 1097 477 1138 527
rect 1131 443 1138 477
rect 1097 409 1138 443
rect 1131 375 1138 409
rect 122 341 180 357
rect 122 307 130 341
rect 164 307 180 341
rect 1097 341 1138 375
rect 122 289 180 307
rect 17 249 87 255
rect 17 215 37 249
rect 71 215 87 249
rect 20 163 70 179
rect 131 173 180 289
rect 224 289 712 323
rect 224 249 437 289
rect 224 215 370 249
rect 404 215 437 249
rect 471 249 602 255
rect 471 215 516 249
rect 550 215 602 249
rect 636 249 712 289
rect 636 215 652 249
rect 686 215 712 249
rect 746 289 1053 323
rect 1131 307 1138 341
rect 1097 291 1138 307
rect 746 249 822 289
rect 1019 255 1053 289
rect 746 215 762 249
rect 796 215 822 249
rect 856 249 975 255
rect 856 215 908 249
rect 942 215 975 249
rect 1019 249 1167 255
rect 1019 215 1044 249
rect 1078 215 1167 249
rect 20 129 36 163
rect 104 163 180 173
rect 104 129 130 163
rect 164 129 180 163
rect 224 163 660 181
rect 258 129 422 163
rect 456 129 610 163
rect 644 129 660 163
rect 704 163 1146 181
rect 704 129 713 163
rect 747 147 908 163
rect 747 129 770 147
rect 20 95 70 129
rect 224 95 274 129
rect 704 95 770 129
rect 882 129 908 147
rect 942 145 1096 163
rect 942 129 958 145
rect 20 61 36 95
rect 70 61 224 95
rect 258 61 274 95
rect 20 51 274 61
rect 312 61 328 95
rect 362 61 516 95
rect 550 61 713 95
rect 747 61 770 95
rect 312 51 770 61
rect 814 95 848 111
rect 814 17 848 61
rect 882 95 958 129
rect 1070 129 1096 145
rect 1130 129 1146 163
rect 882 61 908 95
rect 942 61 958 95
rect 882 51 958 61
rect 1002 95 1036 111
rect 1002 17 1036 61
rect 1070 95 1146 129
rect 1070 61 1096 95
rect 1130 61 1146 95
rect 1070 51 1146 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 303 221 337 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 305 357 339 391 0 FreeSans 400 0 0 0 Y
port 10 nsew signal output
flabel locali s 941 221 975 255 0 FreeSans 400 180 0 0 A2
port 2 nsew signal input
flabel locali s 1019 255 1053 289 0 FreeSans 400 180 0 0 A1
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 C1
port 5 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221ai_2
rlabel locali s 1019 215 1167 255 1 A1
port 1 nsew signal input
rlabel locali s 746 289 1053 323 1 A1
port 1 nsew signal input
rlabel locali s 746 215 822 289 1 A1
port 1 nsew signal input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2519174
string GDS_START 2510028
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
