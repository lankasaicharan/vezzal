magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 4 248 488 258
rect 4 49 959 248
rect 0 0 960 49
<< scpmos >>
rect 89 368 125 592
rect 179 368 215 592
rect 269 368 305 592
rect 359 368 395 592
rect 561 368 597 592
rect 651 368 687 592
rect 741 368 777 592
rect 841 368 877 592
<< nmoslvt >>
rect 87 84 117 232
rect 173 84 203 232
rect 273 84 303 232
rect 373 84 403 232
rect 573 74 603 222
rect 659 74 689 222
rect 746 74 776 222
rect 841 74 871 222
<< ndiff >>
rect 30 220 87 232
rect 30 186 42 220
rect 76 186 87 220
rect 30 130 87 186
rect 30 96 42 130
rect 76 96 87 130
rect 30 84 87 96
rect 117 224 173 232
rect 117 190 128 224
rect 162 190 173 224
rect 117 153 173 190
rect 117 119 128 153
rect 162 119 173 153
rect 117 84 173 119
rect 203 220 273 232
rect 203 186 228 220
rect 262 186 273 220
rect 203 130 273 186
rect 203 96 228 130
rect 262 96 273 130
rect 203 84 273 96
rect 303 217 373 232
rect 303 183 328 217
rect 362 183 373 217
rect 303 84 373 183
rect 403 130 462 232
rect 403 96 415 130
rect 449 96 462 130
rect 403 84 462 96
rect 516 143 573 222
rect 516 109 528 143
rect 562 109 573 143
rect 516 74 573 109
rect 603 210 659 222
rect 603 176 614 210
rect 648 176 659 210
rect 603 120 659 176
rect 603 86 614 120
rect 648 86 659 120
rect 603 74 659 86
rect 689 143 746 222
rect 689 109 700 143
rect 734 109 746 143
rect 689 74 746 109
rect 776 210 841 222
rect 776 176 787 210
rect 821 176 841 210
rect 776 120 841 176
rect 776 86 787 120
rect 821 86 841 120
rect 776 74 841 86
rect 871 199 933 222
rect 871 165 882 199
rect 916 165 933 199
rect 871 120 933 165
rect 871 86 882 120
rect 916 86 933 120
rect 871 74 933 86
<< pdiff >>
rect 33 580 89 592
rect 33 546 45 580
rect 79 546 89 580
rect 33 510 89 546
rect 33 476 45 510
rect 79 476 89 510
rect 33 440 89 476
rect 33 406 45 440
rect 79 406 89 440
rect 33 368 89 406
rect 125 580 179 592
rect 125 546 135 580
rect 169 546 179 580
rect 125 510 179 546
rect 125 476 135 510
rect 169 476 179 510
rect 125 440 179 476
rect 125 406 135 440
rect 169 406 179 440
rect 125 368 179 406
rect 215 580 269 592
rect 215 546 225 580
rect 259 546 269 580
rect 215 508 269 546
rect 215 474 225 508
rect 259 474 269 508
rect 215 368 269 474
rect 305 580 359 592
rect 305 546 315 580
rect 349 546 359 580
rect 305 510 359 546
rect 305 476 315 510
rect 349 476 359 510
rect 305 440 359 476
rect 305 406 315 440
rect 349 406 359 440
rect 305 368 359 406
rect 395 580 451 592
rect 395 546 405 580
rect 439 546 451 580
rect 395 508 451 546
rect 395 474 405 508
rect 439 474 451 508
rect 395 368 451 474
rect 505 580 561 592
rect 505 546 517 580
rect 551 546 561 580
rect 505 508 561 546
rect 505 474 517 508
rect 551 474 561 508
rect 505 368 561 474
rect 597 531 651 592
rect 597 497 607 531
rect 641 497 651 531
rect 597 440 651 497
rect 597 406 607 440
rect 641 406 651 440
rect 597 368 651 406
rect 687 580 741 592
rect 687 546 697 580
rect 731 546 741 580
rect 687 497 741 546
rect 687 463 697 497
rect 731 463 741 497
rect 687 414 741 463
rect 687 380 697 414
rect 731 380 741 414
rect 687 368 741 380
rect 777 580 841 592
rect 777 546 787 580
rect 821 546 841 580
rect 777 482 841 546
rect 777 448 787 482
rect 821 448 841 482
rect 777 368 841 448
rect 877 580 933 592
rect 877 546 887 580
rect 921 546 933 580
rect 877 497 933 546
rect 877 463 887 497
rect 921 463 933 497
rect 877 414 933 463
rect 877 380 887 414
rect 921 380 933 414
rect 877 368 933 380
<< ndiffc >>
rect 42 186 76 220
rect 42 96 76 130
rect 128 190 162 224
rect 128 119 162 153
rect 228 186 262 220
rect 228 96 262 130
rect 328 183 362 217
rect 415 96 449 130
rect 528 109 562 143
rect 614 176 648 210
rect 614 86 648 120
rect 700 109 734 143
rect 787 176 821 210
rect 787 86 821 120
rect 882 165 916 199
rect 882 86 916 120
<< pdiffc >>
rect 45 546 79 580
rect 45 476 79 510
rect 45 406 79 440
rect 135 546 169 580
rect 135 476 169 510
rect 135 406 169 440
rect 225 546 259 580
rect 225 474 259 508
rect 315 546 349 580
rect 315 476 349 510
rect 315 406 349 440
rect 405 546 439 580
rect 405 474 439 508
rect 517 546 551 580
rect 517 474 551 508
rect 607 497 641 531
rect 607 406 641 440
rect 697 546 731 580
rect 697 463 731 497
rect 697 380 731 414
rect 787 546 821 580
rect 787 448 821 482
rect 887 546 921 580
rect 887 463 921 497
rect 887 380 921 414
<< poly >>
rect 89 592 125 618
rect 179 592 215 618
rect 269 592 305 618
rect 359 592 395 618
rect 561 592 597 618
rect 651 592 687 618
rect 741 592 777 618
rect 841 592 877 618
rect 89 336 125 368
rect 44 326 125 336
rect 179 326 215 368
rect 44 320 215 326
rect 44 286 60 320
rect 94 286 215 320
rect 44 270 215 286
rect 269 336 305 368
rect 359 336 395 368
rect 269 320 403 336
rect 561 330 597 368
rect 651 330 687 368
rect 741 330 777 368
rect 841 330 877 368
rect 269 286 285 320
rect 319 286 353 320
rect 387 286 403 320
rect 269 270 403 286
rect 87 232 117 270
rect 173 232 203 270
rect 273 232 303 270
rect 373 232 403 270
rect 487 314 689 330
rect 487 280 503 314
rect 537 280 571 314
rect 605 280 639 314
rect 673 280 689 314
rect 487 264 689 280
rect 573 222 603 264
rect 659 222 689 264
rect 737 326 877 330
rect 737 314 939 326
rect 737 280 753 314
rect 787 280 821 314
rect 855 310 939 314
rect 855 280 889 310
rect 737 276 889 280
rect 923 276 939 310
rect 737 260 939 276
rect 746 222 776 260
rect 841 222 871 260
rect 87 58 117 84
rect 173 58 203 84
rect 273 58 303 84
rect 373 58 403 84
rect 573 48 603 74
rect 659 48 689 74
rect 746 48 776 74
rect 841 48 871 74
<< polycont >>
rect 60 286 94 320
rect 285 286 319 320
rect 353 286 387 320
rect 503 280 537 314
rect 571 280 605 314
rect 639 280 673 314
rect 753 280 787 314
rect 821 280 855 314
rect 889 276 923 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 29 580 79 649
rect 29 546 45 580
rect 29 510 79 546
rect 29 476 45 510
rect 29 440 79 476
rect 29 406 45 440
rect 29 390 79 406
rect 119 580 185 596
rect 119 546 135 580
rect 169 546 185 580
rect 119 510 185 546
rect 119 476 135 510
rect 169 476 185 510
rect 119 440 185 476
rect 225 580 259 649
rect 225 508 259 546
rect 225 458 259 474
rect 299 580 365 596
rect 299 546 315 580
rect 349 546 365 580
rect 299 510 365 546
rect 299 476 315 510
rect 349 476 365 510
rect 119 406 135 440
rect 169 424 185 440
rect 299 440 365 476
rect 405 580 455 649
rect 439 546 455 580
rect 405 508 455 546
rect 439 474 455 508
rect 405 458 455 474
rect 501 581 731 615
rect 501 580 551 581
rect 501 546 517 580
rect 697 580 731 581
rect 501 508 551 546
rect 501 474 517 508
rect 501 458 551 474
rect 591 531 657 547
rect 591 497 607 531
rect 641 497 657 531
rect 299 424 315 440
rect 169 406 315 424
rect 349 424 365 440
rect 591 440 657 497
rect 591 424 607 440
rect 349 406 607 424
rect 641 406 657 440
rect 119 390 657 406
rect 697 497 731 546
rect 697 414 731 463
rect 771 580 837 649
rect 771 546 787 580
rect 821 546 837 580
rect 771 482 837 546
rect 771 448 787 482
rect 821 448 837 482
rect 771 432 837 448
rect 871 580 937 596
rect 871 546 887 580
rect 921 546 937 580
rect 871 497 937 546
rect 871 463 887 497
rect 921 463 937 497
rect 25 320 110 356
rect 25 286 60 320
rect 94 286 110 320
rect 25 270 110 286
rect 144 236 178 390
rect 871 414 937 463
rect 871 398 887 414
rect 731 380 887 398
rect 921 380 937 414
rect 697 364 937 380
rect 217 320 403 356
rect 217 286 285 320
rect 319 286 353 320
rect 387 286 403 320
rect 217 270 403 286
rect 487 330 647 356
rect 487 314 689 330
rect 487 280 503 314
rect 537 280 571 314
rect 605 280 639 314
rect 673 280 689 314
rect 487 264 689 280
rect 737 314 939 330
rect 737 280 753 314
rect 787 280 821 314
rect 855 310 939 314
rect 855 280 889 310
rect 737 276 889 280
rect 923 276 939 310
rect 737 264 939 276
rect 873 236 939 264
rect 26 220 76 236
rect 26 186 42 220
rect 26 130 76 186
rect 26 96 42 130
rect 112 224 178 236
rect 112 190 128 224
rect 162 190 178 224
rect 112 153 178 190
rect 112 119 128 153
rect 162 119 178 153
rect 212 220 278 236
rect 212 186 228 220
rect 262 186 278 220
rect 212 146 278 186
rect 312 230 378 236
rect 312 217 832 230
rect 312 183 328 217
rect 362 210 832 217
rect 362 196 614 210
rect 362 183 378 196
rect 312 180 378 183
rect 648 196 787 210
rect 212 130 466 146
rect 26 85 76 96
rect 212 96 228 130
rect 262 96 415 130
rect 449 96 466 130
rect 212 85 466 96
rect 26 51 466 85
rect 512 143 578 159
rect 512 109 528 143
rect 562 109 578 143
rect 512 17 578 109
rect 614 120 648 176
rect 821 176 832 210
rect 614 70 648 86
rect 684 143 750 159
rect 684 109 700 143
rect 734 109 750 143
rect 684 17 750 109
rect 787 120 832 176
rect 821 86 832 120
rect 787 70 832 86
rect 866 199 937 202
rect 866 165 882 199
rect 916 165 937 199
rect 866 120 937 165
rect 866 86 882 120
rect 916 86 937 120
rect 866 17 937 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o211ai_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 3862434
string GDS_START 3853508
<< end >>
