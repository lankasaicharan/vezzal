magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 572 157 951 241
rect 14 49 951 157
rect 0 0 960 49
<< scnmos >>
rect 93 47 123 131
rect 246 47 276 131
rect 332 47 362 131
rect 462 47 492 131
rect 548 47 578 131
rect 651 47 681 215
rect 737 47 767 215
rect 842 131 872 215
<< scpmoshvt >>
rect 160 403 190 487
rect 246 403 276 487
rect 318 403 348 487
rect 390 403 420 487
rect 462 403 492 487
rect 658 367 688 619
rect 744 367 774 619
rect 849 367 879 451
<< ndiff >>
rect 598 187 651 215
rect 598 153 606 187
rect 640 153 651 187
rect 598 131 651 153
rect 40 106 93 131
rect 40 72 48 106
rect 82 72 93 106
rect 40 47 93 72
rect 123 105 246 131
rect 123 71 201 105
rect 235 71 246 105
rect 123 47 246 71
rect 276 103 332 131
rect 276 69 287 103
rect 321 69 332 103
rect 276 47 332 69
rect 362 81 462 131
rect 362 47 389 81
rect 423 47 462 81
rect 492 106 548 131
rect 492 72 503 106
rect 537 72 548 106
rect 492 47 548 72
rect 578 93 651 131
rect 578 59 606 93
rect 640 59 651 93
rect 578 47 651 59
rect 681 203 737 215
rect 681 169 692 203
rect 726 169 737 203
rect 681 101 737 169
rect 681 67 692 101
rect 726 67 737 101
rect 681 47 737 67
rect 767 163 842 215
rect 767 129 778 163
rect 812 131 842 163
rect 872 190 925 215
rect 872 156 883 190
rect 917 156 925 190
rect 872 131 925 156
rect 812 129 820 131
rect 767 93 820 129
rect 767 59 778 93
rect 812 59 820 93
rect 767 47 820 59
rect 377 39 435 47
<< pdiff >>
rect 107 462 160 487
rect 107 428 115 462
rect 149 428 160 462
rect 107 403 160 428
rect 190 462 246 487
rect 190 428 201 462
rect 235 428 246 462
rect 190 403 246 428
rect 276 403 318 487
rect 348 403 390 487
rect 420 403 462 487
rect 492 449 545 487
rect 492 415 503 449
rect 537 415 545 449
rect 492 403 545 415
rect 605 595 658 619
rect 605 561 613 595
rect 647 561 658 595
rect 605 367 658 561
rect 688 439 744 619
rect 688 405 699 439
rect 733 405 744 439
rect 688 367 744 405
rect 774 595 827 619
rect 774 561 785 595
rect 819 561 827 595
rect 774 451 827 561
rect 774 367 849 451
rect 879 428 932 451
rect 879 394 890 428
rect 924 394 932 428
rect 879 367 932 394
<< ndiffc >>
rect 606 153 640 187
rect 48 72 82 106
rect 201 71 235 105
rect 287 69 321 103
rect 389 47 423 81
rect 503 72 537 106
rect 606 59 640 93
rect 692 169 726 203
rect 692 67 726 101
rect 778 129 812 163
rect 883 156 917 190
rect 778 59 812 93
<< pdiffc >>
rect 115 428 149 462
rect 201 428 235 462
rect 503 415 537 449
rect 613 561 647 595
rect 699 405 733 439
rect 785 561 819 595
rect 890 394 924 428
<< poly >>
rect 495 605 590 621
rect 658 619 688 645
rect 744 619 774 645
rect 495 571 511 605
rect 545 571 590 605
rect 495 555 590 571
rect 160 487 190 513
rect 246 487 276 513
rect 318 487 348 513
rect 390 487 420 513
rect 462 487 492 513
rect 160 367 190 403
rect 93 337 190 367
rect 93 287 123 337
rect 246 289 276 403
rect 93 271 168 287
rect 93 237 118 271
rect 152 237 168 271
rect 93 203 168 237
rect 93 169 118 203
rect 152 169 168 203
rect 93 153 168 169
rect 210 273 276 289
rect 210 239 226 273
rect 260 239 276 273
rect 210 205 276 239
rect 210 171 226 205
rect 260 171 276 205
rect 318 237 348 403
rect 390 309 420 403
rect 462 381 492 403
rect 560 381 590 555
rect 462 351 590 381
rect 849 451 879 477
rect 390 293 492 309
rect 390 279 442 293
rect 426 259 442 279
rect 476 259 492 293
rect 318 221 384 237
rect 318 187 334 221
rect 368 187 384 221
rect 318 171 384 187
rect 426 225 492 259
rect 426 191 442 225
rect 476 191 492 225
rect 426 175 492 191
rect 210 155 276 171
rect 93 131 123 153
rect 246 131 276 155
rect 332 131 362 171
rect 462 131 492 175
rect 534 189 564 351
rect 658 345 688 367
rect 651 315 688 345
rect 651 303 681 315
rect 606 287 681 303
rect 606 253 622 287
rect 656 267 681 287
rect 744 267 774 367
rect 849 335 879 367
rect 656 253 774 267
rect 606 237 774 253
rect 842 319 909 335
rect 842 285 859 319
rect 893 285 909 319
rect 842 269 909 285
rect 651 215 681 237
rect 737 215 767 237
rect 842 215 872 269
rect 534 159 578 189
rect 548 131 578 159
rect 842 105 872 131
rect 93 21 123 47
rect 246 21 276 47
rect 332 21 362 47
rect 462 21 492 47
rect 548 21 578 47
rect 651 21 681 47
rect 737 21 767 47
<< polycont >>
rect 511 571 545 605
rect 118 237 152 271
rect 118 169 152 203
rect 226 239 260 273
rect 226 171 260 205
rect 442 259 476 293
rect 334 187 368 221
rect 442 191 476 225
rect 622 253 656 287
rect 859 285 893 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 99 462 158 478
rect 99 428 115 462
rect 149 428 158 462
rect 99 359 158 428
rect 192 462 251 649
rect 495 605 561 615
rect 495 571 511 605
rect 545 571 561 605
rect 495 523 561 571
rect 597 595 663 649
rect 597 561 613 595
rect 647 561 663 595
rect 597 557 663 561
rect 769 595 835 649
rect 769 561 785 595
rect 819 561 835 595
rect 769 557 835 561
rect 495 489 841 523
rect 192 428 201 462
rect 235 428 251 462
rect 192 409 251 428
rect 487 449 562 455
rect 487 415 503 449
rect 537 415 562 449
rect 487 399 562 415
rect 32 325 492 359
rect 32 106 82 325
rect 426 293 492 325
rect 32 72 48 106
rect 116 271 163 287
rect 116 237 118 271
rect 152 237 163 271
rect 116 203 163 237
rect 116 169 118 203
rect 152 169 163 203
rect 116 94 163 169
rect 207 273 262 289
rect 207 239 226 273
rect 260 239 262 273
rect 207 205 262 239
rect 207 171 226 205
rect 260 171 262 205
rect 300 221 384 291
rect 300 187 334 221
rect 368 187 384 221
rect 300 185 384 187
rect 426 259 442 293
rect 476 259 492 293
rect 426 225 492 259
rect 426 191 442 225
rect 476 191 492 225
rect 426 185 492 191
rect 528 303 562 399
rect 690 439 739 455
rect 690 405 699 439
rect 733 405 739 439
rect 528 287 656 303
rect 528 253 622 287
rect 528 237 656 253
rect 207 155 262 171
rect 528 151 562 237
rect 690 203 739 405
rect 773 452 841 489
rect 773 428 940 452
rect 773 394 890 428
rect 924 394 940 428
rect 773 386 940 394
rect 773 247 807 386
rect 843 319 943 352
rect 843 285 859 319
rect 893 285 943 319
rect 843 281 943 285
rect 773 213 933 247
rect 197 105 249 121
rect 296 119 562 151
rect 32 56 82 72
rect 197 71 201 105
rect 235 71 249 105
rect 197 17 249 71
rect 283 117 562 119
rect 283 103 330 117
rect 283 69 287 103
rect 321 69 330 103
rect 487 106 562 117
rect 283 53 330 69
rect 373 81 439 83
rect 373 47 389 81
rect 423 47 439 81
rect 487 72 503 106
rect 537 72 562 106
rect 487 56 562 72
rect 596 187 656 203
rect 596 153 606 187
rect 640 153 656 187
rect 596 93 656 153
rect 596 59 606 93
rect 640 59 656 93
rect 373 17 439 47
rect 596 17 656 59
rect 690 169 692 203
rect 726 169 739 203
rect 867 190 933 213
rect 690 101 739 169
rect 690 67 692 101
rect 726 67 739 101
rect 690 51 739 67
rect 773 163 828 179
rect 773 129 778 163
rect 812 129 828 163
rect 867 156 883 190
rect 917 156 933 190
rect 867 140 933 156
rect 773 93 828 129
rect 773 59 778 93
rect 812 59 828 93
rect 773 17 828 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or4bb_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6658578
string GDS_START 6650180
<< end >>
