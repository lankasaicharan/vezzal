magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 15 49 855 157
rect 0 0 864 49
<< scnmos >>
rect 98 47 128 131
rect 176 47 206 131
rect 284 47 314 131
rect 398 47 428 131
rect 512 47 542 131
rect 584 47 614 131
rect 670 47 700 131
rect 742 47 772 131
<< scpmoshvt >>
rect 84 409 134 609
rect 190 409 240 609
rect 296 409 346 609
rect 406 409 456 609
rect 512 409 562 609
rect 730 409 780 609
<< ndiff >>
rect 41 103 98 131
rect 41 69 53 103
rect 87 69 98 103
rect 41 47 98 69
rect 128 47 176 131
rect 206 47 284 131
rect 314 47 398 131
rect 428 111 512 131
rect 428 77 467 111
rect 501 77 512 111
rect 428 47 512 77
rect 542 47 584 131
rect 614 93 670 131
rect 614 59 625 93
rect 659 59 670 93
rect 614 47 670 59
rect 700 47 742 131
rect 772 111 829 131
rect 772 77 783 111
rect 817 77 829 111
rect 772 47 829 77
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 190 609
rect 134 563 145 597
rect 179 563 190 597
rect 134 526 190 563
rect 134 492 145 526
rect 179 492 190 526
rect 134 455 190 492
rect 134 421 145 455
rect 179 421 190 455
rect 134 409 190 421
rect 240 597 296 609
rect 240 563 251 597
rect 285 563 296 597
rect 240 526 296 563
rect 240 492 251 526
rect 285 492 296 526
rect 240 455 296 492
rect 240 421 251 455
rect 285 421 296 455
rect 240 409 296 421
rect 346 597 406 609
rect 346 563 357 597
rect 391 563 406 597
rect 346 505 406 563
rect 346 471 357 505
rect 391 471 406 505
rect 346 409 406 471
rect 456 597 512 609
rect 456 563 467 597
rect 501 563 512 597
rect 456 526 512 563
rect 456 492 467 526
rect 501 492 512 526
rect 456 455 512 492
rect 456 421 467 455
rect 501 421 512 455
rect 456 409 512 421
rect 562 597 619 609
rect 562 563 573 597
rect 607 563 619 597
rect 562 526 619 563
rect 562 492 573 526
rect 607 492 619 526
rect 562 455 619 492
rect 562 421 573 455
rect 607 421 619 455
rect 562 409 619 421
rect 673 597 730 609
rect 673 563 685 597
rect 719 563 730 597
rect 673 505 730 563
rect 673 471 685 505
rect 719 471 730 505
rect 673 409 730 471
rect 780 597 837 609
rect 780 563 791 597
rect 825 563 837 597
rect 780 526 837 563
rect 780 492 791 526
rect 825 492 837 526
rect 780 455 837 492
rect 780 421 791 455
rect 825 421 837 455
rect 780 409 837 421
<< ndiffc >>
rect 53 69 87 103
rect 467 77 501 111
rect 625 59 659 93
rect 783 77 817 111
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 492 179 526
rect 145 421 179 455
rect 251 563 285 597
rect 251 492 285 526
rect 251 421 285 455
rect 357 563 391 597
rect 357 471 391 505
rect 467 563 501 597
rect 467 492 501 526
rect 467 421 501 455
rect 573 563 607 597
rect 573 492 607 526
rect 573 421 607 455
rect 685 563 719 597
rect 685 471 719 505
rect 791 563 825 597
rect 791 492 825 526
rect 791 421 825 455
<< poly >>
rect 84 609 134 635
rect 190 609 240 635
rect 296 609 346 635
rect 406 609 456 635
rect 512 609 562 635
rect 730 609 780 635
rect 84 299 134 409
rect 21 283 114 299
rect 190 287 240 409
rect 296 287 346 409
rect 406 349 456 409
rect 512 349 562 409
rect 398 333 464 349
rect 398 299 414 333
rect 448 299 464 333
rect 21 249 37 283
rect 71 249 114 283
rect 21 215 114 249
rect 21 181 37 215
rect 71 195 114 215
rect 176 271 242 287
rect 176 237 192 271
rect 226 237 242 271
rect 176 203 242 237
rect 71 181 128 195
rect 21 165 128 181
rect 98 131 128 165
rect 176 169 192 203
rect 226 169 242 203
rect 176 153 242 169
rect 284 271 350 287
rect 284 237 300 271
rect 334 237 350 271
rect 284 203 350 237
rect 284 169 300 203
rect 334 169 350 203
rect 284 153 350 169
rect 398 265 464 299
rect 398 231 414 265
rect 448 231 464 265
rect 532 333 614 349
rect 532 299 548 333
rect 582 299 614 333
rect 532 265 614 299
rect 730 287 780 409
rect 532 245 548 265
rect 398 215 464 231
rect 512 231 548 245
rect 582 231 614 265
rect 512 215 614 231
rect 176 131 206 153
rect 284 131 314 153
rect 398 131 428 215
rect 512 131 542 215
rect 584 131 614 215
rect 665 271 780 287
rect 665 237 681 271
rect 715 237 780 271
rect 665 203 780 237
rect 665 169 681 203
rect 715 169 780 203
rect 665 153 780 169
rect 670 131 700 153
rect 742 131 772 153
rect 98 21 128 47
rect 176 21 206 47
rect 284 21 314 47
rect 398 21 428 47
rect 512 21 542 47
rect 584 21 614 47
rect 670 21 700 47
rect 742 21 772 47
<< polycont >>
rect 414 299 448 333
rect 37 249 71 283
rect 37 181 71 215
rect 192 237 226 271
rect 192 169 226 203
rect 300 237 334 271
rect 300 169 334 203
rect 414 231 448 265
rect 548 299 582 333
rect 548 231 582 265
rect 681 237 715 271
rect 681 169 715 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 526 89 563
rect 23 492 39 526
rect 73 492 89 526
rect 23 455 89 492
rect 23 421 39 455
rect 73 421 89 455
rect 23 369 89 421
rect 129 597 195 649
rect 129 563 145 597
rect 179 563 195 597
rect 129 526 195 563
rect 129 492 145 526
rect 179 492 195 526
rect 129 455 195 492
rect 129 421 145 455
rect 179 421 195 455
rect 129 405 195 421
rect 235 597 301 613
rect 235 563 251 597
rect 285 563 301 597
rect 235 526 301 563
rect 235 492 251 526
rect 285 492 301 526
rect 235 455 301 492
rect 341 597 407 649
rect 341 563 357 597
rect 391 563 407 597
rect 341 505 407 563
rect 341 471 357 505
rect 391 471 407 505
rect 341 455 407 471
rect 451 597 517 613
rect 451 563 467 597
rect 501 563 517 597
rect 451 526 517 563
rect 451 492 467 526
rect 501 492 517 526
rect 451 455 517 492
rect 235 421 251 455
rect 285 421 301 455
rect 235 419 301 421
rect 451 421 467 455
rect 501 421 517 455
rect 451 419 517 421
rect 235 385 517 419
rect 557 597 623 613
rect 557 563 573 597
rect 607 563 623 597
rect 557 526 623 563
rect 557 492 573 526
rect 607 492 623 526
rect 557 455 623 492
rect 669 597 735 649
rect 669 563 685 597
rect 719 563 735 597
rect 669 505 735 563
rect 669 471 685 505
rect 719 471 735 505
rect 669 455 735 471
rect 775 597 841 613
rect 775 563 791 597
rect 825 563 841 597
rect 775 526 841 563
rect 775 492 791 526
rect 825 492 841 526
rect 775 455 841 492
rect 557 421 573 455
rect 607 421 623 455
rect 557 419 623 421
rect 775 421 791 455
rect 825 421 841 455
rect 557 385 731 419
rect 235 369 301 385
rect 23 335 301 369
rect 398 333 464 349
rect 398 299 414 333
rect 448 299 464 333
rect 21 283 87 299
rect 21 249 37 283
rect 71 249 87 283
rect 21 215 87 249
rect 21 181 37 215
rect 71 181 87 215
rect 21 165 87 181
rect 123 271 242 287
rect 123 237 192 271
rect 226 237 242 271
rect 123 203 242 237
rect 123 169 192 203
rect 226 169 242 203
rect 37 103 87 129
rect 37 69 53 103
rect 123 88 242 169
rect 284 271 359 287
rect 284 237 300 271
rect 334 237 359 271
rect 284 203 359 237
rect 398 265 464 299
rect 398 231 414 265
rect 448 231 464 265
rect 398 215 464 231
rect 505 333 598 349
rect 505 299 548 333
rect 582 299 598 333
rect 505 265 598 299
rect 505 231 548 265
rect 582 231 598 265
rect 505 215 598 231
rect 665 271 731 385
rect 665 237 681 271
rect 715 237 731 271
rect 284 169 300 203
rect 334 169 359 203
rect 665 203 731 237
rect 665 179 681 203
rect 284 88 359 169
rect 451 169 681 179
rect 715 169 731 203
rect 451 145 731 169
rect 451 111 517 145
rect 775 135 841 421
rect 37 17 87 69
rect 451 77 467 111
rect 501 77 517 111
rect 767 111 841 135
rect 451 53 517 77
rect 609 93 675 109
rect 609 59 625 93
rect 659 59 675 93
rect 609 17 675 59
rect 767 77 783 111
rect 817 77 841 111
rect 767 53 841 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a41o_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6634410
string GDS_START 6625596
<< end >>
