magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 693 248 1151 258
rect 206 228 1151 248
rect 1 49 1151 228
rect 0 0 1152 49
<< scnmos >>
rect 84 74 114 202
rect 282 74 312 222
rect 374 74 404 222
rect 460 74 490 222
rect 578 74 608 222
rect 776 84 806 232
rect 862 84 892 232
rect 948 84 978 232
rect 1038 84 1068 232
<< scpmoshvt >>
rect 164 368 194 568
rect 272 368 302 592
rect 362 368 392 592
rect 525 368 555 592
rect 615 368 645 592
rect 725 368 755 592
rect 815 368 845 592
rect 945 368 975 592
rect 1035 368 1065 592
<< ndiff >>
rect 27 153 84 202
rect 27 119 39 153
rect 73 119 84 153
rect 27 74 84 119
rect 114 146 164 202
rect 114 127 171 146
rect 232 138 282 222
rect 114 93 125 127
rect 159 93 171 127
rect 114 74 171 93
rect 225 123 282 138
rect 225 89 237 123
rect 271 89 282 123
rect 225 74 282 89
rect 312 210 374 222
rect 312 176 326 210
rect 360 176 374 210
rect 312 74 374 176
rect 404 136 460 222
rect 404 102 415 136
rect 449 102 460 136
rect 404 74 460 102
rect 490 100 578 222
rect 490 74 517 100
rect 505 66 517 74
rect 551 74 578 100
rect 608 180 658 222
rect 719 194 776 232
rect 608 160 665 180
rect 608 126 619 160
rect 653 126 665 160
rect 608 107 665 126
rect 719 160 731 194
rect 765 160 776 194
rect 719 123 776 160
rect 608 74 658 107
rect 726 84 776 123
rect 806 133 862 232
rect 806 99 817 133
rect 851 99 862 133
rect 806 84 862 99
rect 892 220 948 232
rect 892 186 903 220
rect 937 186 948 220
rect 892 130 948 186
rect 892 96 903 130
rect 937 96 948 130
rect 892 84 948 96
rect 978 133 1038 232
rect 978 99 989 133
rect 1023 99 1038 133
rect 978 84 1038 99
rect 1068 220 1125 232
rect 1068 186 1079 220
rect 1113 186 1125 220
rect 1068 130 1125 186
rect 1068 96 1079 130
rect 1113 96 1125 130
rect 1068 84 1125 96
rect 551 66 563 74
rect 505 54 563 66
<< pdiff >>
rect 212 574 272 592
rect 212 568 224 574
rect 105 556 164 568
rect 105 522 117 556
rect 151 522 164 556
rect 105 485 164 522
rect 105 451 117 485
rect 151 451 164 485
rect 105 414 164 451
rect 105 380 117 414
rect 151 380 164 414
rect 105 368 164 380
rect 194 540 224 568
rect 258 540 272 574
rect 194 506 272 540
rect 194 472 224 506
rect 258 472 272 506
rect 194 438 272 472
rect 194 404 224 438
rect 258 404 272 438
rect 194 368 272 404
rect 302 580 362 592
rect 302 546 315 580
rect 349 546 362 580
rect 302 500 362 546
rect 302 466 315 500
rect 349 466 362 500
rect 302 420 362 466
rect 302 386 315 420
rect 349 386 362 420
rect 302 368 362 386
rect 392 580 525 592
rect 392 546 405 580
rect 439 546 478 580
rect 512 546 525 580
rect 392 508 525 546
rect 392 474 405 508
rect 439 474 478 508
rect 512 474 525 508
rect 392 368 525 474
rect 555 580 615 592
rect 555 546 568 580
rect 602 546 615 580
rect 555 497 615 546
rect 555 463 568 497
rect 602 463 615 497
rect 555 414 615 463
rect 555 380 568 414
rect 602 380 615 414
rect 555 368 615 380
rect 645 580 725 592
rect 645 546 668 580
rect 702 546 725 580
rect 645 500 725 546
rect 645 466 668 500
rect 702 466 725 500
rect 645 368 725 466
rect 755 580 815 592
rect 755 546 768 580
rect 802 546 815 580
rect 755 500 815 546
rect 755 466 768 500
rect 802 466 815 500
rect 755 424 815 466
rect 755 390 768 424
rect 802 390 815 424
rect 755 368 815 390
rect 845 580 945 592
rect 845 546 880 580
rect 914 546 945 580
rect 845 499 945 546
rect 845 465 880 499
rect 914 465 945 499
rect 845 368 945 465
rect 975 580 1035 592
rect 975 546 988 580
rect 1022 546 1035 580
rect 975 500 1035 546
rect 975 466 988 500
rect 1022 466 1035 500
rect 975 424 1035 466
rect 975 390 988 424
rect 1022 390 1035 424
rect 975 368 1035 390
rect 1065 580 1125 592
rect 1065 546 1078 580
rect 1112 546 1125 580
rect 1065 508 1125 546
rect 1065 474 1078 508
rect 1112 474 1125 508
rect 1065 440 1125 474
rect 1065 406 1078 440
rect 1112 406 1125 440
rect 1065 368 1125 406
<< ndiffc >>
rect 39 119 73 153
rect 125 93 159 127
rect 237 89 271 123
rect 326 176 360 210
rect 415 102 449 136
rect 517 66 551 100
rect 619 126 653 160
rect 731 160 765 194
rect 817 99 851 133
rect 903 186 937 220
rect 903 96 937 130
rect 989 99 1023 133
rect 1079 186 1113 220
rect 1079 96 1113 130
<< pdiffc >>
rect 117 522 151 556
rect 117 451 151 485
rect 117 380 151 414
rect 224 540 258 574
rect 224 472 258 506
rect 224 404 258 438
rect 315 546 349 580
rect 315 466 349 500
rect 315 386 349 420
rect 405 546 439 580
rect 478 546 512 580
rect 405 474 439 508
rect 478 474 512 508
rect 568 546 602 580
rect 568 463 602 497
rect 568 380 602 414
rect 668 546 702 580
rect 668 466 702 500
rect 768 546 802 580
rect 768 466 802 500
rect 768 390 802 424
rect 880 546 914 580
rect 880 465 914 499
rect 988 546 1022 580
rect 988 466 1022 500
rect 988 390 1022 424
rect 1078 546 1112 580
rect 1078 474 1112 508
rect 1078 406 1112 440
<< poly >>
rect 164 568 194 594
rect 272 592 302 618
rect 362 592 392 618
rect 525 592 555 618
rect 615 592 645 618
rect 725 592 755 618
rect 815 592 845 618
rect 945 592 975 618
rect 1035 592 1065 618
rect 164 353 194 368
rect 272 353 302 368
rect 362 353 392 368
rect 525 353 555 368
rect 615 353 645 368
rect 725 353 755 368
rect 815 353 845 368
rect 945 353 975 368
rect 1035 353 1065 368
rect 161 302 197 353
rect 63 286 197 302
rect 63 252 79 286
rect 113 252 147 286
rect 181 252 197 286
rect 269 336 305 353
rect 359 336 395 353
rect 522 336 558 353
rect 612 336 648 353
rect 722 336 758 353
rect 812 336 848 353
rect 945 336 978 353
rect 1032 336 1068 353
rect 269 320 404 336
rect 269 286 294 320
rect 328 286 404 320
rect 269 270 404 286
rect 452 320 648 336
rect 452 286 468 320
rect 502 286 648 320
rect 452 270 648 286
rect 705 320 848 336
rect 705 286 721 320
rect 755 286 789 320
rect 823 300 848 320
rect 948 320 1068 336
rect 823 286 892 300
rect 705 270 892 286
rect 63 236 197 252
rect 84 202 114 236
rect 282 222 312 270
rect 374 222 404 270
rect 460 222 490 270
rect 578 222 608 270
rect 776 232 806 270
rect 862 232 892 270
rect 948 286 964 320
rect 998 286 1068 320
rect 948 270 1068 286
rect 948 232 978 270
rect 1038 232 1068 270
rect 84 48 114 74
rect 282 48 312 74
rect 374 48 404 74
rect 460 48 490 74
rect 578 48 608 74
rect 776 58 806 84
rect 862 58 892 84
rect 948 58 978 84
rect 1038 58 1068 84
<< polycont >>
rect 79 252 113 286
rect 147 252 181 286
rect 294 286 328 320
rect 468 286 502 320
rect 721 286 755 320
rect 789 286 823 320
rect 964 286 998 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 208 574 274 649
rect 101 556 167 572
rect 101 522 117 556
rect 151 522 167 556
rect 101 485 167 522
rect 101 451 117 485
rect 151 451 167 485
rect 101 414 167 451
rect 101 380 117 414
rect 151 380 167 414
rect 208 540 224 574
rect 258 540 274 574
rect 208 506 274 540
rect 208 472 224 506
rect 258 472 274 506
rect 208 438 274 472
rect 208 404 224 438
rect 258 404 274 438
rect 310 580 365 596
rect 310 546 315 580
rect 349 546 365 580
rect 310 500 365 546
rect 310 466 315 500
rect 349 466 365 500
rect 310 424 365 466
rect 399 580 518 649
rect 399 546 405 580
rect 439 546 478 580
rect 512 546 518 580
rect 399 508 518 546
rect 399 474 405 508
rect 439 474 478 508
rect 512 474 518 508
rect 399 458 518 474
rect 552 580 618 596
rect 552 546 568 580
rect 602 546 618 580
rect 552 497 618 546
rect 552 463 568 497
rect 602 463 618 497
rect 552 424 618 463
rect 652 580 718 649
rect 652 546 668 580
rect 702 546 718 580
rect 652 500 718 546
rect 652 466 668 500
rect 702 466 718 500
rect 652 458 718 466
rect 752 580 818 596
rect 752 546 768 580
rect 802 546 818 580
rect 752 500 818 546
rect 752 466 768 500
rect 802 466 818 500
rect 752 424 818 466
rect 864 580 930 649
rect 864 546 880 580
rect 914 546 930 580
rect 864 499 930 546
rect 864 465 880 499
rect 914 465 930 499
rect 864 458 930 465
rect 972 580 1038 596
rect 972 546 988 580
rect 1022 546 1038 580
rect 972 500 1038 546
rect 972 466 988 500
rect 1022 466 1038 500
rect 972 424 1038 466
rect 310 420 768 424
rect 101 370 167 380
rect 310 386 315 420
rect 349 414 768 420
rect 349 390 568 414
rect 349 386 365 390
rect 310 370 365 386
rect 552 380 568 390
rect 602 390 768 414
rect 802 390 988 424
rect 1022 390 1038 424
rect 1072 580 1129 649
rect 1072 546 1078 580
rect 1112 546 1129 580
rect 1072 508 1129 546
rect 1072 474 1078 508
rect 1112 474 1129 508
rect 1072 440 1129 474
rect 1072 406 1078 440
rect 1112 406 1129 440
rect 1072 390 1129 406
rect 602 380 647 390
rect 101 336 265 370
rect 552 364 647 380
rect 231 320 344 336
rect 25 286 197 302
rect 25 252 79 286
rect 113 252 147 286
rect 181 252 197 286
rect 25 236 197 252
rect 231 286 294 320
rect 328 286 344 320
rect 231 270 344 286
rect 409 320 518 356
rect 409 286 468 320
rect 502 286 518 320
rect 409 270 518 286
rect 231 202 265 270
rect 601 236 647 364
rect 697 320 839 356
rect 697 286 721 320
rect 755 286 789 320
rect 823 286 839 320
rect 697 270 839 286
rect 889 320 1127 356
rect 889 286 964 320
rect 998 286 1127 320
rect 889 270 1127 286
rect 23 168 265 202
rect 307 210 647 236
rect 307 176 326 210
rect 360 202 647 210
rect 715 220 1129 236
rect 360 176 379 202
rect 23 153 73 168
rect 307 160 379 176
rect 715 194 903 220
rect 415 160 669 168
rect 23 119 39 153
rect 415 136 619 160
rect 23 70 73 119
rect 109 127 175 134
rect 109 93 125 127
rect 159 93 175 127
rect 109 17 175 93
rect 221 123 415 126
rect 221 89 237 123
rect 271 102 415 123
rect 449 134 619 136
rect 449 102 465 134
rect 603 126 619 134
rect 653 126 669 160
rect 603 119 669 126
rect 715 160 731 194
rect 765 186 903 194
rect 937 186 1079 220
rect 1113 186 1129 220
rect 715 119 765 160
rect 801 133 867 152
rect 271 89 465 102
rect 221 70 465 89
rect 501 66 517 100
rect 551 85 567 100
rect 801 99 817 133
rect 851 99 867 133
rect 801 85 867 99
rect 551 66 867 85
rect 901 130 939 186
rect 901 96 903 130
rect 937 96 939 130
rect 901 80 939 96
rect 973 133 1039 152
rect 973 99 989 133
rect 1023 99 1039 133
rect 501 51 867 66
rect 973 17 1039 99
rect 1079 130 1129 186
rect 1113 96 1129 130
rect 1079 80 1129 96
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand4b_2
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 762264
string GDS_START 752122
<< end >>
