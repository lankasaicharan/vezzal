magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 3 259 277 263
rect 3 49 1133 259
rect 0 0 1152 49
<< scnmos >>
rect 82 69 112 237
rect 168 69 198 237
rect 358 65 388 233
rect 458 65 488 233
rect 544 65 574 233
rect 664 65 694 233
rect 750 65 780 233
rect 844 65 874 233
rect 930 65 960 233
rect 1024 65 1054 233
<< scpmoshvt >>
rect 82 367 112 619
rect 168 367 198 619
rect 358 367 388 619
rect 458 367 488 619
rect 544 367 574 619
rect 630 367 660 619
rect 764 367 794 619
rect 866 367 896 619
rect 952 367 982 619
rect 1038 367 1068 619
<< ndiff >>
rect 29 192 82 237
rect 29 158 37 192
rect 71 158 82 192
rect 29 115 82 158
rect 29 81 37 115
rect 71 81 82 115
rect 29 69 82 81
rect 112 229 168 237
rect 112 195 123 229
rect 157 195 168 229
rect 112 153 168 195
rect 112 119 123 153
rect 157 119 168 153
rect 112 69 168 119
rect 198 225 251 237
rect 198 191 209 225
rect 243 191 251 225
rect 198 115 251 191
rect 198 81 209 115
rect 243 81 251 115
rect 198 69 251 81
rect 305 183 358 233
rect 305 149 313 183
rect 347 149 358 183
rect 305 111 358 149
rect 305 77 313 111
rect 347 77 358 111
rect 305 65 358 77
rect 388 225 458 233
rect 388 191 413 225
rect 447 191 458 225
rect 388 153 458 191
rect 388 119 413 153
rect 447 119 458 153
rect 388 65 458 119
rect 488 124 544 233
rect 488 90 499 124
rect 533 90 544 124
rect 488 65 544 90
rect 574 225 664 233
rect 574 191 619 225
rect 653 191 664 225
rect 574 153 664 191
rect 574 119 589 153
rect 623 119 664 153
rect 574 65 664 119
rect 694 192 750 233
rect 694 158 705 192
rect 739 158 750 192
rect 694 111 750 158
rect 694 77 705 111
rect 739 77 750 111
rect 694 65 750 77
rect 780 132 844 233
rect 780 98 795 132
rect 829 98 844 132
rect 780 65 844 98
rect 874 208 930 233
rect 874 174 885 208
rect 919 174 930 208
rect 874 111 930 174
rect 874 77 885 111
rect 919 77 930 111
rect 874 65 930 77
rect 960 132 1024 233
rect 960 98 975 132
rect 1009 98 1024 132
rect 960 65 1024 98
rect 1054 208 1107 233
rect 1054 174 1065 208
rect 1099 174 1107 208
rect 1054 111 1107 174
rect 1054 77 1065 111
rect 1099 77 1107 111
rect 1054 65 1107 77
<< pdiff >>
rect 29 607 82 619
rect 29 573 37 607
rect 71 573 82 607
rect 29 519 82 573
rect 29 485 37 519
rect 71 485 82 519
rect 29 434 82 485
rect 29 400 37 434
rect 71 400 82 434
rect 29 367 82 400
rect 112 599 168 619
rect 112 565 123 599
rect 157 565 168 599
rect 112 504 168 565
rect 112 470 123 504
rect 157 470 168 504
rect 112 413 168 470
rect 112 379 123 413
rect 157 379 168 413
rect 112 367 168 379
rect 198 607 358 619
rect 198 573 209 607
rect 243 573 313 607
rect 347 573 358 607
rect 198 515 358 573
rect 198 481 209 515
rect 243 481 313 515
rect 347 481 358 515
rect 198 367 358 481
rect 388 599 458 619
rect 388 565 406 599
rect 440 565 458 599
rect 388 527 458 565
rect 388 493 406 527
rect 440 493 458 527
rect 388 367 458 493
rect 488 547 544 619
rect 488 513 499 547
rect 533 513 544 547
rect 488 443 544 513
rect 488 409 499 443
rect 533 409 544 443
rect 488 367 544 409
rect 574 599 630 619
rect 574 565 585 599
rect 619 565 630 599
rect 574 527 630 565
rect 574 493 585 527
rect 619 493 630 527
rect 574 367 630 493
rect 660 607 764 619
rect 660 573 695 607
rect 729 573 764 607
rect 660 519 764 573
rect 660 485 695 519
rect 729 485 764 519
rect 660 367 764 485
rect 794 599 866 619
rect 794 565 821 599
rect 855 565 866 599
rect 794 527 866 565
rect 794 493 821 527
rect 855 493 866 527
rect 794 367 866 493
rect 896 545 952 619
rect 896 511 907 545
rect 941 511 952 545
rect 896 443 952 511
rect 896 409 907 443
rect 941 409 952 443
rect 896 367 952 409
rect 982 599 1038 619
rect 982 565 993 599
rect 1027 565 1038 599
rect 982 529 1038 565
rect 982 495 993 529
rect 1027 495 1038 529
rect 982 459 1038 495
rect 982 425 993 459
rect 1027 425 1038 459
rect 982 367 1038 425
rect 1068 607 1121 619
rect 1068 573 1079 607
rect 1113 573 1121 607
rect 1068 530 1121 573
rect 1068 496 1079 530
rect 1113 496 1121 530
rect 1068 443 1121 496
rect 1068 409 1079 443
rect 1113 409 1121 443
rect 1068 367 1121 409
<< ndiffc >>
rect 37 158 71 192
rect 37 81 71 115
rect 123 195 157 229
rect 123 119 157 153
rect 209 191 243 225
rect 209 81 243 115
rect 313 149 347 183
rect 313 77 347 111
rect 413 191 447 225
rect 413 119 447 153
rect 499 90 533 124
rect 619 191 653 225
rect 589 119 623 153
rect 705 158 739 192
rect 705 77 739 111
rect 795 98 829 132
rect 885 174 919 208
rect 885 77 919 111
rect 975 98 1009 132
rect 1065 174 1099 208
rect 1065 77 1099 111
<< pdiffc >>
rect 37 573 71 607
rect 37 485 71 519
rect 37 400 71 434
rect 123 565 157 599
rect 123 470 157 504
rect 123 379 157 413
rect 209 573 243 607
rect 313 573 347 607
rect 209 481 243 515
rect 313 481 347 515
rect 406 565 440 599
rect 406 493 440 527
rect 499 513 533 547
rect 499 409 533 443
rect 585 565 619 599
rect 585 493 619 527
rect 695 573 729 607
rect 695 485 729 519
rect 821 565 855 599
rect 821 493 855 527
rect 907 511 941 545
rect 907 409 941 443
rect 993 565 1027 599
rect 993 495 1027 529
rect 993 425 1027 459
rect 1079 573 1113 607
rect 1079 496 1113 530
rect 1079 409 1113 443
<< poly >>
rect 82 619 112 645
rect 168 619 198 645
rect 358 619 388 645
rect 458 619 488 645
rect 544 619 574 645
rect 630 619 660 645
rect 764 619 794 645
rect 866 619 896 645
rect 952 619 982 645
rect 1038 619 1068 645
rect 82 325 112 367
rect 168 325 198 367
rect 358 335 388 367
rect 21 309 198 325
rect 21 275 37 309
rect 71 275 198 309
rect 21 259 198 275
rect 270 319 404 335
rect 270 285 286 319
rect 320 285 354 319
rect 388 285 404 319
rect 270 269 404 285
rect 458 321 488 367
rect 544 321 574 367
rect 630 335 660 367
rect 764 335 794 367
rect 458 305 574 321
rect 458 271 517 305
rect 551 271 574 305
rect 82 237 112 259
rect 168 237 198 259
rect 358 233 388 269
rect 458 255 574 271
rect 616 319 694 335
rect 616 285 644 319
rect 678 285 694 319
rect 616 269 694 285
rect 736 319 802 335
rect 866 321 896 367
rect 952 321 982 367
rect 1038 321 1068 367
rect 736 285 752 319
rect 786 285 802 319
rect 736 269 802 285
rect 844 305 982 321
rect 844 271 860 305
rect 894 271 932 305
rect 966 271 982 305
rect 458 233 488 255
rect 544 233 574 255
rect 664 233 694 269
rect 750 233 780 269
rect 844 255 982 271
rect 1024 305 1131 321
rect 1024 271 1081 305
rect 1115 271 1131 305
rect 1024 255 1131 271
rect 844 233 874 255
rect 930 233 960 255
rect 1024 233 1054 255
rect 82 43 112 69
rect 168 43 198 69
rect 358 39 388 65
rect 458 39 488 65
rect 544 39 574 65
rect 664 39 694 65
rect 750 39 780 65
rect 844 39 874 65
rect 930 39 960 65
rect 1024 39 1054 65
<< polycont >>
rect 37 275 71 309
rect 286 285 320 319
rect 354 285 388 319
rect 517 271 551 305
rect 644 285 678 319
rect 752 285 786 319
rect 860 271 894 305
rect 932 271 966 305
rect 1081 271 1115 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 21 607 73 649
rect 21 573 37 607
rect 71 573 73 607
rect 21 519 73 573
rect 21 485 37 519
rect 71 485 73 519
rect 21 434 73 485
rect 21 400 37 434
rect 71 400 73 434
rect 21 384 73 400
rect 107 599 159 615
rect 107 565 123 599
rect 157 565 159 599
rect 107 504 159 565
rect 107 470 123 504
rect 157 470 159 504
rect 193 607 363 649
rect 193 573 209 607
rect 243 573 313 607
rect 347 573 363 607
rect 193 515 363 573
rect 193 481 209 515
rect 243 481 313 515
rect 347 481 363 515
rect 193 477 363 481
rect 397 599 635 615
rect 397 565 406 599
rect 440 581 585 599
rect 440 565 449 581
rect 397 527 449 565
rect 583 565 585 581
rect 619 565 635 599
rect 397 493 406 527
rect 440 493 449 527
rect 397 477 449 493
rect 483 513 499 547
rect 533 513 549 547
rect 107 443 159 470
rect 483 443 549 513
rect 583 527 635 565
rect 583 493 585 527
rect 619 493 635 527
rect 583 477 635 493
rect 679 607 745 649
rect 679 573 695 607
rect 729 573 745 607
rect 679 519 745 573
rect 679 485 695 519
rect 729 485 745 519
rect 679 477 745 485
rect 805 599 1029 615
rect 805 565 821 599
rect 855 579 993 599
rect 855 565 857 579
rect 805 527 857 565
rect 991 565 993 579
rect 1027 565 1029 599
rect 805 493 821 527
rect 855 493 857 527
rect 805 477 857 493
rect 891 511 907 545
rect 941 511 957 545
rect 891 443 957 511
rect 107 413 499 443
rect 107 379 123 413
rect 157 409 499 413
rect 533 409 907 443
rect 941 409 957 443
rect 991 529 1029 565
rect 991 495 993 529
rect 1027 495 1029 529
rect 991 459 1029 495
rect 991 425 993 459
rect 1027 425 1029 459
rect 991 409 1029 425
rect 1063 607 1129 649
rect 1063 573 1079 607
rect 1113 573 1129 607
rect 1063 530 1129 573
rect 1063 496 1079 530
rect 1113 496 1129 530
rect 1063 443 1129 496
rect 1063 409 1079 443
rect 1113 409 1129 443
rect 157 379 267 409
rect 107 369 267 379
rect 107 363 236 369
rect 18 309 71 350
rect 18 275 37 309
rect 18 242 71 275
rect 107 229 173 363
rect 301 341 694 375
rect 301 335 463 341
rect 270 319 463 335
rect 270 285 286 319
rect 320 285 354 319
rect 388 285 463 319
rect 628 319 694 341
rect 497 305 567 307
rect 497 271 517 305
rect 551 271 567 305
rect 21 192 73 208
rect 21 158 37 192
rect 71 158 73 192
rect 21 115 73 158
rect 107 195 123 229
rect 157 195 173 229
rect 107 153 173 195
rect 107 119 123 153
rect 157 119 173 153
rect 209 225 463 251
rect 497 242 567 271
rect 628 285 644 319
rect 678 285 694 319
rect 628 269 694 285
rect 736 339 1134 375
rect 736 319 803 339
rect 736 285 752 319
rect 786 285 803 319
rect 1069 305 1134 339
rect 736 269 803 285
rect 844 271 860 305
rect 894 271 932 305
rect 966 271 1035 305
rect 844 242 1035 271
rect 1069 271 1081 305
rect 1115 271 1134 305
rect 1069 242 1134 271
rect 243 217 413 225
rect 243 191 247 217
rect 21 81 37 115
rect 71 85 73 115
rect 209 115 247 191
rect 397 191 413 217
rect 447 208 463 225
rect 601 225 669 229
rect 601 208 619 225
rect 447 191 619 208
rect 653 191 669 225
rect 71 81 209 85
rect 243 81 247 115
rect 21 51 247 81
rect 297 149 313 183
rect 347 149 363 183
rect 297 111 363 149
rect 397 174 669 191
rect 397 153 463 174
rect 397 119 413 153
rect 447 119 463 153
rect 573 153 669 174
rect 497 124 539 140
rect 297 77 313 111
rect 347 85 363 111
rect 497 90 499 124
rect 533 90 539 124
rect 573 119 589 153
rect 623 119 669 153
rect 703 192 885 208
rect 703 158 705 192
rect 739 174 885 192
rect 919 174 1065 208
rect 1099 174 1115 208
rect 739 158 743 174
rect 497 85 539 90
rect 703 111 743 158
rect 703 85 705 111
rect 347 77 705 85
rect 739 77 743 111
rect 297 51 743 77
rect 779 132 845 140
rect 779 98 795 132
rect 829 98 845 132
rect 779 17 845 98
rect 879 111 925 174
rect 879 77 885 111
rect 919 77 925 111
rect 879 61 925 77
rect 959 132 1025 140
rect 959 98 975 132
rect 1009 98 1025 132
rect 959 17 1025 98
rect 1059 111 1115 174
rect 1059 77 1065 111
rect 1099 77 1115 111
rect 1059 61 1115 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221ai_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5825700
string GDS_START 5814850
<< end >>
