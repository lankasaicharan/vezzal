magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
rect 275 329 443 331
<< pwell >>
rect 900 235 1533 241
rect 350 180 1533 235
rect 51 49 1533 180
rect 0 0 1536 49
<< scnmos >>
rect 134 70 164 154
rect 220 70 250 154
rect 429 125 459 209
rect 537 125 567 209
rect 609 125 639 209
rect 695 125 725 209
rect 789 125 819 209
rect 979 47 1009 215
rect 1051 47 1081 215
rect 1166 47 1196 215
rect 1252 47 1282 215
rect 1338 47 1368 215
rect 1424 47 1454 215
<< scpmoshvt >>
rect 80 468 110 596
rect 220 468 250 596
rect 429 447 459 575
rect 537 447 567 575
rect 609 447 639 575
rect 718 447 748 531
rect 790 447 820 531
rect 979 367 1009 619
rect 1065 367 1095 619
rect 1164 367 1194 619
rect 1252 367 1282 619
rect 1338 367 1368 619
rect 1424 367 1454 619
<< ndiff >>
rect 77 116 134 154
rect 77 82 85 116
rect 119 82 134 116
rect 77 70 134 82
rect 164 116 220 154
rect 164 82 175 116
rect 209 82 220 116
rect 164 70 220 82
rect 250 116 303 154
rect 250 82 261 116
rect 295 82 303 116
rect 250 70 303 82
rect 376 197 429 209
rect 376 163 384 197
rect 418 163 429 197
rect 376 125 429 163
rect 459 171 537 209
rect 459 137 474 171
rect 508 137 537 171
rect 459 125 537 137
rect 567 125 609 209
rect 639 173 695 209
rect 639 139 650 173
rect 684 139 695 173
rect 639 125 695 139
rect 725 125 789 209
rect 819 175 872 209
rect 819 141 830 175
rect 864 141 872 175
rect 819 125 872 141
rect 926 171 979 215
rect 926 137 934 171
rect 968 137 979 171
rect 926 101 979 137
rect 926 67 934 101
rect 968 67 979 101
rect 926 47 979 67
rect 1009 47 1051 215
rect 1081 133 1166 215
rect 1081 99 1105 133
rect 1139 99 1166 133
rect 1081 47 1166 99
rect 1196 203 1252 215
rect 1196 169 1207 203
rect 1241 169 1252 203
rect 1196 101 1252 169
rect 1196 67 1207 101
rect 1241 67 1252 101
rect 1196 47 1252 67
rect 1282 183 1338 215
rect 1282 149 1293 183
rect 1327 149 1338 183
rect 1282 93 1338 149
rect 1282 59 1293 93
rect 1327 59 1338 93
rect 1282 47 1338 59
rect 1368 203 1424 215
rect 1368 169 1379 203
rect 1413 169 1424 203
rect 1368 101 1424 169
rect 1368 67 1379 101
rect 1413 67 1424 101
rect 1368 47 1424 67
rect 1454 183 1507 215
rect 1454 149 1465 183
rect 1499 149 1507 183
rect 1454 93 1507 149
rect 1454 59 1465 93
rect 1499 59 1507 93
rect 1454 47 1507 59
<< pdiff >>
rect 27 584 80 596
rect 27 550 35 584
rect 69 550 80 584
rect 27 514 80 550
rect 27 480 35 514
rect 69 480 80 514
rect 27 468 80 480
rect 110 584 220 596
rect 110 550 121 584
rect 155 550 220 584
rect 110 468 220 550
rect 250 514 303 596
rect 250 480 261 514
rect 295 480 303 514
rect 250 468 303 480
rect 357 447 429 575
rect 459 563 537 575
rect 459 529 481 563
rect 515 529 537 563
rect 459 447 537 529
rect 567 447 609 575
rect 639 561 696 575
rect 639 527 654 561
rect 688 531 696 561
rect 926 570 979 619
rect 926 536 934 570
rect 968 536 979 570
rect 926 531 979 536
rect 688 527 718 531
rect 639 493 718 527
rect 639 459 663 493
rect 697 459 718 493
rect 639 447 718 459
rect 748 447 790 531
rect 820 447 979 531
rect 357 411 407 447
rect 357 377 365 411
rect 399 377 407 411
rect 357 365 407 377
rect 926 367 979 447
rect 1009 599 1065 619
rect 1009 565 1020 599
rect 1054 565 1065 599
rect 1009 510 1065 565
rect 1009 476 1020 510
rect 1054 476 1065 510
rect 1009 367 1065 476
rect 1095 570 1164 619
rect 1095 536 1112 570
rect 1146 536 1164 570
rect 1095 367 1164 536
rect 1194 599 1252 619
rect 1194 565 1207 599
rect 1241 565 1252 599
rect 1194 506 1252 565
rect 1194 472 1207 506
rect 1241 472 1252 506
rect 1194 413 1252 472
rect 1194 379 1207 413
rect 1241 379 1252 413
rect 1194 367 1252 379
rect 1282 607 1338 619
rect 1282 573 1293 607
rect 1327 573 1338 607
rect 1282 533 1338 573
rect 1282 499 1293 533
rect 1327 499 1338 533
rect 1282 455 1338 499
rect 1282 421 1293 455
rect 1327 421 1338 455
rect 1282 367 1338 421
rect 1368 599 1424 619
rect 1368 565 1379 599
rect 1413 565 1424 599
rect 1368 506 1424 565
rect 1368 472 1379 506
rect 1413 472 1424 506
rect 1368 413 1424 472
rect 1368 379 1379 413
rect 1413 379 1424 413
rect 1368 367 1424 379
rect 1454 607 1507 619
rect 1454 573 1465 607
rect 1499 573 1507 607
rect 1454 533 1507 573
rect 1454 499 1465 533
rect 1499 499 1507 533
rect 1454 455 1507 499
rect 1454 421 1465 455
rect 1499 421 1507 455
rect 1454 367 1507 421
<< ndiffc >>
rect 85 82 119 116
rect 175 82 209 116
rect 261 82 295 116
rect 384 163 418 197
rect 474 137 508 171
rect 650 139 684 173
rect 830 141 864 175
rect 934 137 968 171
rect 934 67 968 101
rect 1105 99 1139 133
rect 1207 169 1241 203
rect 1207 67 1241 101
rect 1293 149 1327 183
rect 1293 59 1327 93
rect 1379 169 1413 203
rect 1379 67 1413 101
rect 1465 149 1499 183
rect 1465 59 1499 93
<< pdiffc >>
rect 35 550 69 584
rect 35 480 69 514
rect 121 550 155 584
rect 261 480 295 514
rect 481 529 515 563
rect 654 527 688 561
rect 934 536 968 570
rect 663 459 697 493
rect 365 377 399 411
rect 1020 565 1054 599
rect 1020 476 1054 510
rect 1112 536 1146 570
rect 1207 565 1241 599
rect 1207 472 1241 506
rect 1207 379 1241 413
rect 1293 573 1327 607
rect 1293 499 1327 533
rect 1293 421 1327 455
rect 1379 565 1413 599
rect 1379 472 1413 506
rect 1379 379 1413 413
rect 1465 573 1499 607
rect 1465 499 1499 533
rect 1465 421 1499 455
<< poly >>
rect 80 596 110 622
rect 220 596 250 622
rect 979 619 1009 645
rect 1065 619 1095 645
rect 1164 619 1194 645
rect 1252 619 1282 645
rect 1338 619 1368 645
rect 1424 619 1454 645
rect 429 575 459 601
rect 537 575 567 601
rect 609 575 639 601
rect 80 310 110 468
rect 220 436 250 468
rect 158 420 250 436
rect 158 386 174 420
rect 208 386 250 420
rect 158 370 250 386
rect 80 294 164 310
rect 80 260 114 294
rect 148 260 164 294
rect 80 226 164 260
rect 80 192 114 226
rect 148 192 164 226
rect 80 176 164 192
rect 134 154 164 176
rect 220 154 250 370
rect 718 531 748 557
rect 790 531 820 557
rect 429 331 459 447
rect 537 415 567 447
rect 318 315 459 331
rect 318 281 334 315
rect 368 281 459 315
rect 501 399 567 415
rect 501 365 517 399
rect 551 365 567 399
rect 501 331 567 365
rect 609 415 639 447
rect 609 399 675 415
rect 609 365 625 399
rect 659 365 675 399
rect 609 349 675 365
rect 718 337 748 447
rect 501 297 517 331
rect 551 297 567 331
rect 717 307 748 337
rect 790 415 820 447
rect 790 399 856 415
rect 790 365 806 399
rect 840 365 856 399
rect 790 331 856 365
rect 501 281 567 297
rect 318 265 459 281
rect 134 44 164 70
rect 220 44 250 70
rect 318 51 348 265
rect 429 209 459 265
rect 537 209 567 281
rect 609 277 747 307
rect 790 297 806 331
rect 840 297 856 331
rect 979 303 1009 367
rect 1065 308 1095 367
rect 1164 335 1194 367
rect 1252 335 1282 367
rect 1338 335 1368 367
rect 1424 335 1454 367
rect 1164 319 1454 335
rect 790 281 856 297
rect 905 287 1009 303
rect 609 209 639 277
rect 790 265 825 281
rect 789 235 825 265
rect 905 253 921 287
rect 955 253 1009 287
rect 905 237 1009 253
rect 695 209 725 235
rect 789 209 819 235
rect 979 215 1009 237
rect 1051 292 1117 308
rect 1051 258 1067 292
rect 1101 258 1117 292
rect 1164 285 1181 319
rect 1215 285 1249 319
rect 1283 285 1317 319
rect 1351 285 1385 319
rect 1419 285 1454 319
rect 1164 269 1454 285
rect 1051 242 1117 258
rect 1051 215 1081 242
rect 1166 215 1196 269
rect 1252 215 1282 269
rect 1338 215 1368 269
rect 1424 215 1454 269
rect 429 99 459 125
rect 537 99 567 125
rect 609 51 639 125
rect 695 103 725 125
rect 318 21 639 51
rect 681 87 747 103
rect 789 99 819 125
rect 681 53 697 87
rect 731 53 747 87
rect 681 37 747 53
rect 979 21 1009 47
rect 1051 21 1081 47
rect 1166 21 1196 47
rect 1252 21 1282 47
rect 1338 21 1368 47
rect 1424 21 1454 47
<< polycont >>
rect 174 386 208 420
rect 114 260 148 294
rect 114 192 148 226
rect 334 281 368 315
rect 517 365 551 399
rect 625 365 659 399
rect 517 297 551 331
rect 806 365 840 399
rect 806 297 840 331
rect 921 253 955 287
rect 1067 258 1101 292
rect 1181 285 1215 319
rect 1249 285 1283 319
rect 1317 285 1351 319
rect 1385 285 1419 319
rect 697 53 731 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 19 584 73 600
rect 19 550 35 584
rect 69 550 73 584
rect 19 514 73 550
rect 107 584 157 649
rect 107 550 121 584
rect 155 550 157 584
rect 107 532 157 550
rect 191 566 402 600
rect 19 480 35 514
rect 69 498 73 514
rect 191 498 225 566
rect 69 480 225 498
rect 19 464 225 480
rect 259 514 301 532
rect 259 480 261 514
rect 295 480 301 514
rect 19 134 73 464
rect 127 420 225 430
rect 127 386 174 420
rect 208 386 225 420
rect 127 384 225 386
rect 107 294 203 350
rect 107 260 114 294
rect 148 260 203 294
rect 107 226 203 260
rect 107 192 114 226
rect 148 192 203 226
rect 107 168 203 192
rect 259 331 301 480
rect 335 489 402 566
rect 465 563 531 649
rect 465 529 481 563
rect 515 529 531 563
rect 465 523 531 529
rect 638 561 745 577
rect 638 527 654 561
rect 688 527 745 561
rect 918 570 984 649
rect 918 536 934 570
rect 968 536 984 570
rect 918 528 984 536
rect 1018 599 1062 615
rect 1018 565 1020 599
rect 1054 565 1062 599
rect 638 493 745 527
rect 1018 510 1062 565
rect 1096 570 1162 649
rect 1096 536 1112 570
rect 1146 536 1162 570
rect 1096 528 1162 536
rect 1205 599 1243 615
rect 1205 565 1207 599
rect 1241 565 1243 599
rect 1018 494 1020 510
rect 335 455 567 489
rect 349 411 454 421
rect 349 377 365 411
rect 399 377 454 411
rect 349 365 454 377
rect 259 315 384 331
rect 259 281 334 315
rect 368 281 384 315
rect 259 279 384 281
rect 19 116 125 134
rect 19 82 85 116
rect 119 82 125 116
rect 19 66 125 82
rect 159 116 225 134
rect 159 82 175 116
rect 209 82 225 116
rect 159 17 225 82
rect 259 116 299 279
rect 420 245 454 365
rect 501 399 567 455
rect 638 459 663 493
rect 697 459 745 493
rect 638 449 745 459
rect 501 365 517 399
rect 551 365 567 399
rect 501 331 567 365
rect 501 297 517 331
rect 551 297 567 331
rect 501 281 567 297
rect 609 399 675 415
rect 609 365 625 399
rect 659 365 675 399
rect 609 245 675 365
rect 380 211 675 245
rect 709 247 745 449
rect 790 476 1020 494
rect 1054 494 1062 510
rect 1205 506 1243 565
rect 1054 476 1171 494
rect 790 460 1171 476
rect 790 399 856 460
rect 790 365 806 399
rect 840 365 856 399
rect 790 331 856 365
rect 790 297 806 331
rect 840 297 856 331
rect 790 281 856 297
rect 905 287 955 303
rect 905 253 921 287
rect 905 247 955 253
rect 709 213 955 247
rect 989 292 1103 426
rect 989 258 1067 292
rect 1101 258 1103 292
rect 989 242 1103 258
rect 1137 319 1171 460
rect 1205 472 1207 506
rect 1241 472 1243 506
rect 1205 413 1243 472
rect 1277 607 1343 649
rect 1277 573 1293 607
rect 1327 573 1343 607
rect 1277 533 1343 573
rect 1277 499 1293 533
rect 1327 499 1343 533
rect 1277 455 1343 499
rect 1277 421 1293 455
rect 1327 421 1343 455
rect 1377 599 1415 615
rect 1377 565 1379 599
rect 1413 565 1415 599
rect 1377 506 1415 565
rect 1377 472 1379 506
rect 1413 472 1415 506
rect 1205 379 1207 413
rect 1241 387 1243 413
rect 1377 413 1415 472
rect 1449 607 1515 649
rect 1449 573 1465 607
rect 1499 573 1515 607
rect 1449 533 1515 573
rect 1449 499 1465 533
rect 1499 499 1515 533
rect 1449 455 1515 499
rect 1449 421 1465 455
rect 1499 421 1515 455
rect 1377 387 1379 413
rect 1241 379 1379 387
rect 1413 387 1415 413
rect 1413 379 1519 387
rect 1205 353 1519 379
rect 1137 285 1181 319
rect 1215 285 1249 319
rect 1283 285 1317 319
rect 1351 285 1385 319
rect 1419 285 1435 319
rect 380 197 422 211
rect 380 163 384 197
rect 418 163 422 197
rect 380 147 422 163
rect 458 171 524 175
rect 259 82 261 116
rect 295 82 299 116
rect 259 66 299 82
rect 458 137 474 171
rect 508 137 524 171
rect 458 17 524 137
rect 564 99 598 211
rect 709 177 745 213
rect 1137 208 1171 285
rect 1469 251 1519 353
rect 989 179 1171 208
rect 634 173 745 177
rect 634 139 650 173
rect 684 139 745 173
rect 634 133 745 139
rect 814 175 880 179
rect 814 141 830 175
rect 864 141 880 175
rect 564 87 747 99
rect 564 53 697 87
rect 731 53 747 87
rect 564 51 747 53
rect 814 17 880 141
rect 918 174 1171 179
rect 1205 217 1519 251
rect 1205 203 1243 217
rect 918 171 1023 174
rect 918 137 934 171
rect 968 145 1023 171
rect 1205 169 1207 203
rect 1241 169 1243 203
rect 1377 203 1415 217
rect 968 137 984 145
rect 918 101 984 137
rect 918 67 934 101
rect 968 67 984 101
rect 918 51 984 67
rect 1089 133 1155 140
rect 1089 99 1105 133
rect 1139 99 1155 133
rect 1205 117 1243 169
rect 1089 17 1155 99
rect 1191 101 1243 117
rect 1191 67 1207 101
rect 1241 67 1243 101
rect 1191 51 1243 67
rect 1277 149 1293 183
rect 1327 149 1343 183
rect 1277 93 1343 149
rect 1277 59 1293 93
rect 1327 59 1343 93
rect 1277 17 1343 59
rect 1377 169 1379 203
rect 1413 169 1415 203
rect 1377 101 1415 169
rect 1377 67 1379 101
rect 1413 67 1415 101
rect 1377 51 1415 67
rect 1449 149 1465 183
rect 1499 149 1515 183
rect 1449 93 1515 149
rect 1449 59 1465 93
rect 1499 59 1515 93
rect 1449 17 1515 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrtn_4
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2690072
string GDS_START 2678132
<< end >>
