magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 332 2054 704
rect 709 317 961 332
<< pwell >>
rect 1 273 652 279
rect 1 248 1162 273
rect 1 49 1999 248
rect 0 0 2016 49
<< scpmos >>
rect 81 392 117 592
rect 171 392 207 592
rect 261 392 297 592
rect 351 392 387 592
rect 555 379 591 547
rect 645 379 681 547
rect 735 379 771 547
rect 856 410 892 578
rect 946 410 982 578
rect 1051 368 1087 536
rect 1183 368 1219 592
rect 1305 368 1341 592
rect 1395 368 1431 592
rect 1485 368 1521 592
rect 1575 368 1611 592
rect 1665 368 1701 592
rect 1755 368 1791 592
rect 1897 368 1933 592
<< nmoslvt >>
rect 84 125 114 253
rect 171 125 201 253
rect 257 125 287 253
rect 343 125 373 253
rect 435 125 465 253
rect 529 125 559 253
rect 765 119 795 247
rect 851 119 881 247
rect 951 119 981 247
rect 1051 119 1081 247
rect 1245 74 1275 222
rect 1331 74 1361 222
rect 1417 74 1447 222
rect 1503 74 1533 222
rect 1589 74 1619 222
rect 1675 74 1705 222
rect 1775 74 1805 222
rect 1886 74 1916 222
<< ndiff >>
rect 27 241 84 253
rect 27 207 39 241
rect 73 207 84 241
rect 27 171 84 207
rect 27 137 39 171
rect 73 137 84 171
rect 27 125 84 137
rect 114 172 171 253
rect 114 138 125 172
rect 159 138 171 172
rect 114 125 171 138
rect 201 241 257 253
rect 201 207 212 241
rect 246 207 257 241
rect 201 171 257 207
rect 201 137 212 171
rect 246 137 257 171
rect 201 125 257 137
rect 287 172 343 253
rect 287 138 298 172
rect 332 138 343 172
rect 287 125 343 138
rect 373 241 435 253
rect 373 207 384 241
rect 418 207 435 241
rect 373 171 435 207
rect 373 137 384 171
rect 418 137 435 171
rect 373 125 435 137
rect 465 241 529 253
rect 465 207 484 241
rect 518 207 529 241
rect 465 171 529 207
rect 465 137 484 171
rect 518 137 529 171
rect 465 125 529 137
rect 559 239 626 253
rect 559 205 584 239
rect 618 205 626 239
rect 559 171 626 205
rect 559 137 584 171
rect 618 137 626 171
rect 559 125 626 137
rect 707 231 765 247
rect 707 197 720 231
rect 754 197 765 231
rect 707 163 765 197
rect 707 129 720 163
rect 754 129 765 163
rect 707 119 765 129
rect 795 235 851 247
rect 795 201 806 235
rect 840 201 851 235
rect 795 165 851 201
rect 795 131 806 165
rect 840 131 851 165
rect 795 119 851 131
rect 881 235 951 247
rect 881 201 906 235
rect 940 201 951 235
rect 881 165 951 201
rect 881 131 906 165
rect 940 131 951 165
rect 881 119 951 131
rect 981 235 1051 247
rect 981 201 1006 235
rect 1040 201 1051 235
rect 981 165 1051 201
rect 981 131 1006 165
rect 1040 131 1051 165
rect 981 119 1051 131
rect 1081 235 1136 247
rect 1081 201 1092 235
rect 1126 201 1136 235
rect 1081 165 1136 201
rect 1081 131 1092 165
rect 1126 131 1136 165
rect 1081 119 1136 131
rect 1190 210 1245 222
rect 1190 176 1200 210
rect 1234 176 1245 210
rect 1190 120 1245 176
rect 1190 86 1200 120
rect 1234 86 1245 120
rect 1190 74 1245 86
rect 1275 210 1331 222
rect 1275 176 1286 210
rect 1320 176 1331 210
rect 1275 120 1331 176
rect 1275 86 1286 120
rect 1320 86 1331 120
rect 1275 74 1331 86
rect 1361 123 1417 222
rect 1361 89 1372 123
rect 1406 89 1417 123
rect 1361 74 1417 89
rect 1447 210 1503 222
rect 1447 176 1458 210
rect 1492 176 1503 210
rect 1447 74 1503 176
rect 1533 123 1589 222
rect 1533 89 1544 123
rect 1578 89 1589 123
rect 1533 74 1589 89
rect 1619 210 1675 222
rect 1619 176 1630 210
rect 1664 176 1675 210
rect 1619 120 1675 176
rect 1619 86 1630 120
rect 1664 86 1675 120
rect 1619 74 1675 86
rect 1705 133 1775 222
rect 1705 99 1730 133
rect 1764 99 1775 133
rect 1705 74 1775 99
rect 1805 210 1886 222
rect 1805 176 1830 210
rect 1864 176 1886 210
rect 1805 120 1886 176
rect 1805 86 1830 120
rect 1864 86 1886 120
rect 1805 74 1886 86
rect 1916 146 1973 222
rect 1916 112 1927 146
rect 1961 112 1973 146
rect 1916 74 1973 112
<< pdiff >>
rect 27 577 81 592
rect 27 543 37 577
rect 71 543 81 577
rect 27 509 81 543
rect 27 475 37 509
rect 71 475 81 509
rect 27 441 81 475
rect 27 407 37 441
rect 71 407 81 441
rect 27 392 81 407
rect 117 577 171 592
rect 117 543 127 577
rect 161 543 171 577
rect 117 509 171 543
rect 117 475 127 509
rect 161 475 171 509
rect 117 392 171 475
rect 207 580 261 592
rect 207 546 217 580
rect 251 546 261 580
rect 207 510 261 546
rect 207 476 217 510
rect 251 476 261 510
rect 207 441 261 476
rect 207 407 217 441
rect 251 407 261 441
rect 207 392 261 407
rect 297 531 351 592
rect 297 497 307 531
rect 341 497 351 531
rect 297 441 351 497
rect 297 407 307 441
rect 341 407 351 441
rect 297 392 351 407
rect 387 580 441 592
rect 387 546 397 580
rect 431 546 441 580
rect 387 493 441 546
rect 387 459 397 493
rect 431 459 441 493
rect 387 392 441 459
rect 806 547 856 578
rect 501 531 555 547
rect 501 497 511 531
rect 545 497 555 531
rect 501 379 555 497
rect 591 431 645 547
rect 591 397 601 431
rect 635 397 645 431
rect 591 379 645 397
rect 681 535 735 547
rect 681 501 691 535
rect 725 501 735 535
rect 681 379 735 501
rect 771 410 856 547
rect 892 566 946 578
rect 892 532 902 566
rect 936 532 946 566
rect 892 410 946 532
rect 982 536 1032 578
rect 1102 566 1183 592
rect 1102 536 1126 566
rect 982 414 1051 536
rect 982 410 1007 414
rect 771 399 841 410
rect 771 379 796 399
rect 786 365 796 379
rect 830 365 841 399
rect 786 353 841 365
rect 997 380 1007 410
rect 1041 380 1051 414
rect 997 368 1051 380
rect 1087 532 1126 536
rect 1160 532 1183 566
rect 1087 368 1183 532
rect 1219 414 1305 592
rect 1219 380 1260 414
rect 1294 380 1305 414
rect 1219 368 1305 380
rect 1341 573 1395 592
rect 1341 539 1351 573
rect 1385 539 1395 573
rect 1341 368 1395 539
rect 1431 414 1485 592
rect 1431 380 1441 414
rect 1475 380 1485 414
rect 1431 368 1485 380
rect 1521 573 1575 592
rect 1521 539 1531 573
rect 1565 539 1575 573
rect 1521 368 1575 539
rect 1611 580 1665 592
rect 1611 546 1621 580
rect 1655 546 1665 580
rect 1611 503 1665 546
rect 1611 469 1621 503
rect 1655 469 1665 503
rect 1611 414 1665 469
rect 1611 380 1621 414
rect 1655 380 1665 414
rect 1611 368 1665 380
rect 1701 584 1755 592
rect 1701 550 1711 584
rect 1745 550 1755 584
rect 1701 498 1755 550
rect 1701 464 1711 498
rect 1745 464 1755 498
rect 1701 368 1755 464
rect 1791 580 1897 592
rect 1791 546 1831 580
rect 1865 546 1897 580
rect 1791 503 1897 546
rect 1791 469 1831 503
rect 1865 469 1897 503
rect 1791 414 1897 469
rect 1791 380 1831 414
rect 1865 380 1897 414
rect 1791 368 1897 380
rect 1933 580 1989 592
rect 1933 546 1943 580
rect 1977 546 1989 580
rect 1933 500 1989 546
rect 1933 466 1943 500
rect 1977 466 1989 500
rect 1933 368 1989 466
<< ndiffc >>
rect 39 207 73 241
rect 39 137 73 171
rect 125 138 159 172
rect 212 207 246 241
rect 212 137 246 171
rect 298 138 332 172
rect 384 207 418 241
rect 384 137 418 171
rect 484 207 518 241
rect 484 137 518 171
rect 584 205 618 239
rect 584 137 618 171
rect 720 197 754 231
rect 720 129 754 163
rect 806 201 840 235
rect 806 131 840 165
rect 906 201 940 235
rect 906 131 940 165
rect 1006 201 1040 235
rect 1006 131 1040 165
rect 1092 201 1126 235
rect 1092 131 1126 165
rect 1200 176 1234 210
rect 1200 86 1234 120
rect 1286 176 1320 210
rect 1286 86 1320 120
rect 1372 89 1406 123
rect 1458 176 1492 210
rect 1544 89 1578 123
rect 1630 176 1664 210
rect 1630 86 1664 120
rect 1730 99 1764 133
rect 1830 176 1864 210
rect 1830 86 1864 120
rect 1927 112 1961 146
<< pdiffc >>
rect 37 543 71 577
rect 37 475 71 509
rect 37 407 71 441
rect 127 543 161 577
rect 127 475 161 509
rect 217 546 251 580
rect 217 476 251 510
rect 217 407 251 441
rect 307 497 341 531
rect 307 407 341 441
rect 397 546 431 580
rect 397 459 431 493
rect 511 497 545 531
rect 601 397 635 431
rect 691 501 725 535
rect 902 532 936 566
rect 796 365 830 399
rect 1007 380 1041 414
rect 1126 532 1160 566
rect 1260 380 1294 414
rect 1351 539 1385 573
rect 1441 380 1475 414
rect 1531 539 1565 573
rect 1621 546 1655 580
rect 1621 469 1655 503
rect 1621 380 1655 414
rect 1711 550 1745 584
rect 1711 464 1745 498
rect 1831 546 1865 580
rect 1831 469 1865 503
rect 1831 380 1865 414
rect 1943 546 1977 580
rect 1943 466 1977 500
<< poly >>
rect 81 592 117 618
rect 171 592 207 618
rect 261 592 297 618
rect 351 592 387 618
rect 456 615 892 645
rect 81 357 117 392
rect 171 357 207 392
rect 261 376 297 392
rect 351 376 387 392
rect 456 376 486 615
rect 555 547 591 573
rect 645 547 681 573
rect 735 547 771 615
rect 856 578 892 615
rect 946 578 982 604
rect 1183 592 1219 618
rect 1305 592 1341 618
rect 1395 592 1431 618
rect 1485 592 1521 618
rect 1575 592 1611 618
rect 1665 592 1701 618
rect 1755 592 1791 618
rect 1897 592 1933 618
rect 1051 536 1087 562
rect 81 341 201 357
rect 81 307 128 341
rect 162 307 201 341
rect 261 346 486 376
rect 555 347 591 379
rect 645 347 681 379
rect 261 341 387 346
rect 261 321 329 341
rect 81 291 201 307
rect 84 253 114 291
rect 171 253 201 291
rect 257 307 329 321
rect 363 307 387 341
rect 257 291 387 307
rect 555 331 681 347
rect 555 298 631 331
rect 435 297 631 298
rect 665 297 681 331
rect 735 336 771 379
rect 856 384 892 410
rect 735 306 881 336
rect 257 253 287 291
rect 343 253 373 291
rect 435 268 681 297
rect 435 253 465 268
rect 529 253 559 268
rect 765 247 795 306
rect 851 247 881 306
rect 946 326 982 410
rect 1051 326 1087 368
rect 946 292 1087 326
rect 1183 330 1219 368
rect 1305 330 1341 368
rect 1395 330 1431 368
rect 1485 330 1521 368
rect 1183 314 1521 330
rect 1183 300 1205 314
rect 951 262 1081 292
rect 1189 280 1205 300
rect 1239 280 1273 314
rect 1307 280 1341 314
rect 1375 294 1521 314
rect 1575 330 1611 368
rect 1665 330 1701 368
rect 1755 330 1791 368
rect 1897 330 1933 368
rect 1575 314 1945 330
rect 1375 280 1533 294
rect 1189 264 1533 280
rect 1575 280 1591 314
rect 1625 280 1664 314
rect 1698 280 1743 314
rect 1777 280 1822 314
rect 1856 280 1895 314
rect 1929 280 1945 314
rect 1575 264 1945 280
rect 951 247 981 262
rect 1051 247 1081 262
rect 84 99 114 125
rect 171 51 201 125
rect 257 99 287 125
rect 343 99 373 125
rect 435 99 465 125
rect 529 99 559 125
rect 1245 222 1275 264
rect 1331 222 1361 264
rect 1417 222 1447 264
rect 1503 222 1533 264
rect 1589 222 1619 264
rect 1675 222 1705 264
rect 1775 222 1805 264
rect 1886 222 1916 264
rect 765 93 795 119
rect 851 93 881 119
rect 951 51 981 119
rect 1051 93 1081 119
rect 171 21 981 51
rect 1245 48 1275 74
rect 1331 48 1361 74
rect 1417 48 1447 74
rect 1503 48 1533 74
rect 1589 48 1619 74
rect 1675 48 1705 74
rect 1775 48 1805 74
rect 1886 48 1916 74
<< polycont >>
rect 128 307 162 341
rect 329 307 363 341
rect 631 297 665 331
rect 1205 280 1239 314
rect 1273 280 1307 314
rect 1341 280 1375 314
rect 1591 280 1625 314
rect 1664 280 1698 314
rect 1743 280 1777 314
rect 1822 280 1856 314
rect 1895 280 1929 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 21 577 77 593
rect 21 543 37 577
rect 71 543 77 577
rect 21 509 77 543
rect 21 475 37 509
rect 71 475 77 509
rect 21 441 77 475
rect 111 577 161 649
rect 111 543 127 577
rect 111 509 161 543
rect 111 475 127 509
rect 111 459 161 475
rect 201 581 447 615
rect 201 580 251 581
rect 201 546 217 580
rect 381 580 447 581
rect 201 510 251 546
rect 201 476 217 510
rect 21 407 37 441
rect 71 425 77 441
rect 201 441 251 476
rect 201 425 217 441
rect 71 407 217 425
rect 21 391 251 407
rect 291 531 347 547
rect 291 497 307 531
rect 341 497 347 531
rect 291 441 347 497
rect 381 546 397 580
rect 431 546 447 580
rect 381 493 447 546
rect 381 459 397 493
rect 431 459 447 493
rect 495 531 561 649
rect 495 497 511 531
rect 545 497 561 531
rect 675 535 741 649
rect 675 501 691 535
rect 725 501 741 535
rect 886 566 952 649
rect 886 532 902 566
rect 936 532 952 566
rect 1098 566 1189 649
rect 1098 532 1126 566
rect 1160 532 1189 566
rect 1335 573 1401 649
rect 1335 539 1351 573
rect 1385 539 1401 573
rect 1335 532 1401 539
rect 1515 573 1581 649
rect 1515 539 1531 573
rect 1565 539 1581 573
rect 1515 532 1581 539
rect 1615 580 1661 596
rect 1615 546 1621 580
rect 1655 546 1661 580
rect 1615 503 1661 546
rect 495 481 561 497
rect 780 467 1579 498
rect 617 464 1579 467
rect 617 447 814 464
rect 291 407 307 441
rect 341 425 347 441
rect 585 433 814 447
rect 585 431 651 433
rect 585 425 601 431
rect 341 407 601 425
rect 291 397 601 407
rect 635 397 651 431
rect 991 414 1210 430
rect 991 399 1007 414
rect 291 391 651 397
rect 500 381 651 391
rect 25 341 263 357
rect 25 307 128 341
rect 162 307 263 341
rect 25 291 263 307
rect 313 341 455 357
rect 313 307 329 341
rect 363 307 455 341
rect 313 291 455 307
rect 500 257 534 381
rect 780 365 796 399
rect 830 380 1007 399
rect 1041 380 1210 414
rect 830 365 1210 380
rect 780 364 1210 365
rect 1244 414 1511 430
rect 1244 380 1260 414
rect 1294 380 1441 414
rect 1475 380 1511 414
rect 1244 364 1511 380
rect 780 349 846 364
rect 780 347 814 349
rect 615 331 814 347
rect 615 297 631 331
rect 665 315 814 331
rect 1176 330 1210 364
rect 665 297 856 315
rect 615 281 856 297
rect 23 241 434 257
rect 23 207 39 241
rect 73 223 212 241
rect 23 171 73 207
rect 196 207 212 223
rect 246 223 384 241
rect 23 137 39 171
rect 23 121 73 137
rect 109 172 159 189
rect 109 138 125 172
rect 109 17 159 138
rect 196 171 246 207
rect 368 207 384 223
rect 418 207 434 241
rect 196 137 212 171
rect 196 121 246 137
rect 282 172 332 189
rect 282 138 298 172
rect 282 17 332 138
rect 368 171 434 207
rect 368 137 384 171
rect 418 137 434 171
rect 368 87 434 137
rect 468 241 534 257
rect 468 207 484 241
rect 518 207 534 241
rect 468 171 534 207
rect 468 137 484 171
rect 518 137 534 171
rect 468 121 534 137
rect 568 239 634 247
rect 568 205 584 239
rect 618 205 634 239
rect 568 171 634 205
rect 568 137 584 171
rect 618 137 634 171
rect 568 87 634 137
rect 368 53 634 87
rect 704 231 756 247
rect 704 197 720 231
rect 754 197 756 231
rect 704 163 756 197
rect 704 129 720 163
rect 754 129 756 163
rect 790 235 856 281
rect 790 201 806 235
rect 840 201 856 235
rect 790 165 856 201
rect 790 131 806 165
rect 840 131 856 165
rect 890 285 1142 319
rect 890 235 956 285
rect 890 201 906 235
rect 940 201 956 235
rect 890 165 956 201
rect 890 131 906 165
rect 940 131 956 165
rect 704 97 756 129
rect 890 97 956 131
rect 704 63 956 97
rect 990 235 1056 251
rect 990 201 1006 235
rect 1040 201 1056 235
rect 990 165 1056 201
rect 990 131 1006 165
rect 1040 131 1056 165
rect 990 17 1056 131
rect 1092 235 1142 285
rect 1176 314 1391 330
rect 1176 280 1205 314
rect 1239 280 1273 314
rect 1307 280 1341 314
rect 1375 280 1391 314
rect 1176 264 1391 280
rect 1126 201 1142 235
rect 1442 226 1511 364
rect 1545 330 1579 464
rect 1615 469 1621 503
rect 1655 469 1661 503
rect 1615 430 1661 469
rect 1695 584 1761 649
rect 1695 550 1711 584
rect 1745 550 1761 584
rect 1695 498 1761 550
rect 1695 464 1711 498
rect 1745 464 1761 498
rect 1815 580 1881 596
rect 1815 546 1831 580
rect 1865 546 1881 580
rect 1815 503 1881 546
rect 1815 469 1831 503
rect 1865 469 1881 503
rect 1815 430 1881 469
rect 1927 580 1993 649
rect 1927 546 1943 580
rect 1977 546 1993 580
rect 1927 500 1993 546
rect 1927 466 1943 500
rect 1977 466 1993 500
rect 1927 464 1993 466
rect 1615 424 1999 430
rect 1615 414 1759 424
rect 1615 380 1621 414
rect 1655 390 1759 414
rect 1793 414 1951 424
rect 1793 390 1831 414
rect 1655 380 1831 390
rect 1865 390 1951 414
rect 1985 390 1999 424
rect 1865 380 1999 390
rect 1615 364 1999 380
rect 1545 314 1929 330
rect 1545 280 1591 314
rect 1625 280 1664 314
rect 1698 280 1743 314
rect 1777 280 1822 314
rect 1856 280 1895 314
rect 1545 264 1929 280
rect 1965 230 1999 364
rect 1092 165 1142 201
rect 1126 131 1142 165
rect 1092 115 1142 131
rect 1184 210 1234 226
rect 1184 176 1200 210
rect 1184 120 1234 176
rect 1184 86 1200 120
rect 1184 17 1234 86
rect 1270 210 1511 226
rect 1270 176 1286 210
rect 1320 176 1458 210
rect 1492 176 1511 210
rect 1630 210 1999 230
rect 1664 196 1830 210
rect 1664 176 1680 196
rect 1270 120 1320 176
rect 1270 86 1286 120
rect 1270 70 1320 86
rect 1356 123 1422 142
rect 1356 89 1372 123
rect 1406 89 1422 123
rect 1356 17 1422 89
rect 1528 123 1594 142
rect 1528 89 1544 123
rect 1578 89 1594 123
rect 1528 17 1594 89
rect 1630 120 1680 176
rect 1814 176 1830 196
rect 1864 196 1999 210
rect 1864 176 1880 196
rect 1664 86 1680 120
rect 1630 70 1680 86
rect 1714 133 1780 162
rect 1714 99 1730 133
rect 1764 99 1780 133
rect 1714 17 1780 99
rect 1814 120 1880 176
rect 1814 86 1830 120
rect 1864 86 1880 120
rect 1814 70 1880 86
rect 1916 146 1977 162
rect 1916 112 1927 146
rect 1961 112 1977 146
rect 1916 17 1977 112
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 1759 390 1793 424
rect 1951 390 1985 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 1747 424 1805 430
rect 1747 390 1759 424
rect 1793 421 1805 424
rect 1939 424 1997 430
rect 1939 421 1951 424
rect 1793 393 1951 421
rect 1793 390 1805 393
rect 1747 384 1805 390
rect 1939 390 1951 393
rect 1985 390 1997 424
rect 1939 384 1997 390
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ha_4
flabel metal1 s 1951 390 1985 424 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 1471 390 1505 424 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 3833044
string GDS_START 3818516
<< end >>
