magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 331 1958 704
rect 311 313 1121 331
<< pwell >>
rect 11 241 285 245
rect 11 49 1904 241
rect 0 0 1920 49
<< scnmos >>
rect 90 51 120 219
rect 176 51 206 219
rect 380 47 410 215
rect 466 47 496 215
rect 586 47 616 215
rect 672 47 702 215
rect 772 47 802 215
rect 858 47 888 215
rect 944 47 974 215
rect 1030 47 1060 215
rect 1193 47 1223 215
rect 1279 47 1309 215
rect 1365 47 1395 215
rect 1451 47 1481 215
rect 1537 47 1567 215
rect 1623 47 1653 215
rect 1709 47 1739 215
rect 1795 47 1825 215
<< scpmoshvt >>
rect 90 367 120 619
rect 176 367 206 619
rect 400 349 430 601
rect 486 349 516 601
rect 572 349 602 601
rect 658 349 688 601
rect 744 349 774 601
rect 830 349 860 601
rect 916 349 946 601
rect 1002 349 1032 601
rect 1192 367 1222 619
rect 1278 367 1308 619
rect 1364 367 1394 619
rect 1450 367 1480 619
rect 1537 367 1567 619
rect 1623 367 1653 619
rect 1709 367 1739 619
rect 1795 367 1825 619
<< ndiff >>
rect 37 207 90 219
rect 37 173 45 207
rect 79 173 90 207
rect 37 101 90 173
rect 37 67 45 101
rect 79 67 90 101
rect 37 51 90 67
rect 120 171 176 219
rect 120 137 131 171
rect 165 137 176 171
rect 120 97 176 137
rect 120 63 131 97
rect 165 63 176 97
rect 120 51 176 63
rect 206 207 259 219
rect 206 173 217 207
rect 251 173 259 207
rect 206 101 259 173
rect 206 67 217 101
rect 251 67 259 101
rect 206 51 259 67
rect 313 163 380 215
rect 313 129 321 163
rect 355 129 380 163
rect 313 93 380 129
rect 313 59 321 93
rect 355 59 380 93
rect 313 47 380 59
rect 410 157 466 215
rect 410 123 421 157
rect 455 123 466 157
rect 410 89 466 123
rect 410 55 421 89
rect 455 55 466 89
rect 410 47 466 55
rect 496 89 586 215
rect 496 55 523 89
rect 557 55 586 89
rect 496 47 586 55
rect 616 157 672 215
rect 616 123 627 157
rect 661 123 672 157
rect 616 89 672 123
rect 616 55 627 89
rect 661 55 672 89
rect 616 47 672 55
rect 702 89 772 215
rect 702 55 727 89
rect 761 55 772 89
rect 702 47 772 55
rect 802 203 858 215
rect 802 169 813 203
rect 847 169 858 203
rect 802 101 858 169
rect 802 67 813 101
rect 847 67 858 101
rect 802 47 858 67
rect 888 165 944 215
rect 888 131 899 165
rect 933 131 944 165
rect 888 89 944 131
rect 888 55 899 89
rect 933 55 944 89
rect 888 47 944 55
rect 974 203 1030 215
rect 974 169 985 203
rect 1019 169 1030 203
rect 974 101 1030 169
rect 974 67 985 101
rect 1019 67 1030 101
rect 974 47 1030 67
rect 1060 163 1193 215
rect 1060 129 1071 163
rect 1105 129 1148 163
rect 1182 129 1193 163
rect 1060 89 1193 129
rect 1060 55 1071 89
rect 1105 55 1148 89
rect 1182 55 1193 89
rect 1060 47 1193 55
rect 1223 203 1279 215
rect 1223 169 1234 203
rect 1268 169 1279 203
rect 1223 101 1279 169
rect 1223 67 1234 101
rect 1268 67 1279 101
rect 1223 47 1279 67
rect 1309 167 1365 215
rect 1309 133 1320 167
rect 1354 133 1365 167
rect 1309 93 1365 133
rect 1309 59 1320 93
rect 1354 59 1365 93
rect 1309 47 1365 59
rect 1395 203 1451 215
rect 1395 169 1406 203
rect 1440 169 1451 203
rect 1395 101 1451 169
rect 1395 67 1406 101
rect 1440 67 1451 101
rect 1395 47 1451 67
rect 1481 167 1537 215
rect 1481 133 1492 167
rect 1526 133 1537 167
rect 1481 93 1537 133
rect 1481 59 1492 93
rect 1526 59 1537 93
rect 1481 47 1537 59
rect 1567 203 1623 215
rect 1567 169 1578 203
rect 1612 169 1623 203
rect 1567 101 1623 169
rect 1567 67 1578 101
rect 1612 67 1623 101
rect 1567 47 1623 67
rect 1653 167 1709 215
rect 1653 133 1664 167
rect 1698 133 1709 167
rect 1653 93 1709 133
rect 1653 59 1664 93
rect 1698 59 1709 93
rect 1653 47 1709 59
rect 1739 203 1795 215
rect 1739 169 1750 203
rect 1784 169 1795 203
rect 1739 101 1795 169
rect 1739 67 1750 101
rect 1784 67 1795 101
rect 1739 47 1795 67
rect 1825 203 1878 215
rect 1825 169 1836 203
rect 1870 169 1878 203
rect 1825 93 1878 169
rect 1825 59 1836 93
rect 1870 59 1878 93
rect 1825 47 1878 59
<< pdiff >>
rect 37 599 90 619
rect 37 565 45 599
rect 79 565 90 599
rect 37 515 90 565
rect 37 481 45 515
rect 79 481 90 515
rect 37 436 90 481
rect 37 402 45 436
rect 79 402 90 436
rect 37 367 90 402
rect 120 577 176 619
rect 120 543 131 577
rect 165 543 176 577
rect 120 367 176 543
rect 206 424 259 619
rect 206 390 217 424
rect 251 390 259 424
rect 206 367 259 390
rect 347 576 400 601
rect 347 542 355 576
rect 389 542 400 576
rect 347 349 400 542
rect 430 531 486 601
rect 430 497 441 531
rect 475 497 486 531
rect 430 463 486 497
rect 430 429 441 463
rect 475 429 486 463
rect 430 391 486 429
rect 430 357 441 391
rect 475 357 486 391
rect 430 349 486 357
rect 516 593 572 601
rect 516 559 527 593
rect 561 559 572 593
rect 516 518 572 559
rect 516 484 527 518
rect 561 484 572 518
rect 516 439 572 484
rect 516 405 527 439
rect 561 405 572 439
rect 516 349 572 405
rect 602 531 658 601
rect 602 497 613 531
rect 647 497 658 531
rect 602 459 658 497
rect 602 425 613 459
rect 647 425 658 459
rect 602 391 658 425
rect 602 357 613 391
rect 647 357 658 391
rect 602 349 658 357
rect 688 593 744 601
rect 688 559 699 593
rect 733 559 744 593
rect 688 525 744 559
rect 688 491 699 525
rect 733 491 744 525
rect 688 457 744 491
rect 688 423 699 457
rect 733 423 744 457
rect 688 349 744 423
rect 774 589 830 601
rect 774 555 785 589
rect 819 555 830 589
rect 774 513 830 555
rect 774 479 785 513
rect 819 479 830 513
rect 774 349 830 479
rect 860 531 916 601
rect 860 497 871 531
rect 905 497 916 531
rect 860 441 916 497
rect 860 407 871 441
rect 905 407 916 441
rect 860 349 916 407
rect 946 589 1002 601
rect 946 555 957 589
rect 991 555 1002 589
rect 946 513 1002 555
rect 946 479 957 513
rect 991 479 1002 513
rect 946 349 1002 479
rect 1032 527 1085 601
rect 1032 493 1043 527
rect 1077 493 1085 527
rect 1032 457 1085 493
rect 1032 423 1043 457
rect 1077 423 1085 457
rect 1032 349 1085 423
rect 1139 525 1192 619
rect 1139 491 1147 525
rect 1181 491 1192 525
rect 1139 441 1192 491
rect 1139 407 1147 441
rect 1181 407 1192 441
rect 1139 367 1192 407
rect 1222 599 1278 619
rect 1222 565 1233 599
rect 1267 565 1278 599
rect 1222 515 1278 565
rect 1222 481 1233 515
rect 1267 481 1278 515
rect 1222 367 1278 481
rect 1308 527 1364 619
rect 1308 493 1319 527
rect 1353 493 1364 527
rect 1308 413 1364 493
rect 1308 379 1319 413
rect 1353 379 1364 413
rect 1308 367 1364 379
rect 1394 599 1450 619
rect 1394 565 1405 599
rect 1439 565 1450 599
rect 1394 523 1450 565
rect 1394 489 1405 523
rect 1439 489 1450 523
rect 1394 445 1450 489
rect 1394 411 1405 445
rect 1439 411 1450 445
rect 1394 367 1450 411
rect 1480 599 1537 619
rect 1480 565 1491 599
rect 1525 565 1537 599
rect 1480 510 1537 565
rect 1480 476 1491 510
rect 1525 476 1537 510
rect 1480 413 1537 476
rect 1480 379 1491 413
rect 1525 379 1537 413
rect 1480 367 1537 379
rect 1567 607 1623 619
rect 1567 573 1578 607
rect 1612 573 1623 607
rect 1567 493 1623 573
rect 1567 459 1578 493
rect 1612 459 1623 493
rect 1567 367 1623 459
rect 1653 599 1709 619
rect 1653 565 1664 599
rect 1698 565 1709 599
rect 1653 515 1709 565
rect 1653 481 1664 515
rect 1698 481 1709 515
rect 1653 420 1709 481
rect 1653 386 1664 420
rect 1698 386 1709 420
rect 1653 367 1709 386
rect 1739 607 1795 619
rect 1739 573 1750 607
rect 1784 573 1795 607
rect 1739 493 1795 573
rect 1739 459 1750 493
rect 1784 459 1795 493
rect 1739 367 1795 459
rect 1825 599 1878 619
rect 1825 565 1836 599
rect 1870 565 1878 599
rect 1825 515 1878 565
rect 1825 481 1836 515
rect 1870 481 1878 515
rect 1825 420 1878 481
rect 1825 386 1836 420
rect 1870 386 1878 420
rect 1825 367 1878 386
<< ndiffc >>
rect 45 173 79 207
rect 45 67 79 101
rect 131 137 165 171
rect 131 63 165 97
rect 217 173 251 207
rect 217 67 251 101
rect 321 129 355 163
rect 321 59 355 93
rect 421 123 455 157
rect 421 55 455 89
rect 523 55 557 89
rect 627 123 661 157
rect 627 55 661 89
rect 727 55 761 89
rect 813 169 847 203
rect 813 67 847 101
rect 899 131 933 165
rect 899 55 933 89
rect 985 169 1019 203
rect 985 67 1019 101
rect 1071 129 1105 163
rect 1148 129 1182 163
rect 1071 55 1105 89
rect 1148 55 1182 89
rect 1234 169 1268 203
rect 1234 67 1268 101
rect 1320 133 1354 167
rect 1320 59 1354 93
rect 1406 169 1440 203
rect 1406 67 1440 101
rect 1492 133 1526 167
rect 1492 59 1526 93
rect 1578 169 1612 203
rect 1578 67 1612 101
rect 1664 133 1698 167
rect 1664 59 1698 93
rect 1750 169 1784 203
rect 1750 67 1784 101
rect 1836 169 1870 203
rect 1836 59 1870 93
<< pdiffc >>
rect 45 565 79 599
rect 45 481 79 515
rect 45 402 79 436
rect 131 543 165 577
rect 217 390 251 424
rect 355 542 389 576
rect 441 497 475 531
rect 441 429 475 463
rect 441 357 475 391
rect 527 559 561 593
rect 527 484 561 518
rect 527 405 561 439
rect 613 497 647 531
rect 613 425 647 459
rect 613 357 647 391
rect 699 559 733 593
rect 699 491 733 525
rect 699 423 733 457
rect 785 555 819 589
rect 785 479 819 513
rect 871 497 905 531
rect 871 407 905 441
rect 957 555 991 589
rect 957 479 991 513
rect 1043 493 1077 527
rect 1043 423 1077 457
rect 1147 491 1181 525
rect 1147 407 1181 441
rect 1233 565 1267 599
rect 1233 481 1267 515
rect 1319 493 1353 527
rect 1319 379 1353 413
rect 1405 565 1439 599
rect 1405 489 1439 523
rect 1405 411 1439 445
rect 1491 565 1525 599
rect 1491 476 1525 510
rect 1491 379 1525 413
rect 1578 573 1612 607
rect 1578 459 1612 493
rect 1664 565 1698 599
rect 1664 481 1698 515
rect 1664 386 1698 420
rect 1750 573 1784 607
rect 1750 459 1784 493
rect 1836 565 1870 599
rect 1836 481 1870 515
rect 1836 386 1870 420
<< poly >>
rect 90 619 120 645
rect 176 619 206 645
rect 400 601 430 627
rect 486 601 516 627
rect 572 601 602 627
rect 658 601 688 627
rect 744 601 774 627
rect 830 601 860 627
rect 916 601 946 627
rect 1002 601 1032 627
rect 1192 619 1222 645
rect 1278 619 1308 645
rect 1364 619 1394 645
rect 1450 619 1480 645
rect 1537 619 1567 645
rect 1623 619 1653 645
rect 1709 619 1739 645
rect 1795 619 1825 645
rect 90 325 120 367
rect 29 309 120 325
rect 29 275 45 309
rect 79 275 120 309
rect 29 259 120 275
rect 90 219 120 259
rect 176 335 206 367
rect 176 319 251 335
rect 176 285 201 319
rect 235 285 251 319
rect 400 317 430 349
rect 486 317 516 349
rect 572 317 602 349
rect 658 317 688 349
rect 744 317 774 349
rect 830 317 860 349
rect 916 317 946 349
rect 1002 317 1032 349
rect 1192 321 1222 367
rect 1278 321 1308 367
rect 1364 321 1394 367
rect 1450 321 1480 367
rect 1537 325 1567 367
rect 1623 325 1653 367
rect 1709 325 1739 367
rect 1795 325 1825 367
rect 176 269 251 285
rect 364 301 702 317
rect 176 219 206 269
rect 364 267 380 301
rect 414 267 448 301
rect 482 267 516 301
rect 550 267 584 301
rect 618 267 652 301
rect 686 267 702 301
rect 364 251 702 267
rect 744 301 1060 317
rect 744 267 760 301
rect 794 267 828 301
rect 862 267 896 301
rect 930 267 964 301
rect 998 267 1060 301
rect 744 251 1060 267
rect 1157 305 1495 321
rect 1157 271 1173 305
rect 1207 271 1241 305
rect 1275 271 1309 305
rect 1343 271 1377 305
rect 1411 271 1445 305
rect 1479 271 1495 305
rect 1157 255 1495 271
rect 1537 309 1899 325
rect 1537 275 1577 309
rect 1611 275 1645 309
rect 1679 275 1713 309
rect 1747 275 1781 309
rect 1815 275 1849 309
rect 1883 275 1899 309
rect 1537 259 1899 275
rect 380 215 410 251
rect 466 215 496 251
rect 586 215 616 251
rect 672 215 702 251
rect 772 215 802 251
rect 858 215 888 251
rect 944 215 974 251
rect 1030 215 1060 251
rect 1193 215 1223 255
rect 1279 215 1309 255
rect 1365 215 1395 255
rect 1451 215 1481 255
rect 1537 215 1567 259
rect 1623 215 1653 259
rect 1709 215 1739 259
rect 1795 215 1825 259
rect 90 25 120 51
rect 176 25 206 51
rect 380 21 410 47
rect 466 21 496 47
rect 586 21 616 47
rect 672 21 702 47
rect 772 21 802 47
rect 858 21 888 47
rect 944 21 974 47
rect 1030 21 1060 47
rect 1193 21 1223 47
rect 1279 21 1309 47
rect 1365 21 1395 47
rect 1451 21 1481 47
rect 1537 21 1567 47
rect 1623 21 1653 47
rect 1709 21 1739 47
rect 1795 21 1825 47
<< polycont >>
rect 45 275 79 309
rect 201 285 235 319
rect 380 267 414 301
rect 448 267 482 301
rect 516 267 550 301
rect 584 267 618 301
rect 652 267 686 301
rect 760 267 794 301
rect 828 267 862 301
rect 896 267 930 301
rect 964 267 998 301
rect 1173 271 1207 305
rect 1241 271 1275 305
rect 1309 271 1343 305
rect 1377 271 1411 305
rect 1445 271 1479 305
rect 1577 275 1611 309
rect 1645 275 1679 309
rect 1713 275 1747 309
rect 1781 275 1815 309
rect 1849 275 1883 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 29 599 81 615
rect 29 565 45 599
rect 79 565 81 599
rect 29 515 81 565
rect 115 577 181 649
rect 115 543 131 577
rect 165 543 181 577
rect 115 530 181 543
rect 339 593 735 615
rect 339 581 527 593
rect 339 576 405 581
rect 339 542 355 576
rect 389 542 405 576
rect 511 559 527 581
rect 561 581 699 593
rect 561 559 577 581
rect 339 530 405 542
rect 439 531 477 547
rect 29 481 45 515
rect 79 496 81 515
rect 439 497 441 531
rect 475 497 477 531
rect 79 481 405 496
rect 29 462 405 481
rect 29 436 165 462
rect 29 402 45 436
rect 79 402 165 436
rect 29 386 165 402
rect 201 424 327 428
rect 201 390 217 424
rect 251 390 327 424
rect 201 386 327 390
rect 17 309 95 352
rect 17 275 45 309
rect 79 275 95 309
rect 129 239 165 386
rect 199 319 257 352
rect 199 285 201 319
rect 235 285 257 319
rect 199 269 257 285
rect 29 207 165 239
rect 291 235 327 386
rect 364 303 405 462
rect 439 463 477 497
rect 439 429 441 463
rect 475 429 477 463
rect 439 391 477 429
rect 511 518 577 559
rect 691 559 699 581
rect 733 559 735 593
rect 511 484 527 518
rect 561 484 577 518
rect 511 439 577 484
rect 511 405 527 439
rect 561 405 577 439
rect 611 531 657 547
rect 611 497 613 531
rect 647 497 657 531
rect 611 459 657 497
rect 611 425 613 459
rect 647 425 657 459
rect 439 357 441 391
rect 475 371 477 391
rect 611 391 657 425
rect 691 525 735 559
rect 691 491 699 525
rect 733 491 735 525
rect 691 457 735 491
rect 769 599 1455 615
rect 769 589 1233 599
rect 769 555 785 589
rect 819 581 957 589
rect 819 555 835 581
rect 769 513 835 555
rect 941 555 957 581
rect 991 577 1233 589
rect 991 555 1007 577
rect 769 479 785 513
rect 819 479 835 513
rect 769 475 835 479
rect 869 531 907 547
rect 869 497 871 531
rect 905 497 907 531
rect 691 423 699 457
rect 733 441 735 457
rect 869 441 907 497
rect 941 513 1007 555
rect 1217 565 1233 577
rect 1267 577 1405 599
rect 1267 565 1283 577
rect 941 479 957 513
rect 991 479 1007 513
rect 941 475 1007 479
rect 1041 527 1093 543
rect 1041 493 1043 527
rect 1077 493 1093 527
rect 1041 457 1093 493
rect 1041 441 1043 457
rect 733 423 871 441
rect 691 407 871 423
rect 905 423 1043 441
rect 1077 423 1093 457
rect 905 407 1093 423
rect 1131 525 1183 543
rect 1131 491 1147 525
rect 1181 491 1183 525
rect 1131 441 1183 491
rect 1217 515 1283 565
rect 1389 565 1405 577
rect 1439 565 1455 599
rect 1217 481 1233 515
rect 1267 481 1283 515
rect 1217 475 1283 481
rect 1317 527 1355 543
rect 1317 493 1319 527
rect 1353 493 1355 527
rect 1317 441 1355 493
rect 1131 407 1147 441
rect 1181 413 1355 441
rect 1181 407 1319 413
rect 611 371 613 391
rect 475 357 613 371
rect 647 373 657 391
rect 1303 379 1319 407
rect 1353 379 1355 413
rect 1389 523 1455 565
rect 1389 489 1405 523
rect 1439 489 1455 523
rect 1389 445 1455 489
rect 1389 411 1405 445
rect 1439 411 1455 445
rect 1489 599 1528 615
rect 1489 565 1491 599
rect 1525 565 1528 599
rect 1489 510 1528 565
rect 1489 476 1491 510
rect 1525 476 1528 510
rect 1489 420 1528 476
rect 1562 607 1628 649
rect 1562 573 1578 607
rect 1612 573 1628 607
rect 1562 493 1628 573
rect 1562 459 1578 493
rect 1612 459 1628 493
rect 1562 454 1628 459
rect 1662 599 1700 615
rect 1662 565 1664 599
rect 1698 565 1700 599
rect 1662 515 1700 565
rect 1662 481 1664 515
rect 1698 481 1700 515
rect 1662 420 1700 481
rect 1734 607 1800 649
rect 1734 573 1750 607
rect 1784 573 1800 607
rect 1734 493 1800 573
rect 1734 459 1750 493
rect 1784 459 1800 493
rect 1734 454 1800 459
rect 1834 599 1886 615
rect 1834 565 1836 599
rect 1870 565 1886 599
rect 1834 515 1886 565
rect 1834 481 1836 515
rect 1870 481 1886 515
rect 1834 420 1886 481
rect 1489 413 1664 420
rect 1303 375 1355 379
rect 1489 379 1491 413
rect 1525 386 1664 413
rect 1698 386 1836 420
rect 1870 386 1886 420
rect 1489 375 1525 379
rect 647 357 1123 373
rect 439 337 1123 357
rect 364 301 702 303
rect 364 267 380 301
rect 414 267 448 301
rect 482 267 516 301
rect 550 267 584 301
rect 618 267 652 301
rect 686 267 702 301
rect 744 301 1014 303
rect 744 267 760 301
rect 794 267 828 301
rect 862 267 896 301
rect 930 267 964 301
rect 998 267 1014 301
rect 29 173 45 207
rect 79 205 165 207
rect 215 233 327 235
rect 744 233 778 267
rect 1050 235 1123 337
rect 1157 305 1241 366
rect 1303 341 1525 375
rect 1559 309 1899 352
rect 1157 271 1173 305
rect 1207 271 1241 305
rect 1275 271 1309 305
rect 1343 271 1377 305
rect 1411 271 1445 305
rect 1479 271 1495 305
rect 1559 275 1577 309
rect 1611 275 1645 309
rect 1679 275 1713 309
rect 1747 275 1781 309
rect 1815 275 1849 309
rect 1883 275 1899 309
rect 1050 233 1793 235
rect 215 207 778 233
rect 29 101 79 173
rect 215 173 217 207
rect 251 199 778 207
rect 812 203 1793 233
rect 251 173 267 199
rect 29 67 45 101
rect 29 51 79 67
rect 115 137 131 171
rect 165 137 181 171
rect 115 97 181 137
rect 115 63 131 97
rect 165 63 181 97
rect 115 17 181 63
rect 215 101 267 173
rect 812 169 813 203
rect 847 199 985 203
rect 847 169 849 199
rect 812 165 849 169
rect 983 169 985 199
rect 1019 197 1234 203
rect 1019 169 1021 197
rect 215 67 217 101
rect 251 67 267 101
rect 215 51 267 67
rect 305 129 321 163
rect 355 129 371 163
rect 305 93 371 129
rect 305 59 321 93
rect 355 59 371 93
rect 305 17 371 59
rect 405 157 849 165
rect 405 123 421 157
rect 455 131 627 157
rect 455 123 473 131
rect 405 89 473 123
rect 611 123 627 131
rect 661 131 849 157
rect 661 123 677 131
rect 405 55 421 89
rect 455 55 473 89
rect 405 51 473 55
rect 507 89 573 97
rect 507 55 523 89
rect 557 55 573 89
rect 507 17 573 55
rect 611 89 677 123
rect 811 101 849 131
rect 611 55 627 89
rect 661 55 677 89
rect 611 51 677 55
rect 711 89 777 97
rect 711 55 727 89
rect 761 55 777 89
rect 711 17 777 55
rect 811 67 813 101
rect 847 67 849 101
rect 811 51 849 67
rect 883 131 899 165
rect 933 131 949 165
rect 883 89 949 131
rect 883 55 899 89
rect 933 55 949 89
rect 883 17 949 55
rect 983 101 1021 169
rect 1232 169 1234 197
rect 1268 201 1406 203
rect 1268 169 1270 201
rect 983 67 985 101
rect 1019 67 1021 101
rect 983 51 1021 67
rect 1055 129 1071 163
rect 1105 129 1148 163
rect 1182 129 1198 163
rect 1055 89 1198 129
rect 1055 55 1071 89
rect 1105 55 1148 89
rect 1182 55 1198 89
rect 1055 17 1198 55
rect 1232 101 1270 169
rect 1404 169 1406 201
rect 1440 201 1578 203
rect 1440 169 1442 201
rect 1232 67 1234 101
rect 1268 67 1270 101
rect 1232 51 1270 67
rect 1304 133 1320 167
rect 1354 133 1370 167
rect 1304 93 1370 133
rect 1304 59 1320 93
rect 1354 59 1370 93
rect 1304 17 1370 59
rect 1404 101 1442 169
rect 1576 169 1578 201
rect 1612 201 1750 203
rect 1612 169 1614 201
rect 1404 67 1406 101
rect 1440 67 1442 101
rect 1404 51 1442 67
rect 1476 133 1492 167
rect 1526 133 1542 167
rect 1476 93 1542 133
rect 1476 59 1492 93
rect 1526 59 1542 93
rect 1476 17 1542 59
rect 1576 101 1614 169
rect 1748 169 1750 201
rect 1784 169 1793 203
rect 1576 67 1578 101
rect 1612 67 1614 101
rect 1576 51 1614 67
rect 1648 133 1664 167
rect 1698 133 1714 167
rect 1648 93 1714 133
rect 1648 59 1664 93
rect 1698 59 1714 93
rect 1648 17 1714 59
rect 1748 101 1793 169
rect 1748 67 1750 101
rect 1784 67 1793 101
rect 1748 51 1793 67
rect 1827 203 1886 219
rect 1827 169 1836 203
rect 1870 169 1886 203
rect 1827 93 1886 169
rect 1827 59 1836 93
rect 1870 59 1886 93
rect 1827 17 1886 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4bb_4
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3376264
string GDS_START 3360376
<< end >>
