magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 187 49 977 180
rect 0 0 1152 49
<< scnmos >>
rect 266 70 296 154
rect 352 70 382 154
rect 438 70 468 154
rect 524 70 554 154
rect 610 70 640 154
rect 696 70 726 154
rect 782 70 812 154
rect 868 70 898 154
<< scpmoshvt >>
rect 94 367 124 619
rect 180 367 210 619
rect 266 367 296 619
rect 352 367 382 619
rect 438 367 468 619
rect 524 367 554 619
rect 610 367 640 619
rect 696 367 726 619
rect 782 367 812 619
rect 868 367 898 619
rect 954 367 984 619
rect 1040 367 1070 619
<< ndiff >>
rect 213 118 266 154
rect 213 84 221 118
rect 255 84 266 118
rect 213 70 266 84
rect 296 129 352 154
rect 296 95 307 129
rect 341 95 352 129
rect 296 70 352 95
rect 382 118 438 154
rect 382 84 393 118
rect 427 84 438 118
rect 382 70 438 84
rect 468 129 524 154
rect 468 95 479 129
rect 513 95 524 129
rect 468 70 524 95
rect 554 118 610 154
rect 554 84 565 118
rect 599 84 610 118
rect 554 70 610 84
rect 640 129 696 154
rect 640 95 651 129
rect 685 95 696 129
rect 640 70 696 95
rect 726 118 782 154
rect 726 84 737 118
rect 771 84 782 118
rect 726 70 782 84
rect 812 129 868 154
rect 812 95 823 129
rect 857 95 868 129
rect 812 70 868 95
rect 898 118 951 154
rect 898 84 909 118
rect 943 84 951 118
rect 898 70 951 84
<< pdiff >>
rect 41 599 94 619
rect 41 565 49 599
rect 83 565 94 599
rect 41 529 94 565
rect 41 495 49 529
rect 83 495 94 529
rect 41 461 94 495
rect 41 427 49 461
rect 83 427 94 461
rect 41 367 94 427
rect 124 593 180 619
rect 124 559 135 593
rect 169 559 180 593
rect 124 505 180 559
rect 124 471 135 505
rect 169 471 180 505
rect 124 417 180 471
rect 124 383 135 417
rect 169 383 180 417
rect 124 367 180 383
rect 210 599 266 619
rect 210 565 221 599
rect 255 565 266 599
rect 210 529 266 565
rect 210 495 221 529
rect 255 495 266 529
rect 210 461 266 495
rect 210 427 221 461
rect 255 427 266 461
rect 210 367 266 427
rect 296 593 352 619
rect 296 559 307 593
rect 341 559 352 593
rect 296 505 352 559
rect 296 471 307 505
rect 341 471 352 505
rect 296 417 352 471
rect 296 383 307 417
rect 341 383 352 417
rect 296 367 352 383
rect 382 599 438 619
rect 382 565 393 599
rect 427 565 438 599
rect 382 529 438 565
rect 382 495 393 529
rect 427 495 438 529
rect 382 461 438 495
rect 382 427 393 461
rect 427 427 438 461
rect 382 367 438 427
rect 468 593 524 619
rect 468 559 479 593
rect 513 559 524 593
rect 468 505 524 559
rect 468 471 479 505
rect 513 471 524 505
rect 468 417 524 471
rect 468 383 479 417
rect 513 383 524 417
rect 468 367 524 383
rect 554 599 610 619
rect 554 565 565 599
rect 599 565 610 599
rect 554 529 610 565
rect 554 495 565 529
rect 599 495 610 529
rect 554 461 610 495
rect 554 427 565 461
rect 599 427 610 461
rect 554 367 610 427
rect 640 593 696 619
rect 640 559 651 593
rect 685 559 696 593
rect 640 505 696 559
rect 640 471 651 505
rect 685 471 696 505
rect 640 417 696 471
rect 640 383 651 417
rect 685 383 696 417
rect 640 367 696 383
rect 726 599 782 619
rect 726 565 737 599
rect 771 565 782 599
rect 726 529 782 565
rect 726 495 737 529
rect 771 495 782 529
rect 726 461 782 495
rect 726 427 737 461
rect 771 427 782 461
rect 726 367 782 427
rect 812 593 868 619
rect 812 559 823 593
rect 857 559 868 593
rect 812 505 868 559
rect 812 471 823 505
rect 857 471 868 505
rect 812 417 868 471
rect 812 383 823 417
rect 857 383 868 417
rect 812 367 868 383
rect 898 599 954 619
rect 898 565 909 599
rect 943 565 954 599
rect 898 529 954 565
rect 898 495 909 529
rect 943 495 954 529
rect 898 461 954 495
rect 898 427 909 461
rect 943 427 954 461
rect 898 367 954 427
rect 984 593 1040 619
rect 984 559 995 593
rect 1029 559 1040 593
rect 984 505 1040 559
rect 984 471 995 505
rect 1029 471 1040 505
rect 984 417 1040 471
rect 984 383 995 417
rect 1029 383 1040 417
rect 984 367 1040 383
rect 1070 599 1123 619
rect 1070 565 1081 599
rect 1115 565 1123 599
rect 1070 529 1123 565
rect 1070 495 1081 529
rect 1115 495 1123 529
rect 1070 461 1123 495
rect 1070 427 1081 461
rect 1115 427 1123 461
rect 1070 367 1123 427
<< ndiffc >>
rect 221 84 255 118
rect 307 95 341 129
rect 393 84 427 118
rect 479 95 513 129
rect 565 84 599 118
rect 651 95 685 129
rect 737 84 771 118
rect 823 95 857 129
rect 909 84 943 118
<< pdiffc >>
rect 49 565 83 599
rect 49 495 83 529
rect 49 427 83 461
rect 135 559 169 593
rect 135 471 169 505
rect 135 383 169 417
rect 221 565 255 599
rect 221 495 255 529
rect 221 427 255 461
rect 307 559 341 593
rect 307 471 341 505
rect 307 383 341 417
rect 393 565 427 599
rect 393 495 427 529
rect 393 427 427 461
rect 479 559 513 593
rect 479 471 513 505
rect 479 383 513 417
rect 565 565 599 599
rect 565 495 599 529
rect 565 427 599 461
rect 651 559 685 593
rect 651 471 685 505
rect 651 383 685 417
rect 737 565 771 599
rect 737 495 771 529
rect 737 427 771 461
rect 823 559 857 593
rect 823 471 857 505
rect 823 383 857 417
rect 909 565 943 599
rect 909 495 943 529
rect 909 427 943 461
rect 995 559 1029 593
rect 995 471 1029 505
rect 995 383 1029 417
rect 1081 565 1115 599
rect 1081 495 1115 529
rect 1081 427 1115 461
<< poly >>
rect 94 619 124 645
rect 180 619 210 645
rect 266 619 296 645
rect 352 619 382 645
rect 438 619 468 645
rect 524 619 554 645
rect 610 619 640 645
rect 696 619 726 645
rect 782 619 812 645
rect 868 619 898 645
rect 954 619 984 645
rect 1040 619 1070 645
rect 94 308 124 367
rect 180 308 210 367
rect 266 308 296 367
rect 352 308 382 367
rect 438 308 468 367
rect 524 308 554 367
rect 610 308 640 367
rect 696 308 726 367
rect 782 308 812 367
rect 868 308 898 367
rect 954 308 984 367
rect 1040 308 1070 367
rect 94 292 1070 308
rect 94 258 119 292
rect 153 258 187 292
rect 221 258 255 292
rect 289 258 323 292
rect 357 258 391 292
rect 425 258 459 292
rect 493 258 527 292
rect 561 258 595 292
rect 629 258 663 292
rect 697 258 731 292
rect 765 258 799 292
rect 833 258 867 292
rect 901 258 935 292
rect 969 258 1003 292
rect 1037 258 1070 292
rect 94 242 1070 258
rect 266 154 296 242
rect 352 154 382 242
rect 438 154 468 242
rect 524 154 554 242
rect 610 154 640 242
rect 696 154 726 242
rect 782 154 812 242
rect 868 154 898 242
rect 266 44 296 70
rect 352 44 382 70
rect 438 44 468 70
rect 524 44 554 70
rect 610 44 640 70
rect 696 44 726 70
rect 782 44 812 70
rect 868 44 898 70
<< polycont >>
rect 119 258 153 292
rect 187 258 221 292
rect 255 258 289 292
rect 323 258 357 292
rect 391 258 425 292
rect 459 258 493 292
rect 527 258 561 292
rect 595 258 629 292
rect 663 258 697 292
rect 731 258 765 292
rect 799 258 833 292
rect 867 258 901 292
rect 935 258 969 292
rect 1003 258 1037 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 40 599 92 615
rect 40 545 49 599
rect 83 545 92 599
rect 40 529 92 545
rect 40 495 49 529
rect 83 495 92 529
rect 40 461 92 495
rect 40 427 49 461
rect 83 427 92 461
rect 40 411 92 427
rect 127 593 178 609
rect 127 559 135 593
rect 169 559 178 593
rect 127 505 178 559
rect 127 471 135 505
rect 169 471 178 505
rect 127 417 178 471
rect 127 383 135 417
rect 169 383 178 417
rect 212 599 264 615
rect 212 579 221 599
rect 212 545 220 579
rect 255 565 264 599
rect 254 545 264 565
rect 212 529 264 545
rect 212 495 221 529
rect 255 495 264 529
rect 212 461 264 495
rect 212 427 221 461
rect 255 427 264 461
rect 212 411 264 427
rect 299 593 350 609
rect 299 559 307 593
rect 341 559 350 593
rect 299 505 350 559
rect 299 471 307 505
rect 341 471 350 505
rect 299 417 350 471
rect 127 377 178 383
rect 299 383 307 417
rect 341 383 350 417
rect 384 599 436 615
rect 384 565 393 599
rect 427 579 436 599
rect 384 545 394 565
rect 428 545 436 579
rect 384 529 436 545
rect 384 495 393 529
rect 427 495 436 529
rect 384 461 436 495
rect 384 427 393 461
rect 427 427 436 461
rect 384 411 436 427
rect 471 593 522 609
rect 471 559 479 593
rect 513 559 522 593
rect 471 505 522 559
rect 471 471 479 505
rect 513 471 522 505
rect 471 417 522 471
rect 299 377 350 383
rect 471 383 479 417
rect 513 383 522 417
rect 556 599 608 615
rect 556 545 565 599
rect 599 545 608 599
rect 556 529 608 545
rect 556 495 565 529
rect 599 495 608 529
rect 556 461 608 495
rect 556 427 565 461
rect 599 427 608 461
rect 556 411 608 427
rect 643 593 694 609
rect 643 559 651 593
rect 685 559 694 593
rect 643 505 694 559
rect 643 471 651 505
rect 685 471 694 505
rect 643 417 694 471
rect 471 377 522 383
rect 643 383 651 417
rect 685 383 694 417
rect 728 599 780 615
rect 728 565 737 599
rect 771 579 780 599
rect 728 545 738 565
rect 772 545 780 579
rect 728 529 780 545
rect 728 495 737 529
rect 771 495 780 529
rect 728 461 780 495
rect 728 427 737 461
rect 771 427 780 461
rect 728 411 780 427
rect 815 593 866 609
rect 815 559 823 593
rect 857 559 866 593
rect 815 505 866 559
rect 815 471 823 505
rect 857 471 866 505
rect 815 417 866 471
rect 643 377 694 383
rect 815 383 823 417
rect 857 383 866 417
rect 900 599 952 615
rect 900 565 909 599
rect 943 579 952 599
rect 900 545 910 565
rect 944 545 952 579
rect 900 529 952 545
rect 900 495 909 529
rect 943 495 952 529
rect 900 461 952 495
rect 900 427 909 461
rect 943 427 952 461
rect 900 411 952 427
rect 986 593 1038 609
rect 986 559 995 593
rect 1029 559 1038 593
rect 986 505 1038 559
rect 986 471 995 505
rect 1029 471 1038 505
rect 986 417 1038 471
rect 815 377 866 383
rect 986 383 995 417
rect 1029 383 1038 417
rect 1072 599 1123 615
rect 1072 565 1081 599
rect 1115 579 1123 599
rect 1072 545 1082 565
rect 1116 545 1123 579
rect 1072 529 1123 545
rect 1072 495 1081 529
rect 1115 495 1123 529
rect 1072 461 1123 495
rect 1072 427 1081 461
rect 1115 427 1123 461
rect 1072 411 1123 427
rect 986 377 1038 383
rect 35 342 1124 377
rect 35 208 69 342
rect 103 292 1053 308
rect 103 258 119 292
rect 153 258 187 292
rect 221 258 255 292
rect 289 258 323 292
rect 357 258 391 292
rect 425 258 459 292
rect 493 258 527 292
rect 561 258 595 292
rect 629 258 663 292
rect 697 258 731 292
rect 765 258 799 292
rect 833 258 867 292
rect 901 258 935 292
rect 969 258 1003 292
rect 1037 258 1053 292
rect 103 242 1053 258
rect 1087 208 1124 342
rect 35 168 1124 208
rect 205 118 264 134
rect 205 84 221 118
rect 255 84 264 118
rect 205 17 264 84
rect 298 129 350 168
rect 298 95 307 129
rect 341 95 350 129
rect 298 79 350 95
rect 384 118 436 134
rect 384 84 393 118
rect 427 84 436 118
rect 384 17 436 84
rect 470 129 522 168
rect 470 95 479 129
rect 513 95 522 129
rect 470 79 522 95
rect 556 118 608 134
rect 556 84 565 118
rect 599 84 608 118
rect 556 17 608 84
rect 642 129 694 168
rect 642 95 651 129
rect 685 95 694 129
rect 642 79 694 95
rect 728 118 780 134
rect 728 84 737 118
rect 771 84 780 118
rect 728 17 780 84
rect 814 129 866 168
rect 814 95 823 129
rect 857 95 866 129
rect 814 79 866 95
rect 900 118 959 134
rect 900 84 909 118
rect 943 84 959 118
rect 900 17 959 84
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 49 565 83 579
rect 49 545 83 565
rect 220 565 221 579
rect 221 565 254 579
rect 220 545 254 565
rect 394 565 427 579
rect 427 565 428 579
rect 394 545 428 565
rect 565 565 599 579
rect 565 545 599 565
rect 738 565 771 579
rect 771 565 772 579
rect 738 545 772 565
rect 910 565 943 579
rect 943 565 944 579
rect 910 545 944 565
rect 1082 565 1115 579
rect 1115 565 1116 579
rect 1082 545 1116 565
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 14 579 1138 589
rect 14 545 49 579
rect 83 545 220 579
rect 254 545 394 579
rect 428 545 565 579
rect 599 545 738 579
rect 772 545 910 579
rect 944 545 1082 579
rect 1116 545 1138 579
rect 14 538 1138 545
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 invkapwr_8
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 14 538 1138 589 0 FreeSans 200 0 0 0 KAPWR
port 2 nsew power bidirectional
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y
string GDS_END 3700086
string GDS_START 3689228
<< end >>
