magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 337 710 704
rect -38 331 150 337
rect 441 331 710 337
<< pwell >>
rect 192 289 399 295
rect 1 157 399 289
rect 1 49 671 157
rect 0 0 672 49
<< scnmos >>
rect 80 179 110 263
rect 166 179 196 263
rect 290 185 320 269
rect 390 47 420 131
rect 476 47 506 131
rect 562 47 592 131
<< scpmoshvt >>
rect 89 535 119 619
rect 208 535 238 619
rect 280 535 310 619
rect 366 535 396 619
rect 460 535 490 619
rect 553 535 583 619
<< ndiff >>
rect 218 263 290 269
rect 27 251 80 263
rect 27 217 35 251
rect 69 217 80 251
rect 27 179 80 217
rect 110 251 166 263
rect 110 217 121 251
rect 155 217 166 251
rect 110 179 166 217
rect 196 225 290 263
rect 196 191 226 225
rect 260 191 290 225
rect 196 185 290 191
rect 320 257 373 269
rect 320 223 331 257
rect 365 223 373 257
rect 320 185 373 223
rect 196 179 268 185
rect 333 93 390 131
rect 333 59 341 93
rect 375 59 390 93
rect 333 47 390 59
rect 420 119 476 131
rect 420 85 431 119
rect 465 85 476 119
rect 420 47 476 85
rect 506 93 562 131
rect 506 59 517 93
rect 551 59 562 93
rect 506 47 562 59
rect 592 119 645 131
rect 592 85 603 119
rect 637 85 645 119
rect 592 47 645 85
<< pdiff >>
rect 36 581 89 619
rect 36 547 44 581
rect 78 547 89 581
rect 36 535 89 547
rect 119 607 208 619
rect 119 573 146 607
rect 180 573 208 607
rect 119 535 208 573
rect 238 535 280 619
rect 310 589 366 619
rect 310 555 321 589
rect 355 555 366 589
rect 310 535 366 555
rect 396 535 460 619
rect 490 607 553 619
rect 490 573 508 607
rect 542 573 553 607
rect 490 535 553 573
rect 583 581 636 619
rect 583 547 594 581
rect 628 547 636 581
rect 583 535 636 547
<< ndiffc >>
rect 35 217 69 251
rect 121 217 155 251
rect 226 191 260 225
rect 331 223 365 257
rect 341 59 375 93
rect 431 85 465 119
rect 517 59 551 93
rect 603 85 637 119
<< pdiffc >>
rect 44 547 78 581
rect 146 573 180 607
rect 321 555 355 589
rect 508 573 542 607
rect 594 547 628 581
<< poly >>
rect 89 619 119 645
rect 208 619 238 645
rect 280 619 310 645
rect 366 619 396 645
rect 460 619 490 645
rect 553 619 583 645
rect 89 513 119 535
rect 41 483 119 513
rect 208 507 238 535
rect 41 321 71 483
rect 161 477 238 507
rect 161 435 191 477
rect 119 419 191 435
rect 280 429 310 535
rect 366 503 396 535
rect 119 385 135 419
rect 169 385 191 419
rect 119 369 191 385
rect 233 413 310 429
rect 233 379 249 413
rect 283 379 310 413
rect 41 291 110 321
rect 80 263 110 291
rect 155 315 185 369
rect 233 363 310 379
rect 352 487 418 503
rect 352 453 368 487
rect 402 453 418 487
rect 352 419 418 453
rect 352 385 368 419
rect 402 385 418 419
rect 352 369 418 385
rect 280 321 310 363
rect 155 285 196 315
rect 280 291 320 321
rect 166 263 196 285
rect 290 269 320 291
rect 80 144 110 179
rect 166 153 196 179
rect 290 159 320 185
rect 388 183 418 369
rect 460 352 490 535
rect 553 460 583 535
rect 532 444 604 460
rect 532 410 548 444
rect 582 410 604 444
rect 532 394 604 410
rect 460 336 526 352
rect 460 302 476 336
rect 510 302 526 336
rect 460 268 526 302
rect 460 234 476 268
rect 510 234 526 268
rect 460 218 526 234
rect 388 153 420 183
rect 58 128 124 144
rect 390 131 420 153
rect 476 131 506 218
rect 574 176 604 394
rect 562 146 604 176
rect 562 131 592 146
rect 58 94 74 128
rect 108 94 124 128
rect 58 78 124 94
rect 390 21 420 47
rect 476 21 506 47
rect 562 21 592 47
<< polycont >>
rect 135 385 169 419
rect 249 379 283 413
rect 368 453 402 487
rect 368 385 402 419
rect 548 410 582 444
rect 476 302 510 336
rect 476 234 510 268
rect 74 94 108 128
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 130 607 196 649
rect 28 581 94 585
rect 28 547 44 581
rect 78 547 94 581
rect 130 573 146 607
rect 180 573 196 607
rect 508 607 546 649
rect 130 569 196 573
rect 249 589 472 605
rect 28 533 94 547
rect 249 555 321 589
rect 355 555 472 589
rect 542 573 546 607
rect 508 557 546 573
rect 590 581 652 597
rect 249 539 472 555
rect 249 533 283 539
rect 28 499 283 533
rect 28 251 73 499
rect 319 487 402 503
rect 319 453 368 487
rect 119 419 185 424
rect 119 385 135 419
rect 169 385 185 419
rect 223 413 283 429
rect 223 379 249 413
rect 223 363 283 379
rect 319 419 402 453
rect 319 385 368 419
rect 438 460 472 539
rect 590 547 594 581
rect 628 547 652 581
rect 590 531 652 547
rect 438 444 582 460
rect 438 410 548 444
rect 438 394 582 410
rect 319 369 402 385
rect 460 336 555 352
rect 618 350 652 531
rect 460 302 476 336
rect 510 302 555 336
rect 28 217 35 251
rect 69 217 73 251
rect 28 201 73 217
rect 117 265 369 299
rect 117 251 159 265
rect 117 217 121 251
rect 155 217 159 251
rect 327 257 369 265
rect 117 201 159 217
rect 210 225 276 229
rect 210 191 226 225
rect 260 191 276 225
rect 327 223 331 257
rect 365 223 369 257
rect 327 207 369 223
rect 460 268 555 302
rect 460 234 476 268
rect 510 234 555 268
rect 460 218 555 234
rect 210 167 276 191
rect 21 128 171 144
rect 210 133 469 167
rect 21 94 74 128
rect 108 94 171 128
rect 427 119 469 133
rect 21 78 171 94
rect 325 93 391 97
rect 325 59 341 93
rect 375 59 391 93
rect 427 85 431 119
rect 465 85 469 119
rect 599 119 652 350
rect 427 69 469 85
rect 513 93 555 109
rect 325 17 391 59
rect 513 59 517 93
rect 551 59 555 93
rect 599 85 603 119
rect 637 85 652 119
rect 599 69 652 85
rect 513 17 555 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221a_m
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4866088
string GDS_START 4858706
<< end >>
