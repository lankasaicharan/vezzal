magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 318 161 863 241
rect 1 49 863 161
rect 0 0 864 49
<< scnmos >>
rect 80 51 110 135
rect 166 51 196 135
rect 397 131 427 215
rect 469 131 499 215
rect 577 131 607 215
rect 649 131 679 215
rect 754 47 784 215
<< scpmoshvt >>
rect 100 531 130 615
rect 186 531 216 615
rect 383 393 413 477
rect 469 393 499 477
rect 563 393 593 477
rect 649 393 679 477
rect 754 367 784 619
<< ndiff >>
rect 344 181 397 215
rect 344 147 352 181
rect 386 147 397 181
rect 27 107 80 135
rect 27 73 35 107
rect 69 73 80 107
rect 27 51 80 73
rect 110 107 166 135
rect 110 73 121 107
rect 155 73 166 107
rect 110 51 166 73
rect 196 107 249 135
rect 344 131 397 147
rect 427 131 469 215
rect 499 131 577 215
rect 607 131 649 215
rect 679 203 754 215
rect 679 169 697 203
rect 731 169 754 203
rect 679 131 754 169
rect 196 73 207 107
rect 241 73 249 107
rect 196 51 249 73
rect 701 93 754 131
rect 701 59 709 93
rect 743 59 754 93
rect 701 47 754 59
rect 784 203 837 215
rect 784 169 795 203
rect 829 169 837 203
rect 784 101 837 169
rect 784 67 795 101
rect 829 67 837 101
rect 784 47 837 67
<< pdiff >>
rect 47 590 100 615
rect 47 556 55 590
rect 89 556 100 590
rect 47 531 100 556
rect 130 590 186 615
rect 130 556 141 590
rect 175 556 186 590
rect 130 531 186 556
rect 216 590 269 615
rect 216 556 227 590
rect 261 556 269 590
rect 216 531 269 556
rect 701 607 754 619
rect 701 573 709 607
rect 743 573 754 607
rect 701 539 754 573
rect 701 505 709 539
rect 743 505 754 539
rect 701 477 754 505
rect 330 463 383 477
rect 330 429 338 463
rect 372 429 383 463
rect 330 393 383 429
rect 413 452 469 477
rect 413 418 424 452
rect 458 418 469 452
rect 413 393 469 418
rect 499 452 563 477
rect 499 418 513 452
rect 547 418 563 452
rect 499 393 563 418
rect 593 452 649 477
rect 593 418 604 452
rect 638 418 649 452
rect 593 393 649 418
rect 679 459 754 477
rect 679 425 690 459
rect 724 425 754 459
rect 679 393 754 425
rect 701 367 754 393
rect 784 599 837 619
rect 784 565 795 599
rect 829 565 837 599
rect 784 529 837 565
rect 784 495 795 529
rect 829 495 837 529
rect 784 457 837 495
rect 784 423 795 457
rect 829 423 837 457
rect 784 367 837 423
<< ndiffc >>
rect 352 147 386 181
rect 35 73 69 107
rect 121 73 155 107
rect 697 169 731 203
rect 207 73 241 107
rect 709 59 743 93
rect 795 169 829 203
rect 795 67 829 101
<< pdiffc >>
rect 55 556 89 590
rect 141 556 175 590
rect 227 556 261 590
rect 709 573 743 607
rect 709 505 743 539
rect 338 429 372 463
rect 424 418 458 452
rect 513 418 547 452
rect 604 418 638 452
rect 690 425 724 459
rect 795 565 829 599
rect 795 495 829 529
rect 795 423 829 457
<< poly >>
rect 100 615 130 641
rect 186 615 216 641
rect 754 619 784 645
rect 603 601 679 617
rect 603 567 619 601
rect 653 567 679 601
rect 603 551 679 567
rect 100 498 130 531
rect 100 468 138 498
rect 72 452 138 468
rect 72 418 88 452
rect 122 418 138 452
rect 72 384 138 418
rect 186 415 216 531
rect 383 477 413 503
rect 469 477 499 503
rect 563 477 593 503
rect 649 477 679 551
rect 72 350 88 384
rect 122 350 138 384
rect 72 334 138 350
rect 180 385 216 415
rect 80 135 110 334
rect 180 223 210 385
rect 252 321 318 337
rect 252 287 268 321
rect 302 301 318 321
rect 383 301 413 393
rect 302 287 427 301
rect 252 271 427 287
rect 166 207 232 223
rect 397 215 427 271
rect 469 215 499 393
rect 563 303 593 393
rect 541 287 607 303
rect 541 253 557 287
rect 591 253 607 287
rect 541 237 607 253
rect 577 215 607 237
rect 649 215 679 393
rect 754 335 784 367
rect 721 319 787 335
rect 721 285 737 319
rect 771 285 787 319
rect 721 269 787 285
rect 754 215 784 269
rect 166 173 182 207
rect 216 173 232 207
rect 166 157 232 173
rect 166 135 196 157
rect 397 105 427 131
rect 469 109 499 131
rect 469 93 535 109
rect 577 105 607 131
rect 649 105 679 131
rect 469 59 485 93
rect 519 59 535 93
rect 80 25 110 51
rect 166 25 196 51
rect 469 43 535 59
rect 754 21 784 47
<< polycont >>
rect 619 567 653 601
rect 88 418 122 452
rect 88 350 122 384
rect 268 287 302 321
rect 557 253 591 287
rect 737 285 771 319
rect 182 173 216 207
rect 485 59 519 93
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 18 590 91 606
rect 18 556 55 590
rect 89 556 91 590
rect 18 540 91 556
rect 125 590 191 649
rect 125 556 141 590
rect 175 556 191 590
rect 125 540 191 556
rect 225 590 277 606
rect 225 556 227 590
rect 261 556 277 590
rect 18 300 52 540
rect 88 452 176 506
rect 122 418 176 452
rect 88 384 176 418
rect 122 357 176 384
rect 225 391 277 556
rect 322 463 388 649
rect 322 429 338 463
rect 372 429 388 463
rect 322 425 388 429
rect 422 452 463 468
rect 422 418 424 452
rect 458 418 463 452
rect 225 357 388 391
rect 122 350 138 357
rect 88 334 138 350
rect 185 321 318 323
rect 185 300 268 321
rect 18 287 268 300
rect 302 287 318 321
rect 18 285 318 287
rect 18 266 219 285
rect 18 107 78 266
rect 354 251 388 357
rect 112 207 216 223
rect 112 173 182 207
rect 112 157 216 173
rect 266 217 388 251
rect 422 375 463 418
rect 497 452 563 649
rect 597 601 669 615
rect 597 567 619 601
rect 653 567 669 601
rect 597 525 669 567
rect 703 607 751 649
rect 703 573 709 607
rect 743 573 751 607
rect 703 539 751 573
rect 703 505 709 539
rect 743 505 751 539
rect 703 475 751 505
rect 497 418 513 452
rect 547 418 563 452
rect 497 409 563 418
rect 597 452 648 468
rect 597 418 604 452
rect 638 418 648 452
rect 597 375 648 418
rect 682 459 751 475
rect 682 425 690 459
rect 724 425 751 459
rect 682 409 751 425
rect 785 599 847 615
rect 785 565 795 599
rect 829 565 847 599
rect 785 529 847 565
rect 785 495 795 529
rect 829 495 847 529
rect 785 457 847 495
rect 785 423 795 457
rect 829 423 847 457
rect 785 407 847 423
rect 422 341 771 375
rect 266 123 300 217
rect 422 183 462 341
rect 721 319 771 341
rect 336 181 462 183
rect 336 147 352 181
rect 386 147 462 181
rect 511 287 653 303
rect 511 253 557 287
rect 591 253 653 287
rect 721 285 737 319
rect 721 269 771 285
rect 511 150 653 253
rect 805 219 847 407
rect 687 203 751 219
rect 687 169 697 203
rect 731 169 751 203
rect 336 135 462 147
rect 18 73 35 107
rect 69 73 78 107
rect 18 57 78 73
rect 112 107 164 123
rect 112 73 121 107
rect 155 73 164 107
rect 112 17 164 73
rect 198 107 300 123
rect 198 73 207 107
rect 241 101 300 107
rect 241 93 535 101
rect 241 73 485 93
rect 198 59 485 73
rect 519 59 535 93
rect 198 51 535 59
rect 687 93 751 169
rect 687 59 709 93
rect 743 59 751 93
rect 687 17 751 59
rect 785 203 847 219
rect 785 169 795 203
rect 829 169 847 203
rect 785 101 847 169
rect 785 67 795 101
rect 829 67 847 101
rect 785 51 847 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4bb_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5234594
string GDS_START 5226482
<< end >>
