magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 75 49 707 241
rect 0 0 768 49
<< scnmos >>
rect 154 47 184 215
rect 244 47 274 215
rect 330 47 360 215
rect 426 47 456 215
rect 512 47 542 215
rect 598 47 628 215
<< scpmoshvt >>
rect 89 367 119 619
rect 244 367 274 619
rect 330 367 360 619
rect 426 367 456 619
rect 512 367 542 619
rect 658 367 688 619
<< ndiff >>
rect 101 203 154 215
rect 101 169 109 203
rect 143 169 154 203
rect 101 93 154 169
rect 101 59 109 93
rect 143 59 154 93
rect 101 47 154 59
rect 184 186 244 215
rect 184 152 195 186
rect 229 152 244 186
rect 184 101 244 152
rect 184 67 195 101
rect 229 67 244 101
rect 184 47 244 67
rect 274 126 330 215
rect 274 92 285 126
rect 319 92 330 126
rect 274 47 330 92
rect 360 202 426 215
rect 360 168 376 202
rect 410 168 426 202
rect 360 101 426 168
rect 360 67 376 101
rect 410 67 426 101
rect 360 47 426 67
rect 456 126 512 215
rect 456 92 467 126
rect 501 92 512 126
rect 456 47 512 92
rect 542 186 598 215
rect 542 152 553 186
rect 587 152 598 186
rect 542 101 598 152
rect 542 67 553 101
rect 587 67 598 101
rect 542 47 598 67
rect 628 203 681 215
rect 628 169 639 203
rect 673 169 681 203
rect 628 93 681 169
rect 628 59 639 93
rect 673 59 681 93
rect 628 47 681 59
<< pdiff >>
rect 36 599 89 619
rect 36 565 44 599
rect 78 565 89 599
rect 36 510 89 565
rect 36 476 44 510
rect 78 476 89 510
rect 36 413 89 476
rect 36 379 44 413
rect 78 379 89 413
rect 36 367 89 379
rect 119 607 244 619
rect 119 573 130 607
rect 164 573 199 607
rect 233 573 244 607
rect 119 529 244 573
rect 119 495 130 529
rect 164 495 244 529
rect 119 455 244 495
rect 119 421 130 455
rect 164 421 244 455
rect 119 367 244 421
rect 274 599 330 619
rect 274 565 285 599
rect 319 565 330 599
rect 274 527 330 565
rect 274 493 285 527
rect 319 493 330 527
rect 274 367 330 493
rect 360 607 426 619
rect 360 573 371 607
rect 405 573 426 607
rect 360 367 426 573
rect 456 443 512 619
rect 456 409 467 443
rect 501 409 512 443
rect 456 367 512 409
rect 542 605 658 619
rect 542 571 553 605
rect 587 571 658 605
rect 542 509 658 571
rect 542 475 613 509
rect 647 475 658 509
rect 542 367 658 475
rect 688 599 741 619
rect 688 565 699 599
rect 733 565 741 599
rect 688 516 741 565
rect 688 482 699 516
rect 733 482 741 516
rect 688 425 741 482
rect 688 391 699 425
rect 733 391 741 425
rect 688 367 741 391
<< ndiffc >>
rect 109 169 143 203
rect 109 59 143 93
rect 195 152 229 186
rect 195 67 229 101
rect 285 92 319 126
rect 376 168 410 202
rect 376 67 410 101
rect 467 92 501 126
rect 553 152 587 186
rect 553 67 587 101
rect 639 169 673 203
rect 639 59 673 93
<< pdiffc >>
rect 44 565 78 599
rect 44 476 78 510
rect 44 379 78 413
rect 130 573 164 607
rect 199 573 233 607
rect 130 495 164 529
rect 130 421 164 455
rect 285 565 319 599
rect 285 493 319 527
rect 371 573 405 607
rect 467 409 501 443
rect 553 571 587 605
rect 613 475 647 509
rect 699 565 733 599
rect 699 482 733 516
rect 699 391 733 425
<< poly >>
rect 89 619 119 645
rect 244 619 274 645
rect 330 619 360 645
rect 426 619 456 645
rect 512 619 542 645
rect 658 619 688 645
rect 89 303 119 367
rect 244 303 274 367
rect 330 335 360 367
rect 426 345 456 367
rect 512 345 542 367
rect 89 287 274 303
rect 89 253 127 287
rect 161 253 198 287
rect 232 253 274 287
rect 316 319 384 335
rect 316 285 334 319
rect 368 285 384 319
rect 316 269 384 285
rect 426 287 542 345
rect 658 323 688 367
rect 89 237 274 253
rect 154 215 184 237
rect 244 215 274 237
rect 330 215 360 269
rect 426 253 461 287
rect 495 253 542 287
rect 426 237 542 253
rect 426 215 456 237
rect 512 215 542 237
rect 598 307 747 323
rect 598 273 614 307
rect 648 273 697 307
rect 731 273 747 307
rect 598 237 747 273
rect 598 215 628 237
rect 154 21 184 47
rect 244 21 274 47
rect 330 21 360 47
rect 426 21 456 47
rect 512 21 542 47
rect 598 21 628 47
<< polycont >>
rect 127 253 161 287
rect 198 253 232 287
rect 334 285 368 319
rect 461 253 495 287
rect 614 273 648 307
rect 697 273 731 307
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 28 599 82 615
rect 28 565 44 599
rect 78 565 82 599
rect 28 510 82 565
rect 28 476 44 510
rect 78 476 82 510
rect 28 413 82 476
rect 28 379 44 413
rect 78 379 82 413
rect 116 607 249 649
rect 116 573 130 607
rect 164 573 199 607
rect 233 573 249 607
rect 116 563 249 573
rect 283 599 321 615
rect 283 565 285 599
rect 319 565 321 599
rect 116 529 164 563
rect 283 529 321 565
rect 355 607 663 615
rect 355 573 371 607
rect 405 605 663 607
rect 405 573 553 605
rect 355 571 553 573
rect 587 571 663 605
rect 355 563 663 571
rect 116 495 130 529
rect 116 455 164 495
rect 116 421 130 455
rect 116 405 164 421
rect 198 527 569 529
rect 198 493 285 527
rect 319 493 569 527
rect 28 371 82 379
rect 198 371 232 493
rect 28 337 232 371
rect 266 443 501 459
rect 266 409 467 443
rect 266 393 501 409
rect 535 425 569 493
rect 603 509 663 563
rect 603 475 613 509
rect 647 475 663 509
rect 603 459 663 475
rect 697 599 749 615
rect 697 565 699 599
rect 733 565 749 599
rect 697 516 749 565
rect 697 482 699 516
rect 733 482 749 516
rect 697 425 749 482
rect 31 287 232 303
rect 31 253 127 287
rect 161 253 198 287
rect 31 237 232 253
rect 266 208 300 393
rect 535 391 699 425
rect 733 391 749 425
rect 334 321 749 357
rect 334 319 374 321
rect 368 285 374 319
rect 588 307 749 321
rect 334 269 374 285
rect 408 253 461 287
rect 495 253 552 287
rect 588 273 614 307
rect 648 273 697 307
rect 731 273 749 307
rect 588 257 749 273
rect 408 242 552 253
rect 266 203 596 208
rect 93 169 109 203
rect 143 169 159 203
rect 93 93 159 169
rect 93 59 109 93
rect 143 59 159 93
rect 93 17 159 59
rect 193 202 596 203
rect 193 186 376 202
rect 193 152 195 186
rect 229 168 376 186
rect 410 186 596 202
rect 410 168 553 186
rect 229 152 235 168
rect 193 101 235 152
rect 193 67 195 101
rect 229 67 235 101
rect 193 51 235 67
rect 269 126 335 134
rect 269 92 285 126
rect 319 92 335 126
rect 269 17 335 92
rect 369 101 417 168
rect 551 152 553 168
rect 587 152 596 186
rect 369 67 376 101
rect 410 67 417 101
rect 369 51 417 67
rect 451 126 517 134
rect 451 92 467 126
rect 501 92 517 126
rect 451 17 517 92
rect 551 101 596 152
rect 551 67 553 101
rect 587 67 596 101
rect 551 51 596 67
rect 630 203 689 219
rect 630 169 639 203
rect 673 169 689 203
rect 630 93 689 169
rect 630 59 639 93
rect 673 59 689 93
rect 630 17 689 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor3_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2639272
string GDS_START 2632062
<< end >>
