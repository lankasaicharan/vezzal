magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3794 1975
<< nwell >>
rect -38 331 2534 704
<< pwell >>
rect 1 49 2319 183
rect 0 0 2496 49
<< scnmos >>
rect 80 47 110 157
rect 152 47 182 157
rect 238 47 268 157
rect 310 47 340 157
rect 396 47 426 157
rect 468 47 498 157
rect 554 47 584 157
rect 626 47 656 157
rect 716 47 746 157
rect 788 47 818 157
rect 874 47 904 157
rect 946 47 976 157
rect 1032 47 1062 157
rect 1104 47 1134 157
rect 1190 47 1220 157
rect 1262 47 1292 157
rect 1348 47 1378 157
rect 1420 47 1450 157
rect 1506 47 1536 157
rect 1578 47 1608 157
rect 1664 47 1694 157
rect 1736 47 1766 157
rect 1822 47 1852 157
rect 1894 47 1924 157
rect 1980 47 2010 157
rect 2052 47 2082 157
rect 2138 47 2168 157
rect 2210 47 2240 157
<< scpmoshvt >>
rect 80 417 130 617
rect 186 417 236 617
rect 292 417 342 617
rect 398 417 448 617
rect 504 417 554 617
rect 610 417 660 617
rect 716 417 766 617
rect 822 417 872 617
rect 928 417 978 617
rect 1034 417 1084 617
rect 1140 417 1190 617
rect 1246 417 1296 617
rect 1352 417 1402 617
rect 1458 417 1508 617
rect 1564 417 1614 617
rect 1670 417 1720 617
rect 1776 417 1826 617
rect 1882 417 1932 617
rect 1988 417 2038 617
rect 2094 417 2144 617
rect 2200 417 2250 617
rect 2306 417 2356 617
<< ndiff >>
rect 27 105 80 157
rect 27 71 35 105
rect 69 71 80 105
rect 27 47 80 71
rect 110 47 152 157
rect 182 105 238 157
rect 182 71 193 105
rect 227 71 238 105
rect 182 47 238 71
rect 268 47 310 157
rect 340 105 396 157
rect 340 71 351 105
rect 385 71 396 105
rect 340 47 396 71
rect 426 47 468 157
rect 498 105 554 157
rect 498 71 509 105
rect 543 71 554 105
rect 498 47 554 71
rect 584 47 626 157
rect 656 105 716 157
rect 656 71 667 105
rect 701 71 716 105
rect 656 47 716 71
rect 746 47 788 157
rect 818 105 874 157
rect 818 71 829 105
rect 863 71 874 105
rect 818 47 874 71
rect 904 47 946 157
rect 976 105 1032 157
rect 976 71 987 105
rect 1021 71 1032 105
rect 976 47 1032 71
rect 1062 47 1104 157
rect 1134 105 1190 157
rect 1134 71 1145 105
rect 1179 71 1190 105
rect 1134 47 1190 71
rect 1220 47 1262 157
rect 1292 105 1348 157
rect 1292 71 1303 105
rect 1337 71 1348 105
rect 1292 47 1348 71
rect 1378 47 1420 157
rect 1450 105 1506 157
rect 1450 71 1461 105
rect 1495 71 1506 105
rect 1450 47 1506 71
rect 1536 47 1578 157
rect 1608 105 1664 157
rect 1608 71 1619 105
rect 1653 71 1664 105
rect 1608 47 1664 71
rect 1694 47 1736 157
rect 1766 105 1822 157
rect 1766 71 1777 105
rect 1811 71 1822 105
rect 1766 47 1822 71
rect 1852 47 1894 157
rect 1924 105 1980 157
rect 1924 71 1935 105
rect 1969 71 1980 105
rect 1924 47 1980 71
rect 2010 47 2052 157
rect 2082 105 2138 157
rect 2082 71 2093 105
rect 2127 71 2138 105
rect 2082 47 2138 71
rect 2168 47 2210 157
rect 2240 105 2293 157
rect 2240 71 2251 105
rect 2285 71 2293 105
rect 2240 47 2293 71
<< pdiff >>
rect 27 599 80 617
rect 27 565 35 599
rect 69 565 80 599
rect 27 531 80 565
rect 27 497 35 531
rect 69 497 80 531
rect 27 463 80 497
rect 27 429 35 463
rect 69 429 80 463
rect 27 417 80 429
rect 130 599 186 617
rect 130 565 141 599
rect 175 565 186 599
rect 130 531 186 565
rect 130 497 141 531
rect 175 497 186 531
rect 130 463 186 497
rect 130 429 141 463
rect 175 429 186 463
rect 130 417 186 429
rect 236 599 292 617
rect 236 565 247 599
rect 281 565 292 599
rect 236 531 292 565
rect 236 497 247 531
rect 281 497 292 531
rect 236 463 292 497
rect 236 429 247 463
rect 281 429 292 463
rect 236 417 292 429
rect 342 599 398 617
rect 342 565 353 599
rect 387 565 398 599
rect 342 531 398 565
rect 342 497 353 531
rect 387 497 398 531
rect 342 463 398 497
rect 342 429 353 463
rect 387 429 398 463
rect 342 417 398 429
rect 448 599 504 617
rect 448 565 459 599
rect 493 565 504 599
rect 448 531 504 565
rect 448 497 459 531
rect 493 497 504 531
rect 448 463 504 497
rect 448 429 459 463
rect 493 429 504 463
rect 448 417 504 429
rect 554 599 610 617
rect 554 565 565 599
rect 599 565 610 599
rect 554 531 610 565
rect 554 497 565 531
rect 599 497 610 531
rect 554 463 610 497
rect 554 429 565 463
rect 599 429 610 463
rect 554 417 610 429
rect 660 599 716 617
rect 660 565 671 599
rect 705 565 716 599
rect 660 531 716 565
rect 660 497 671 531
rect 705 497 716 531
rect 660 463 716 497
rect 660 429 671 463
rect 705 429 716 463
rect 660 417 716 429
rect 766 599 822 617
rect 766 565 777 599
rect 811 565 822 599
rect 766 531 822 565
rect 766 497 777 531
rect 811 497 822 531
rect 766 463 822 497
rect 766 429 777 463
rect 811 429 822 463
rect 766 417 822 429
rect 872 599 928 617
rect 872 565 883 599
rect 917 565 928 599
rect 872 531 928 565
rect 872 497 883 531
rect 917 497 928 531
rect 872 463 928 497
rect 872 429 883 463
rect 917 429 928 463
rect 872 417 928 429
rect 978 599 1034 617
rect 978 565 989 599
rect 1023 565 1034 599
rect 978 531 1034 565
rect 978 497 989 531
rect 1023 497 1034 531
rect 978 463 1034 497
rect 978 429 989 463
rect 1023 429 1034 463
rect 978 417 1034 429
rect 1084 599 1140 617
rect 1084 565 1095 599
rect 1129 565 1140 599
rect 1084 531 1140 565
rect 1084 497 1095 531
rect 1129 497 1140 531
rect 1084 463 1140 497
rect 1084 429 1095 463
rect 1129 429 1140 463
rect 1084 417 1140 429
rect 1190 599 1246 617
rect 1190 565 1201 599
rect 1235 565 1246 599
rect 1190 531 1246 565
rect 1190 497 1201 531
rect 1235 497 1246 531
rect 1190 463 1246 497
rect 1190 429 1201 463
rect 1235 429 1246 463
rect 1190 417 1246 429
rect 1296 599 1352 617
rect 1296 565 1307 599
rect 1341 565 1352 599
rect 1296 531 1352 565
rect 1296 497 1307 531
rect 1341 497 1352 531
rect 1296 463 1352 497
rect 1296 429 1307 463
rect 1341 429 1352 463
rect 1296 417 1352 429
rect 1402 599 1458 617
rect 1402 565 1413 599
rect 1447 565 1458 599
rect 1402 531 1458 565
rect 1402 497 1413 531
rect 1447 497 1458 531
rect 1402 463 1458 497
rect 1402 429 1413 463
rect 1447 429 1458 463
rect 1402 417 1458 429
rect 1508 599 1564 617
rect 1508 565 1519 599
rect 1553 565 1564 599
rect 1508 531 1564 565
rect 1508 497 1519 531
rect 1553 497 1564 531
rect 1508 463 1564 497
rect 1508 429 1519 463
rect 1553 429 1564 463
rect 1508 417 1564 429
rect 1614 599 1670 617
rect 1614 565 1625 599
rect 1659 565 1670 599
rect 1614 531 1670 565
rect 1614 497 1625 531
rect 1659 497 1670 531
rect 1614 463 1670 497
rect 1614 429 1625 463
rect 1659 429 1670 463
rect 1614 417 1670 429
rect 1720 599 1776 617
rect 1720 565 1731 599
rect 1765 565 1776 599
rect 1720 531 1776 565
rect 1720 497 1731 531
rect 1765 497 1776 531
rect 1720 463 1776 497
rect 1720 429 1731 463
rect 1765 429 1776 463
rect 1720 417 1776 429
rect 1826 599 1882 617
rect 1826 565 1837 599
rect 1871 565 1882 599
rect 1826 531 1882 565
rect 1826 497 1837 531
rect 1871 497 1882 531
rect 1826 463 1882 497
rect 1826 429 1837 463
rect 1871 429 1882 463
rect 1826 417 1882 429
rect 1932 599 1988 617
rect 1932 565 1943 599
rect 1977 565 1988 599
rect 1932 531 1988 565
rect 1932 497 1943 531
rect 1977 497 1988 531
rect 1932 463 1988 497
rect 1932 429 1943 463
rect 1977 429 1988 463
rect 1932 417 1988 429
rect 2038 599 2094 617
rect 2038 565 2049 599
rect 2083 565 2094 599
rect 2038 531 2094 565
rect 2038 497 2049 531
rect 2083 497 2094 531
rect 2038 463 2094 497
rect 2038 429 2049 463
rect 2083 429 2094 463
rect 2038 417 2094 429
rect 2144 599 2200 617
rect 2144 565 2155 599
rect 2189 565 2200 599
rect 2144 531 2200 565
rect 2144 497 2155 531
rect 2189 497 2200 531
rect 2144 463 2200 497
rect 2144 429 2155 463
rect 2189 429 2200 463
rect 2144 417 2200 429
rect 2250 599 2306 617
rect 2250 565 2261 599
rect 2295 565 2306 599
rect 2250 531 2306 565
rect 2250 497 2261 531
rect 2295 497 2306 531
rect 2250 463 2306 497
rect 2250 429 2261 463
rect 2295 429 2306 463
rect 2250 417 2306 429
rect 2356 599 2409 617
rect 2356 565 2367 599
rect 2401 565 2409 599
rect 2356 531 2409 565
rect 2356 497 2367 531
rect 2401 497 2409 531
rect 2356 463 2409 497
rect 2356 429 2367 463
rect 2401 429 2409 463
rect 2356 417 2409 429
<< ndiffc >>
rect 35 71 69 105
rect 193 71 227 105
rect 351 71 385 105
rect 509 71 543 105
rect 667 71 701 105
rect 829 71 863 105
rect 987 71 1021 105
rect 1145 71 1179 105
rect 1303 71 1337 105
rect 1461 71 1495 105
rect 1619 71 1653 105
rect 1777 71 1811 105
rect 1935 71 1969 105
rect 2093 71 2127 105
rect 2251 71 2285 105
<< pdiffc >>
rect 35 565 69 599
rect 35 497 69 531
rect 35 429 69 463
rect 141 565 175 599
rect 141 497 175 531
rect 141 429 175 463
rect 247 565 281 599
rect 247 497 281 531
rect 247 429 281 463
rect 353 565 387 599
rect 353 497 387 531
rect 353 429 387 463
rect 459 565 493 599
rect 459 497 493 531
rect 459 429 493 463
rect 565 565 599 599
rect 565 497 599 531
rect 565 429 599 463
rect 671 565 705 599
rect 671 497 705 531
rect 671 429 705 463
rect 777 565 811 599
rect 777 497 811 531
rect 777 429 811 463
rect 883 565 917 599
rect 883 497 917 531
rect 883 429 917 463
rect 989 565 1023 599
rect 989 497 1023 531
rect 989 429 1023 463
rect 1095 565 1129 599
rect 1095 497 1129 531
rect 1095 429 1129 463
rect 1201 565 1235 599
rect 1201 497 1235 531
rect 1201 429 1235 463
rect 1307 565 1341 599
rect 1307 497 1341 531
rect 1307 429 1341 463
rect 1413 565 1447 599
rect 1413 497 1447 531
rect 1413 429 1447 463
rect 1519 565 1553 599
rect 1519 497 1553 531
rect 1519 429 1553 463
rect 1625 565 1659 599
rect 1625 497 1659 531
rect 1625 429 1659 463
rect 1731 565 1765 599
rect 1731 497 1765 531
rect 1731 429 1765 463
rect 1837 565 1871 599
rect 1837 497 1871 531
rect 1837 429 1871 463
rect 1943 565 1977 599
rect 1943 497 1977 531
rect 1943 429 1977 463
rect 2049 565 2083 599
rect 2049 497 2083 531
rect 2049 429 2083 463
rect 2155 565 2189 599
rect 2155 497 2189 531
rect 2155 429 2189 463
rect 2261 565 2295 599
rect 2261 497 2295 531
rect 2261 429 2295 463
rect 2367 565 2401 599
rect 2367 497 2401 531
rect 2367 429 2401 463
<< poly >>
rect 80 617 130 645
rect 186 617 236 645
rect 292 617 342 645
rect 398 617 448 645
rect 504 617 554 645
rect 610 617 660 645
rect 716 617 766 645
rect 822 617 872 645
rect 928 617 978 645
rect 1034 617 1084 645
rect 1140 617 1190 645
rect 1246 617 1296 645
rect 1352 617 1402 645
rect 1458 617 1508 645
rect 1564 617 1614 645
rect 1670 617 1720 645
rect 1776 617 1826 645
rect 1882 617 1932 645
rect 1988 617 2038 645
rect 2094 617 2144 645
rect 2200 617 2250 645
rect 2306 617 2356 645
rect 80 313 130 417
rect 186 313 236 417
rect 292 313 342 417
rect 398 313 448 417
rect 504 313 554 417
rect 610 313 660 417
rect 80 297 660 313
rect 80 263 96 297
rect 130 263 660 297
rect 80 229 660 263
rect 80 195 96 229
rect 130 195 660 229
rect 80 179 660 195
rect 716 309 766 417
rect 822 309 872 417
rect 928 309 978 417
rect 1034 309 1084 417
rect 1140 309 1190 417
rect 1246 309 1296 417
rect 1352 309 1402 417
rect 1458 309 1508 417
rect 1564 309 1614 417
rect 1670 309 1720 417
rect 1776 309 1826 417
rect 1882 309 1932 417
rect 1988 309 2038 417
rect 2094 309 2144 417
rect 2200 309 2250 417
rect 2306 309 2356 417
rect 716 291 2384 309
rect 716 257 732 291
rect 766 257 933 291
rect 967 257 1028 291
rect 1062 257 1310 291
rect 1344 257 1566 291
rect 1600 257 1661 291
rect 1695 257 1946 291
rect 1980 257 2198 291
rect 2232 257 2266 291
rect 2300 257 2334 291
rect 2368 257 2384 291
rect 716 241 2384 257
rect 80 157 110 179
rect 152 157 182 179
rect 238 157 268 179
rect 310 157 340 179
rect 396 157 426 179
rect 468 157 498 179
rect 554 157 584 179
rect 626 157 656 179
rect 716 157 746 241
rect 788 157 818 241
rect 874 157 904 241
rect 946 157 976 241
rect 1032 157 1062 241
rect 1104 157 1134 241
rect 1190 157 1220 241
rect 1262 157 1292 241
rect 1348 157 1378 241
rect 1420 157 1450 241
rect 1506 157 1536 241
rect 1578 157 1608 241
rect 1664 157 1694 241
rect 1736 157 1766 241
rect 1822 157 1852 241
rect 1894 157 1924 241
rect 1980 157 2010 241
rect 2052 157 2082 241
rect 2138 157 2168 241
rect 2210 157 2240 241
rect 80 21 110 47
rect 152 21 182 47
rect 238 21 268 47
rect 310 21 340 47
rect 396 21 426 47
rect 468 21 498 47
rect 554 21 584 47
rect 626 21 656 47
rect 716 21 746 47
rect 788 21 818 47
rect 874 21 904 47
rect 946 21 976 47
rect 1032 21 1062 47
rect 1104 21 1134 47
rect 1190 21 1220 47
rect 1262 21 1292 47
rect 1348 21 1378 47
rect 1420 21 1450 47
rect 1506 21 1536 47
rect 1578 21 1608 47
rect 1664 21 1694 47
rect 1736 21 1766 47
rect 1822 21 1852 47
rect 1894 21 1924 47
rect 1980 21 2010 47
rect 2052 21 2082 47
rect 2138 21 2168 47
rect 2210 21 2240 47
<< polycont >>
rect 96 263 130 297
rect 96 195 130 229
rect 732 257 766 291
rect 933 257 967 291
rect 1028 257 1062 291
rect 1310 257 1344 291
rect 1566 257 1600 291
rect 1661 257 1695 291
rect 1946 257 1980 291
rect 2198 257 2232 291
rect 2266 257 2300 291
rect 2334 257 2368 291
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 19 599 85 649
rect 19 565 35 599
rect 69 565 85 599
rect 19 531 85 565
rect 19 497 35 531
rect 69 497 85 531
rect 19 463 85 497
rect 19 429 35 463
rect 69 429 85 463
rect 19 413 85 429
rect 119 599 211 615
rect 119 565 141 599
rect 175 565 211 599
rect 119 531 211 565
rect 119 497 141 531
rect 175 497 211 531
rect 119 463 211 497
rect 119 429 141 463
rect 175 429 211 463
rect 119 403 211 429
rect 245 599 297 649
rect 245 565 247 599
rect 281 565 297 599
rect 245 531 297 565
rect 245 497 247 531
rect 281 497 297 531
rect 245 463 297 497
rect 245 429 247 463
rect 281 429 297 463
rect 245 413 297 429
rect 337 599 403 615
rect 337 565 353 599
rect 387 565 403 599
rect 337 531 403 565
rect 337 497 353 531
rect 387 497 403 531
rect 337 463 403 497
rect 337 429 353 463
rect 387 429 403 463
rect 25 313 74 361
rect 25 297 139 313
rect 25 263 96 297
rect 130 263 139 297
rect 25 229 139 263
rect 25 195 96 229
rect 130 195 139 229
rect 25 155 139 195
rect 177 307 211 403
rect 337 307 403 429
rect 443 599 509 649
rect 443 565 459 599
rect 493 565 509 599
rect 443 531 509 565
rect 443 497 459 531
rect 493 497 509 531
rect 443 463 509 497
rect 443 429 459 463
rect 493 429 509 463
rect 443 417 509 429
rect 549 599 615 615
rect 549 565 565 599
rect 599 565 615 599
rect 549 531 615 565
rect 549 497 565 531
rect 599 497 615 531
rect 549 463 615 497
rect 549 429 565 463
rect 599 429 615 463
rect 549 307 615 429
rect 655 599 721 649
rect 655 565 671 599
rect 705 565 721 599
rect 655 531 721 565
rect 655 497 671 531
rect 705 497 721 531
rect 655 463 721 497
rect 655 429 671 463
rect 705 429 721 463
rect 655 417 721 429
rect 761 599 827 615
rect 761 565 777 599
rect 811 565 827 599
rect 761 531 827 565
rect 761 497 777 531
rect 811 497 827 531
rect 761 463 827 497
rect 761 429 777 463
rect 811 429 827 463
rect 761 424 827 429
rect 761 390 777 424
rect 811 390 827 424
rect 867 599 933 649
rect 867 565 883 599
rect 917 565 933 599
rect 867 531 933 565
rect 867 497 883 531
rect 917 497 933 531
rect 867 463 933 497
rect 867 429 883 463
rect 917 429 933 463
rect 867 417 933 429
rect 973 599 1039 615
rect 973 565 989 599
rect 1023 565 1039 599
rect 973 531 1039 565
rect 973 497 989 531
rect 1023 497 1039 531
rect 973 463 1039 497
rect 973 429 989 463
rect 1023 429 1039 463
rect 973 424 1039 429
rect 761 375 827 390
rect 973 390 991 424
rect 1025 390 1039 424
rect 1079 599 1145 649
rect 1079 565 1095 599
rect 1129 565 1145 599
rect 1079 531 1145 565
rect 1079 497 1095 531
rect 1129 497 1145 531
rect 1079 463 1145 497
rect 1079 429 1095 463
rect 1129 429 1145 463
rect 1079 417 1145 429
rect 1185 599 1251 615
rect 1185 565 1201 599
rect 1235 565 1251 599
rect 1185 531 1251 565
rect 1185 497 1201 531
rect 1235 497 1251 531
rect 1185 463 1251 497
rect 1185 429 1201 463
rect 1235 429 1251 463
rect 1185 424 1251 429
rect 973 384 1039 390
rect 1185 390 1201 424
rect 1235 390 1251 424
rect 1291 599 1357 649
rect 1291 565 1307 599
rect 1341 565 1357 599
rect 1291 531 1357 565
rect 1291 497 1307 531
rect 1341 497 1357 531
rect 1291 463 1357 497
rect 1291 429 1307 463
rect 1341 429 1357 463
rect 1291 417 1357 429
rect 1397 599 1463 615
rect 1397 565 1413 599
rect 1447 565 1463 599
rect 1397 531 1463 565
rect 1397 497 1413 531
rect 1447 497 1463 531
rect 1397 463 1463 497
rect 1397 429 1413 463
rect 1447 429 1463 463
rect 1397 424 1463 429
rect 761 341 879 375
rect 1185 358 1251 390
rect 177 291 782 307
rect 177 276 732 291
rect 177 242 607 276
rect 641 242 703 276
rect 766 257 782 291
rect 737 242 782 257
rect 177 241 782 242
rect 25 105 85 121
rect 25 71 35 105
rect 69 71 85 105
rect 25 17 85 71
rect 177 105 246 241
rect 490 236 782 241
rect 177 71 193 105
rect 227 71 246 105
rect 177 53 246 71
rect 335 105 401 121
rect 335 71 351 105
rect 385 71 401 105
rect 335 17 401 71
rect 490 105 559 236
rect 816 207 879 341
rect 917 291 1078 302
rect 917 257 933 291
rect 967 276 1028 291
rect 967 257 991 276
rect 917 242 991 257
rect 1025 257 1028 276
rect 1062 257 1078 291
rect 1025 242 1078 257
rect 917 236 1078 242
rect 490 71 509 105
rect 543 71 559 105
rect 490 53 559 71
rect 651 105 717 121
rect 651 71 667 105
rect 701 71 717 105
rect 651 17 717 71
rect 813 105 879 207
rect 1129 234 1251 358
rect 1397 390 1414 424
rect 1448 390 1463 424
rect 1503 599 1569 649
rect 1503 565 1519 599
rect 1553 565 1569 599
rect 1503 531 1569 565
rect 1503 497 1519 531
rect 1553 497 1569 531
rect 1503 463 1569 497
rect 1503 429 1519 463
rect 1553 429 1569 463
rect 1503 417 1569 429
rect 1609 599 1675 615
rect 1609 565 1625 599
rect 1659 565 1675 599
rect 1609 531 1675 565
rect 1609 497 1625 531
rect 1659 497 1675 531
rect 1609 463 1675 497
rect 1609 429 1625 463
rect 1659 429 1675 463
rect 1609 424 1675 429
rect 1397 358 1463 390
rect 1609 390 1626 424
rect 1660 390 1675 424
rect 1715 599 1781 649
rect 1715 565 1731 599
rect 1765 565 1781 599
rect 1715 531 1781 565
rect 1715 497 1731 531
rect 1765 497 1781 531
rect 1715 463 1781 497
rect 1715 429 1731 463
rect 1765 429 1781 463
rect 1715 417 1781 429
rect 1821 599 1887 615
rect 1821 565 1837 599
rect 1871 565 1887 599
rect 1821 531 1887 565
rect 1821 497 1837 531
rect 1871 497 1887 531
rect 1821 463 1887 497
rect 1821 429 1837 463
rect 1871 429 1887 463
rect 1821 424 1887 429
rect 1609 384 1675 390
rect 1821 390 1838 424
rect 1872 390 1887 424
rect 1927 599 1993 649
rect 1927 565 1943 599
rect 1977 565 1993 599
rect 1927 531 1993 565
rect 1927 497 1943 531
rect 1977 497 1993 531
rect 1927 463 1993 497
rect 1927 429 1943 463
rect 1977 429 1993 463
rect 1927 417 1993 429
rect 2033 599 2099 615
rect 2033 565 2049 599
rect 2083 565 2099 599
rect 2033 531 2099 565
rect 2033 497 2049 531
rect 2083 497 2099 531
rect 2033 463 2099 497
rect 2033 429 2049 463
rect 2083 429 2099 463
rect 2033 424 2099 429
rect 1821 358 1887 390
rect 1294 291 1360 302
rect 1294 242 1310 291
rect 1344 242 1360 291
rect 1294 236 1360 242
rect 1397 234 1511 358
rect 1550 291 1711 302
rect 1550 257 1566 291
rect 1600 276 1661 291
rect 1695 276 1711 291
rect 1601 257 1661 276
rect 1550 242 1567 257
rect 1601 242 1663 257
rect 1697 242 1711 276
rect 1550 236 1711 242
rect 813 71 829 105
rect 863 71 879 105
rect 813 53 879 71
rect 971 105 1037 121
rect 971 71 987 105
rect 1021 71 1037 105
rect 971 17 1037 71
rect 1129 105 1195 234
rect 1129 71 1145 105
rect 1179 71 1195 105
rect 1129 53 1195 71
rect 1287 105 1353 121
rect 1287 71 1303 105
rect 1337 71 1353 105
rect 1287 17 1353 71
rect 1445 105 1511 234
rect 1761 234 1887 358
rect 2033 390 2047 424
rect 2081 390 2099 424
rect 2139 599 2205 649
rect 2139 565 2155 599
rect 2189 565 2205 599
rect 2139 531 2205 565
rect 2139 497 2155 531
rect 2189 497 2205 531
rect 2139 463 2205 497
rect 2139 429 2155 463
rect 2189 429 2205 463
rect 2139 417 2205 429
rect 2245 599 2311 615
rect 2245 565 2261 599
rect 2295 565 2311 599
rect 2245 531 2311 565
rect 2245 497 2261 531
rect 2295 497 2311 531
rect 2245 463 2311 497
rect 2245 429 2261 463
rect 2295 429 2311 463
rect 2245 424 2311 429
rect 2033 358 2099 390
rect 2245 390 2261 424
rect 2295 390 2311 424
rect 2351 599 2417 649
rect 2351 565 2367 599
rect 2401 565 2417 599
rect 2351 531 2417 565
rect 2351 497 2367 531
rect 2401 497 2417 531
rect 2351 463 2417 497
rect 2351 429 2367 463
rect 2401 429 2417 463
rect 2351 417 2417 429
rect 2245 384 2311 390
rect 1930 291 1996 302
rect 1930 257 1946 291
rect 1980 276 1996 291
rect 1930 242 1951 257
rect 1985 242 1996 276
rect 1930 236 1996 242
rect 2033 234 2143 358
rect 2182 291 2384 302
rect 2182 257 2198 291
rect 2232 276 2266 291
rect 2232 257 2239 276
rect 2300 257 2334 291
rect 2368 276 2384 291
rect 2182 242 2239 257
rect 2273 242 2335 257
rect 2369 242 2384 276
rect 2182 236 2384 242
rect 1445 71 1461 105
rect 1495 71 1511 105
rect 1445 53 1511 71
rect 1603 105 1669 121
rect 1603 71 1619 105
rect 1653 71 1669 105
rect 1603 17 1669 71
rect 1761 105 1827 234
rect 1761 71 1777 105
rect 1811 71 1827 105
rect 1761 53 1827 71
rect 1919 105 1985 121
rect 1919 71 1935 105
rect 1969 71 1985 105
rect 1919 17 1985 71
rect 2077 105 2143 234
rect 2077 71 2093 105
rect 2127 71 2143 105
rect 2077 53 2143 71
rect 2235 105 2301 121
rect 2235 71 2251 105
rect 2285 71 2301 105
rect 2235 17 2301 71
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 777 390 811 424
rect 991 390 1025 424
rect 1201 390 1235 424
rect 607 242 641 276
rect 703 257 732 276
rect 732 257 737 276
rect 703 242 737 257
rect 991 242 1025 276
rect 1414 390 1448 424
rect 1626 390 1660 424
rect 1838 390 1872 424
rect 1310 257 1344 276
rect 1310 242 1344 257
rect 1567 257 1600 276
rect 1600 257 1601 276
rect 1663 257 1695 276
rect 1695 257 1697 276
rect 1567 242 1601 257
rect 1663 242 1697 257
rect 2047 390 2081 424
rect 2261 390 2295 424
rect 1951 257 1980 276
rect 1980 257 1985 276
rect 1951 242 1985 257
rect 2239 257 2266 276
rect 2266 257 2273 276
rect 2335 257 2368 276
rect 2368 257 2369 276
rect 2239 242 2273 257
rect 2335 242 2369 257
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 683 2496 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 0 617 2496 649
rect 761 424 2311 430
rect 761 390 777 424
rect 811 390 991 424
rect 1025 390 1201 424
rect 1235 390 1414 424
rect 1448 390 1626 424
rect 1660 390 1838 424
rect 1872 390 2047 424
rect 2081 390 2261 424
rect 2295 390 2311 424
rect 761 384 2311 390
rect 595 276 2381 282
rect 595 242 607 276
rect 641 242 703 276
rect 737 242 991 276
rect 1025 242 1310 276
rect 1344 242 1567 276
rect 1601 242 1663 276
rect 1697 242 1951 276
rect 1985 242 2239 276
rect 2273 242 2335 276
rect 2369 242 2381 276
rect 595 236 2381 242
rect 0 17 2496 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
rect 0 -49 2496 -17
<< labels >>
flabel pwell s 0 0 2496 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 2496 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkbuflp_16
flabel metal1 s 761 384 2311 430 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel metal1 s 0 617 2496 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 2496 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2496 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5421446
string GDS_START 5405212
<< end >>
