magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 3 49 671 166
rect 0 0 672 49
<< scnmos >>
rect 86 56 116 140
rect 158 56 188 140
rect 244 56 274 140
rect 322 56 352 140
rect 400 56 430 140
rect 486 56 516 140
rect 558 56 588 140
<< scpmoshvt >>
rect 105 409 155 609
rect 211 409 261 609
rect 317 409 367 609
rect 423 409 473 609
rect 529 409 579 609
<< ndiff >>
rect 29 106 86 140
rect 29 72 41 106
rect 75 72 86 106
rect 29 56 86 72
rect 116 56 158 140
rect 188 115 244 140
rect 188 81 199 115
rect 233 81 244 115
rect 188 56 244 81
rect 274 56 322 140
rect 352 56 400 140
rect 430 115 486 140
rect 430 81 441 115
rect 475 81 486 115
rect 430 56 486 81
rect 516 56 558 140
rect 588 115 645 140
rect 588 81 599 115
rect 633 81 645 115
rect 588 56 645 81
<< pdiff >>
rect 48 597 105 609
rect 48 563 60 597
rect 94 563 105 597
rect 48 526 105 563
rect 48 492 60 526
rect 94 492 105 526
rect 48 455 105 492
rect 48 421 60 455
rect 94 421 105 455
rect 48 409 105 421
rect 155 597 211 609
rect 155 563 166 597
rect 200 563 211 597
rect 155 526 211 563
rect 155 492 166 526
rect 200 492 211 526
rect 155 455 211 492
rect 155 421 166 455
rect 200 421 211 455
rect 155 409 211 421
rect 261 597 317 609
rect 261 563 272 597
rect 306 563 317 597
rect 261 525 317 563
rect 261 491 272 525
rect 306 491 317 525
rect 261 409 317 491
rect 367 597 423 609
rect 367 563 378 597
rect 412 563 423 597
rect 367 526 423 563
rect 367 492 378 526
rect 412 492 423 526
rect 367 455 423 492
rect 367 421 378 455
rect 412 421 423 455
rect 367 409 423 421
rect 473 597 529 609
rect 473 563 484 597
rect 518 563 529 597
rect 473 526 529 563
rect 473 492 484 526
rect 518 492 529 526
rect 473 455 529 492
rect 473 421 484 455
rect 518 421 529 455
rect 473 409 529 421
rect 579 597 636 609
rect 579 563 590 597
rect 624 563 636 597
rect 579 526 636 563
rect 579 492 590 526
rect 624 492 636 526
rect 579 455 636 492
rect 579 421 590 455
rect 624 421 636 455
rect 579 409 636 421
<< ndiffc >>
rect 41 72 75 106
rect 199 81 233 115
rect 441 81 475 115
rect 599 81 633 115
<< pdiffc >>
rect 60 563 94 597
rect 60 492 94 526
rect 60 421 94 455
rect 166 563 200 597
rect 166 492 200 526
rect 166 421 200 455
rect 272 563 306 597
rect 272 491 306 525
rect 378 563 412 597
rect 378 492 412 526
rect 378 421 412 455
rect 484 563 518 597
rect 484 492 518 526
rect 484 421 518 455
rect 590 563 624 597
rect 590 492 624 526
rect 590 421 624 455
<< poly >>
rect 105 609 155 635
rect 211 609 261 635
rect 317 609 367 635
rect 423 609 473 635
rect 529 609 579 635
rect 105 299 155 409
rect 211 299 261 409
rect 317 299 367 409
rect 423 299 473 409
rect 529 369 579 409
rect 521 353 587 369
rect 521 319 537 353
rect 571 319 587 353
rect 86 283 155 299
rect 86 249 105 283
rect 139 249 155 283
rect 86 185 155 249
rect 197 283 263 299
rect 197 249 213 283
rect 247 249 263 283
rect 197 233 263 249
rect 305 283 371 299
rect 305 249 321 283
rect 355 249 371 283
rect 305 233 371 249
rect 413 283 479 299
rect 413 249 429 283
rect 463 249 479 283
rect 413 233 479 249
rect 521 285 587 319
rect 521 251 537 285
rect 571 251 587 285
rect 521 235 587 251
rect 233 185 263 233
rect 86 155 188 185
rect 233 155 274 185
rect 86 140 116 155
rect 158 140 188 155
rect 244 140 274 155
rect 322 140 352 233
rect 413 185 443 233
rect 557 185 587 235
rect 400 155 443 185
rect 486 155 588 185
rect 400 140 430 155
rect 486 140 516 155
rect 558 140 588 155
rect 86 30 116 56
rect 158 30 188 56
rect 244 30 274 56
rect 322 30 352 56
rect 400 30 430 56
rect 486 30 516 56
rect 558 30 588 56
<< polycont >>
rect 537 319 571 353
rect 105 249 139 283
rect 213 249 247 283
rect 321 249 355 283
rect 429 249 463 283
rect 537 251 571 285
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 19 597 110 613
rect 19 563 60 597
rect 94 563 110 597
rect 19 526 110 563
rect 19 492 60 526
rect 94 492 110 526
rect 19 455 110 492
rect 19 421 60 455
rect 94 421 110 455
rect 19 369 110 421
rect 150 597 216 613
rect 150 563 166 597
rect 200 563 216 597
rect 150 526 216 563
rect 150 492 166 526
rect 200 492 216 526
rect 150 455 216 492
rect 256 597 322 649
rect 256 563 272 597
rect 306 563 322 597
rect 256 525 322 563
rect 256 491 272 525
rect 306 491 322 525
rect 256 475 322 491
rect 362 597 428 613
rect 362 563 378 597
rect 412 563 428 597
rect 362 526 428 563
rect 362 492 378 526
rect 412 492 428 526
rect 150 421 166 455
rect 200 439 216 455
rect 362 455 428 492
rect 362 439 378 455
rect 200 421 378 439
rect 412 421 428 455
rect 150 405 428 421
rect 468 597 534 649
rect 468 563 484 597
rect 518 563 534 597
rect 468 526 534 563
rect 468 492 484 526
rect 518 492 534 526
rect 468 455 534 492
rect 468 421 484 455
rect 518 421 534 455
rect 468 405 534 421
rect 574 597 654 613
rect 574 563 590 597
rect 624 563 654 597
rect 574 526 654 563
rect 574 492 590 526
rect 624 492 654 526
rect 574 455 654 492
rect 574 421 590 455
rect 624 421 654 455
rect 574 405 654 421
rect 19 353 584 369
rect 19 335 537 353
rect 19 197 53 335
rect 521 319 537 335
rect 571 319 584 353
rect 89 283 161 299
rect 89 249 105 283
rect 139 249 161 283
rect 89 233 161 249
rect 197 283 263 299
rect 197 249 213 283
rect 247 249 263 283
rect 197 233 263 249
rect 305 283 371 299
rect 305 249 321 283
rect 355 249 371 283
rect 19 163 249 197
rect 25 106 91 127
rect 25 72 41 106
rect 75 72 91 106
rect 25 17 91 72
rect 183 115 249 163
rect 183 81 199 115
rect 233 81 249 115
rect 305 88 371 249
rect 409 283 479 299
rect 409 249 429 283
rect 463 249 479 283
rect 409 233 479 249
rect 521 285 584 319
rect 521 251 537 285
rect 571 251 584 285
rect 521 235 584 251
rect 620 144 654 405
rect 425 115 491 144
rect 183 53 249 81
rect 425 81 441 115
rect 475 81 491 115
rect 425 17 491 81
rect 583 115 654 144
rect 583 81 599 115
rect 633 81 654 115
rect 583 53 654 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a31o_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2765118
string GDS_START 2758480
<< end >>
