magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 1 49 634 241
rect 0 0 672 49
<< scnmos >>
rect 80 47 110 215
rect 152 47 182 215
rect 267 47 297 215
rect 353 47 383 215
rect 439 47 469 215
rect 525 47 555 215
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 267 367 297 619
rect 353 367 383 619
rect 439 367 469 619
rect 525 367 555 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 101 80 169
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 47 152 215
rect 182 163 267 215
rect 182 129 207 163
rect 241 129 267 163
rect 182 89 267 129
rect 182 55 207 89
rect 241 55 267 89
rect 182 47 267 55
rect 297 203 353 215
rect 297 169 308 203
rect 342 169 353 203
rect 297 101 353 169
rect 297 67 308 101
rect 342 67 353 101
rect 297 47 353 67
rect 383 177 439 215
rect 383 143 394 177
rect 428 143 439 177
rect 383 93 439 143
rect 383 59 394 93
rect 428 59 439 93
rect 383 47 439 59
rect 469 203 525 215
rect 469 169 480 203
rect 514 169 525 203
rect 469 101 525 169
rect 469 67 480 101
rect 514 67 525 101
rect 469 47 525 67
rect 555 177 608 215
rect 555 143 566 177
rect 600 143 608 177
rect 555 93 608 143
rect 555 59 566 93
rect 600 59 608 93
rect 555 47 608 59
<< pdiff >>
rect 27 607 80 619
rect 27 573 35 607
rect 69 573 80 607
rect 27 511 80 573
rect 27 477 35 511
rect 69 477 80 511
rect 27 418 80 477
rect 27 384 35 418
rect 69 384 80 418
rect 27 367 80 384
rect 110 599 166 619
rect 110 565 121 599
rect 155 565 166 599
rect 110 517 166 565
rect 110 483 121 517
rect 155 483 166 517
rect 110 436 166 483
rect 110 402 121 436
rect 155 402 166 436
rect 110 367 166 402
rect 196 607 267 619
rect 196 573 214 607
rect 248 573 267 607
rect 196 494 267 573
rect 196 460 214 494
rect 248 460 267 494
rect 196 367 267 460
rect 297 599 353 619
rect 297 565 308 599
rect 342 565 353 599
rect 297 511 353 565
rect 297 477 308 511
rect 342 477 353 511
rect 297 413 353 477
rect 297 379 308 413
rect 342 379 353 413
rect 297 367 353 379
rect 383 611 439 619
rect 383 577 394 611
rect 428 577 439 611
rect 383 532 439 577
rect 383 498 394 532
rect 428 498 439 532
rect 383 457 439 498
rect 383 423 394 457
rect 428 423 439 457
rect 383 367 439 423
rect 469 599 525 619
rect 469 565 480 599
rect 514 565 525 599
rect 469 511 525 565
rect 469 477 480 511
rect 514 477 525 511
rect 469 413 525 477
rect 469 379 480 413
rect 514 379 525 413
rect 469 367 525 379
rect 555 607 608 619
rect 555 573 566 607
rect 600 573 608 607
rect 555 532 608 573
rect 555 498 566 532
rect 600 498 608 532
rect 555 457 608 498
rect 555 423 566 457
rect 600 423 608 457
rect 555 367 608 423
<< ndiffc >>
rect 35 169 69 203
rect 35 67 69 101
rect 207 129 241 163
rect 207 55 241 89
rect 308 169 342 203
rect 308 67 342 101
rect 394 143 428 177
rect 394 59 428 93
rect 480 169 514 203
rect 480 67 514 101
rect 566 143 600 177
rect 566 59 600 93
<< pdiffc >>
rect 35 573 69 607
rect 35 477 69 511
rect 35 384 69 418
rect 121 565 155 599
rect 121 483 155 517
rect 121 402 155 436
rect 214 573 248 607
rect 214 460 248 494
rect 308 565 342 599
rect 308 477 342 511
rect 308 379 342 413
rect 394 577 428 611
rect 394 498 428 532
rect 394 423 428 457
rect 480 565 514 599
rect 480 477 514 511
rect 480 379 514 413
rect 566 573 600 607
rect 566 498 600 532
rect 566 423 600 457
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 267 619 297 645
rect 353 619 383 645
rect 439 619 469 645
rect 525 619 555 645
rect 80 345 110 367
rect 25 315 110 345
rect 166 335 196 367
rect 152 319 218 335
rect 25 309 91 315
rect 25 275 41 309
rect 75 275 91 309
rect 25 267 91 275
rect 152 285 168 319
rect 202 285 218 319
rect 152 269 218 285
rect 267 333 297 367
rect 353 333 383 367
rect 439 333 469 367
rect 525 333 555 367
rect 267 317 555 333
rect 267 283 283 317
rect 317 283 351 317
rect 385 283 419 317
rect 453 283 487 317
rect 521 283 555 317
rect 25 237 110 267
rect 80 215 110 237
rect 152 215 182 269
rect 267 267 555 283
rect 267 215 297 267
rect 353 215 383 267
rect 439 215 469 267
rect 525 215 555 267
rect 80 21 110 47
rect 152 21 182 47
rect 267 21 297 47
rect 353 21 383 47
rect 439 21 469 47
rect 525 21 555 47
<< polycont >>
rect 41 275 75 309
rect 168 285 202 319
rect 283 283 317 317
rect 351 283 385 317
rect 419 283 453 317
rect 487 283 521 317
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 19 607 85 649
rect 19 573 35 607
rect 69 573 85 607
rect 19 511 85 573
rect 19 477 35 511
rect 69 477 85 511
rect 19 418 85 477
rect 19 384 35 418
rect 69 384 85 418
rect 119 599 157 615
rect 119 565 121 599
rect 155 565 157 599
rect 119 517 157 565
rect 119 483 121 517
rect 155 483 157 517
rect 119 436 157 483
rect 198 607 264 649
rect 198 573 214 607
rect 248 573 264 607
rect 198 494 264 573
rect 198 460 214 494
rect 248 460 264 494
rect 198 454 264 460
rect 306 599 344 615
rect 306 565 308 599
rect 342 565 344 599
rect 306 511 344 565
rect 306 477 308 511
rect 342 477 344 511
rect 119 402 121 436
rect 155 420 157 436
rect 155 402 272 420
rect 119 386 272 402
rect 25 309 91 350
rect 25 275 41 309
rect 75 275 91 309
rect 25 265 91 275
rect 127 319 204 350
rect 127 285 168 319
rect 202 285 204 319
rect 127 265 204 285
rect 238 321 272 386
rect 306 413 344 477
rect 378 611 444 649
rect 378 577 394 611
rect 428 577 444 611
rect 378 532 444 577
rect 378 498 394 532
rect 428 498 444 532
rect 378 457 444 498
rect 378 423 394 457
rect 428 423 444 457
rect 478 599 516 615
rect 478 565 480 599
rect 514 565 516 599
rect 478 511 516 565
rect 478 477 480 511
rect 514 477 516 511
rect 306 379 308 413
rect 342 389 344 413
rect 478 413 516 477
rect 550 607 616 649
rect 550 573 566 607
rect 600 573 616 607
rect 550 532 616 573
rect 550 498 566 532
rect 600 498 616 532
rect 550 457 616 498
rect 550 423 566 457
rect 600 423 616 457
rect 478 389 480 413
rect 342 379 480 389
rect 514 389 516 413
rect 514 379 652 389
rect 306 355 652 379
rect 238 317 537 321
rect 238 283 283 317
rect 317 283 351 317
rect 385 283 419 317
rect 453 283 487 317
rect 521 283 537 317
rect 238 281 537 283
rect 238 231 272 281
rect 571 247 652 355
rect 19 203 272 231
rect 19 169 35 203
rect 69 197 272 203
rect 306 213 652 247
rect 306 203 344 213
rect 69 169 85 197
rect 19 101 85 169
rect 306 169 308 203
rect 342 169 344 203
rect 478 203 516 213
rect 19 67 35 101
rect 69 67 85 101
rect 19 51 85 67
rect 191 129 207 163
rect 241 129 257 163
rect 191 89 257 129
rect 191 55 207 89
rect 241 55 257 89
rect 191 17 257 55
rect 306 101 344 169
rect 306 67 308 101
rect 342 67 344 101
rect 306 51 344 67
rect 378 143 394 177
rect 428 143 444 177
rect 378 93 444 143
rect 378 59 394 93
rect 428 59 444 93
rect 378 17 444 59
rect 478 169 480 203
rect 514 169 516 203
rect 478 101 516 169
rect 478 67 480 101
rect 514 67 516 101
rect 478 51 516 67
rect 550 143 566 177
rect 600 143 616 177
rect 550 93 616 143
rect 550 59 566 93
rect 600 59 616 93
rect 550 17 616 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and2_4
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3532380
string GDS_START 3525880
<< end >>
