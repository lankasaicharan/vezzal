magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1345 2586 1852
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 1 21 1235 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 177 47 207 177
rect 271 47 301 177
rect 375 47 405 177
rect 459 47 489 177
rect 553 47 583 177
rect 657 47 687 177
rect 741 47 771 177
rect 835 47 865 177
rect 929 47 959 177
rect 1033 47 1063 177
rect 1127 47 1157 177
<< scpmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 461 297 497 497
rect 555 297 591 497
rect 649 297 685 497
rect 743 297 779 497
rect 837 297 873 497
rect 931 297 967 497
rect 1025 297 1061 497
rect 1119 297 1155 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 177 177
rect 113 129 133 163
rect 167 129 177 163
rect 113 95 177 129
rect 113 61 133 95
rect 167 61 177 95
rect 113 47 177 61
rect 207 95 271 177
rect 207 61 227 95
rect 261 61 271 95
rect 207 47 271 61
rect 301 163 375 177
rect 301 129 321 163
rect 355 129 375 163
rect 301 95 375 129
rect 301 61 321 95
rect 355 61 375 95
rect 301 47 375 61
rect 405 95 459 177
rect 405 61 415 95
rect 449 61 459 95
rect 405 47 459 61
rect 489 163 553 177
rect 489 129 509 163
rect 543 129 553 163
rect 489 95 553 129
rect 489 61 509 95
rect 543 61 553 95
rect 489 47 553 61
rect 583 95 657 177
rect 583 61 603 95
rect 637 61 657 95
rect 583 47 657 61
rect 687 163 741 177
rect 687 129 697 163
rect 731 129 741 163
rect 687 95 741 129
rect 687 61 697 95
rect 731 61 741 95
rect 687 47 741 61
rect 771 95 835 177
rect 771 61 791 95
rect 825 61 835 95
rect 771 47 835 61
rect 865 163 929 177
rect 865 129 885 163
rect 919 129 929 163
rect 865 95 929 129
rect 865 61 885 95
rect 919 61 929 95
rect 865 47 929 61
rect 959 95 1033 177
rect 959 61 979 95
rect 1013 61 1033 95
rect 959 47 1033 61
rect 1063 163 1127 177
rect 1063 129 1073 163
rect 1107 129 1127 163
rect 1063 95 1127 129
rect 1063 61 1073 95
rect 1107 61 1127 95
rect 1063 47 1127 61
rect 1157 95 1209 177
rect 1157 61 1167 95
rect 1201 61 1209 95
rect 1157 47 1209 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 297 179 375
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 477 367 497
rect 309 443 321 477
rect 355 443 367 477
rect 309 409 367 443
rect 309 375 321 409
rect 355 375 367 409
rect 309 297 367 375
rect 403 477 461 497
rect 403 443 415 477
rect 449 443 461 477
rect 403 409 461 443
rect 403 375 415 409
rect 449 375 461 409
rect 403 341 461 375
rect 403 307 415 341
rect 449 307 461 341
rect 403 297 461 307
rect 497 341 555 497
rect 497 307 509 341
rect 543 307 555 341
rect 497 297 555 307
rect 591 477 649 497
rect 591 443 603 477
rect 637 443 649 477
rect 591 409 649 443
rect 591 375 603 409
rect 637 375 649 409
rect 591 297 649 375
rect 685 477 743 497
rect 685 443 697 477
rect 731 443 743 477
rect 685 409 743 443
rect 685 375 697 409
rect 731 375 743 409
rect 685 341 743 375
rect 685 307 697 341
rect 731 307 743 341
rect 685 297 743 307
rect 779 409 837 497
rect 779 375 791 409
rect 825 375 837 409
rect 779 297 837 375
rect 873 477 931 497
rect 873 443 885 477
rect 919 443 931 477
rect 873 297 931 443
rect 967 409 1025 497
rect 967 375 979 409
rect 1013 375 1025 409
rect 967 297 1025 375
rect 1061 477 1119 497
rect 1061 443 1073 477
rect 1107 443 1119 477
rect 1061 297 1119 443
rect 1155 477 1209 497
rect 1155 443 1167 477
rect 1201 443 1209 477
rect 1155 297 1209 443
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 415 61 449 95
rect 509 129 543 163
rect 509 61 543 95
rect 603 61 637 95
rect 697 129 731 163
rect 697 61 731 95
rect 791 61 825 95
rect 885 129 919 163
rect 885 61 919 95
rect 979 61 1013 95
rect 1073 129 1107 163
rect 1073 61 1107 95
rect 1167 61 1201 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 443 167 477
rect 133 375 167 409
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 443 355 477
rect 321 375 355 409
rect 415 443 449 477
rect 415 375 449 409
rect 415 307 449 341
rect 509 307 543 341
rect 603 443 637 477
rect 603 375 637 409
rect 697 443 731 477
rect 697 375 731 409
rect 697 307 731 341
rect 791 375 825 409
rect 885 443 919 477
rect 979 375 1013 409
rect 1073 443 1107 477
rect 1167 443 1201 477
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 461 497 497 523
rect 555 497 591 523
rect 649 497 685 523
rect 743 497 779 523
rect 837 497 873 523
rect 931 497 967 523
rect 1025 497 1061 523
rect 1119 497 1155 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 461 282 497 297
rect 555 282 591 297
rect 649 282 685 297
rect 743 282 779 297
rect 837 282 873 297
rect 931 282 967 297
rect 1025 282 1061 297
rect 1119 282 1155 297
rect 83 265 123 282
rect 177 265 217 282
rect 271 265 311 282
rect 365 265 405 282
rect 83 249 405 265
rect 83 215 99 249
rect 133 215 177 249
rect 211 215 255 249
rect 289 215 333 249
rect 367 215 405 249
rect 83 199 405 215
rect 83 177 113 199
rect 177 177 207 199
rect 271 177 301 199
rect 375 177 405 199
rect 459 265 499 282
rect 553 265 593 282
rect 647 265 687 282
rect 459 249 687 265
rect 459 215 475 249
rect 509 215 553 249
rect 587 215 687 249
rect 459 199 687 215
rect 459 177 489 199
rect 553 177 583 199
rect 657 177 687 199
rect 741 265 781 282
rect 835 265 875 282
rect 929 265 969 282
rect 1023 265 1063 282
rect 1117 265 1157 282
rect 741 249 1063 265
rect 741 215 913 249
rect 947 215 991 249
rect 1025 215 1063 249
rect 741 199 1063 215
rect 1109 249 1185 265
rect 1109 215 1125 249
rect 1159 215 1185 249
rect 1109 199 1185 215
rect 741 177 771 199
rect 835 177 865 199
rect 929 177 959 199
rect 1033 177 1063 199
rect 1127 177 1157 199
rect 83 21 113 47
rect 177 21 207 47
rect 271 21 301 47
rect 375 21 405 47
rect 459 21 489 47
rect 553 21 583 47
rect 657 21 687 47
rect 741 21 771 47
rect 835 21 865 47
rect 929 21 959 47
rect 1033 21 1063 47
rect 1127 21 1157 47
<< polycont >>
rect 99 215 133 249
rect 177 215 211 249
rect 255 215 289 249
rect 333 215 367 249
rect 475 215 509 249
rect 553 215 587 249
rect 913 215 947 249
rect 991 215 1025 249
rect 1125 215 1159 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 30 477 81 493
rect 30 443 39 477
rect 73 443 81 477
rect 30 409 81 443
rect 30 375 39 409
rect 73 375 81 409
rect 30 341 81 375
rect 125 477 175 527
rect 125 443 133 477
rect 167 443 175 477
rect 125 409 175 443
rect 125 375 133 409
rect 167 375 175 409
rect 125 359 175 375
rect 219 477 269 493
rect 219 443 227 477
rect 261 443 269 477
rect 219 409 269 443
rect 219 375 227 409
rect 261 375 269 409
rect 30 307 39 341
rect 73 325 81 341
rect 219 341 269 375
rect 313 477 363 527
rect 313 443 321 477
rect 355 443 363 477
rect 313 409 363 443
rect 313 375 321 409
rect 355 375 363 409
rect 313 359 363 375
rect 407 477 645 493
rect 407 443 415 477
rect 449 459 603 477
rect 449 443 539 459
rect 407 425 539 443
rect 573 443 603 459
rect 637 443 645 477
rect 573 425 645 443
rect 407 417 645 425
rect 407 409 457 417
rect 407 375 415 409
rect 449 375 457 409
rect 595 409 645 417
rect 219 325 227 341
rect 73 307 227 325
rect 261 325 269 341
rect 407 341 457 375
rect 407 325 415 341
rect 261 307 415 325
rect 449 307 457 341
rect 30 291 457 307
rect 501 341 551 383
rect 595 375 603 409
rect 637 375 645 409
rect 595 359 645 375
rect 689 477 1115 493
rect 689 443 697 477
rect 731 459 885 477
rect 731 443 739 459
rect 689 409 739 443
rect 877 443 885 459
rect 919 459 1073 477
rect 919 443 927 459
rect 877 427 927 443
rect 1065 443 1073 459
rect 1107 443 1115 477
rect 1065 427 1115 443
rect 1159 477 1209 493
rect 1159 459 1167 477
rect 1159 425 1161 459
rect 1201 443 1209 477
rect 1195 425 1209 443
rect 689 375 697 409
rect 731 375 739 409
rect 501 307 509 341
rect 543 325 551 341
rect 689 341 739 375
rect 783 409 833 425
rect 783 375 791 409
rect 825 393 833 409
rect 971 409 1021 425
rect 971 393 979 409
rect 825 375 979 393
rect 1013 391 1021 409
rect 1013 375 1269 391
rect 783 357 1269 375
rect 689 325 697 341
rect 543 307 697 325
rect 731 307 739 341
rect 501 291 739 307
rect 783 289 1143 323
rect 783 257 817 289
rect 18 249 405 257
rect 18 215 99 249
rect 133 215 177 249
rect 211 215 255 249
rect 289 215 333 249
rect 367 215 405 249
rect 459 249 817 257
rect 1109 257 1143 289
rect 459 215 475 249
rect 509 215 553 249
rect 587 215 817 249
rect 851 249 1063 255
rect 851 215 913 249
rect 947 215 991 249
rect 1025 215 1063 249
rect 1109 249 1177 257
rect 1109 215 1125 249
rect 1159 215 1177 249
rect 1211 181 1269 357
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 1269 181
rect 107 129 133 163
rect 167 145 321 163
rect 167 129 183 145
rect 107 95 183 129
rect 295 129 321 145
rect 355 145 509 163
rect 355 129 371 145
rect 107 61 133 95
rect 167 61 183 95
rect 107 51 183 61
rect 227 95 261 111
rect 227 17 261 61
rect 295 95 371 129
rect 483 129 509 145
rect 543 145 697 163
rect 543 129 559 145
rect 295 61 321 95
rect 355 61 371 95
rect 295 51 371 61
rect 415 95 449 111
rect 415 17 449 61
rect 483 95 559 129
rect 671 129 697 145
rect 731 145 885 163
rect 731 129 747 145
rect 483 61 509 95
rect 543 61 559 95
rect 483 51 559 61
rect 603 95 637 111
rect 603 17 637 61
rect 671 95 747 129
rect 859 129 885 145
rect 919 145 1073 163
rect 919 129 935 145
rect 671 61 697 95
rect 731 61 747 95
rect 671 51 747 61
rect 791 95 825 111
rect 791 17 825 61
rect 859 95 935 129
rect 1047 129 1073 145
rect 1107 145 1269 163
rect 1107 129 1123 145
rect 859 61 885 95
rect 919 61 935 95
rect 859 51 935 61
rect 979 95 1013 111
rect 979 17 1013 61
rect 1047 95 1123 129
rect 1047 61 1073 95
rect 1107 61 1123 95
rect 1047 51 1123 61
rect 1167 95 1201 111
rect 1167 17 1201 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 539 425 573 459
rect 1161 443 1167 459
rect 1167 443 1195 459
rect 1161 425 1195 443
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 527 459 596 467
rect 527 425 539 459
rect 573 456 596 459
rect 1139 459 1208 467
rect 1139 456 1161 459
rect 573 428 1161 456
rect 573 425 596 428
rect 527 413 596 425
rect 1139 425 1161 428
rect 1195 425 1208 459
rect 1139 413 1208 425
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< comment >>
rect 846 -85 847 -84
<< labels >>
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 580 221 614 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 1225 289 1259 323 0 FreeSans 400 0 0 0 Y
port 8 nsew signal output
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor3_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1307502
string GDS_START 1297610
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
