magic
tech sky130A
magscale 1 2
timestamp 1627201166
<< checkpaint >>
rect -1260 -1260 3542 3598
<< pwell >>
rect 1178 1416 1199 1465
<< poly >>
rect 0 2322 2282 2338
rect 0 2288 97 2322
rect 131 2288 165 2322
rect 199 2288 233 2322
rect 267 2288 301 2322
rect 335 2288 369 2322
rect 403 2288 437 2322
rect 471 2288 505 2322
rect 539 2288 573 2322
rect 607 2288 641 2322
rect 675 2288 709 2322
rect 743 2288 777 2322
rect 811 2288 845 2322
rect 879 2288 913 2322
rect 947 2288 981 2322
rect 1015 2288 1049 2322
rect 1083 2288 1199 2322
rect 1233 2288 1267 2322
rect 1301 2288 1335 2322
rect 1369 2288 1403 2322
rect 1437 2288 1471 2322
rect 1505 2288 1539 2322
rect 1573 2288 1607 2322
rect 1641 2288 1675 2322
rect 1709 2288 1743 2322
rect 1777 2288 1811 2322
rect 1845 2288 1879 2322
rect 1913 2288 1947 2322
rect 1981 2288 2015 2322
rect 2049 2288 2083 2322
rect 2117 2288 2151 2322
rect 2185 2288 2282 2322
rect 0 2274 2282 2288
rect 0 2240 16 2274
rect 50 2240 2232 2274
rect 2266 2240 2282 2274
rect 0 2206 2282 2240
rect 0 2172 16 2206
rect 50 2172 2232 2206
rect 2266 2172 2282 2206
rect 0 2138 2282 2172
rect 0 2104 16 2138
rect 50 2104 2232 2138
rect 2266 2104 2282 2138
rect 0 2070 2282 2104
rect 0 2036 16 2070
rect 50 2036 2232 2070
rect 2266 2036 2282 2070
rect 0 2002 2282 2036
rect 0 1968 16 2002
rect 50 1968 2232 2002
rect 2266 1968 2282 2002
rect 0 1934 2282 1968
rect 0 1900 16 1934
rect 50 1900 2232 1934
rect 2266 1900 2282 1934
rect 0 1866 2282 1900
rect 0 1832 16 1866
rect 50 1832 2232 1866
rect 2266 1832 2282 1866
rect 0 1798 2282 1832
rect 0 1764 16 1798
rect 50 1764 2232 1798
rect 2266 1764 2282 1798
rect 0 1730 2282 1764
rect 0 1696 16 1730
rect 50 1696 2232 1730
rect 2266 1696 2282 1730
rect 0 1662 2282 1696
rect 0 1628 16 1662
rect 50 1628 2232 1662
rect 2266 1628 2282 1662
rect 0 1594 2282 1628
rect 0 1560 16 1594
rect 50 1560 2232 1594
rect 2266 1560 2282 1594
rect 0 1526 2282 1560
rect 0 1492 16 1526
rect 50 1492 2232 1526
rect 2266 1492 2282 1526
rect 0 1458 2282 1492
rect 0 1424 16 1458
rect 50 1424 2232 1458
rect 2266 1424 2282 1458
rect 0 1390 2282 1424
rect 0 1356 16 1390
rect 50 1356 2232 1390
rect 2266 1356 2282 1390
rect 0 1322 2282 1356
rect 0 1288 16 1322
rect 50 1288 2232 1322
rect 2266 1288 2282 1322
rect 0 1254 2282 1288
rect 0 1220 16 1254
rect 50 1220 2232 1254
rect 2266 1220 2282 1254
rect 0 1186 2282 1220
rect 0 1152 16 1186
rect 50 1152 2232 1186
rect 2266 1152 2282 1186
rect 0 1118 2282 1152
rect 0 1084 16 1118
rect 50 1084 2232 1118
rect 2266 1084 2282 1118
rect 0 1050 2282 1084
rect 0 1016 16 1050
rect 50 1016 2232 1050
rect 2266 1016 2282 1050
rect 0 982 2282 1016
rect 0 948 16 982
rect 50 948 2232 982
rect 2266 948 2282 982
rect 0 914 2282 948
rect 0 880 16 914
rect 50 880 2232 914
rect 2266 880 2282 914
rect 0 846 2282 880
rect 0 812 16 846
rect 50 812 2232 846
rect 2266 812 2282 846
rect 0 778 2282 812
rect 0 744 16 778
rect 50 744 2232 778
rect 2266 744 2282 778
rect 0 710 2282 744
rect 0 676 16 710
rect 50 676 2232 710
rect 2266 676 2282 710
rect 0 642 2282 676
rect 0 608 16 642
rect 50 608 2232 642
rect 2266 608 2282 642
rect 0 574 2282 608
rect 0 540 16 574
rect 50 540 2232 574
rect 2266 540 2282 574
rect 0 506 2282 540
rect 0 472 16 506
rect 50 472 2232 506
rect 2266 472 2282 506
rect 0 438 2282 472
rect 0 404 16 438
rect 50 404 2232 438
rect 2266 404 2282 438
rect 0 370 2282 404
rect 0 336 16 370
rect 50 336 2232 370
rect 2266 336 2282 370
rect 0 302 2282 336
rect 0 268 16 302
rect 50 268 2232 302
rect 2266 268 2282 302
rect 0 234 2282 268
rect 0 200 16 234
rect 50 200 2232 234
rect 2266 200 2282 234
rect 0 166 2282 200
rect 0 132 16 166
rect 50 132 2232 166
rect 2266 132 2282 166
rect 0 98 2282 132
rect 0 64 16 98
rect 50 64 2232 98
rect 2266 64 2282 98
rect 0 50 2282 64
rect 0 16 97 50
rect 131 16 165 50
rect 199 16 233 50
rect 267 16 301 50
rect 335 16 369 50
rect 403 16 437 50
rect 471 16 505 50
rect 539 16 573 50
rect 607 16 641 50
rect 675 16 709 50
rect 743 16 777 50
rect 811 16 845 50
rect 879 16 913 50
rect 947 16 981 50
rect 1015 16 1049 50
rect 1083 16 1199 50
rect 1233 16 1267 50
rect 1301 16 1335 50
rect 1369 16 1403 50
rect 1437 16 1471 50
rect 1505 16 1539 50
rect 1573 16 1607 50
rect 1641 16 1675 50
rect 1709 16 1743 50
rect 1777 16 1811 50
rect 1845 16 1879 50
rect 1913 16 1947 50
rect 1981 16 2015 50
rect 2049 16 2083 50
rect 2117 16 2151 50
rect 2185 16 2282 50
rect 0 0 2282 16
<< polycont >>
rect 97 2288 131 2322
rect 165 2288 199 2322
rect 233 2288 267 2322
rect 301 2288 335 2322
rect 369 2288 403 2322
rect 437 2288 471 2322
rect 505 2288 539 2322
rect 573 2288 607 2322
rect 641 2288 675 2322
rect 709 2288 743 2322
rect 777 2288 811 2322
rect 845 2288 879 2322
rect 913 2288 947 2322
rect 981 2288 1015 2322
rect 1049 2288 1083 2322
rect 1199 2288 1233 2322
rect 1267 2288 1301 2322
rect 1335 2288 1369 2322
rect 1403 2288 1437 2322
rect 1471 2288 1505 2322
rect 1539 2288 1573 2322
rect 1607 2288 1641 2322
rect 1675 2288 1709 2322
rect 1743 2288 1777 2322
rect 1811 2288 1845 2322
rect 1879 2288 1913 2322
rect 1947 2288 1981 2322
rect 2015 2288 2049 2322
rect 2083 2288 2117 2322
rect 2151 2288 2185 2322
rect 16 2240 50 2274
rect 2232 2240 2266 2274
rect 16 2172 50 2206
rect 2232 2172 2266 2206
rect 16 2104 50 2138
rect 2232 2104 2266 2138
rect 16 2036 50 2070
rect 2232 2036 2266 2070
rect 16 1968 50 2002
rect 2232 1968 2266 2002
rect 16 1900 50 1934
rect 2232 1900 2266 1934
rect 16 1832 50 1866
rect 2232 1832 2266 1866
rect 16 1764 50 1798
rect 2232 1764 2266 1798
rect 16 1696 50 1730
rect 2232 1696 2266 1730
rect 16 1628 50 1662
rect 2232 1628 2266 1662
rect 16 1560 50 1594
rect 2232 1560 2266 1594
rect 16 1492 50 1526
rect 2232 1492 2266 1526
rect 16 1424 50 1458
rect 2232 1424 2266 1458
rect 16 1356 50 1390
rect 2232 1356 2266 1390
rect 16 1288 50 1322
rect 2232 1288 2266 1322
rect 16 1220 50 1254
rect 2232 1220 2266 1254
rect 16 1152 50 1186
rect 2232 1152 2266 1186
rect 16 1084 50 1118
rect 2232 1084 2266 1118
rect 16 1016 50 1050
rect 2232 1016 2266 1050
rect 16 948 50 982
rect 2232 948 2266 982
rect 16 880 50 914
rect 2232 880 2266 914
rect 16 812 50 846
rect 2232 812 2266 846
rect 16 744 50 778
rect 2232 744 2266 778
rect 16 676 50 710
rect 2232 676 2266 710
rect 16 608 50 642
rect 2232 608 2266 642
rect 16 540 50 574
rect 2232 540 2266 574
rect 16 472 50 506
rect 2232 472 2266 506
rect 16 404 50 438
rect 2232 404 2266 438
rect 16 336 50 370
rect 2232 336 2266 370
rect 16 268 50 302
rect 2232 268 2266 302
rect 16 200 50 234
rect 2232 200 2266 234
rect 16 132 50 166
rect 2232 132 2266 166
rect 16 64 50 98
rect 2232 64 2266 98
rect 97 16 131 50
rect 165 16 199 50
rect 233 16 267 50
rect 301 16 335 50
rect 369 16 403 50
rect 437 16 471 50
rect 505 16 539 50
rect 573 16 607 50
rect 641 16 675 50
rect 709 16 743 50
rect 777 16 811 50
rect 845 16 879 50
rect 913 16 947 50
rect 981 16 1015 50
rect 1049 16 1083 50
rect 1199 16 1233 50
rect 1267 16 1301 50
rect 1335 16 1369 50
rect 1403 16 1437 50
rect 1471 16 1505 50
rect 1539 16 1573 50
rect 1607 16 1641 50
rect 1675 16 1709 50
rect 1743 16 1777 50
rect 1811 16 1845 50
rect 1879 16 1913 50
rect 1947 16 1981 50
rect 2015 16 2049 50
rect 2083 16 2117 50
rect 2151 16 2185 50
<< locali >>
rect 0 2322 2282 2338
rect 0 2288 80 2322
rect 131 2288 152 2322
rect 199 2288 224 2322
rect 267 2288 296 2322
rect 335 2288 368 2322
rect 403 2288 437 2322
rect 474 2288 505 2322
rect 546 2288 573 2322
rect 618 2288 641 2322
rect 690 2288 709 2322
rect 762 2288 777 2322
rect 834 2288 845 2322
rect 906 2288 913 2322
rect 978 2288 981 2322
rect 1015 2288 1016 2322
rect 1083 2288 1088 2322
rect 1122 2288 1160 2322
rect 1194 2288 1199 2322
rect 1266 2288 1267 2322
rect 1301 2288 1304 2322
rect 1369 2288 1376 2322
rect 1437 2288 1448 2322
rect 1505 2288 1520 2322
rect 1573 2288 1592 2322
rect 1641 2288 1664 2322
rect 1709 2288 1736 2322
rect 1777 2288 1808 2322
rect 1845 2288 1879 2322
rect 1914 2288 1947 2322
rect 1986 2288 2015 2322
rect 2058 2288 2083 2322
rect 2130 2288 2151 2322
rect 2202 2288 2282 2322
rect 0 2274 2282 2288
rect 0 2240 16 2274
rect 50 2272 2232 2274
rect 50 2240 66 2272
rect 0 2222 66 2240
rect 2216 2240 2232 2272
rect 2266 2240 2282 2274
rect 0 2172 16 2222
rect 50 2172 66 2222
rect 100 2220 2181 2238
rect 100 2200 1124 2220
rect 0 2166 66 2172
rect 1114 2186 1124 2200
rect 1158 2200 2181 2220
rect 2216 2222 2282 2240
rect 1158 2186 1168 2200
rect 0 2150 1080 2166
rect 0 2104 16 2150
rect 50 2132 1080 2150
rect 1114 2148 1168 2186
rect 2216 2172 2232 2222
rect 2266 2172 2282 2222
rect 2216 2166 2282 2172
rect 50 2104 66 2132
rect 0 2078 66 2104
rect 1114 2114 1124 2148
rect 1158 2114 1168 2148
rect 1202 2150 2282 2166
rect 1202 2132 2232 2150
rect 1114 2098 1168 2114
rect 2216 2104 2232 2132
rect 2266 2104 2282 2150
rect 0 2036 16 2078
rect 50 2036 66 2078
rect 100 2076 2181 2098
rect 100 2060 1124 2076
rect 0 2026 66 2036
rect 1114 2042 1124 2060
rect 1158 2060 2181 2076
rect 2216 2078 2282 2104
rect 1158 2042 1168 2060
rect 0 2006 1080 2026
rect 0 1968 16 2006
rect 50 1992 1080 2006
rect 1114 2004 1168 2042
rect 2216 2036 2232 2078
rect 2266 2036 2282 2078
rect 2216 2026 2282 2036
rect 50 1968 66 1992
rect 0 1934 66 1968
rect 1114 1970 1124 2004
rect 1158 1970 1168 2004
rect 1202 2006 2282 2026
rect 1202 1992 2232 2006
rect 1114 1958 1168 1970
rect 2216 1968 2232 1992
rect 2266 1968 2282 2006
rect 0 1900 16 1934
rect 50 1900 66 1934
rect 100 1932 2181 1958
rect 100 1920 1124 1932
rect 0 1886 66 1900
rect 1114 1898 1124 1920
rect 1158 1920 2181 1932
rect 2216 1934 2282 1968
rect 1158 1898 1168 1920
rect 0 1866 1080 1886
rect 0 1828 16 1866
rect 50 1852 1080 1866
rect 1114 1860 1168 1898
rect 2216 1900 2232 1934
rect 2266 1900 2282 1934
rect 2216 1886 2282 1900
rect 50 1828 66 1852
rect 0 1798 66 1828
rect 1114 1826 1124 1860
rect 1158 1826 1168 1860
rect 1202 1866 2282 1886
rect 1202 1852 2232 1866
rect 1114 1818 1168 1826
rect 2216 1828 2232 1852
rect 2266 1828 2282 1866
rect 0 1756 16 1798
rect 50 1756 66 1798
rect 100 1788 2181 1818
rect 100 1780 1124 1788
rect 0 1746 66 1756
rect 1114 1754 1124 1780
rect 1158 1780 2181 1788
rect 2216 1798 2282 1828
rect 1158 1754 1168 1780
rect 0 1730 1080 1746
rect 0 1684 16 1730
rect 50 1712 1080 1730
rect 1114 1716 1168 1754
rect 2216 1756 2232 1798
rect 2266 1756 2282 1798
rect 2216 1746 2282 1756
rect 50 1684 66 1712
rect 0 1662 66 1684
rect 1114 1682 1124 1716
rect 1158 1682 1168 1716
rect 1202 1730 2282 1746
rect 1202 1712 2232 1730
rect 1114 1678 1168 1682
rect 2216 1684 2232 1712
rect 2266 1684 2282 1730
rect 0 1612 16 1662
rect 50 1612 66 1662
rect 100 1644 2181 1678
rect 100 1640 1124 1644
rect 0 1606 66 1612
rect 1114 1610 1124 1640
rect 1158 1640 2181 1644
rect 2216 1662 2282 1684
rect 1158 1610 1168 1640
rect 0 1594 1080 1606
rect 0 1540 16 1594
rect 50 1572 1080 1594
rect 1114 1572 1168 1610
rect 2216 1612 2232 1662
rect 2266 1612 2282 1662
rect 2216 1606 2282 1612
rect 1202 1594 2282 1606
rect 1202 1572 2232 1594
rect 50 1540 66 1572
rect 0 1526 66 1540
rect 1114 1538 1124 1572
rect 1158 1538 1168 1572
rect 2216 1540 2232 1572
rect 2266 1540 2282 1594
rect 0 1468 16 1526
rect 50 1468 66 1526
rect 100 1500 2181 1538
rect 2216 1526 2282 1540
rect 0 1466 66 1468
rect 1114 1466 1124 1500
rect 1158 1466 1168 1500
rect 2216 1468 2232 1526
rect 2266 1468 2282 1526
rect 2216 1466 2282 1468
rect 0 1458 1080 1466
rect 0 1396 16 1458
rect 50 1430 1080 1458
rect 50 1396 66 1430
rect 1114 1428 1168 1466
rect 1202 1458 2282 1466
rect 1202 1432 2232 1458
rect 1114 1396 1124 1428
rect 0 1390 66 1396
rect 0 1324 16 1390
rect 50 1326 66 1390
rect 100 1394 1124 1396
rect 1158 1398 1168 1428
rect 1158 1394 2181 1398
rect 100 1360 2181 1394
rect 2216 1396 2232 1432
rect 2266 1396 2282 1458
rect 2216 1390 2282 1396
rect 1114 1356 1168 1360
rect 50 1324 1080 1326
rect 0 1322 1080 1324
rect 0 1288 16 1322
rect 50 1292 1080 1322
rect 1114 1322 1124 1356
rect 1158 1322 1168 1356
rect 2216 1326 2232 1390
rect 50 1288 66 1292
rect 0 1286 66 1288
rect 0 1220 16 1286
rect 50 1220 66 1286
rect 1114 1284 1168 1322
rect 1202 1324 2232 1326
rect 2266 1324 2282 1390
rect 1202 1322 2282 1324
rect 1202 1292 2232 1322
rect 1114 1258 1124 1284
rect 100 1250 1124 1258
rect 1158 1258 1168 1284
rect 2216 1288 2232 1292
rect 2266 1288 2282 1322
rect 2216 1286 2282 1288
rect 1158 1250 2181 1258
rect 100 1220 2181 1250
rect 2216 1220 2232 1286
rect 2266 1220 2282 1286
rect 0 1186 66 1220
rect 0 1152 16 1186
rect 50 1152 1080 1186
rect 0 1118 66 1152
rect 1114 1118 1168 1220
rect 2216 1186 2282 1220
rect 1202 1152 2232 1186
rect 2266 1152 2282 1186
rect 2216 1118 2282 1152
rect 0 1052 16 1118
rect 50 1052 66 1118
rect 100 1088 2181 1118
rect 100 1080 1124 1088
rect 0 1050 66 1052
rect 0 1016 16 1050
rect 50 1046 66 1050
rect 1114 1054 1124 1080
rect 1158 1080 2181 1088
rect 1158 1054 1168 1080
rect 50 1016 1080 1046
rect 0 1014 1080 1016
rect 0 948 16 1014
rect 50 1012 1080 1014
rect 1114 1016 1168 1054
rect 2216 1052 2232 1118
rect 2266 1052 2282 1118
rect 2216 1050 2282 1052
rect 2216 1046 2232 1050
rect 50 948 66 1012
rect 1114 982 1124 1016
rect 1158 982 1168 1016
rect 1202 1016 2232 1046
rect 2266 1016 2282 1050
rect 1202 1014 2282 1016
rect 1202 1012 2232 1014
rect 1114 978 1168 982
rect 0 942 66 948
rect 0 880 16 942
rect 50 906 66 942
rect 100 944 2181 978
rect 100 940 1124 944
rect 1114 910 1124 940
rect 1158 940 2181 944
rect 2216 948 2232 1012
rect 2266 948 2282 1014
rect 2216 942 2282 948
rect 1158 910 1168 940
rect 50 880 1080 906
rect 0 872 1080 880
rect 1114 872 1168 910
rect 2216 906 2232 942
rect 1202 880 2232 906
rect 2266 880 2282 942
rect 1202 872 2282 880
rect 0 870 66 872
rect 0 812 16 870
rect 50 812 66 870
rect 1114 838 1124 872
rect 1158 838 1168 872
rect 2216 870 2282 872
rect 0 798 66 812
rect 100 800 2181 838
rect 2216 812 2232 870
rect 2266 812 2282 870
rect 0 744 16 798
rect 50 766 66 798
rect 1114 766 1124 800
rect 1158 766 1168 800
rect 2216 798 2282 812
rect 2216 766 2232 798
rect 50 744 1080 766
rect 0 732 1080 744
rect 0 726 66 732
rect 0 676 16 726
rect 50 676 66 726
rect 1114 728 1168 766
rect 1202 744 2232 766
rect 2266 744 2282 798
rect 1202 732 2282 744
rect 1114 698 1124 728
rect 0 654 66 676
rect 100 694 1124 698
rect 1158 698 1168 728
rect 2216 726 2282 732
rect 1158 694 2181 698
rect 100 660 2181 694
rect 2216 676 2232 726
rect 2266 676 2282 726
rect 0 608 16 654
rect 50 626 66 654
rect 1114 656 1168 660
rect 50 608 1080 626
rect 0 592 1080 608
rect 1114 622 1124 656
rect 1158 622 1168 656
rect 2216 654 2282 676
rect 2216 626 2232 654
rect 0 582 66 592
rect 0 540 16 582
rect 50 540 66 582
rect 1114 584 1168 622
rect 1202 608 2232 626
rect 2266 608 2282 654
rect 1202 592 2282 608
rect 1114 558 1124 584
rect 0 510 66 540
rect 100 550 1124 558
rect 1158 558 1168 584
rect 2216 582 2282 592
rect 1158 550 2181 558
rect 100 520 2181 550
rect 2216 540 2232 582
rect 2266 540 2282 582
rect 0 472 16 510
rect 50 486 66 510
rect 1114 512 1168 520
rect 50 472 1080 486
rect 0 452 1080 472
rect 1114 478 1124 512
rect 1158 478 1168 512
rect 2216 510 2282 540
rect 2216 486 2232 510
rect 0 438 66 452
rect 0 404 16 438
rect 50 404 66 438
rect 1114 440 1168 478
rect 1202 472 2232 486
rect 2266 472 2282 510
rect 1202 452 2282 472
rect 1114 418 1124 440
rect 0 370 66 404
rect 100 406 1124 418
rect 1158 418 1168 440
rect 2216 438 2282 452
rect 1158 406 2181 418
rect 100 380 2181 406
rect 2216 404 2232 438
rect 2266 404 2282 438
rect 0 332 16 370
rect 50 346 66 370
rect 1114 368 1168 380
rect 50 332 1080 346
rect 0 312 1080 332
rect 1114 334 1124 368
rect 1158 334 1168 368
rect 2216 370 2282 404
rect 2216 346 2232 370
rect 0 302 66 312
rect 0 260 16 302
rect 50 260 66 302
rect 1114 296 1168 334
rect 1202 332 2232 346
rect 2266 332 2282 370
rect 1202 312 2282 332
rect 1114 278 1124 296
rect 0 234 66 260
rect 100 262 1124 278
rect 1158 278 1168 296
rect 2216 302 2282 312
rect 1158 262 2181 278
rect 100 240 2181 262
rect 2216 260 2232 302
rect 2266 260 2282 302
rect 0 188 16 234
rect 50 206 66 234
rect 1114 224 1168 240
rect 50 188 1080 206
rect 0 172 1080 188
rect 1114 190 1124 224
rect 1158 190 1168 224
rect 2216 234 2282 260
rect 2216 206 2232 234
rect 0 166 66 172
rect 0 116 16 166
rect 50 116 66 166
rect 1114 152 1168 190
rect 1202 188 2232 206
rect 2266 188 2282 234
rect 1202 172 2282 188
rect 1114 138 1124 152
rect 0 98 66 116
rect 100 118 1124 138
rect 1158 138 1168 152
rect 2216 166 2282 172
rect 1158 118 2181 138
rect 100 100 2181 118
rect 2216 116 2232 166
rect 2266 116 2282 166
rect 0 64 16 98
rect 50 66 66 98
rect 2216 98 2282 116
rect 2216 66 2232 98
rect 50 64 2232 66
rect 2266 64 2282 98
rect 0 50 2282 64
rect 0 16 80 50
rect 131 16 152 50
rect 199 16 224 50
rect 267 16 296 50
rect 335 16 368 50
rect 403 16 437 50
rect 474 16 505 50
rect 546 16 573 50
rect 618 16 641 50
rect 690 16 709 50
rect 762 16 777 50
rect 834 16 845 50
rect 906 16 913 50
rect 978 16 981 50
rect 1015 16 1016 50
rect 1083 16 1088 50
rect 1122 16 1160 50
rect 1194 16 1199 50
rect 1266 16 1267 50
rect 1301 16 1304 50
rect 1369 16 1376 50
rect 1437 16 1448 50
rect 1505 16 1520 50
rect 1573 16 1592 50
rect 1641 16 1664 50
rect 1709 16 1736 50
rect 1777 16 1808 50
rect 1845 16 1879 50
rect 1914 16 1947 50
rect 1986 16 2015 50
rect 2058 16 2083 50
rect 2130 16 2151 50
rect 2202 16 2282 50
rect 0 0 2282 16
<< viali >>
rect 80 2288 97 2322
rect 97 2288 114 2322
rect 152 2288 165 2322
rect 165 2288 186 2322
rect 224 2288 233 2322
rect 233 2288 258 2322
rect 296 2288 301 2322
rect 301 2288 330 2322
rect 368 2288 369 2322
rect 369 2288 402 2322
rect 440 2288 471 2322
rect 471 2288 474 2322
rect 512 2288 539 2322
rect 539 2288 546 2322
rect 584 2288 607 2322
rect 607 2288 618 2322
rect 656 2288 675 2322
rect 675 2288 690 2322
rect 728 2288 743 2322
rect 743 2288 762 2322
rect 800 2288 811 2322
rect 811 2288 834 2322
rect 872 2288 879 2322
rect 879 2288 906 2322
rect 944 2288 947 2322
rect 947 2288 978 2322
rect 1016 2288 1049 2322
rect 1049 2288 1050 2322
rect 1088 2288 1122 2322
rect 1160 2288 1194 2322
rect 1232 2288 1233 2322
rect 1233 2288 1266 2322
rect 1304 2288 1335 2322
rect 1335 2288 1338 2322
rect 1376 2288 1403 2322
rect 1403 2288 1410 2322
rect 1448 2288 1471 2322
rect 1471 2288 1482 2322
rect 1520 2288 1539 2322
rect 1539 2288 1554 2322
rect 1592 2288 1607 2322
rect 1607 2288 1626 2322
rect 1664 2288 1675 2322
rect 1675 2288 1698 2322
rect 1736 2288 1743 2322
rect 1743 2288 1770 2322
rect 1808 2288 1811 2322
rect 1811 2288 1842 2322
rect 1880 2288 1913 2322
rect 1913 2288 1914 2322
rect 1952 2288 1981 2322
rect 1981 2288 1986 2322
rect 2024 2288 2049 2322
rect 2049 2288 2058 2322
rect 2096 2288 2117 2322
rect 2117 2288 2130 2322
rect 2168 2288 2185 2322
rect 2185 2288 2202 2322
rect 16 2206 50 2222
rect 16 2188 50 2206
rect 1124 2186 1158 2220
rect 16 2138 50 2150
rect 16 2116 50 2138
rect 2232 2206 2266 2222
rect 2232 2188 2266 2206
rect 1124 2114 1158 2148
rect 2232 2138 2266 2150
rect 2232 2116 2266 2138
rect 16 2070 50 2078
rect 16 2044 50 2070
rect 1124 2042 1158 2076
rect 16 2002 50 2006
rect 16 1972 50 2002
rect 2232 2070 2266 2078
rect 2232 2044 2266 2070
rect 1124 1970 1158 2004
rect 2232 2002 2266 2006
rect 2232 1972 2266 2002
rect 16 1900 50 1934
rect 1124 1898 1158 1932
rect 16 1832 50 1862
rect 2232 1900 2266 1934
rect 16 1828 50 1832
rect 1124 1826 1158 1860
rect 2232 1832 2266 1862
rect 2232 1828 2266 1832
rect 16 1764 50 1790
rect 16 1756 50 1764
rect 1124 1754 1158 1788
rect 16 1696 50 1718
rect 2232 1764 2266 1790
rect 2232 1756 2266 1764
rect 16 1684 50 1696
rect 1124 1682 1158 1716
rect 2232 1696 2266 1718
rect 2232 1684 2266 1696
rect 16 1628 50 1646
rect 16 1612 50 1628
rect 1124 1610 1158 1644
rect 16 1560 50 1574
rect 2232 1628 2266 1646
rect 2232 1612 2266 1628
rect 16 1540 50 1560
rect 1124 1538 1158 1572
rect 2232 1560 2266 1574
rect 2232 1540 2266 1560
rect 16 1492 50 1502
rect 16 1468 50 1492
rect 1124 1466 1158 1500
rect 2232 1492 2266 1502
rect 2232 1468 2266 1492
rect 16 1424 50 1430
rect 16 1396 50 1424
rect 16 1356 50 1358
rect 16 1324 50 1356
rect 1124 1394 1158 1428
rect 2232 1424 2266 1430
rect 2232 1396 2266 1424
rect 1124 1322 1158 1356
rect 2232 1356 2266 1358
rect 16 1254 50 1286
rect 16 1252 50 1254
rect 2232 1324 2266 1356
rect 1124 1250 1158 1284
rect 2232 1254 2266 1286
rect 2232 1252 2266 1254
rect 16 1084 50 1086
rect 16 1052 50 1084
rect 1124 1054 1158 1088
rect 16 982 50 1014
rect 2232 1084 2266 1086
rect 2232 1052 2266 1084
rect 16 980 50 982
rect 1124 982 1158 1016
rect 16 914 50 942
rect 16 908 50 914
rect 1124 910 1158 944
rect 2232 982 2266 1014
rect 2232 980 2266 982
rect 2232 914 2266 942
rect 2232 908 2266 914
rect 16 846 50 870
rect 16 836 50 846
rect 1124 838 1158 872
rect 2232 846 2266 870
rect 2232 836 2266 846
rect 16 778 50 798
rect 16 764 50 778
rect 1124 766 1158 800
rect 2232 778 2266 798
rect 16 710 50 726
rect 16 692 50 710
rect 2232 764 2266 778
rect 1124 694 1158 728
rect 2232 710 2266 726
rect 2232 692 2266 710
rect 16 642 50 654
rect 16 620 50 642
rect 1124 622 1158 656
rect 2232 642 2266 654
rect 16 574 50 582
rect 16 548 50 574
rect 2232 620 2266 642
rect 1124 550 1158 584
rect 2232 574 2266 582
rect 2232 548 2266 574
rect 16 506 50 510
rect 16 476 50 506
rect 1124 478 1158 512
rect 2232 506 2266 510
rect 16 404 50 438
rect 2232 476 2266 506
rect 1124 406 1158 440
rect 2232 404 2266 438
rect 16 336 50 366
rect 16 332 50 336
rect 1124 334 1158 368
rect 16 268 50 294
rect 16 260 50 268
rect 2232 336 2266 366
rect 2232 332 2266 336
rect 1124 262 1158 296
rect 2232 268 2266 294
rect 2232 260 2266 268
rect 16 200 50 222
rect 16 188 50 200
rect 1124 190 1158 224
rect 16 132 50 150
rect 16 116 50 132
rect 2232 200 2266 222
rect 2232 188 2266 200
rect 1124 118 1158 152
rect 2232 132 2266 150
rect 2232 116 2266 132
rect 80 16 97 50
rect 97 16 114 50
rect 152 16 165 50
rect 165 16 186 50
rect 224 16 233 50
rect 233 16 258 50
rect 296 16 301 50
rect 301 16 330 50
rect 368 16 369 50
rect 369 16 402 50
rect 440 16 471 50
rect 471 16 474 50
rect 512 16 539 50
rect 539 16 546 50
rect 584 16 607 50
rect 607 16 618 50
rect 656 16 675 50
rect 675 16 690 50
rect 728 16 743 50
rect 743 16 762 50
rect 800 16 811 50
rect 811 16 834 50
rect 872 16 879 50
rect 879 16 906 50
rect 944 16 947 50
rect 947 16 978 50
rect 1016 16 1049 50
rect 1049 16 1050 50
rect 1088 16 1122 50
rect 1160 16 1194 50
rect 1232 16 1233 50
rect 1233 16 1266 50
rect 1304 16 1335 50
rect 1335 16 1338 50
rect 1376 16 1403 50
rect 1403 16 1410 50
rect 1448 16 1471 50
rect 1471 16 1482 50
rect 1520 16 1539 50
rect 1539 16 1554 50
rect 1592 16 1607 50
rect 1607 16 1626 50
rect 1664 16 1675 50
rect 1675 16 1698 50
rect 1736 16 1743 50
rect 1743 16 1770 50
rect 1808 16 1811 50
rect 1811 16 1842 50
rect 1880 16 1913 50
rect 1913 16 1914 50
rect 1952 16 1981 50
rect 1981 16 1986 50
rect 2024 16 2049 50
rect 2049 16 2058 50
rect 2096 16 2117 50
rect 2117 16 2130 50
rect 2168 16 2185 50
rect 2185 16 2202 50
<< metal1 >>
rect 0 2331 2282 2338
rect 0 2322 88 2331
rect 0 2288 80 2322
rect 0 2282 88 2288
rect 0 2230 7 2282
rect 59 2279 88 2282
rect 140 2279 152 2331
rect 204 2279 216 2331
rect 268 2279 280 2331
rect 332 2279 344 2331
rect 396 2322 408 2331
rect 460 2322 472 2331
rect 524 2322 536 2331
rect 588 2322 600 2331
rect 652 2322 664 2331
rect 402 2288 408 2322
rect 652 2288 656 2322
rect 396 2279 408 2288
rect 460 2279 472 2288
rect 524 2279 536 2288
rect 588 2279 600 2288
rect 652 2279 664 2288
rect 716 2279 728 2331
rect 780 2279 792 2331
rect 844 2279 856 2331
rect 908 2279 920 2331
rect 972 2322 984 2331
rect 1036 2322 1246 2331
rect 1298 2322 1310 2331
rect 978 2288 984 2322
rect 1050 2288 1088 2322
rect 1122 2288 1160 2322
rect 1194 2288 1232 2322
rect 1298 2288 1304 2322
rect 972 2279 984 2288
rect 1036 2279 1246 2288
rect 1298 2279 1310 2288
rect 1362 2279 1374 2331
rect 1426 2279 1438 2331
rect 1490 2279 1502 2331
rect 1554 2279 1566 2331
rect 1618 2322 1630 2331
rect 1682 2322 1694 2331
rect 1746 2322 1758 2331
rect 1810 2322 1822 2331
rect 1874 2322 1886 2331
rect 1626 2288 1630 2322
rect 1874 2288 1880 2322
rect 1618 2279 1630 2288
rect 1682 2279 1694 2288
rect 1746 2279 1758 2288
rect 1810 2279 1822 2288
rect 1874 2279 1886 2288
rect 1938 2279 1950 2331
rect 2002 2279 2014 2331
rect 2066 2279 2078 2331
rect 2130 2279 2142 2331
rect 2194 2322 2282 2331
rect 2202 2288 2282 2322
rect 2194 2282 2282 2288
rect 2194 2279 2223 2282
rect 59 2272 2223 2279
rect 59 2230 66 2272
rect 0 2222 66 2230
rect 0 2218 16 2222
rect 50 2218 66 2222
rect 0 2166 7 2218
rect 59 2166 66 2218
rect 0 2154 66 2166
rect 0 2102 7 2154
rect 59 2102 66 2154
rect 0 2090 66 2102
rect 0 2038 7 2090
rect 59 2038 66 2090
rect 0 2026 66 2038
rect 0 1974 7 2026
rect 59 1974 66 2026
rect 0 1972 16 1974
rect 50 1972 66 1974
rect 0 1962 66 1972
rect 0 1910 7 1962
rect 59 1910 66 1962
rect 0 1900 16 1910
rect 50 1900 66 1910
rect 0 1898 66 1900
rect 0 1846 7 1898
rect 59 1846 66 1898
rect 0 1834 16 1846
rect 50 1834 66 1846
rect 0 1782 7 1834
rect 59 1782 66 1834
rect 0 1770 16 1782
rect 50 1770 66 1782
rect 0 1718 7 1770
rect 59 1718 66 1770
rect 0 1706 16 1718
rect 50 1706 66 1718
rect 0 1654 7 1706
rect 59 1654 66 1706
rect 0 1646 66 1654
rect 0 1642 16 1646
rect 50 1642 66 1646
rect 0 1590 7 1642
rect 59 1590 66 1642
rect 0 1578 66 1590
rect 0 1526 7 1578
rect 59 1526 66 1578
rect 0 1514 66 1526
rect 0 1462 7 1514
rect 59 1462 66 1514
rect 0 1450 66 1462
rect 0 1398 7 1450
rect 59 1398 66 1450
rect 0 1396 16 1398
rect 50 1396 66 1398
rect 0 1386 66 1396
rect 0 1334 7 1386
rect 59 1334 66 1386
rect 0 1324 16 1334
rect 50 1324 66 1334
rect 0 1322 66 1324
rect 0 1270 7 1322
rect 59 1270 66 1322
rect 0 1252 16 1270
rect 50 1252 66 1270
rect 0 1086 66 1252
rect 0 1068 16 1086
rect 50 1068 66 1086
rect 0 1016 7 1068
rect 59 1016 66 1068
rect 0 1014 66 1016
rect 0 1004 16 1014
rect 50 1004 66 1014
rect 0 952 7 1004
rect 59 952 66 1004
rect 0 942 66 952
rect 0 940 16 942
rect 50 940 66 942
rect 0 888 7 940
rect 59 888 66 940
rect 0 876 66 888
rect 0 824 7 876
rect 59 824 66 876
rect 0 812 66 824
rect 0 760 7 812
rect 59 760 66 812
rect 0 748 66 760
rect 0 696 7 748
rect 59 696 66 748
rect 0 692 16 696
rect 50 692 66 696
rect 0 684 66 692
rect 0 632 7 684
rect 59 632 66 684
rect 0 620 16 632
rect 50 620 66 632
rect 0 568 7 620
rect 59 568 66 620
rect 0 556 16 568
rect 50 556 66 568
rect 0 504 7 556
rect 59 504 66 556
rect 0 492 16 504
rect 50 492 66 504
rect 0 440 7 492
rect 59 440 66 492
rect 0 438 66 440
rect 0 428 16 438
rect 50 428 66 438
rect 0 376 7 428
rect 59 376 66 428
rect 0 366 66 376
rect 0 364 16 366
rect 50 364 66 366
rect 0 312 7 364
rect 59 312 66 364
rect 0 300 66 312
rect 0 248 7 300
rect 59 248 66 300
rect 0 236 66 248
rect 0 184 7 236
rect 59 184 66 236
rect 0 172 66 184
rect 0 120 7 172
rect 59 120 66 172
rect 0 116 16 120
rect 50 116 66 120
rect 0 108 66 116
rect 0 56 7 108
rect 59 66 66 108
rect 100 1201 128 2244
rect 156 1229 184 2272
rect 212 1201 240 2244
rect 268 1229 296 2272
rect 324 1201 352 2244
rect 380 1229 408 2272
rect 436 1201 464 2244
rect 492 1229 520 2272
rect 548 1201 576 2244
rect 604 1229 632 2272
rect 660 1201 688 2244
rect 716 1229 744 2272
rect 772 1201 800 2244
rect 828 1229 856 2272
rect 884 1201 912 2244
rect 940 1229 968 2272
rect 996 1201 1024 2244
rect 1052 1229 1080 2272
rect 1114 2237 1168 2244
rect 1114 2185 1115 2237
rect 1167 2185 1168 2237
rect 1114 2173 1168 2185
rect 1114 2121 1115 2173
rect 1167 2121 1168 2173
rect 1114 2114 1124 2121
rect 1158 2114 1168 2121
rect 1114 2109 1168 2114
rect 1114 2057 1115 2109
rect 1167 2057 1168 2109
rect 1114 2045 1124 2057
rect 1158 2045 1168 2057
rect 1114 1993 1115 2045
rect 1167 1993 1168 2045
rect 1114 1981 1124 1993
rect 1158 1981 1168 1993
rect 1114 1929 1115 1981
rect 1167 1929 1168 1981
rect 1114 1917 1124 1929
rect 1158 1917 1168 1929
rect 1114 1865 1115 1917
rect 1167 1865 1168 1917
rect 1114 1860 1168 1865
rect 1114 1853 1124 1860
rect 1158 1853 1168 1860
rect 1114 1801 1115 1853
rect 1167 1801 1168 1853
rect 1114 1789 1168 1801
rect 1114 1737 1115 1789
rect 1167 1737 1168 1789
rect 1114 1725 1168 1737
rect 1114 1673 1115 1725
rect 1167 1673 1168 1725
rect 1114 1661 1168 1673
rect 1114 1609 1115 1661
rect 1167 1609 1168 1661
rect 1114 1597 1168 1609
rect 1114 1545 1115 1597
rect 1167 1545 1168 1597
rect 1114 1538 1124 1545
rect 1158 1538 1168 1545
rect 1114 1533 1168 1538
rect 1114 1481 1115 1533
rect 1167 1481 1168 1533
rect 1114 1469 1124 1481
rect 1158 1469 1168 1481
rect 1114 1417 1115 1469
rect 1167 1417 1168 1469
rect 1114 1405 1124 1417
rect 1158 1405 1168 1417
rect 1114 1353 1115 1405
rect 1167 1353 1168 1405
rect 1114 1341 1124 1353
rect 1158 1341 1168 1353
rect 1114 1289 1115 1341
rect 1167 1289 1168 1341
rect 1114 1284 1168 1289
rect 1114 1277 1124 1284
rect 1158 1277 1168 1284
rect 1114 1225 1115 1277
rect 1167 1225 1168 1277
rect 1202 1229 1230 2272
rect 1114 1201 1168 1225
rect 1258 1201 1286 2244
rect 1314 1229 1342 2272
rect 1370 1201 1398 2244
rect 1426 1229 1454 2272
rect 1482 1201 1510 2244
rect 1538 1229 1566 2272
rect 1594 1201 1622 2244
rect 1650 1229 1678 2272
rect 1706 1201 1734 2244
rect 1762 1229 1790 2272
rect 1818 1201 1846 2244
rect 1874 1229 1902 2272
rect 1930 1201 1958 2244
rect 1986 1229 2014 2272
rect 2042 1201 2070 2244
rect 2098 1229 2126 2272
rect 2154 1201 2182 2244
rect 100 1195 2182 1201
rect 100 1143 152 1195
rect 204 1143 216 1195
rect 268 1143 280 1195
rect 332 1143 344 1195
rect 396 1143 408 1195
rect 460 1143 472 1195
rect 524 1143 536 1195
rect 588 1143 600 1195
rect 652 1143 664 1195
rect 716 1143 728 1195
rect 780 1143 792 1195
rect 844 1143 856 1195
rect 908 1143 920 1195
rect 972 1143 984 1195
rect 1036 1143 1048 1195
rect 1100 1143 1182 1195
rect 1234 1143 1246 1195
rect 1298 1143 1310 1195
rect 1362 1143 1374 1195
rect 1426 1143 1438 1195
rect 1490 1143 1502 1195
rect 1554 1143 1566 1195
rect 1618 1143 1630 1195
rect 1682 1143 1694 1195
rect 1746 1143 1758 1195
rect 1810 1143 1822 1195
rect 1874 1143 1886 1195
rect 1938 1143 1950 1195
rect 2002 1143 2014 1195
rect 2066 1143 2078 1195
rect 2130 1143 2182 1195
rect 100 1137 2182 1143
rect 100 94 128 1137
rect 156 66 184 1109
rect 212 94 240 1137
rect 268 66 296 1109
rect 324 94 352 1137
rect 380 66 408 1109
rect 436 94 464 1137
rect 492 66 520 1109
rect 548 94 576 1137
rect 604 66 632 1109
rect 660 94 688 1137
rect 716 66 744 1109
rect 772 94 800 1137
rect 828 66 856 1109
rect 884 94 912 1137
rect 940 66 968 1109
rect 996 94 1024 1137
rect 1114 1113 1168 1137
rect 1052 66 1080 1109
rect 1114 1061 1115 1113
rect 1167 1061 1168 1113
rect 1114 1054 1124 1061
rect 1158 1054 1168 1061
rect 1114 1049 1168 1054
rect 1114 997 1115 1049
rect 1167 997 1168 1049
rect 1114 985 1124 997
rect 1158 985 1168 997
rect 1114 933 1115 985
rect 1167 933 1168 985
rect 1114 921 1124 933
rect 1158 921 1168 933
rect 1114 869 1115 921
rect 1167 869 1168 921
rect 1114 857 1124 869
rect 1158 857 1168 869
rect 1114 805 1115 857
rect 1167 805 1168 857
rect 1114 800 1168 805
rect 1114 793 1124 800
rect 1158 793 1168 800
rect 1114 741 1115 793
rect 1167 741 1168 793
rect 1114 729 1168 741
rect 1114 677 1115 729
rect 1167 677 1168 729
rect 1114 665 1168 677
rect 1114 613 1115 665
rect 1167 613 1168 665
rect 1114 601 1168 613
rect 1114 549 1115 601
rect 1167 549 1168 601
rect 1114 537 1168 549
rect 1114 485 1115 537
rect 1167 485 1168 537
rect 1114 478 1124 485
rect 1158 478 1168 485
rect 1114 473 1168 478
rect 1114 421 1115 473
rect 1167 421 1168 473
rect 1114 409 1124 421
rect 1158 409 1168 421
rect 1114 357 1115 409
rect 1167 357 1168 409
rect 1114 345 1124 357
rect 1158 345 1168 357
rect 1114 293 1115 345
rect 1167 293 1168 345
rect 1114 281 1124 293
rect 1158 281 1168 293
rect 1114 229 1115 281
rect 1167 229 1168 281
rect 1114 224 1168 229
rect 1114 217 1124 224
rect 1158 217 1168 224
rect 1114 165 1115 217
rect 1167 165 1168 217
rect 1114 153 1168 165
rect 1114 101 1115 153
rect 1167 101 1168 153
rect 1114 94 1168 101
rect 1202 66 1230 1109
rect 1258 94 1286 1137
rect 1314 66 1342 1109
rect 1370 94 1398 1137
rect 1426 66 1454 1109
rect 1482 94 1510 1137
rect 1538 66 1566 1109
rect 1594 94 1622 1137
rect 1650 66 1678 1109
rect 1706 94 1734 1137
rect 1762 66 1790 1109
rect 1818 94 1846 1137
rect 1874 66 1902 1109
rect 1930 94 1958 1137
rect 1986 66 2014 1109
rect 2042 94 2070 1137
rect 2098 66 2126 1109
rect 2154 94 2182 1137
rect 2216 2230 2223 2272
rect 2275 2230 2282 2282
rect 2216 2222 2282 2230
rect 2216 2218 2232 2222
rect 2266 2218 2282 2222
rect 2216 2166 2223 2218
rect 2275 2166 2282 2218
rect 2216 2154 2282 2166
rect 2216 2102 2223 2154
rect 2275 2102 2282 2154
rect 2216 2090 2282 2102
rect 2216 2038 2223 2090
rect 2275 2038 2282 2090
rect 2216 2026 2282 2038
rect 2216 1974 2223 2026
rect 2275 1974 2282 2026
rect 2216 1972 2232 1974
rect 2266 1972 2282 1974
rect 2216 1962 2282 1972
rect 2216 1910 2223 1962
rect 2275 1910 2282 1962
rect 2216 1900 2232 1910
rect 2266 1900 2282 1910
rect 2216 1898 2282 1900
rect 2216 1846 2223 1898
rect 2275 1846 2282 1898
rect 2216 1834 2232 1846
rect 2266 1834 2282 1846
rect 2216 1782 2223 1834
rect 2275 1782 2282 1834
rect 2216 1770 2232 1782
rect 2266 1770 2282 1782
rect 2216 1718 2223 1770
rect 2275 1718 2282 1770
rect 2216 1706 2232 1718
rect 2266 1706 2282 1718
rect 2216 1654 2223 1706
rect 2275 1654 2282 1706
rect 2216 1646 2282 1654
rect 2216 1642 2232 1646
rect 2266 1642 2282 1646
rect 2216 1590 2223 1642
rect 2275 1590 2282 1642
rect 2216 1578 2282 1590
rect 2216 1526 2223 1578
rect 2275 1526 2282 1578
rect 2216 1514 2282 1526
rect 2216 1462 2223 1514
rect 2275 1462 2282 1514
rect 2216 1450 2282 1462
rect 2216 1398 2223 1450
rect 2275 1398 2282 1450
rect 2216 1396 2232 1398
rect 2266 1396 2282 1398
rect 2216 1386 2282 1396
rect 2216 1334 2223 1386
rect 2275 1334 2282 1386
rect 2216 1324 2232 1334
rect 2266 1324 2282 1334
rect 2216 1322 2282 1324
rect 2216 1270 2223 1322
rect 2275 1270 2282 1322
rect 2216 1252 2232 1270
rect 2266 1252 2282 1270
rect 2216 1086 2282 1252
rect 2216 1068 2232 1086
rect 2266 1068 2282 1086
rect 2216 1016 2223 1068
rect 2275 1016 2282 1068
rect 2216 1014 2282 1016
rect 2216 1004 2232 1014
rect 2266 1004 2282 1014
rect 2216 952 2223 1004
rect 2275 952 2282 1004
rect 2216 942 2282 952
rect 2216 940 2232 942
rect 2266 940 2282 942
rect 2216 888 2223 940
rect 2275 888 2282 940
rect 2216 876 2282 888
rect 2216 824 2223 876
rect 2275 824 2282 876
rect 2216 812 2282 824
rect 2216 760 2223 812
rect 2275 760 2282 812
rect 2216 748 2282 760
rect 2216 696 2223 748
rect 2275 696 2282 748
rect 2216 692 2232 696
rect 2266 692 2282 696
rect 2216 684 2282 692
rect 2216 632 2223 684
rect 2275 632 2282 684
rect 2216 620 2232 632
rect 2266 620 2282 632
rect 2216 568 2223 620
rect 2275 568 2282 620
rect 2216 556 2232 568
rect 2266 556 2282 568
rect 2216 504 2223 556
rect 2275 504 2282 556
rect 2216 492 2232 504
rect 2266 492 2282 504
rect 2216 440 2223 492
rect 2275 440 2282 492
rect 2216 438 2282 440
rect 2216 428 2232 438
rect 2266 428 2282 438
rect 2216 376 2223 428
rect 2275 376 2282 428
rect 2216 366 2282 376
rect 2216 364 2232 366
rect 2266 364 2282 366
rect 2216 312 2223 364
rect 2275 312 2282 364
rect 2216 300 2282 312
rect 2216 248 2223 300
rect 2275 248 2282 300
rect 2216 236 2282 248
rect 2216 184 2223 236
rect 2275 184 2282 236
rect 2216 172 2282 184
rect 2216 120 2223 172
rect 2275 120 2282 172
rect 2216 116 2232 120
rect 2266 116 2282 120
rect 2216 108 2282 116
rect 2216 66 2223 108
rect 59 59 2223 66
rect 59 56 88 59
rect 0 50 88 56
rect 0 16 80 50
rect 0 7 88 16
rect 140 7 152 59
rect 204 7 216 59
rect 268 7 280 59
rect 332 7 344 59
rect 396 50 408 59
rect 460 50 472 59
rect 524 50 536 59
rect 588 50 600 59
rect 652 50 664 59
rect 402 16 408 50
rect 652 16 656 50
rect 396 7 408 16
rect 460 7 472 16
rect 524 7 536 16
rect 588 7 600 16
rect 652 7 664 16
rect 716 7 728 59
rect 780 7 792 59
rect 844 7 856 59
rect 908 7 920 59
rect 972 50 984 59
rect 1036 50 1246 59
rect 1298 50 1310 59
rect 978 16 984 50
rect 1050 16 1088 50
rect 1122 16 1160 50
rect 1194 16 1232 50
rect 1298 16 1304 50
rect 972 7 984 16
rect 1036 7 1246 16
rect 1298 7 1310 16
rect 1362 7 1374 59
rect 1426 7 1438 59
rect 1490 7 1502 59
rect 1554 7 1566 59
rect 1618 50 1630 59
rect 1682 50 1694 59
rect 1746 50 1758 59
rect 1810 50 1822 59
rect 1874 50 1886 59
rect 1626 16 1630 50
rect 1874 16 1880 50
rect 1618 7 1630 16
rect 1682 7 1694 16
rect 1746 7 1758 16
rect 1810 7 1822 16
rect 1874 7 1886 16
rect 1938 7 1950 59
rect 2002 7 2014 59
rect 2066 7 2078 59
rect 2130 7 2142 59
rect 2194 56 2223 59
rect 2275 56 2282 108
rect 2194 50 2282 56
rect 2202 16 2282 50
rect 2194 7 2282 16
rect 0 0 2282 7
<< via1 >>
rect 88 2322 140 2331
rect 88 2288 114 2322
rect 114 2288 140 2322
rect 7 2230 59 2282
rect 88 2279 140 2288
rect 152 2322 204 2331
rect 152 2288 186 2322
rect 186 2288 204 2322
rect 152 2279 204 2288
rect 216 2322 268 2331
rect 216 2288 224 2322
rect 224 2288 258 2322
rect 258 2288 268 2322
rect 216 2279 268 2288
rect 280 2322 332 2331
rect 280 2288 296 2322
rect 296 2288 330 2322
rect 330 2288 332 2322
rect 280 2279 332 2288
rect 344 2322 396 2331
rect 408 2322 460 2331
rect 472 2322 524 2331
rect 536 2322 588 2331
rect 600 2322 652 2331
rect 664 2322 716 2331
rect 344 2288 368 2322
rect 368 2288 396 2322
rect 408 2288 440 2322
rect 440 2288 460 2322
rect 472 2288 474 2322
rect 474 2288 512 2322
rect 512 2288 524 2322
rect 536 2288 546 2322
rect 546 2288 584 2322
rect 584 2288 588 2322
rect 600 2288 618 2322
rect 618 2288 652 2322
rect 664 2288 690 2322
rect 690 2288 716 2322
rect 344 2279 396 2288
rect 408 2279 460 2288
rect 472 2279 524 2288
rect 536 2279 588 2288
rect 600 2279 652 2288
rect 664 2279 716 2288
rect 728 2322 780 2331
rect 728 2288 762 2322
rect 762 2288 780 2322
rect 728 2279 780 2288
rect 792 2322 844 2331
rect 792 2288 800 2322
rect 800 2288 834 2322
rect 834 2288 844 2322
rect 792 2279 844 2288
rect 856 2322 908 2331
rect 856 2288 872 2322
rect 872 2288 906 2322
rect 906 2288 908 2322
rect 856 2279 908 2288
rect 920 2322 972 2331
rect 984 2322 1036 2331
rect 1246 2322 1298 2331
rect 1310 2322 1362 2331
rect 920 2288 944 2322
rect 944 2288 972 2322
rect 984 2288 1016 2322
rect 1016 2288 1036 2322
rect 1246 2288 1266 2322
rect 1266 2288 1298 2322
rect 1310 2288 1338 2322
rect 1338 2288 1362 2322
rect 920 2279 972 2288
rect 984 2279 1036 2288
rect 1246 2279 1298 2288
rect 1310 2279 1362 2288
rect 1374 2322 1426 2331
rect 1374 2288 1376 2322
rect 1376 2288 1410 2322
rect 1410 2288 1426 2322
rect 1374 2279 1426 2288
rect 1438 2322 1490 2331
rect 1438 2288 1448 2322
rect 1448 2288 1482 2322
rect 1482 2288 1490 2322
rect 1438 2279 1490 2288
rect 1502 2322 1554 2331
rect 1502 2288 1520 2322
rect 1520 2288 1554 2322
rect 1502 2279 1554 2288
rect 1566 2322 1618 2331
rect 1630 2322 1682 2331
rect 1694 2322 1746 2331
rect 1758 2322 1810 2331
rect 1822 2322 1874 2331
rect 1886 2322 1938 2331
rect 1566 2288 1592 2322
rect 1592 2288 1618 2322
rect 1630 2288 1664 2322
rect 1664 2288 1682 2322
rect 1694 2288 1698 2322
rect 1698 2288 1736 2322
rect 1736 2288 1746 2322
rect 1758 2288 1770 2322
rect 1770 2288 1808 2322
rect 1808 2288 1810 2322
rect 1822 2288 1842 2322
rect 1842 2288 1874 2322
rect 1886 2288 1914 2322
rect 1914 2288 1938 2322
rect 1566 2279 1618 2288
rect 1630 2279 1682 2288
rect 1694 2279 1746 2288
rect 1758 2279 1810 2288
rect 1822 2279 1874 2288
rect 1886 2279 1938 2288
rect 1950 2322 2002 2331
rect 1950 2288 1952 2322
rect 1952 2288 1986 2322
rect 1986 2288 2002 2322
rect 1950 2279 2002 2288
rect 2014 2322 2066 2331
rect 2014 2288 2024 2322
rect 2024 2288 2058 2322
rect 2058 2288 2066 2322
rect 2014 2279 2066 2288
rect 2078 2322 2130 2331
rect 2078 2288 2096 2322
rect 2096 2288 2130 2322
rect 2078 2279 2130 2288
rect 2142 2322 2194 2331
rect 2142 2288 2168 2322
rect 2168 2288 2194 2322
rect 2142 2279 2194 2288
rect 7 2188 16 2218
rect 16 2188 50 2218
rect 50 2188 59 2218
rect 7 2166 59 2188
rect 7 2150 59 2154
rect 7 2116 16 2150
rect 16 2116 50 2150
rect 50 2116 59 2150
rect 7 2102 59 2116
rect 7 2078 59 2090
rect 7 2044 16 2078
rect 16 2044 50 2078
rect 50 2044 59 2078
rect 7 2038 59 2044
rect 7 2006 59 2026
rect 7 1974 16 2006
rect 16 1974 50 2006
rect 50 1974 59 2006
rect 7 1934 59 1962
rect 7 1910 16 1934
rect 16 1910 50 1934
rect 50 1910 59 1934
rect 7 1862 59 1898
rect 7 1846 16 1862
rect 16 1846 50 1862
rect 50 1846 59 1862
rect 7 1828 16 1834
rect 16 1828 50 1834
rect 50 1828 59 1834
rect 7 1790 59 1828
rect 7 1782 16 1790
rect 16 1782 50 1790
rect 50 1782 59 1790
rect 7 1756 16 1770
rect 16 1756 50 1770
rect 50 1756 59 1770
rect 7 1718 59 1756
rect 7 1684 16 1706
rect 16 1684 50 1706
rect 50 1684 59 1706
rect 7 1654 59 1684
rect 7 1612 16 1642
rect 16 1612 50 1642
rect 50 1612 59 1642
rect 7 1590 59 1612
rect 7 1574 59 1578
rect 7 1540 16 1574
rect 16 1540 50 1574
rect 50 1540 59 1574
rect 7 1526 59 1540
rect 7 1502 59 1514
rect 7 1468 16 1502
rect 16 1468 50 1502
rect 50 1468 59 1502
rect 7 1462 59 1468
rect 7 1430 59 1450
rect 7 1398 16 1430
rect 16 1398 50 1430
rect 50 1398 59 1430
rect 7 1358 59 1386
rect 7 1334 16 1358
rect 16 1334 50 1358
rect 50 1334 59 1358
rect 7 1286 59 1322
rect 7 1270 16 1286
rect 16 1270 50 1286
rect 50 1270 59 1286
rect 7 1052 16 1068
rect 16 1052 50 1068
rect 50 1052 59 1068
rect 7 1016 59 1052
rect 7 980 16 1004
rect 16 980 50 1004
rect 50 980 59 1004
rect 7 952 59 980
rect 7 908 16 940
rect 16 908 50 940
rect 50 908 59 940
rect 7 888 59 908
rect 7 870 59 876
rect 7 836 16 870
rect 16 836 50 870
rect 50 836 59 870
rect 7 824 59 836
rect 7 798 59 812
rect 7 764 16 798
rect 16 764 50 798
rect 50 764 59 798
rect 7 760 59 764
rect 7 726 59 748
rect 7 696 16 726
rect 16 696 50 726
rect 50 696 59 726
rect 7 654 59 684
rect 7 632 16 654
rect 16 632 50 654
rect 50 632 59 654
rect 7 582 59 620
rect 7 568 16 582
rect 16 568 50 582
rect 50 568 59 582
rect 7 548 16 556
rect 16 548 50 556
rect 50 548 59 556
rect 7 510 59 548
rect 7 504 16 510
rect 16 504 50 510
rect 50 504 59 510
rect 7 476 16 492
rect 16 476 50 492
rect 50 476 59 492
rect 7 440 59 476
rect 7 404 16 428
rect 16 404 50 428
rect 50 404 59 428
rect 7 376 59 404
rect 7 332 16 364
rect 16 332 50 364
rect 50 332 59 364
rect 7 312 59 332
rect 7 294 59 300
rect 7 260 16 294
rect 16 260 50 294
rect 50 260 59 294
rect 7 248 59 260
rect 7 222 59 236
rect 7 188 16 222
rect 16 188 50 222
rect 50 188 59 222
rect 7 184 59 188
rect 7 150 59 172
rect 7 120 16 150
rect 16 120 50 150
rect 50 120 59 150
rect 7 56 59 108
rect 1115 2220 1167 2237
rect 1115 2186 1124 2220
rect 1124 2186 1158 2220
rect 1158 2186 1167 2220
rect 1115 2185 1167 2186
rect 1115 2148 1167 2173
rect 1115 2121 1124 2148
rect 1124 2121 1158 2148
rect 1158 2121 1167 2148
rect 1115 2076 1167 2109
rect 1115 2057 1124 2076
rect 1124 2057 1158 2076
rect 1158 2057 1167 2076
rect 1115 2042 1124 2045
rect 1124 2042 1158 2045
rect 1158 2042 1167 2045
rect 1115 2004 1167 2042
rect 1115 1993 1124 2004
rect 1124 1993 1158 2004
rect 1158 1993 1167 2004
rect 1115 1970 1124 1981
rect 1124 1970 1158 1981
rect 1158 1970 1167 1981
rect 1115 1932 1167 1970
rect 1115 1929 1124 1932
rect 1124 1929 1158 1932
rect 1158 1929 1167 1932
rect 1115 1898 1124 1917
rect 1124 1898 1158 1917
rect 1158 1898 1167 1917
rect 1115 1865 1167 1898
rect 1115 1826 1124 1853
rect 1124 1826 1158 1853
rect 1158 1826 1167 1853
rect 1115 1801 1167 1826
rect 1115 1788 1167 1789
rect 1115 1754 1124 1788
rect 1124 1754 1158 1788
rect 1158 1754 1167 1788
rect 1115 1737 1167 1754
rect 1115 1716 1167 1725
rect 1115 1682 1124 1716
rect 1124 1682 1158 1716
rect 1158 1682 1167 1716
rect 1115 1673 1167 1682
rect 1115 1644 1167 1661
rect 1115 1610 1124 1644
rect 1124 1610 1158 1644
rect 1158 1610 1167 1644
rect 1115 1609 1167 1610
rect 1115 1572 1167 1597
rect 1115 1545 1124 1572
rect 1124 1545 1158 1572
rect 1158 1545 1167 1572
rect 1115 1500 1167 1533
rect 1115 1481 1124 1500
rect 1124 1481 1158 1500
rect 1158 1481 1167 1500
rect 1115 1466 1124 1469
rect 1124 1466 1158 1469
rect 1158 1466 1167 1469
rect 1115 1428 1167 1466
rect 1115 1417 1124 1428
rect 1124 1417 1158 1428
rect 1158 1417 1167 1428
rect 1115 1394 1124 1405
rect 1124 1394 1158 1405
rect 1158 1394 1167 1405
rect 1115 1356 1167 1394
rect 1115 1353 1124 1356
rect 1124 1353 1158 1356
rect 1158 1353 1167 1356
rect 1115 1322 1124 1341
rect 1124 1322 1158 1341
rect 1158 1322 1167 1341
rect 1115 1289 1167 1322
rect 1115 1250 1124 1277
rect 1124 1250 1158 1277
rect 1158 1250 1167 1277
rect 1115 1225 1167 1250
rect 152 1143 204 1195
rect 216 1143 268 1195
rect 280 1143 332 1195
rect 344 1143 396 1195
rect 408 1143 460 1195
rect 472 1143 524 1195
rect 536 1143 588 1195
rect 600 1143 652 1195
rect 664 1143 716 1195
rect 728 1143 780 1195
rect 792 1143 844 1195
rect 856 1143 908 1195
rect 920 1143 972 1195
rect 984 1143 1036 1195
rect 1048 1143 1100 1195
rect 1182 1143 1234 1195
rect 1246 1143 1298 1195
rect 1310 1143 1362 1195
rect 1374 1143 1426 1195
rect 1438 1143 1490 1195
rect 1502 1143 1554 1195
rect 1566 1143 1618 1195
rect 1630 1143 1682 1195
rect 1694 1143 1746 1195
rect 1758 1143 1810 1195
rect 1822 1143 1874 1195
rect 1886 1143 1938 1195
rect 1950 1143 2002 1195
rect 2014 1143 2066 1195
rect 2078 1143 2130 1195
rect 1115 1088 1167 1113
rect 1115 1061 1124 1088
rect 1124 1061 1158 1088
rect 1158 1061 1167 1088
rect 1115 1016 1167 1049
rect 1115 997 1124 1016
rect 1124 997 1158 1016
rect 1158 997 1167 1016
rect 1115 982 1124 985
rect 1124 982 1158 985
rect 1158 982 1167 985
rect 1115 944 1167 982
rect 1115 933 1124 944
rect 1124 933 1158 944
rect 1158 933 1167 944
rect 1115 910 1124 921
rect 1124 910 1158 921
rect 1158 910 1167 921
rect 1115 872 1167 910
rect 1115 869 1124 872
rect 1124 869 1158 872
rect 1158 869 1167 872
rect 1115 838 1124 857
rect 1124 838 1158 857
rect 1158 838 1167 857
rect 1115 805 1167 838
rect 1115 766 1124 793
rect 1124 766 1158 793
rect 1158 766 1167 793
rect 1115 741 1167 766
rect 1115 728 1167 729
rect 1115 694 1124 728
rect 1124 694 1158 728
rect 1158 694 1167 728
rect 1115 677 1167 694
rect 1115 656 1167 665
rect 1115 622 1124 656
rect 1124 622 1158 656
rect 1158 622 1167 656
rect 1115 613 1167 622
rect 1115 584 1167 601
rect 1115 550 1124 584
rect 1124 550 1158 584
rect 1158 550 1167 584
rect 1115 549 1167 550
rect 1115 512 1167 537
rect 1115 485 1124 512
rect 1124 485 1158 512
rect 1158 485 1167 512
rect 1115 440 1167 473
rect 1115 421 1124 440
rect 1124 421 1158 440
rect 1158 421 1167 440
rect 1115 406 1124 409
rect 1124 406 1158 409
rect 1158 406 1167 409
rect 1115 368 1167 406
rect 1115 357 1124 368
rect 1124 357 1158 368
rect 1158 357 1167 368
rect 1115 334 1124 345
rect 1124 334 1158 345
rect 1158 334 1167 345
rect 1115 296 1167 334
rect 1115 293 1124 296
rect 1124 293 1158 296
rect 1158 293 1167 296
rect 1115 262 1124 281
rect 1124 262 1158 281
rect 1158 262 1167 281
rect 1115 229 1167 262
rect 1115 190 1124 217
rect 1124 190 1158 217
rect 1158 190 1167 217
rect 1115 165 1167 190
rect 1115 152 1167 153
rect 1115 118 1124 152
rect 1124 118 1158 152
rect 1158 118 1167 152
rect 1115 101 1167 118
rect 2223 2230 2275 2282
rect 2223 2188 2232 2218
rect 2232 2188 2266 2218
rect 2266 2188 2275 2218
rect 2223 2166 2275 2188
rect 2223 2150 2275 2154
rect 2223 2116 2232 2150
rect 2232 2116 2266 2150
rect 2266 2116 2275 2150
rect 2223 2102 2275 2116
rect 2223 2078 2275 2090
rect 2223 2044 2232 2078
rect 2232 2044 2266 2078
rect 2266 2044 2275 2078
rect 2223 2038 2275 2044
rect 2223 2006 2275 2026
rect 2223 1974 2232 2006
rect 2232 1974 2266 2006
rect 2266 1974 2275 2006
rect 2223 1934 2275 1962
rect 2223 1910 2232 1934
rect 2232 1910 2266 1934
rect 2266 1910 2275 1934
rect 2223 1862 2275 1898
rect 2223 1846 2232 1862
rect 2232 1846 2266 1862
rect 2266 1846 2275 1862
rect 2223 1828 2232 1834
rect 2232 1828 2266 1834
rect 2266 1828 2275 1834
rect 2223 1790 2275 1828
rect 2223 1782 2232 1790
rect 2232 1782 2266 1790
rect 2266 1782 2275 1790
rect 2223 1756 2232 1770
rect 2232 1756 2266 1770
rect 2266 1756 2275 1770
rect 2223 1718 2275 1756
rect 2223 1684 2232 1706
rect 2232 1684 2266 1706
rect 2266 1684 2275 1706
rect 2223 1654 2275 1684
rect 2223 1612 2232 1642
rect 2232 1612 2266 1642
rect 2266 1612 2275 1642
rect 2223 1590 2275 1612
rect 2223 1574 2275 1578
rect 2223 1540 2232 1574
rect 2232 1540 2266 1574
rect 2266 1540 2275 1574
rect 2223 1526 2275 1540
rect 2223 1502 2275 1514
rect 2223 1468 2232 1502
rect 2232 1468 2266 1502
rect 2266 1468 2275 1502
rect 2223 1462 2275 1468
rect 2223 1430 2275 1450
rect 2223 1398 2232 1430
rect 2232 1398 2266 1430
rect 2266 1398 2275 1430
rect 2223 1358 2275 1386
rect 2223 1334 2232 1358
rect 2232 1334 2266 1358
rect 2266 1334 2275 1358
rect 2223 1286 2275 1322
rect 2223 1270 2232 1286
rect 2232 1270 2266 1286
rect 2266 1270 2275 1286
rect 2223 1052 2232 1068
rect 2232 1052 2266 1068
rect 2266 1052 2275 1068
rect 2223 1016 2275 1052
rect 2223 980 2232 1004
rect 2232 980 2266 1004
rect 2266 980 2275 1004
rect 2223 952 2275 980
rect 2223 908 2232 940
rect 2232 908 2266 940
rect 2266 908 2275 940
rect 2223 888 2275 908
rect 2223 870 2275 876
rect 2223 836 2232 870
rect 2232 836 2266 870
rect 2266 836 2275 870
rect 2223 824 2275 836
rect 2223 798 2275 812
rect 2223 764 2232 798
rect 2232 764 2266 798
rect 2266 764 2275 798
rect 2223 760 2275 764
rect 2223 726 2275 748
rect 2223 696 2232 726
rect 2232 696 2266 726
rect 2266 696 2275 726
rect 2223 654 2275 684
rect 2223 632 2232 654
rect 2232 632 2266 654
rect 2266 632 2275 654
rect 2223 582 2275 620
rect 2223 568 2232 582
rect 2232 568 2266 582
rect 2266 568 2275 582
rect 2223 548 2232 556
rect 2232 548 2266 556
rect 2266 548 2275 556
rect 2223 510 2275 548
rect 2223 504 2232 510
rect 2232 504 2266 510
rect 2266 504 2275 510
rect 2223 476 2232 492
rect 2232 476 2266 492
rect 2266 476 2275 492
rect 2223 440 2275 476
rect 2223 404 2232 428
rect 2232 404 2266 428
rect 2266 404 2275 428
rect 2223 376 2275 404
rect 2223 332 2232 364
rect 2232 332 2266 364
rect 2266 332 2275 364
rect 2223 312 2275 332
rect 2223 294 2275 300
rect 2223 260 2232 294
rect 2232 260 2266 294
rect 2266 260 2275 294
rect 2223 248 2275 260
rect 2223 222 2275 236
rect 2223 188 2232 222
rect 2232 188 2266 222
rect 2266 188 2275 222
rect 2223 184 2275 188
rect 2223 150 2275 172
rect 2223 120 2232 150
rect 2232 120 2266 150
rect 2266 120 2275 150
rect 88 50 140 59
rect 88 16 114 50
rect 114 16 140 50
rect 88 7 140 16
rect 152 50 204 59
rect 152 16 186 50
rect 186 16 204 50
rect 152 7 204 16
rect 216 50 268 59
rect 216 16 224 50
rect 224 16 258 50
rect 258 16 268 50
rect 216 7 268 16
rect 280 50 332 59
rect 280 16 296 50
rect 296 16 330 50
rect 330 16 332 50
rect 280 7 332 16
rect 344 50 396 59
rect 408 50 460 59
rect 472 50 524 59
rect 536 50 588 59
rect 600 50 652 59
rect 664 50 716 59
rect 344 16 368 50
rect 368 16 396 50
rect 408 16 440 50
rect 440 16 460 50
rect 472 16 474 50
rect 474 16 512 50
rect 512 16 524 50
rect 536 16 546 50
rect 546 16 584 50
rect 584 16 588 50
rect 600 16 618 50
rect 618 16 652 50
rect 664 16 690 50
rect 690 16 716 50
rect 344 7 396 16
rect 408 7 460 16
rect 472 7 524 16
rect 536 7 588 16
rect 600 7 652 16
rect 664 7 716 16
rect 728 50 780 59
rect 728 16 762 50
rect 762 16 780 50
rect 728 7 780 16
rect 792 50 844 59
rect 792 16 800 50
rect 800 16 834 50
rect 834 16 844 50
rect 792 7 844 16
rect 856 50 908 59
rect 856 16 872 50
rect 872 16 906 50
rect 906 16 908 50
rect 856 7 908 16
rect 920 50 972 59
rect 984 50 1036 59
rect 1246 50 1298 59
rect 1310 50 1362 59
rect 920 16 944 50
rect 944 16 972 50
rect 984 16 1016 50
rect 1016 16 1036 50
rect 1246 16 1266 50
rect 1266 16 1298 50
rect 1310 16 1338 50
rect 1338 16 1362 50
rect 920 7 972 16
rect 984 7 1036 16
rect 1246 7 1298 16
rect 1310 7 1362 16
rect 1374 50 1426 59
rect 1374 16 1376 50
rect 1376 16 1410 50
rect 1410 16 1426 50
rect 1374 7 1426 16
rect 1438 50 1490 59
rect 1438 16 1448 50
rect 1448 16 1482 50
rect 1482 16 1490 50
rect 1438 7 1490 16
rect 1502 50 1554 59
rect 1502 16 1520 50
rect 1520 16 1554 50
rect 1502 7 1554 16
rect 1566 50 1618 59
rect 1630 50 1682 59
rect 1694 50 1746 59
rect 1758 50 1810 59
rect 1822 50 1874 59
rect 1886 50 1938 59
rect 1566 16 1592 50
rect 1592 16 1618 50
rect 1630 16 1664 50
rect 1664 16 1682 50
rect 1694 16 1698 50
rect 1698 16 1736 50
rect 1736 16 1746 50
rect 1758 16 1770 50
rect 1770 16 1808 50
rect 1808 16 1810 50
rect 1822 16 1842 50
rect 1842 16 1874 50
rect 1886 16 1914 50
rect 1914 16 1938 50
rect 1566 7 1618 16
rect 1630 7 1682 16
rect 1694 7 1746 16
rect 1758 7 1810 16
rect 1822 7 1874 16
rect 1886 7 1938 16
rect 1950 50 2002 59
rect 1950 16 1952 50
rect 1952 16 1986 50
rect 1986 16 2002 50
rect 1950 7 2002 16
rect 2014 50 2066 59
rect 2014 16 2024 50
rect 2024 16 2058 50
rect 2058 16 2066 50
rect 2014 7 2066 16
rect 2078 50 2130 59
rect 2078 16 2096 50
rect 2096 16 2130 50
rect 2078 7 2130 16
rect 2142 50 2194 59
rect 2223 56 2275 108
rect 2142 16 2168 50
rect 2168 16 2194 50
rect 2142 7 2194 16
<< metal2 >>
rect 0 2333 1086 2338
rect 0 2282 61 2333
rect 117 2331 141 2333
rect 197 2331 221 2333
rect 277 2331 301 2333
rect 357 2331 381 2333
rect 437 2331 461 2333
rect 517 2331 541 2333
rect 597 2331 621 2333
rect 677 2331 701 2333
rect 757 2331 781 2333
rect 837 2331 861 2333
rect 917 2331 941 2333
rect 997 2331 1021 2333
rect 0 2249 7 2282
rect 59 2277 61 2282
rect 140 2279 141 2331
rect 204 2279 216 2331
rect 277 2279 280 2331
rect 460 2279 461 2331
rect 524 2279 536 2331
rect 597 2279 600 2331
rect 780 2279 781 2331
rect 844 2279 856 2331
rect 917 2279 920 2331
rect 117 2277 141 2279
rect 197 2277 221 2279
rect 277 2277 301 2279
rect 357 2277 381 2279
rect 437 2277 461 2279
rect 517 2277 541 2279
rect 597 2277 621 2279
rect 677 2277 701 2279
rect 757 2277 781 2279
rect 837 2277 861 2279
rect 917 2277 941 2279
rect 997 2277 1021 2279
rect 1077 2277 1086 2333
rect 59 2272 1086 2277
rect 59 2249 66 2272
rect 0 2193 5 2249
rect 61 2193 66 2249
rect 1114 2244 1168 2338
rect 1196 2333 2282 2338
rect 1196 2277 1205 2333
rect 1261 2331 1285 2333
rect 1341 2331 1365 2333
rect 1421 2331 1445 2333
rect 1501 2331 1525 2333
rect 1581 2331 1605 2333
rect 1661 2331 1685 2333
rect 1741 2331 1765 2333
rect 1821 2331 1845 2333
rect 1901 2331 1925 2333
rect 1981 2331 2005 2333
rect 2061 2331 2085 2333
rect 2141 2331 2165 2333
rect 1362 2279 1365 2331
rect 1426 2279 1438 2331
rect 1501 2279 1502 2331
rect 1682 2279 1685 2331
rect 1746 2279 1758 2331
rect 1821 2279 1822 2331
rect 2002 2279 2005 2331
rect 2066 2279 2078 2331
rect 2141 2279 2142 2331
rect 2221 2282 2282 2333
rect 1261 2277 1285 2279
rect 1341 2277 1365 2279
rect 1421 2277 1445 2279
rect 1501 2277 1525 2279
rect 1581 2277 1605 2279
rect 1661 2277 1685 2279
rect 1741 2277 1765 2279
rect 1821 2277 1845 2279
rect 1901 2277 1925 2279
rect 1981 2277 2005 2279
rect 2061 2277 2085 2279
rect 2141 2277 2165 2279
rect 2221 2277 2223 2282
rect 1196 2272 2223 2277
rect 2216 2249 2223 2272
rect 2275 2249 2282 2282
rect 94 2237 2188 2244
rect 94 2216 1115 2237
rect 0 2169 7 2193
rect 59 2188 66 2193
rect 59 2169 1085 2188
rect 0 2113 5 2169
rect 61 2160 1085 2169
rect 1113 2185 1115 2216
rect 1167 2216 2188 2237
rect 1167 2185 1169 2216
rect 2216 2193 2221 2249
rect 2277 2193 2282 2249
rect 2216 2188 2223 2193
rect 1113 2173 1169 2185
rect 61 2113 66 2160
rect 1113 2157 1115 2173
rect 1167 2157 1169 2173
rect 1197 2169 2223 2188
rect 2275 2169 2282 2193
rect 1197 2160 2221 2169
rect 0 2102 7 2113
rect 59 2102 66 2113
rect 94 2104 1113 2132
rect 0 2090 66 2102
rect 0 2089 7 2090
rect 59 2089 66 2090
rect 0 2033 5 2089
rect 61 2076 66 2089
rect 1169 2104 2188 2132
rect 2216 2113 2221 2160
rect 2277 2113 2282 2169
rect 1113 2077 1115 2101
rect 1167 2077 1169 2101
rect 61 2048 1085 2076
rect 2216 2102 2223 2113
rect 2275 2102 2282 2113
rect 2216 2090 2282 2102
rect 2216 2089 2223 2090
rect 2275 2089 2282 2090
rect 2216 2076 2221 2089
rect 61 2033 66 2048
rect 0 2026 66 2033
rect 0 2009 7 2026
rect 59 2009 66 2026
rect 1197 2048 2221 2076
rect 1113 2020 1115 2021
rect 0 1953 5 2009
rect 61 1964 66 2009
rect 94 1997 1115 2020
rect 1167 2020 1169 2021
rect 2216 2033 2221 2048
rect 2277 2033 2282 2089
rect 2216 2026 2282 2033
rect 1167 1997 2188 2020
rect 94 1992 1113 1997
rect 1169 1992 2188 1997
rect 2216 2009 2223 2026
rect 2275 2009 2282 2026
rect 61 1953 1085 1964
rect 0 1929 7 1953
rect 59 1936 1085 1953
rect 2216 1964 2221 2009
rect 59 1929 66 1936
rect 0 1873 5 1929
rect 61 1873 66 1929
rect 1113 1929 1115 1941
rect 1167 1929 1169 1941
rect 1197 1953 2221 1964
rect 2277 1953 2282 2009
rect 1197 1936 2223 1953
rect 1113 1917 1169 1929
rect 94 1880 1113 1908
rect 0 1849 7 1873
rect 59 1852 66 1873
rect 2216 1929 2223 1936
rect 2275 1929 2282 1953
rect 1169 1880 2188 1908
rect 1113 1853 1169 1861
rect 59 1849 1085 1852
rect 0 1793 5 1849
rect 61 1824 1085 1849
rect 1113 1837 1115 1853
rect 1167 1837 1169 1853
rect 2216 1873 2221 1929
rect 2277 1873 2282 1929
rect 2216 1852 2223 1873
rect 61 1793 66 1824
rect 1197 1849 2223 1852
rect 2275 1849 2282 1873
rect 1197 1824 2221 1849
rect 0 1782 7 1793
rect 59 1782 66 1793
rect 0 1770 66 1782
rect 0 1769 7 1770
rect 59 1769 66 1770
rect 0 1713 5 1769
rect 61 1740 66 1769
rect 94 1781 1113 1796
rect 1169 1781 2188 1796
rect 94 1768 1115 1781
rect 1113 1757 1115 1768
rect 1167 1768 2188 1781
rect 2216 1793 2221 1824
rect 2277 1793 2282 1849
rect 2216 1782 2223 1793
rect 2275 1782 2282 1793
rect 2216 1770 2282 1782
rect 2216 1769 2223 1770
rect 2275 1769 2282 1770
rect 1167 1757 1169 1768
rect 61 1713 1085 1740
rect 0 1712 1085 1713
rect 2216 1740 2221 1769
rect 0 1706 66 1712
rect 0 1689 7 1706
rect 59 1689 66 1706
rect 0 1633 5 1689
rect 61 1633 66 1689
rect 1197 1713 2221 1740
rect 2277 1713 2282 1769
rect 1197 1712 2282 1713
rect 1113 1684 1115 1701
rect 94 1677 1115 1684
rect 1167 1684 1169 1701
rect 2216 1706 2282 1712
rect 2216 1689 2223 1706
rect 2275 1689 2282 1706
rect 1167 1677 2188 1684
rect 94 1656 1113 1677
rect 0 1609 7 1633
rect 59 1628 66 1633
rect 59 1609 1085 1628
rect 0 1553 5 1609
rect 61 1600 1085 1609
rect 1169 1656 2188 1677
rect 2216 1633 2221 1689
rect 2277 1633 2282 1689
rect 2216 1628 2223 1633
rect 1113 1609 1115 1621
rect 1167 1609 1169 1621
rect 61 1553 66 1600
rect 1113 1597 1169 1609
rect 1197 1609 2223 1628
rect 2275 1609 2282 1633
rect 1197 1600 2221 1609
rect 0 1529 7 1553
rect 59 1529 66 1553
rect 94 1544 1113 1572
rect 0 1473 5 1529
rect 61 1516 66 1529
rect 1169 1544 2188 1572
rect 2216 1553 2221 1600
rect 2277 1553 2282 1609
rect 1113 1533 1169 1541
rect 1113 1517 1115 1533
rect 1167 1517 1169 1533
rect 61 1488 1085 1516
rect 61 1473 66 1488
rect 0 1462 7 1473
rect 59 1462 66 1473
rect 0 1450 66 1462
rect 2216 1529 2223 1553
rect 2275 1529 2282 1553
rect 2216 1516 2221 1529
rect 1197 1488 2221 1516
rect 1113 1460 1115 1461
rect 0 1449 7 1450
rect 59 1449 66 1450
rect 0 1393 5 1449
rect 61 1404 66 1449
rect 94 1437 1115 1460
rect 1167 1460 1169 1461
rect 2216 1473 2221 1488
rect 2277 1473 2282 1529
rect 2216 1462 2223 1473
rect 2275 1462 2282 1473
rect 1167 1437 2188 1460
rect 94 1432 1113 1437
rect 1169 1432 2188 1437
rect 2216 1450 2282 1462
rect 2216 1449 2223 1450
rect 2275 1449 2282 1450
rect 61 1393 1085 1404
rect 0 1386 1085 1393
rect 0 1369 7 1386
rect 59 1376 1085 1386
rect 2216 1404 2221 1449
rect 59 1369 66 1376
rect 0 1313 5 1369
rect 61 1313 66 1369
rect 1113 1357 1115 1381
rect 1167 1357 1169 1381
rect 1197 1393 2221 1404
rect 2277 1393 2282 1449
rect 1197 1386 2282 1393
rect 1197 1376 2223 1386
rect 94 1320 1113 1348
rect 2216 1369 2223 1376
rect 2275 1369 2282 1386
rect 0 1289 7 1313
rect 59 1292 66 1313
rect 1169 1320 2188 1348
rect 59 1289 1085 1292
rect 0 1233 5 1289
rect 61 1233 1085 1289
rect 0 1225 1085 1233
rect 1113 1289 1115 1301
rect 1167 1289 1169 1301
rect 2216 1313 2221 1369
rect 2277 1313 2282 1369
rect 2216 1292 2223 1313
rect 1113 1277 1169 1289
rect 1197 1289 2223 1292
rect 2275 1289 2282 1313
rect 1197 1233 2221 1289
rect 2277 1233 2282 1289
rect 1197 1225 2282 1233
rect 0 1224 66 1225
rect 2216 1224 2282 1225
rect 1113 1197 1169 1221
rect 74 1196 153 1197
rect 0 1195 153 1196
rect 209 1195 233 1197
rect 289 1195 313 1197
rect 369 1195 393 1197
rect 449 1195 473 1197
rect 529 1195 553 1197
rect 609 1195 633 1197
rect 689 1195 713 1197
rect 769 1195 793 1197
rect 849 1195 873 1197
rect 929 1195 953 1197
rect 1009 1195 1033 1197
rect 1089 1195 1113 1197
rect 0 1143 152 1195
rect 209 1143 216 1195
rect 460 1143 472 1195
rect 529 1143 536 1195
rect 780 1143 792 1195
rect 849 1143 856 1195
rect 1100 1143 1113 1195
rect 0 1142 153 1143
rect 74 1141 153 1142
rect 209 1141 233 1143
rect 289 1141 313 1143
rect 369 1141 393 1143
rect 449 1141 473 1143
rect 529 1141 553 1143
rect 609 1141 633 1143
rect 689 1141 713 1143
rect 769 1141 793 1143
rect 849 1141 873 1143
rect 929 1141 953 1143
rect 1009 1141 1033 1143
rect 1089 1141 1113 1143
rect 1169 1195 1193 1197
rect 1249 1195 1273 1197
rect 1329 1195 1353 1197
rect 1409 1195 1433 1197
rect 1489 1195 1513 1197
rect 1569 1195 1593 1197
rect 1649 1195 1673 1197
rect 1729 1195 1753 1197
rect 1809 1195 1833 1197
rect 1889 1195 1913 1197
rect 1969 1195 1993 1197
rect 2049 1195 2073 1197
rect 2129 1196 2208 1197
rect 2129 1195 2282 1196
rect 1169 1143 1182 1195
rect 1426 1143 1433 1195
rect 1490 1143 1502 1195
rect 1746 1143 1753 1195
rect 1810 1143 1822 1195
rect 2066 1143 2073 1195
rect 2130 1143 2282 1195
rect 1169 1141 1193 1143
rect 1249 1141 1273 1143
rect 1329 1141 1353 1143
rect 1409 1141 1433 1143
rect 1489 1141 1513 1143
rect 1569 1141 1593 1143
rect 1649 1141 1673 1143
rect 1729 1141 1753 1143
rect 1809 1141 1833 1143
rect 1889 1141 1913 1143
rect 1969 1141 1993 1143
rect 2049 1141 2073 1143
rect 2129 1142 2282 1143
rect 2129 1141 2208 1142
rect 1113 1117 1169 1141
rect 0 1113 66 1114
rect 2216 1113 2282 1114
rect 0 1105 1085 1113
rect 0 1049 5 1105
rect 61 1049 1085 1105
rect 0 1025 7 1049
rect 59 1046 1085 1049
rect 1113 1049 1169 1061
rect 59 1025 66 1046
rect 0 969 5 1025
rect 61 969 66 1025
rect 1113 1037 1115 1049
rect 1167 1037 1169 1049
rect 1197 1105 2282 1113
rect 1197 1049 2221 1105
rect 2277 1049 2282 1105
rect 1197 1046 2223 1049
rect 94 990 1113 1018
rect 2216 1025 2223 1046
rect 2275 1025 2282 1049
rect 0 952 7 969
rect 59 962 66 969
rect 1169 990 2188 1018
rect 59 952 1085 962
rect 0 945 1085 952
rect 0 889 5 945
rect 61 934 1085 945
rect 1113 957 1115 981
rect 1167 957 1169 981
rect 2216 969 2221 1025
rect 2277 969 2282 1025
rect 2216 962 2223 969
rect 61 889 66 934
rect 1197 952 2223 962
rect 2275 952 2282 969
rect 1197 945 2282 952
rect 1197 934 2221 945
rect 0 888 7 889
rect 59 888 66 889
rect 0 876 66 888
rect 94 901 1113 906
rect 1169 901 2188 906
rect 94 878 1115 901
rect 0 865 7 876
rect 59 865 66 876
rect 0 809 5 865
rect 61 850 66 865
rect 1113 877 1115 878
rect 1167 878 2188 901
rect 2216 889 2221 934
rect 2277 889 2282 945
rect 2216 888 2223 889
rect 2275 888 2282 889
rect 1167 877 1169 878
rect 61 822 1085 850
rect 61 809 66 822
rect 0 785 7 809
rect 59 785 66 809
rect 2216 876 2282 888
rect 2216 865 2223 876
rect 2275 865 2282 876
rect 2216 850 2221 865
rect 1197 822 2221 850
rect 1113 805 1115 821
rect 1167 805 1169 821
rect 1113 797 1169 805
rect 0 729 5 785
rect 61 738 66 785
rect 94 766 1113 794
rect 2216 809 2221 822
rect 2277 809 2282 865
rect 1169 766 2188 794
rect 2216 785 2223 809
rect 2275 785 2282 809
rect 61 729 1085 738
rect 0 705 7 729
rect 59 710 1085 729
rect 1113 729 1169 741
rect 2216 738 2221 785
rect 1113 717 1115 729
rect 1167 717 1169 729
rect 59 705 66 710
rect 0 649 5 705
rect 61 649 66 705
rect 94 661 1113 682
rect 1197 729 2221 738
rect 2277 729 2282 785
rect 1197 710 2223 729
rect 2216 705 2223 710
rect 2275 705 2282 729
rect 1169 661 2188 682
rect 94 654 1115 661
rect 0 632 7 649
rect 59 632 66 649
rect 0 626 66 632
rect 1113 637 1115 654
rect 1167 654 2188 661
rect 1167 637 1169 654
rect 0 625 1085 626
rect 0 569 5 625
rect 61 598 1085 625
rect 2216 649 2221 705
rect 2277 649 2282 705
rect 2216 632 2223 649
rect 2275 632 2282 649
rect 2216 626 2282 632
rect 61 569 66 598
rect 1197 625 2282 626
rect 1197 598 2221 625
rect 1113 570 1115 581
rect 0 568 7 569
rect 59 568 66 569
rect 0 556 66 568
rect 0 545 7 556
rect 59 545 66 556
rect 0 489 5 545
rect 61 514 66 545
rect 94 557 1115 570
rect 1167 570 1169 581
rect 1167 557 2188 570
rect 94 542 1113 557
rect 1169 542 2188 557
rect 2216 569 2221 598
rect 2277 569 2282 625
rect 2216 568 2223 569
rect 2275 568 2282 569
rect 2216 556 2282 568
rect 2216 545 2223 556
rect 2275 545 2282 556
rect 61 489 1085 514
rect 0 465 7 489
rect 59 486 1085 489
rect 2216 514 2221 545
rect 59 465 66 486
rect 0 409 5 465
rect 61 409 66 465
rect 1113 485 1115 501
rect 1167 485 1169 501
rect 1197 489 2221 514
rect 2277 489 2282 545
rect 1197 486 2223 489
rect 1113 477 1169 485
rect 94 430 1113 458
rect 0 385 7 409
rect 59 402 66 409
rect 2216 465 2223 486
rect 2275 465 2282 489
rect 1169 430 2188 458
rect 1113 409 1169 421
rect 59 385 1085 402
rect 0 329 5 385
rect 61 374 1085 385
rect 1113 397 1115 409
rect 1167 397 1169 409
rect 2216 409 2221 465
rect 2277 409 2282 465
rect 2216 402 2223 409
rect 61 329 66 374
rect 1197 385 2223 402
rect 2275 385 2282 409
rect 1197 374 2221 385
rect 0 312 7 329
rect 59 312 66 329
rect 94 341 1113 346
rect 1169 341 2188 346
rect 94 318 1115 341
rect 0 305 66 312
rect 0 249 5 305
rect 61 290 66 305
rect 1113 317 1115 318
rect 1167 318 2188 341
rect 2216 329 2221 374
rect 2277 329 2282 385
rect 1167 317 1169 318
rect 61 262 1085 290
rect 2216 312 2223 329
rect 2275 312 2282 329
rect 2216 305 2282 312
rect 2216 290 2221 305
rect 61 249 66 262
rect 0 248 7 249
rect 59 248 66 249
rect 0 236 66 248
rect 0 225 7 236
rect 59 225 66 236
rect 1197 262 2221 290
rect 1113 237 1115 261
rect 1167 237 1169 261
rect 0 169 5 225
rect 61 178 66 225
rect 94 206 1113 234
rect 2216 249 2221 262
rect 2277 249 2282 305
rect 2216 248 2223 249
rect 2275 248 2282 249
rect 2216 236 2282 248
rect 1169 206 2188 234
rect 2216 225 2223 236
rect 2275 225 2282 236
rect 61 169 1085 178
rect 0 145 7 169
rect 59 150 1085 169
rect 1113 165 1115 181
rect 1167 165 1169 181
rect 2216 178 2221 225
rect 1113 153 1169 165
rect 59 145 66 150
rect 0 89 5 145
rect 61 89 66 145
rect 1113 122 1115 153
rect 94 101 1115 122
rect 1167 122 1169 153
rect 1197 169 2221 178
rect 2277 169 2282 225
rect 1197 150 2223 169
rect 2216 145 2223 150
rect 2275 145 2282 169
rect 1167 101 2188 122
rect 94 94 2188 101
rect 0 56 7 89
rect 59 66 66 89
rect 59 61 1086 66
rect 59 56 61 61
rect 117 59 141 61
rect 197 59 221 61
rect 277 59 301 61
rect 357 59 381 61
rect 437 59 461 61
rect 517 59 541 61
rect 597 59 621 61
rect 677 59 701 61
rect 757 59 781 61
rect 837 59 861 61
rect 917 59 941 61
rect 997 59 1021 61
rect 0 5 61 56
rect 140 7 141 59
rect 204 7 216 59
rect 277 7 280 59
rect 460 7 461 59
rect 524 7 536 59
rect 597 7 600 59
rect 780 7 781 59
rect 844 7 856 59
rect 917 7 920 59
rect 117 5 141 7
rect 197 5 221 7
rect 277 5 301 7
rect 357 5 381 7
rect 437 5 461 7
rect 517 5 541 7
rect 597 5 621 7
rect 677 5 701 7
rect 757 5 781 7
rect 837 5 861 7
rect 917 5 941 7
rect 997 5 1021 7
rect 1077 5 1086 61
rect 0 0 1086 5
rect 1114 0 1168 94
rect 2216 89 2221 145
rect 2277 89 2282 145
rect 2216 66 2223 89
rect 1196 61 2223 66
rect 1196 5 1205 61
rect 1261 59 1285 61
rect 1341 59 1365 61
rect 1421 59 1445 61
rect 1501 59 1525 61
rect 1581 59 1605 61
rect 1661 59 1685 61
rect 1741 59 1765 61
rect 1821 59 1845 61
rect 1901 59 1925 61
rect 1981 59 2005 61
rect 2061 59 2085 61
rect 2141 59 2165 61
rect 1362 7 1365 59
rect 1426 7 1438 59
rect 1501 7 1502 59
rect 1682 7 1685 59
rect 1746 7 1758 59
rect 1821 7 1822 59
rect 2002 7 2005 59
rect 2066 7 2078 59
rect 2141 7 2142 59
rect 2221 56 2223 61
rect 2275 56 2282 89
rect 1261 5 1285 7
rect 1341 5 1365 7
rect 1421 5 1445 7
rect 1501 5 1525 7
rect 1581 5 1605 7
rect 1661 5 1685 7
rect 1741 5 1765 7
rect 1821 5 1845 7
rect 1901 5 1925 7
rect 1981 5 2005 7
rect 2061 5 2085 7
rect 2141 5 2165 7
rect 2221 5 2282 56
rect 1196 0 2282 5
<< via2 >>
rect 61 2331 117 2333
rect 141 2331 197 2333
rect 221 2331 277 2333
rect 301 2331 357 2333
rect 381 2331 437 2333
rect 461 2331 517 2333
rect 541 2331 597 2333
rect 621 2331 677 2333
rect 701 2331 757 2333
rect 781 2331 837 2333
rect 861 2331 917 2333
rect 941 2331 997 2333
rect 1021 2331 1077 2333
rect 61 2279 88 2331
rect 88 2279 117 2331
rect 141 2279 152 2331
rect 152 2279 197 2331
rect 221 2279 268 2331
rect 268 2279 277 2331
rect 301 2279 332 2331
rect 332 2279 344 2331
rect 344 2279 357 2331
rect 381 2279 396 2331
rect 396 2279 408 2331
rect 408 2279 437 2331
rect 461 2279 472 2331
rect 472 2279 517 2331
rect 541 2279 588 2331
rect 588 2279 597 2331
rect 621 2279 652 2331
rect 652 2279 664 2331
rect 664 2279 677 2331
rect 701 2279 716 2331
rect 716 2279 728 2331
rect 728 2279 757 2331
rect 781 2279 792 2331
rect 792 2279 837 2331
rect 861 2279 908 2331
rect 908 2279 917 2331
rect 941 2279 972 2331
rect 972 2279 984 2331
rect 984 2279 997 2331
rect 1021 2279 1036 2331
rect 1036 2279 1077 2331
rect 61 2277 117 2279
rect 141 2277 197 2279
rect 221 2277 277 2279
rect 301 2277 357 2279
rect 381 2277 437 2279
rect 461 2277 517 2279
rect 541 2277 597 2279
rect 621 2277 677 2279
rect 701 2277 757 2279
rect 781 2277 837 2279
rect 861 2277 917 2279
rect 941 2277 997 2279
rect 1021 2277 1077 2279
rect 5 2230 7 2249
rect 7 2230 59 2249
rect 59 2230 61 2249
rect 5 2218 61 2230
rect 5 2193 7 2218
rect 7 2193 59 2218
rect 59 2193 61 2218
rect 1205 2331 1261 2333
rect 1285 2331 1341 2333
rect 1365 2331 1421 2333
rect 1445 2331 1501 2333
rect 1525 2331 1581 2333
rect 1605 2331 1661 2333
rect 1685 2331 1741 2333
rect 1765 2331 1821 2333
rect 1845 2331 1901 2333
rect 1925 2331 1981 2333
rect 2005 2331 2061 2333
rect 2085 2331 2141 2333
rect 2165 2331 2221 2333
rect 1205 2279 1246 2331
rect 1246 2279 1261 2331
rect 1285 2279 1298 2331
rect 1298 2279 1310 2331
rect 1310 2279 1341 2331
rect 1365 2279 1374 2331
rect 1374 2279 1421 2331
rect 1445 2279 1490 2331
rect 1490 2279 1501 2331
rect 1525 2279 1554 2331
rect 1554 2279 1566 2331
rect 1566 2279 1581 2331
rect 1605 2279 1618 2331
rect 1618 2279 1630 2331
rect 1630 2279 1661 2331
rect 1685 2279 1694 2331
rect 1694 2279 1741 2331
rect 1765 2279 1810 2331
rect 1810 2279 1821 2331
rect 1845 2279 1874 2331
rect 1874 2279 1886 2331
rect 1886 2279 1901 2331
rect 1925 2279 1938 2331
rect 1938 2279 1950 2331
rect 1950 2279 1981 2331
rect 2005 2279 2014 2331
rect 2014 2279 2061 2331
rect 2085 2279 2130 2331
rect 2130 2279 2141 2331
rect 2165 2279 2194 2331
rect 2194 2279 2221 2331
rect 1205 2277 1261 2279
rect 1285 2277 1341 2279
rect 1365 2277 1421 2279
rect 1445 2277 1501 2279
rect 1525 2277 1581 2279
rect 1605 2277 1661 2279
rect 1685 2277 1741 2279
rect 1765 2277 1821 2279
rect 1845 2277 1901 2279
rect 1925 2277 1981 2279
rect 2005 2277 2061 2279
rect 2085 2277 2141 2279
rect 2165 2277 2221 2279
rect 5 2166 7 2169
rect 7 2166 59 2169
rect 59 2166 61 2169
rect 5 2154 61 2166
rect 2221 2230 2223 2249
rect 2223 2230 2275 2249
rect 2275 2230 2277 2249
rect 2221 2218 2277 2230
rect 2221 2193 2223 2218
rect 2223 2193 2275 2218
rect 2275 2193 2277 2218
rect 5 2113 7 2154
rect 7 2113 59 2154
rect 59 2113 61 2154
rect 2221 2166 2223 2169
rect 2223 2166 2275 2169
rect 2275 2166 2277 2169
rect 1113 2121 1115 2157
rect 1115 2121 1167 2157
rect 1167 2121 1169 2157
rect 1113 2109 1169 2121
rect 5 2038 7 2089
rect 7 2038 59 2089
rect 59 2038 61 2089
rect 1113 2101 1115 2109
rect 1115 2101 1167 2109
rect 1167 2101 1169 2109
rect 2221 2154 2277 2166
rect 2221 2113 2223 2154
rect 2223 2113 2275 2154
rect 2275 2113 2277 2154
rect 1113 2057 1115 2077
rect 1115 2057 1167 2077
rect 1167 2057 1169 2077
rect 5 2033 61 2038
rect 1113 2045 1169 2057
rect 1113 2021 1115 2045
rect 1115 2021 1167 2045
rect 1167 2021 1169 2045
rect 5 1974 7 2009
rect 7 1974 59 2009
rect 59 1974 61 2009
rect 5 1962 61 1974
rect 2221 2038 2223 2089
rect 2223 2038 2275 2089
rect 2275 2038 2277 2089
rect 2221 2033 2277 2038
rect 1113 1993 1115 1997
rect 1115 1993 1167 1997
rect 1167 1993 1169 1997
rect 1113 1981 1169 1993
rect 5 1953 7 1962
rect 7 1953 59 1962
rect 59 1953 61 1962
rect 1113 1941 1115 1981
rect 1115 1941 1167 1981
rect 1167 1941 1169 1981
rect 2221 1974 2223 2009
rect 2223 1974 2275 2009
rect 2275 1974 2277 2009
rect 5 1910 7 1929
rect 7 1910 59 1929
rect 59 1910 61 1929
rect 5 1898 61 1910
rect 5 1873 7 1898
rect 7 1873 59 1898
rect 59 1873 61 1898
rect 2221 1962 2277 1974
rect 2221 1953 2223 1962
rect 2223 1953 2275 1962
rect 2275 1953 2277 1962
rect 1113 1865 1115 1917
rect 1115 1865 1167 1917
rect 1167 1865 1169 1917
rect 1113 1861 1169 1865
rect 5 1846 7 1849
rect 7 1846 59 1849
rect 59 1846 61 1849
rect 5 1834 61 1846
rect 5 1793 7 1834
rect 7 1793 59 1834
rect 59 1793 61 1834
rect 2221 1910 2223 1929
rect 2223 1910 2275 1929
rect 2275 1910 2277 1929
rect 2221 1898 2277 1910
rect 2221 1873 2223 1898
rect 2223 1873 2275 1898
rect 2275 1873 2277 1898
rect 1113 1801 1115 1837
rect 1115 1801 1167 1837
rect 1167 1801 1169 1837
rect 2221 1846 2223 1849
rect 2223 1846 2275 1849
rect 2275 1846 2277 1849
rect 2221 1834 2277 1846
rect 5 1718 7 1769
rect 7 1718 59 1769
rect 59 1718 61 1769
rect 1113 1789 1169 1801
rect 1113 1781 1115 1789
rect 1115 1781 1167 1789
rect 1167 1781 1169 1789
rect 2221 1793 2223 1834
rect 2223 1793 2275 1834
rect 2275 1793 2277 1834
rect 5 1713 61 1718
rect 1113 1737 1115 1757
rect 1115 1737 1167 1757
rect 1167 1737 1169 1757
rect 1113 1725 1169 1737
rect 5 1654 7 1689
rect 7 1654 59 1689
rect 59 1654 61 1689
rect 5 1642 61 1654
rect 5 1633 7 1642
rect 7 1633 59 1642
rect 59 1633 61 1642
rect 1113 1701 1115 1725
rect 1115 1701 1167 1725
rect 1167 1701 1169 1725
rect 2221 1718 2223 1769
rect 2223 1718 2275 1769
rect 2275 1718 2277 1769
rect 2221 1713 2277 1718
rect 1113 1673 1115 1677
rect 1115 1673 1167 1677
rect 1167 1673 1169 1677
rect 1113 1661 1169 1673
rect 5 1590 7 1609
rect 7 1590 59 1609
rect 59 1590 61 1609
rect 1113 1621 1115 1661
rect 1115 1621 1167 1661
rect 1167 1621 1169 1661
rect 2221 1654 2223 1689
rect 2223 1654 2275 1689
rect 2275 1654 2277 1689
rect 2221 1642 2277 1654
rect 2221 1633 2223 1642
rect 2223 1633 2275 1642
rect 2275 1633 2277 1642
rect 5 1578 61 1590
rect 5 1553 7 1578
rect 7 1553 59 1578
rect 59 1553 61 1578
rect 1113 1545 1115 1597
rect 1115 1545 1167 1597
rect 1167 1545 1169 1597
rect 5 1526 7 1529
rect 7 1526 59 1529
rect 59 1526 61 1529
rect 5 1514 61 1526
rect 1113 1541 1169 1545
rect 2221 1590 2223 1609
rect 2223 1590 2275 1609
rect 2275 1590 2277 1609
rect 2221 1578 2277 1590
rect 2221 1553 2223 1578
rect 2223 1553 2275 1578
rect 2275 1553 2277 1578
rect 5 1473 7 1514
rect 7 1473 59 1514
rect 59 1473 61 1514
rect 1113 1481 1115 1517
rect 1115 1481 1167 1517
rect 1167 1481 1169 1517
rect 2221 1526 2223 1529
rect 2223 1526 2275 1529
rect 2275 1526 2277 1529
rect 2221 1514 2277 1526
rect 1113 1469 1169 1481
rect 1113 1461 1115 1469
rect 1115 1461 1167 1469
rect 1167 1461 1169 1469
rect 5 1398 7 1449
rect 7 1398 59 1449
rect 59 1398 61 1449
rect 2221 1473 2223 1514
rect 2223 1473 2275 1514
rect 2275 1473 2277 1514
rect 1113 1417 1115 1437
rect 1115 1417 1167 1437
rect 1167 1417 1169 1437
rect 1113 1405 1169 1417
rect 5 1393 61 1398
rect 1113 1381 1115 1405
rect 1115 1381 1167 1405
rect 1167 1381 1169 1405
rect 5 1334 7 1369
rect 7 1334 59 1369
rect 59 1334 61 1369
rect 5 1322 61 1334
rect 5 1313 7 1322
rect 7 1313 59 1322
rect 59 1313 61 1322
rect 2221 1398 2223 1449
rect 2223 1398 2275 1449
rect 2275 1398 2277 1449
rect 2221 1393 2277 1398
rect 1113 1353 1115 1357
rect 1115 1353 1167 1357
rect 1167 1353 1169 1357
rect 1113 1341 1169 1353
rect 1113 1301 1115 1341
rect 1115 1301 1167 1341
rect 1167 1301 1169 1341
rect 5 1270 7 1289
rect 7 1270 59 1289
rect 59 1270 61 1289
rect 5 1233 61 1270
rect 2221 1334 2223 1369
rect 2223 1334 2275 1369
rect 2275 1334 2277 1369
rect 2221 1322 2277 1334
rect 2221 1313 2223 1322
rect 2223 1313 2275 1322
rect 2275 1313 2277 1322
rect 1113 1225 1115 1277
rect 1115 1225 1167 1277
rect 1167 1225 1169 1277
rect 2221 1270 2223 1289
rect 2223 1270 2275 1289
rect 2275 1270 2277 1289
rect 2221 1233 2277 1270
rect 1113 1221 1169 1225
rect 153 1195 209 1197
rect 233 1195 289 1197
rect 313 1195 369 1197
rect 393 1195 449 1197
rect 473 1195 529 1197
rect 553 1195 609 1197
rect 633 1195 689 1197
rect 713 1195 769 1197
rect 793 1195 849 1197
rect 873 1195 929 1197
rect 953 1195 1009 1197
rect 1033 1195 1089 1197
rect 153 1143 204 1195
rect 204 1143 209 1195
rect 233 1143 268 1195
rect 268 1143 280 1195
rect 280 1143 289 1195
rect 313 1143 332 1195
rect 332 1143 344 1195
rect 344 1143 369 1195
rect 393 1143 396 1195
rect 396 1143 408 1195
rect 408 1143 449 1195
rect 473 1143 524 1195
rect 524 1143 529 1195
rect 553 1143 588 1195
rect 588 1143 600 1195
rect 600 1143 609 1195
rect 633 1143 652 1195
rect 652 1143 664 1195
rect 664 1143 689 1195
rect 713 1143 716 1195
rect 716 1143 728 1195
rect 728 1143 769 1195
rect 793 1143 844 1195
rect 844 1143 849 1195
rect 873 1143 908 1195
rect 908 1143 920 1195
rect 920 1143 929 1195
rect 953 1143 972 1195
rect 972 1143 984 1195
rect 984 1143 1009 1195
rect 1033 1143 1036 1195
rect 1036 1143 1048 1195
rect 1048 1143 1089 1195
rect 153 1141 209 1143
rect 233 1141 289 1143
rect 313 1141 369 1143
rect 393 1141 449 1143
rect 473 1141 529 1143
rect 553 1141 609 1143
rect 633 1141 689 1143
rect 713 1141 769 1143
rect 793 1141 849 1143
rect 873 1141 929 1143
rect 953 1141 1009 1143
rect 1033 1141 1089 1143
rect 1113 1141 1169 1197
rect 1193 1195 1249 1197
rect 1273 1195 1329 1197
rect 1353 1195 1409 1197
rect 1433 1195 1489 1197
rect 1513 1195 1569 1197
rect 1593 1195 1649 1197
rect 1673 1195 1729 1197
rect 1753 1195 1809 1197
rect 1833 1195 1889 1197
rect 1913 1195 1969 1197
rect 1993 1195 2049 1197
rect 2073 1195 2129 1197
rect 1193 1143 1234 1195
rect 1234 1143 1246 1195
rect 1246 1143 1249 1195
rect 1273 1143 1298 1195
rect 1298 1143 1310 1195
rect 1310 1143 1329 1195
rect 1353 1143 1362 1195
rect 1362 1143 1374 1195
rect 1374 1143 1409 1195
rect 1433 1143 1438 1195
rect 1438 1143 1489 1195
rect 1513 1143 1554 1195
rect 1554 1143 1566 1195
rect 1566 1143 1569 1195
rect 1593 1143 1618 1195
rect 1618 1143 1630 1195
rect 1630 1143 1649 1195
rect 1673 1143 1682 1195
rect 1682 1143 1694 1195
rect 1694 1143 1729 1195
rect 1753 1143 1758 1195
rect 1758 1143 1809 1195
rect 1833 1143 1874 1195
rect 1874 1143 1886 1195
rect 1886 1143 1889 1195
rect 1913 1143 1938 1195
rect 1938 1143 1950 1195
rect 1950 1143 1969 1195
rect 1993 1143 2002 1195
rect 2002 1143 2014 1195
rect 2014 1143 2049 1195
rect 2073 1143 2078 1195
rect 2078 1143 2129 1195
rect 1193 1141 1249 1143
rect 1273 1141 1329 1143
rect 1353 1141 1409 1143
rect 1433 1141 1489 1143
rect 1513 1141 1569 1143
rect 1593 1141 1649 1143
rect 1673 1141 1729 1143
rect 1753 1141 1809 1143
rect 1833 1141 1889 1143
rect 1913 1141 1969 1143
rect 1993 1141 2049 1143
rect 2073 1141 2129 1143
rect 1113 1113 1169 1117
rect 5 1068 61 1105
rect 5 1049 7 1068
rect 7 1049 59 1068
rect 59 1049 61 1068
rect 1113 1061 1115 1113
rect 1115 1061 1167 1113
rect 1167 1061 1169 1113
rect 5 1016 7 1025
rect 7 1016 59 1025
rect 59 1016 61 1025
rect 5 1004 61 1016
rect 5 969 7 1004
rect 7 969 59 1004
rect 59 969 61 1004
rect 2221 1068 2277 1105
rect 2221 1049 2223 1068
rect 2223 1049 2275 1068
rect 2275 1049 2277 1068
rect 1113 997 1115 1037
rect 1115 997 1167 1037
rect 1167 997 1169 1037
rect 1113 985 1169 997
rect 1113 981 1115 985
rect 1115 981 1167 985
rect 1167 981 1169 985
rect 5 940 61 945
rect 5 889 7 940
rect 7 889 59 940
rect 59 889 61 940
rect 2221 1016 2223 1025
rect 2223 1016 2275 1025
rect 2275 1016 2277 1025
rect 2221 1004 2277 1016
rect 2221 969 2223 1004
rect 2223 969 2275 1004
rect 2275 969 2277 1004
rect 1113 933 1115 957
rect 1115 933 1167 957
rect 1167 933 1169 957
rect 2221 940 2277 945
rect 1113 921 1169 933
rect 1113 901 1115 921
rect 1115 901 1167 921
rect 1167 901 1169 921
rect 5 824 7 865
rect 7 824 59 865
rect 59 824 61 865
rect 2221 889 2223 940
rect 2223 889 2275 940
rect 2275 889 2277 940
rect 1113 869 1115 877
rect 1115 869 1167 877
rect 1167 869 1169 877
rect 1113 857 1169 869
rect 5 812 61 824
rect 5 809 7 812
rect 7 809 59 812
rect 59 809 61 812
rect 1113 821 1115 857
rect 1115 821 1167 857
rect 1167 821 1169 857
rect 2221 824 2223 865
rect 2223 824 2275 865
rect 2275 824 2277 865
rect 5 760 7 785
rect 7 760 59 785
rect 59 760 61 785
rect 5 748 61 760
rect 5 729 7 748
rect 7 729 59 748
rect 59 729 61 748
rect 1113 793 1169 797
rect 2221 812 2277 824
rect 2221 809 2223 812
rect 2223 809 2275 812
rect 2275 809 2277 812
rect 1113 741 1115 793
rect 1115 741 1167 793
rect 1167 741 1169 793
rect 2221 760 2223 785
rect 2223 760 2275 785
rect 2275 760 2277 785
rect 2221 748 2277 760
rect 5 696 7 705
rect 7 696 59 705
rect 59 696 61 705
rect 5 684 61 696
rect 5 649 7 684
rect 7 649 59 684
rect 59 649 61 684
rect 1113 677 1115 717
rect 1115 677 1167 717
rect 1167 677 1169 717
rect 2221 729 2223 748
rect 2223 729 2275 748
rect 2275 729 2277 748
rect 1113 665 1169 677
rect 1113 661 1115 665
rect 1115 661 1167 665
rect 1167 661 1169 665
rect 5 620 61 625
rect 5 569 7 620
rect 7 569 59 620
rect 59 569 61 620
rect 1113 613 1115 637
rect 1115 613 1167 637
rect 1167 613 1169 637
rect 2221 696 2223 705
rect 2223 696 2275 705
rect 2275 696 2277 705
rect 2221 684 2277 696
rect 2221 649 2223 684
rect 2223 649 2275 684
rect 2275 649 2277 684
rect 1113 601 1169 613
rect 1113 581 1115 601
rect 1115 581 1167 601
rect 1167 581 1169 601
rect 2221 620 2277 625
rect 5 504 7 545
rect 7 504 59 545
rect 59 504 61 545
rect 1113 549 1115 557
rect 1115 549 1167 557
rect 1167 549 1169 557
rect 1113 537 1169 549
rect 2221 569 2223 620
rect 2223 569 2275 620
rect 2275 569 2277 620
rect 5 492 61 504
rect 5 489 7 492
rect 7 489 59 492
rect 59 489 61 492
rect 1113 501 1115 537
rect 1115 501 1167 537
rect 1167 501 1169 537
rect 5 440 7 465
rect 7 440 59 465
rect 59 440 61 465
rect 5 428 61 440
rect 5 409 7 428
rect 7 409 59 428
rect 59 409 61 428
rect 2221 504 2223 545
rect 2223 504 2275 545
rect 2275 504 2277 545
rect 2221 492 2277 504
rect 2221 489 2223 492
rect 2223 489 2275 492
rect 2275 489 2277 492
rect 1113 473 1169 477
rect 1113 421 1115 473
rect 1115 421 1167 473
rect 1167 421 1169 473
rect 5 376 7 385
rect 7 376 59 385
rect 59 376 61 385
rect 5 364 61 376
rect 2221 440 2223 465
rect 2223 440 2275 465
rect 2275 440 2277 465
rect 2221 428 2277 440
rect 2221 409 2223 428
rect 2223 409 2275 428
rect 2275 409 2277 428
rect 5 329 7 364
rect 7 329 59 364
rect 59 329 61 364
rect 1113 357 1115 397
rect 1115 357 1167 397
rect 1167 357 1169 397
rect 2221 376 2223 385
rect 2223 376 2275 385
rect 2275 376 2277 385
rect 1113 345 1169 357
rect 1113 341 1115 345
rect 1115 341 1167 345
rect 1167 341 1169 345
rect 5 300 61 305
rect 5 249 7 300
rect 7 249 59 300
rect 59 249 61 300
rect 2221 364 2277 376
rect 2221 329 2223 364
rect 2223 329 2275 364
rect 2275 329 2277 364
rect 1113 293 1115 317
rect 1115 293 1167 317
rect 1167 293 1169 317
rect 1113 281 1169 293
rect 2221 300 2277 305
rect 1113 261 1115 281
rect 1115 261 1167 281
rect 1167 261 1169 281
rect 5 184 7 225
rect 7 184 59 225
rect 59 184 61 225
rect 5 172 61 184
rect 1113 229 1115 237
rect 1115 229 1167 237
rect 1167 229 1169 237
rect 2221 249 2223 300
rect 2223 249 2275 300
rect 2275 249 2277 300
rect 1113 217 1169 229
rect 1113 181 1115 217
rect 1115 181 1167 217
rect 1167 181 1169 217
rect 5 169 7 172
rect 7 169 59 172
rect 59 169 61 172
rect 2221 184 2223 225
rect 2223 184 2275 225
rect 2275 184 2277 225
rect 5 120 7 145
rect 7 120 59 145
rect 59 120 61 145
rect 5 108 61 120
rect 5 89 7 108
rect 7 89 59 108
rect 59 89 61 108
rect 2221 172 2277 184
rect 2221 169 2223 172
rect 2223 169 2275 172
rect 2275 169 2277 172
rect 61 59 117 61
rect 141 59 197 61
rect 221 59 277 61
rect 301 59 357 61
rect 381 59 437 61
rect 461 59 517 61
rect 541 59 597 61
rect 621 59 677 61
rect 701 59 757 61
rect 781 59 837 61
rect 861 59 917 61
rect 941 59 997 61
rect 1021 59 1077 61
rect 61 7 88 59
rect 88 7 117 59
rect 141 7 152 59
rect 152 7 197 59
rect 221 7 268 59
rect 268 7 277 59
rect 301 7 332 59
rect 332 7 344 59
rect 344 7 357 59
rect 381 7 396 59
rect 396 7 408 59
rect 408 7 437 59
rect 461 7 472 59
rect 472 7 517 59
rect 541 7 588 59
rect 588 7 597 59
rect 621 7 652 59
rect 652 7 664 59
rect 664 7 677 59
rect 701 7 716 59
rect 716 7 728 59
rect 728 7 757 59
rect 781 7 792 59
rect 792 7 837 59
rect 861 7 908 59
rect 908 7 917 59
rect 941 7 972 59
rect 972 7 984 59
rect 984 7 997 59
rect 1021 7 1036 59
rect 1036 7 1077 59
rect 61 5 117 7
rect 141 5 197 7
rect 221 5 277 7
rect 301 5 357 7
rect 381 5 437 7
rect 461 5 517 7
rect 541 5 597 7
rect 621 5 677 7
rect 701 5 757 7
rect 781 5 837 7
rect 861 5 917 7
rect 941 5 997 7
rect 1021 5 1077 7
rect 2221 120 2223 145
rect 2223 120 2275 145
rect 2275 120 2277 145
rect 2221 108 2277 120
rect 2221 89 2223 108
rect 2223 89 2275 108
rect 2275 89 2277 108
rect 1205 59 1261 61
rect 1285 59 1341 61
rect 1365 59 1421 61
rect 1445 59 1501 61
rect 1525 59 1581 61
rect 1605 59 1661 61
rect 1685 59 1741 61
rect 1765 59 1821 61
rect 1845 59 1901 61
rect 1925 59 1981 61
rect 2005 59 2061 61
rect 2085 59 2141 61
rect 2165 59 2221 61
rect 1205 7 1246 59
rect 1246 7 1261 59
rect 1285 7 1298 59
rect 1298 7 1310 59
rect 1310 7 1341 59
rect 1365 7 1374 59
rect 1374 7 1421 59
rect 1445 7 1490 59
rect 1490 7 1501 59
rect 1525 7 1554 59
rect 1554 7 1566 59
rect 1566 7 1581 59
rect 1605 7 1618 59
rect 1618 7 1630 59
rect 1630 7 1661 59
rect 1685 7 1694 59
rect 1694 7 1741 59
rect 1765 7 1810 59
rect 1810 7 1821 59
rect 1845 7 1874 59
rect 1874 7 1886 59
rect 1886 7 1901 59
rect 1925 7 1938 59
rect 1938 7 1950 59
rect 1950 7 1981 59
rect 2005 7 2014 59
rect 2014 7 2061 59
rect 2085 7 2130 59
rect 2130 7 2141 59
rect 2165 7 2194 59
rect 2194 7 2221 59
rect 1205 5 1261 7
rect 1285 5 1341 7
rect 1365 5 1421 7
rect 1445 5 1501 7
rect 1525 5 1581 7
rect 1605 5 1661 7
rect 1685 5 1741 7
rect 1765 5 1821 7
rect 1845 5 1901 7
rect 1925 5 1981 7
rect 2005 5 2061 7
rect 2085 5 2141 7
rect 2165 5 2221 7
<< metal3 >>
rect 0 2333 2282 2338
rect 0 2277 61 2333
rect 117 2277 141 2333
rect 197 2277 221 2333
rect 277 2277 301 2333
rect 357 2277 381 2333
rect 437 2277 461 2333
rect 517 2277 541 2333
rect 597 2277 621 2333
rect 677 2277 701 2333
rect 757 2277 781 2333
rect 837 2277 861 2333
rect 917 2277 941 2333
rect 997 2277 1021 2333
rect 1077 2277 1205 2333
rect 1261 2277 1285 2333
rect 1341 2277 1365 2333
rect 1421 2277 1445 2333
rect 1501 2277 1525 2333
rect 1581 2277 1605 2333
rect 1661 2277 1685 2333
rect 1741 2277 1765 2333
rect 1821 2277 1845 2333
rect 1901 2277 1925 2333
rect 1981 2277 2005 2333
rect 2061 2277 2085 2333
rect 2141 2277 2165 2333
rect 2221 2277 2282 2333
rect 0 2272 2282 2277
rect 0 2249 66 2272
rect 0 2193 5 2249
rect 61 2193 66 2249
rect 0 2169 66 2193
rect 0 2113 5 2169
rect 61 2113 66 2169
rect 0 2089 66 2113
rect 0 2033 5 2089
rect 61 2033 66 2089
rect 0 2009 66 2033
rect 0 1953 5 2009
rect 61 1953 66 2009
rect 0 1929 66 1953
rect 0 1873 5 1929
rect 61 1873 66 1929
rect 0 1849 66 1873
rect 0 1793 5 1849
rect 61 1793 66 1849
rect 0 1769 66 1793
rect 0 1713 5 1769
rect 61 1713 66 1769
rect 0 1689 66 1713
rect 0 1633 5 1689
rect 61 1633 66 1689
rect 0 1609 66 1633
rect 0 1553 5 1609
rect 61 1553 66 1609
rect 0 1529 66 1553
rect 0 1473 5 1529
rect 61 1473 66 1529
rect 0 1449 66 1473
rect 0 1393 5 1449
rect 61 1393 66 1449
rect 0 1369 66 1393
rect 0 1313 5 1369
rect 61 1313 66 1369
rect 0 1289 66 1313
rect 0 1233 5 1289
rect 61 1233 66 1289
rect 0 1105 66 1233
rect 0 1049 5 1105
rect 61 1049 66 1105
rect 0 1025 66 1049
rect 0 969 5 1025
rect 61 969 66 1025
rect 0 945 66 969
rect 0 889 5 945
rect 61 889 66 945
rect 0 865 66 889
rect 0 809 5 865
rect 61 809 66 865
rect 0 785 66 809
rect 0 729 5 785
rect 61 729 66 785
rect 0 705 66 729
rect 0 649 5 705
rect 61 649 66 705
rect 0 625 66 649
rect 0 569 5 625
rect 61 569 66 625
rect 0 545 66 569
rect 0 489 5 545
rect 61 489 66 545
rect 0 465 66 489
rect 0 409 5 465
rect 61 409 66 465
rect 0 385 66 409
rect 0 329 5 385
rect 61 329 66 385
rect 0 305 66 329
rect 0 249 5 305
rect 61 249 66 305
rect 0 225 66 249
rect 0 169 5 225
rect 61 169 66 225
rect 0 145 66 169
rect 0 89 5 145
rect 61 89 66 145
rect 126 1202 186 2212
rect 246 1262 306 2272
rect 366 1202 426 2212
rect 486 1262 546 2272
rect 606 1202 666 2212
rect 726 1262 786 2272
rect 846 1202 906 2212
rect 966 1262 1048 2272
rect 1108 2157 1174 2212
rect 1108 2101 1113 2157
rect 1169 2101 1174 2157
rect 1108 2077 1174 2101
rect 1108 2021 1113 2077
rect 1169 2021 1174 2077
rect 1108 1997 1174 2021
rect 1108 1941 1113 1997
rect 1169 1941 1174 1997
rect 1108 1917 1174 1941
rect 1108 1861 1113 1917
rect 1169 1861 1174 1917
rect 1108 1837 1174 1861
rect 1108 1781 1113 1837
rect 1169 1781 1174 1837
rect 1108 1757 1174 1781
rect 1108 1701 1113 1757
rect 1169 1701 1174 1757
rect 1108 1677 1174 1701
rect 1108 1621 1113 1677
rect 1169 1621 1174 1677
rect 1108 1597 1174 1621
rect 1108 1541 1113 1597
rect 1169 1541 1174 1597
rect 1108 1517 1174 1541
rect 1108 1461 1113 1517
rect 1169 1461 1174 1517
rect 1108 1437 1174 1461
rect 1108 1381 1113 1437
rect 1169 1381 1174 1437
rect 1108 1357 1174 1381
rect 1108 1301 1113 1357
rect 1169 1301 1174 1357
rect 1108 1277 1174 1301
rect 1108 1221 1113 1277
rect 1169 1221 1174 1277
rect 1234 1262 1316 2272
rect 1108 1202 1174 1221
rect 1376 1202 1436 2212
rect 1496 1262 1556 2272
rect 1616 1202 1676 2212
rect 1736 1262 1796 2272
rect 1856 1202 1916 2212
rect 1976 1262 2036 2272
rect 2216 2249 2282 2272
rect 2096 1202 2156 2212
rect 126 1197 2156 1202
rect 126 1141 153 1197
rect 209 1141 233 1197
rect 289 1141 313 1197
rect 369 1141 393 1197
rect 449 1141 473 1197
rect 529 1141 553 1197
rect 609 1141 633 1197
rect 689 1141 713 1197
rect 769 1141 793 1197
rect 849 1141 873 1197
rect 929 1141 953 1197
rect 1009 1141 1033 1197
rect 1089 1141 1113 1197
rect 1169 1141 1193 1197
rect 1249 1141 1273 1197
rect 1329 1141 1353 1197
rect 1409 1141 1433 1197
rect 1489 1141 1513 1197
rect 1569 1141 1593 1197
rect 1649 1141 1673 1197
rect 1729 1141 1753 1197
rect 1809 1141 1833 1197
rect 1889 1141 1913 1197
rect 1969 1141 1993 1197
rect 2049 1141 2073 1197
rect 2129 1141 2156 1197
rect 126 1136 2156 1141
rect 126 126 186 1136
rect 0 66 66 89
rect 246 66 306 1076
rect 366 126 426 1136
rect 486 66 546 1076
rect 606 126 666 1136
rect 726 66 786 1076
rect 846 126 906 1136
rect 1108 1117 1174 1136
rect 966 66 1048 1076
rect 1108 1061 1113 1117
rect 1169 1061 1174 1117
rect 1108 1037 1174 1061
rect 1108 981 1113 1037
rect 1169 981 1174 1037
rect 1108 957 1174 981
rect 1108 901 1113 957
rect 1169 901 1174 957
rect 1108 877 1174 901
rect 1108 821 1113 877
rect 1169 821 1174 877
rect 1108 797 1174 821
rect 1108 741 1113 797
rect 1169 741 1174 797
rect 1108 717 1174 741
rect 1108 661 1113 717
rect 1169 661 1174 717
rect 1108 637 1174 661
rect 1108 581 1113 637
rect 1169 581 1174 637
rect 1108 557 1174 581
rect 1108 501 1113 557
rect 1169 501 1174 557
rect 1108 477 1174 501
rect 1108 421 1113 477
rect 1169 421 1174 477
rect 1108 397 1174 421
rect 1108 341 1113 397
rect 1169 341 1174 397
rect 1108 317 1174 341
rect 1108 261 1113 317
rect 1169 261 1174 317
rect 1108 237 1174 261
rect 1108 181 1113 237
rect 1169 181 1174 237
rect 1108 126 1174 181
rect 1234 66 1316 1076
rect 1376 126 1436 1136
rect 1496 66 1556 1076
rect 1616 126 1676 1136
rect 1736 66 1796 1076
rect 1856 126 1916 1136
rect 1976 66 2036 1076
rect 2096 126 2156 1136
rect 2216 2193 2221 2249
rect 2277 2193 2282 2249
rect 2216 2169 2282 2193
rect 2216 2113 2221 2169
rect 2277 2113 2282 2169
rect 2216 2089 2282 2113
rect 2216 2033 2221 2089
rect 2277 2033 2282 2089
rect 2216 2009 2282 2033
rect 2216 1953 2221 2009
rect 2277 1953 2282 2009
rect 2216 1929 2282 1953
rect 2216 1873 2221 1929
rect 2277 1873 2282 1929
rect 2216 1849 2282 1873
rect 2216 1793 2221 1849
rect 2277 1793 2282 1849
rect 2216 1769 2282 1793
rect 2216 1713 2221 1769
rect 2277 1713 2282 1769
rect 2216 1689 2282 1713
rect 2216 1633 2221 1689
rect 2277 1633 2282 1689
rect 2216 1609 2282 1633
rect 2216 1553 2221 1609
rect 2277 1553 2282 1609
rect 2216 1529 2282 1553
rect 2216 1473 2221 1529
rect 2277 1473 2282 1529
rect 2216 1449 2282 1473
rect 2216 1393 2221 1449
rect 2277 1393 2282 1449
rect 2216 1369 2282 1393
rect 2216 1313 2221 1369
rect 2277 1313 2282 1369
rect 2216 1289 2282 1313
rect 2216 1233 2221 1289
rect 2277 1233 2282 1289
rect 2216 1105 2282 1233
rect 2216 1049 2221 1105
rect 2277 1049 2282 1105
rect 2216 1025 2282 1049
rect 2216 969 2221 1025
rect 2277 969 2282 1025
rect 2216 945 2282 969
rect 2216 889 2221 945
rect 2277 889 2282 945
rect 2216 865 2282 889
rect 2216 809 2221 865
rect 2277 809 2282 865
rect 2216 785 2282 809
rect 2216 729 2221 785
rect 2277 729 2282 785
rect 2216 705 2282 729
rect 2216 649 2221 705
rect 2277 649 2282 705
rect 2216 625 2282 649
rect 2216 569 2221 625
rect 2277 569 2282 625
rect 2216 545 2282 569
rect 2216 489 2221 545
rect 2277 489 2282 545
rect 2216 465 2282 489
rect 2216 409 2221 465
rect 2277 409 2282 465
rect 2216 385 2282 409
rect 2216 329 2221 385
rect 2277 329 2282 385
rect 2216 305 2282 329
rect 2216 249 2221 305
rect 2277 249 2282 305
rect 2216 225 2282 249
rect 2216 169 2221 225
rect 2277 169 2282 225
rect 2216 145 2282 169
rect 2216 89 2221 145
rect 2277 89 2282 145
rect 2216 66 2282 89
rect 0 61 2282 66
rect 0 5 61 61
rect 117 5 141 61
rect 197 5 221 61
rect 277 5 301 61
rect 357 5 381 61
rect 437 5 461 61
rect 517 5 541 61
rect 597 5 621 61
rect 677 5 701 61
rect 757 5 781 61
rect 837 5 861 61
rect 917 5 941 61
rect 997 5 1021 61
rect 1077 5 1205 61
rect 1261 5 1285 61
rect 1341 5 1365 61
rect 1421 5 1445 61
rect 1501 5 1525 61
rect 1581 5 1605 61
rect 1661 5 1685 61
rect 1741 5 1765 61
rect 1821 5 1845 61
rect 1901 5 1925 61
rect 1981 5 2005 61
rect 2061 5 2085 61
rect 2141 5 2165 61
rect 2221 5 2282 61
rect 0 0 2282 5
<< metal4 >>
rect 0 0 2282 2338
<< labels >>
flabel metal2 s 1120 2288 1162 2324 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel metal2 s 1018 2297 1048 2325 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal4 s 1776 530 1863 625 0 FreeSans 200 0 0 0 MET4
port 3 nsew
flabel pwell s 1178 1416 1199 1465 0 FreeSans 2000 0 0 0 SUB
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 715040
string GDS_START 656130
<< end >>
