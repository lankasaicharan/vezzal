magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 191 157 568 241
rect 1 49 568 157
rect 0 0 576 49
<< scnmos >>
rect 270 131 300 215
rect 342 131 372 215
rect 80 47 110 131
rect 459 47 489 215
<< scpmoshvt >>
rect 112 367 142 451
rect 231 367 261 451
rect 342 367 372 451
rect 454 367 484 619
<< ndiff >>
rect 217 189 270 215
rect 217 155 225 189
rect 259 155 270 189
rect 217 131 270 155
rect 300 131 342 215
rect 372 187 459 215
rect 372 153 383 187
rect 417 153 459 187
rect 372 131 459 153
rect 27 106 80 131
rect 27 72 35 106
rect 69 72 80 106
rect 27 47 80 72
rect 110 103 163 131
rect 110 69 121 103
rect 155 69 163 103
rect 110 47 163 69
rect 406 93 459 131
rect 406 59 414 93
rect 448 59 459 93
rect 406 47 459 59
rect 489 203 542 215
rect 489 169 500 203
rect 534 169 542 203
rect 489 101 542 169
rect 489 67 500 101
rect 534 67 542 101
rect 489 47 542 67
<< pdiff >>
rect 401 607 454 619
rect 401 573 409 607
rect 443 573 454 607
rect 401 503 454 573
rect 401 469 409 503
rect 443 469 454 503
rect 401 451 454 469
rect 59 426 112 451
rect 59 392 67 426
rect 101 392 112 426
rect 59 367 112 392
rect 142 424 231 451
rect 142 390 169 424
rect 203 390 231 424
rect 142 367 231 390
rect 261 414 342 451
rect 261 380 289 414
rect 323 380 342 414
rect 261 367 342 380
rect 372 414 454 451
rect 372 380 383 414
rect 417 380 454 414
rect 372 367 454 380
rect 484 599 537 619
rect 484 565 495 599
rect 529 565 537 599
rect 484 502 537 565
rect 484 468 495 502
rect 529 468 537 502
rect 484 413 537 468
rect 484 379 495 413
rect 529 379 537 413
rect 484 367 537 379
<< ndiffc >>
rect 225 155 259 189
rect 383 153 417 187
rect 35 72 69 106
rect 121 69 155 103
rect 414 59 448 93
rect 500 169 534 203
rect 500 67 534 101
<< pdiffc >>
rect 409 573 443 607
rect 409 469 443 503
rect 67 392 101 426
rect 169 390 203 424
rect 289 380 323 414
rect 383 380 417 414
rect 495 565 529 599
rect 495 468 529 502
rect 495 379 529 413
<< poly >>
rect 454 619 484 645
rect 303 601 372 617
rect 303 567 319 601
rect 353 567 372 601
rect 303 533 372 567
rect 303 499 319 533
rect 353 499 372 533
rect 303 483 372 499
rect 112 451 142 477
rect 231 451 261 477
rect 342 451 372 483
rect 112 219 142 367
rect 231 333 261 367
rect 195 317 261 333
rect 195 283 211 317
rect 245 283 261 317
rect 195 267 261 283
rect 231 237 300 267
rect 80 203 171 219
rect 270 215 300 237
rect 342 215 372 367
rect 454 303 484 367
rect 414 287 489 303
rect 414 253 430 287
rect 464 253 489 287
rect 414 237 489 253
rect 459 215 489 237
rect 80 169 121 203
rect 155 169 171 203
rect 80 153 171 169
rect 80 131 110 153
rect 270 105 300 131
rect 342 105 372 131
rect 80 21 110 47
rect 459 21 489 47
<< polycont >>
rect 319 567 353 601
rect 319 499 353 533
rect 211 283 245 317
rect 430 253 464 287
rect 121 169 155 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 19 426 108 442
rect 19 392 67 426
rect 101 392 108 426
rect 19 333 108 392
rect 142 430 177 649
rect 211 601 369 615
rect 211 567 319 601
rect 353 567 369 601
rect 211 533 369 567
rect 211 499 319 533
rect 353 499 369 533
rect 211 464 369 499
rect 403 607 457 649
rect 403 573 409 607
rect 443 573 457 607
rect 403 503 457 573
rect 403 469 409 503
rect 443 469 457 503
rect 403 430 457 469
rect 142 424 219 430
rect 142 390 169 424
rect 203 390 219 424
rect 142 374 219 390
rect 279 414 339 430
rect 279 380 289 414
rect 323 380 339 414
rect 19 317 245 333
rect 19 283 211 317
rect 19 267 245 283
rect 279 303 339 380
rect 373 414 457 430
rect 373 380 383 414
rect 417 380 457 414
rect 373 353 457 380
rect 491 599 559 615
rect 491 565 495 599
rect 529 565 559 599
rect 491 502 559 565
rect 491 468 495 502
rect 529 468 559 502
rect 491 413 559 468
rect 491 379 495 413
rect 529 379 559 413
rect 491 339 559 379
rect 279 287 464 303
rect 19 106 77 267
rect 279 253 430 287
rect 279 237 464 253
rect 111 203 175 219
rect 279 205 315 237
rect 111 169 121 203
rect 155 169 175 203
rect 111 153 175 169
rect 209 189 315 205
rect 498 203 559 339
rect 209 155 225 189
rect 259 155 315 189
rect 209 139 315 155
rect 367 187 464 203
rect 367 153 383 187
rect 417 153 464 187
rect 19 72 35 106
rect 69 72 77 106
rect 19 56 77 72
rect 111 103 171 119
rect 111 69 121 103
rect 155 69 171 103
rect 111 17 171 69
rect 367 93 464 153
rect 367 59 414 93
rect 448 59 464 93
rect 367 17 464 59
rect 498 169 500 203
rect 534 169 559 203
rect 498 101 559 169
rect 498 67 500 101
rect 534 67 559 101
rect 498 51 559 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and2b_1
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5120350
string GDS_START 5113958
<< end >>
