magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 29 171 1317 229
rect 29 49 1508 171
rect 0 0 1536 49
<< scnmos >>
rect 108 119 138 203
rect 194 119 224 203
rect 266 119 296 203
rect 352 119 382 203
rect 446 119 476 203
rect 556 119 586 203
rect 751 119 781 203
rect 837 119 867 203
rect 943 119 973 203
rect 1029 119 1059 203
rect 1115 119 1145 203
rect 1209 119 1239 203
rect 1313 61 1343 145
rect 1399 61 1429 145
<< scpmoshvt >>
rect 80 488 110 616
rect 188 532 218 616
rect 266 532 296 616
rect 374 532 404 616
rect 460 532 490 616
rect 554 532 584 616
rect 751 457 781 541
rect 837 457 867 541
rect 943 457 973 541
rect 1029 457 1059 541
rect 1131 457 1161 541
rect 1209 457 1239 541
rect 1317 457 1347 541
rect 1426 457 1456 585
<< ndiff >>
rect 55 175 108 203
rect 55 141 63 175
rect 97 141 108 175
rect 55 119 108 141
rect 138 178 194 203
rect 138 144 149 178
rect 183 144 194 178
rect 138 119 194 144
rect 224 119 266 203
rect 296 178 352 203
rect 296 144 307 178
rect 341 144 352 178
rect 296 119 352 144
rect 382 178 446 203
rect 382 144 399 178
rect 433 144 446 178
rect 382 119 446 144
rect 476 140 556 203
rect 476 119 499 140
rect 491 106 499 119
rect 533 119 556 140
rect 586 178 639 203
rect 586 144 597 178
rect 631 144 639 178
rect 586 119 639 144
rect 698 176 751 203
rect 698 142 706 176
rect 740 142 751 176
rect 698 119 751 142
rect 781 176 837 203
rect 781 142 792 176
rect 826 142 837 176
rect 781 119 837 142
rect 867 165 943 203
rect 867 131 888 165
rect 922 131 943 165
rect 867 119 943 131
rect 973 176 1029 203
rect 973 142 984 176
rect 1018 142 1029 176
rect 973 119 1029 142
rect 1059 176 1115 203
rect 1059 142 1070 176
rect 1104 142 1115 176
rect 1059 119 1115 142
rect 1145 119 1209 203
rect 1239 145 1291 203
rect 1239 119 1313 145
rect 533 106 541 119
rect 491 90 541 106
rect 1261 61 1313 119
rect 1343 120 1399 145
rect 1343 86 1354 120
rect 1388 86 1399 120
rect 1343 61 1399 86
rect 1429 120 1482 145
rect 1429 86 1440 120
rect 1474 86 1482 120
rect 1429 61 1482 86
<< pdiff >>
rect 27 604 80 616
rect 27 570 35 604
rect 69 570 80 604
rect 27 534 80 570
rect 27 500 35 534
rect 69 500 80 534
rect 27 488 80 500
rect 110 582 188 616
rect 110 548 132 582
rect 166 548 188 582
rect 110 532 188 548
rect 218 532 266 616
rect 296 591 374 616
rect 296 557 320 591
rect 354 557 374 591
rect 296 532 374 557
rect 404 591 460 616
rect 404 557 415 591
rect 449 557 460 591
rect 404 532 460 557
rect 490 603 554 616
rect 490 569 505 603
rect 539 569 554 603
rect 490 532 554 569
rect 584 591 637 616
rect 584 557 595 591
rect 629 557 637 591
rect 584 532 637 557
rect 110 488 163 532
rect 1369 566 1426 585
rect 1369 541 1377 566
rect 698 515 751 541
rect 698 481 706 515
rect 740 481 751 515
rect 698 457 751 481
rect 781 517 837 541
rect 781 483 792 517
rect 826 483 837 517
rect 781 457 837 483
rect 867 525 943 541
rect 867 491 888 525
rect 922 491 943 525
rect 867 457 943 491
rect 973 517 1029 541
rect 973 483 984 517
rect 1018 483 1029 517
rect 973 457 1029 483
rect 1059 517 1131 541
rect 1059 483 1079 517
rect 1113 483 1131 517
rect 1059 457 1131 483
rect 1161 457 1209 541
rect 1239 457 1317 541
rect 1347 532 1377 541
rect 1411 532 1426 566
rect 1347 457 1426 532
rect 1456 573 1509 585
rect 1456 539 1467 573
rect 1501 539 1509 573
rect 1456 503 1509 539
rect 1456 469 1467 503
rect 1501 469 1509 503
rect 1456 457 1509 469
<< ndiffc >>
rect 63 141 97 175
rect 149 144 183 178
rect 307 144 341 178
rect 399 144 433 178
rect 499 106 533 140
rect 597 144 631 178
rect 706 142 740 176
rect 792 142 826 176
rect 888 131 922 165
rect 984 142 1018 176
rect 1070 142 1104 176
rect 1354 86 1388 120
rect 1440 86 1474 120
<< pdiffc >>
rect 35 570 69 604
rect 35 500 69 534
rect 132 548 166 582
rect 320 557 354 591
rect 415 557 449 591
rect 505 569 539 603
rect 595 557 629 591
rect 706 481 740 515
rect 792 483 826 517
rect 888 491 922 525
rect 984 483 1018 517
rect 1079 483 1113 517
rect 1377 532 1411 566
rect 1467 539 1501 573
rect 1467 469 1501 503
<< poly >>
rect 80 616 110 642
rect 188 616 218 642
rect 266 616 296 642
rect 374 616 404 642
rect 460 616 490 642
rect 554 616 584 642
rect 653 615 1347 645
rect 80 291 110 488
rect 188 405 218 532
rect 266 464 296 532
rect 266 448 332 464
rect 266 414 282 448
rect 316 414 332 448
rect 158 389 224 405
rect 158 355 174 389
rect 208 355 224 389
rect 158 339 224 355
rect 80 275 151 291
rect 80 241 101 275
rect 135 241 151 275
rect 80 225 151 241
rect 108 203 138 225
rect 194 203 224 339
rect 266 398 332 414
rect 266 203 296 398
rect 374 296 404 532
rect 460 480 490 532
rect 554 510 584 532
rect 653 510 683 615
rect 751 541 781 567
rect 837 541 867 567
rect 943 541 973 615
rect 1029 541 1059 567
rect 1131 541 1161 567
rect 1209 541 1239 567
rect 1317 541 1347 615
rect 1426 585 1456 611
rect 554 480 683 510
rect 446 464 512 480
rect 446 430 462 464
rect 496 430 512 464
rect 446 414 512 430
rect 338 280 404 296
rect 338 246 354 280
rect 388 246 404 280
rect 452 255 482 414
rect 554 366 584 480
rect 524 350 590 366
rect 524 316 540 350
rect 574 316 590 350
rect 524 300 590 316
rect 751 308 781 457
rect 837 401 867 457
rect 829 385 895 401
rect 829 351 845 385
rect 879 351 895 385
rect 829 335 895 351
rect 338 230 404 246
rect 352 203 382 230
rect 446 225 482 255
rect 446 203 476 225
rect 556 203 586 300
rect 687 292 781 308
rect 687 258 703 292
rect 737 258 781 292
rect 687 242 781 258
rect 751 203 781 242
rect 837 203 867 335
rect 943 203 973 457
rect 1029 255 1059 457
rect 1131 325 1161 457
rect 1209 425 1239 457
rect 1209 409 1275 425
rect 1209 375 1225 409
rect 1259 375 1275 409
rect 1209 359 1275 375
rect 1101 309 1167 325
rect 1101 275 1117 309
rect 1151 275 1167 309
rect 1101 259 1167 275
rect 1209 317 1245 359
rect 1023 225 1059 255
rect 1029 203 1059 225
rect 1115 203 1145 259
rect 1209 203 1239 317
rect 1317 311 1347 457
rect 1313 281 1353 311
rect 108 51 138 119
rect 194 93 224 119
rect 266 93 296 119
rect 352 93 382 119
rect 446 93 476 119
rect 1313 145 1343 281
rect 1426 239 1456 457
rect 1385 223 1456 239
rect 1385 189 1401 223
rect 1435 189 1456 223
rect 1385 167 1456 189
rect 1399 145 1429 167
rect 556 93 586 119
rect 751 93 781 119
rect 837 93 867 119
rect 943 93 973 119
rect 1029 51 1059 119
rect 1115 93 1145 119
rect 1209 93 1239 119
rect 108 21 1059 51
rect 1313 35 1343 61
rect 1399 35 1429 61
<< polycont >>
rect 282 414 316 448
rect 174 355 208 389
rect 101 241 135 275
rect 462 430 496 464
rect 354 246 388 280
rect 540 316 574 350
rect 845 351 879 385
rect 703 258 737 292
rect 1225 375 1259 409
rect 1117 275 1151 309
rect 1401 189 1435 223
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 17 604 85 615
rect 17 570 35 604
rect 69 570 85 604
rect 17 534 85 570
rect 17 500 35 534
rect 69 500 85 534
rect 119 582 178 649
rect 119 548 132 582
rect 166 548 178 582
rect 119 532 178 548
rect 212 591 365 607
rect 212 557 320 591
rect 354 557 365 591
rect 212 541 365 557
rect 399 591 455 607
rect 399 557 415 591
rect 449 557 455 591
rect 489 603 555 649
rect 489 569 505 603
rect 539 569 555 603
rect 489 566 555 569
rect 589 591 645 607
rect 17 191 65 500
rect 212 473 246 541
rect 399 532 455 557
rect 589 557 595 591
rect 629 557 645 591
rect 589 532 645 557
rect 399 498 645 532
rect 694 515 749 649
rect 106 439 246 473
rect 694 481 706 515
rect 740 481 749 515
rect 694 465 749 481
rect 783 517 838 533
rect 783 483 792 517
rect 826 483 838 517
rect 872 525 938 649
rect 1361 566 1427 649
rect 872 491 888 525
rect 922 491 938 525
rect 872 487 938 491
rect 972 517 1029 533
rect 280 448 462 464
rect 106 291 140 439
rect 280 414 282 448
rect 316 430 462 448
rect 496 430 660 464
rect 316 414 660 430
rect 783 453 838 483
rect 972 483 984 517
rect 1018 483 1029 517
rect 972 453 1029 483
rect 1063 517 1129 533
rect 1361 532 1377 566
rect 1411 532 1427 566
rect 1361 527 1427 532
rect 1461 573 1519 589
rect 1461 539 1467 573
rect 1501 539 1519 573
rect 1063 483 1079 517
rect 1113 493 1129 517
rect 1461 503 1519 539
rect 1113 483 1391 493
rect 1063 459 1391 483
rect 783 419 1029 453
rect 174 389 224 405
rect 280 398 660 414
rect 208 364 224 389
rect 626 385 660 398
rect 1202 409 1315 425
rect 1202 385 1225 409
rect 208 355 590 364
rect 174 350 590 355
rect 626 351 845 385
rect 879 375 1225 385
rect 1259 375 1315 409
rect 879 351 1315 375
rect 174 316 540 350
rect 574 316 590 350
rect 174 314 590 316
rect 99 275 140 291
rect 687 309 1167 317
rect 687 292 1117 309
rect 687 280 703 292
rect 99 241 101 275
rect 135 259 140 275
rect 135 241 304 259
rect 338 246 354 280
rect 388 258 703 280
rect 737 275 1117 292
rect 1151 275 1167 309
rect 737 273 1167 275
rect 737 258 758 273
rect 1101 259 1167 273
rect 388 246 758 258
rect 99 225 304 241
rect 690 226 758 246
rect 251 194 304 225
rect 17 175 99 191
rect 17 141 63 175
rect 97 141 99 175
rect 17 125 99 141
rect 133 178 199 191
rect 133 144 149 178
rect 183 144 199 178
rect 133 17 199 144
rect 251 178 349 194
rect 251 144 307 178
rect 341 144 349 178
rect 251 128 349 144
rect 383 178 647 212
rect 792 205 1028 239
rect 1225 238 1315 351
rect 1349 239 1391 459
rect 1461 469 1467 503
rect 1501 469 1519 503
rect 1461 281 1519 469
rect 383 144 399 178
rect 433 144 449 178
rect 583 144 597 178
rect 631 144 647 178
rect 383 128 449 144
rect 483 140 549 144
rect 483 106 499 140
rect 533 106 549 140
rect 583 128 647 144
rect 690 176 756 192
rect 690 142 706 176
rect 740 142 756 176
rect 483 17 549 106
rect 690 17 756 142
rect 792 176 838 205
rect 826 142 838 176
rect 972 176 1028 205
rect 1349 223 1435 239
rect 1349 204 1401 223
rect 792 126 838 142
rect 872 165 938 171
rect 872 131 888 165
rect 922 131 938 165
rect 872 17 938 131
rect 972 142 984 176
rect 1018 142 1028 176
rect 972 126 1028 142
rect 1062 189 1401 204
rect 1062 176 1435 189
rect 1062 142 1070 176
rect 1104 170 1435 176
rect 1104 167 1304 170
rect 1104 142 1120 167
rect 1062 126 1120 142
rect 1469 136 1519 281
rect 1338 120 1397 136
rect 1338 86 1354 120
rect 1388 86 1397 120
rect 1338 17 1397 86
rect 1431 120 1519 136
rect 1431 86 1440 120
rect 1474 86 1519 120
rect 1431 70 1519 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fa_0
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 1471 168 1505 202 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1471 390 1505 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1471 464 1505 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1471 538 1505 572 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2445140
string GDS_START 2433158
<< end >>
