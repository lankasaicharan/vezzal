magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 877 241 1151 263
rect 9 49 1151 241
rect 0 0 1152 49
<< scnmos >>
rect 88 47 118 215
rect 174 47 204 215
rect 260 47 290 215
rect 346 47 376 215
rect 440 47 470 215
rect 594 47 624 215
rect 680 47 710 215
rect 766 47 796 215
rect 956 69 986 237
rect 1042 69 1072 237
<< scpmoshvt >>
rect 88 367 118 619
rect 174 367 204 619
rect 260 367 290 619
rect 346 367 376 619
rect 536 367 566 619
rect 622 367 652 619
rect 708 367 738 619
rect 870 367 900 619
rect 956 367 986 619
rect 1042 367 1072 619
<< ndiff >>
rect 903 225 956 237
rect 35 203 88 215
rect 35 169 43 203
rect 77 169 88 203
rect 35 101 88 169
rect 35 67 43 101
rect 77 67 88 101
rect 35 47 88 67
rect 118 127 174 215
rect 118 93 129 127
rect 163 93 174 127
rect 118 47 174 93
rect 204 203 260 215
rect 204 169 215 203
rect 249 169 260 203
rect 204 101 260 169
rect 204 67 215 101
rect 249 67 260 101
rect 204 47 260 67
rect 290 127 346 215
rect 290 93 301 127
rect 335 93 346 127
rect 290 47 346 93
rect 376 203 440 215
rect 376 169 390 203
rect 424 169 440 203
rect 376 101 440 169
rect 376 67 390 101
rect 424 67 440 101
rect 376 47 440 67
rect 470 127 594 215
rect 470 93 481 127
rect 515 93 549 127
rect 583 93 594 127
rect 470 47 594 93
rect 624 203 680 215
rect 624 169 635 203
rect 669 169 680 203
rect 624 101 680 169
rect 624 67 635 101
rect 669 67 680 101
rect 624 47 680 67
rect 710 127 766 215
rect 710 93 721 127
rect 755 93 766 127
rect 710 47 766 93
rect 796 169 849 215
rect 796 135 807 169
rect 841 135 849 169
rect 796 47 849 135
rect 903 191 911 225
rect 945 191 956 225
rect 903 153 956 191
rect 903 119 911 153
rect 945 119 956 153
rect 903 69 956 119
rect 986 124 1042 237
rect 986 90 997 124
rect 1031 90 1042 124
rect 986 69 1042 90
rect 1072 208 1125 237
rect 1072 174 1083 208
rect 1117 174 1125 208
rect 1072 117 1125 174
rect 1072 83 1083 117
rect 1117 83 1125 117
rect 1072 69 1125 83
<< pdiff >>
rect 35 599 88 619
rect 35 565 43 599
rect 77 565 88 599
rect 35 510 88 565
rect 35 476 43 510
rect 77 476 88 510
rect 35 413 88 476
rect 35 379 43 413
rect 77 379 88 413
rect 35 367 88 379
rect 118 607 174 619
rect 118 573 129 607
rect 163 573 174 607
rect 118 518 174 573
rect 118 484 129 518
rect 163 484 174 518
rect 118 423 174 484
rect 118 389 129 423
rect 163 389 174 423
rect 118 367 174 389
rect 204 599 260 619
rect 204 565 215 599
rect 249 565 260 599
rect 204 510 260 565
rect 204 476 215 510
rect 249 476 260 510
rect 204 413 260 476
rect 204 379 215 413
rect 249 379 260 413
rect 204 367 260 379
rect 290 597 346 619
rect 290 563 301 597
rect 335 563 346 597
rect 290 511 346 563
rect 290 477 301 511
rect 335 477 346 511
rect 290 423 346 477
rect 290 389 301 423
rect 335 389 346 423
rect 290 367 346 389
rect 376 531 429 619
rect 376 497 387 531
rect 421 497 429 531
rect 376 413 429 497
rect 376 379 387 413
rect 421 379 429 413
rect 376 367 429 379
rect 483 531 536 619
rect 483 497 491 531
rect 525 497 536 531
rect 483 413 536 497
rect 483 379 491 413
rect 525 379 536 413
rect 483 367 536 379
rect 566 597 622 619
rect 566 563 577 597
rect 611 563 622 597
rect 566 521 622 563
rect 566 487 577 521
rect 611 487 622 521
rect 566 441 622 487
rect 566 407 577 441
rect 611 407 622 441
rect 566 367 622 407
rect 652 599 708 619
rect 652 565 663 599
rect 697 565 708 599
rect 652 510 708 565
rect 652 476 663 510
rect 697 476 708 510
rect 652 413 708 476
rect 652 379 663 413
rect 697 379 708 413
rect 652 367 708 379
rect 738 607 870 619
rect 738 573 749 607
rect 783 573 825 607
rect 859 573 870 607
rect 738 526 870 573
rect 738 492 749 526
rect 783 492 825 526
rect 859 492 870 526
rect 738 441 870 492
rect 738 407 749 441
rect 783 407 825 441
rect 859 407 870 441
rect 738 367 870 407
rect 900 599 956 619
rect 900 565 911 599
rect 945 565 956 599
rect 900 510 956 565
rect 900 476 911 510
rect 945 476 956 510
rect 900 413 956 476
rect 900 379 911 413
rect 945 379 956 413
rect 900 367 956 379
rect 986 607 1042 619
rect 986 573 997 607
rect 1031 573 1042 607
rect 986 526 1042 573
rect 986 492 997 526
rect 1031 492 1042 526
rect 986 445 1042 492
rect 986 411 997 445
rect 1031 411 1042 445
rect 986 367 1042 411
rect 1072 599 1125 619
rect 1072 565 1083 599
rect 1117 565 1125 599
rect 1072 510 1125 565
rect 1072 476 1083 510
rect 1117 476 1125 510
rect 1072 413 1125 476
rect 1072 379 1083 413
rect 1117 379 1125 413
rect 1072 367 1125 379
<< ndiffc >>
rect 43 169 77 203
rect 43 67 77 101
rect 129 93 163 127
rect 215 169 249 203
rect 215 67 249 101
rect 301 93 335 127
rect 390 169 424 203
rect 390 67 424 101
rect 481 93 515 127
rect 549 93 583 127
rect 635 169 669 203
rect 635 67 669 101
rect 721 93 755 127
rect 807 135 841 169
rect 911 191 945 225
rect 911 119 945 153
rect 997 90 1031 124
rect 1083 174 1117 208
rect 1083 83 1117 117
<< pdiffc >>
rect 43 565 77 599
rect 43 476 77 510
rect 43 379 77 413
rect 129 573 163 607
rect 129 484 163 518
rect 129 389 163 423
rect 215 565 249 599
rect 215 476 249 510
rect 215 379 249 413
rect 301 563 335 597
rect 301 477 335 511
rect 301 389 335 423
rect 387 497 421 531
rect 387 379 421 413
rect 491 497 525 531
rect 491 379 525 413
rect 577 563 611 597
rect 577 487 611 521
rect 577 407 611 441
rect 663 565 697 599
rect 663 476 697 510
rect 663 379 697 413
rect 749 573 783 607
rect 825 573 859 607
rect 749 492 783 526
rect 825 492 859 526
rect 749 407 783 441
rect 825 407 859 441
rect 911 565 945 599
rect 911 476 945 510
rect 911 379 945 413
rect 997 573 1031 607
rect 997 492 1031 526
rect 997 411 1031 445
rect 1083 565 1117 599
rect 1083 476 1117 510
rect 1083 379 1117 413
<< poly >>
rect 88 619 118 645
rect 174 619 204 645
rect 260 619 290 645
rect 346 619 376 645
rect 536 619 566 645
rect 622 619 652 645
rect 708 619 738 645
rect 870 619 900 645
rect 956 619 986 645
rect 1042 619 1072 645
rect 88 303 118 367
rect 174 303 204 367
rect 260 303 290 367
rect 346 303 376 367
rect 536 345 566 367
rect 622 345 652 367
rect 708 345 738 367
rect 870 345 900 367
rect 536 321 652 345
rect 440 315 652 321
rect 440 305 624 315
rect 55 287 204 303
rect 55 253 71 287
rect 105 253 139 287
rect 173 253 204 287
rect 55 237 204 253
rect 246 287 380 303
rect 246 253 262 287
rect 296 253 330 287
rect 364 253 380 287
rect 246 237 380 253
rect 440 271 484 305
rect 518 271 574 305
rect 608 271 624 305
rect 440 255 624 271
rect 694 287 900 345
rect 694 267 710 287
rect 88 215 118 237
rect 174 215 204 237
rect 260 215 290 237
rect 346 215 376 237
rect 440 215 470 255
rect 594 215 624 255
rect 680 253 710 267
rect 744 253 778 287
rect 812 270 900 287
rect 956 325 986 367
rect 1042 325 1072 367
rect 956 309 1127 325
rect 956 275 1077 309
rect 1111 275 1127 309
rect 812 253 868 270
rect 680 237 868 253
rect 956 259 1127 275
rect 956 237 986 259
rect 1042 237 1072 259
rect 680 215 710 237
rect 766 215 796 237
rect 88 21 118 47
rect 174 21 204 47
rect 260 21 290 47
rect 346 21 376 47
rect 440 21 470 47
rect 594 21 624 47
rect 680 21 710 47
rect 766 21 796 47
rect 956 43 986 69
rect 1042 43 1072 69
<< polycont >>
rect 71 253 105 287
rect 139 253 173 287
rect 262 253 296 287
rect 330 253 364 287
rect 484 271 518 305
rect 574 271 608 305
rect 710 253 744 287
rect 778 253 812 287
rect 1077 275 1111 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 27 599 79 615
rect 27 565 43 599
rect 77 565 79 599
rect 27 510 79 565
rect 27 476 43 510
rect 77 476 79 510
rect 27 413 79 476
rect 27 379 43 413
rect 77 379 79 413
rect 113 607 179 649
rect 113 573 129 607
rect 163 573 179 607
rect 113 518 179 573
rect 113 484 129 518
rect 163 484 179 518
rect 113 423 179 484
rect 113 389 129 423
rect 163 389 179 423
rect 213 599 251 615
rect 213 565 215 599
rect 249 565 251 599
rect 213 510 251 565
rect 213 476 215 510
rect 249 476 251 510
rect 213 413 251 476
rect 27 355 79 379
rect 213 379 215 413
rect 249 379 251 413
rect 285 597 627 615
rect 285 563 301 597
rect 335 581 577 597
rect 335 563 351 581
rect 285 511 351 563
rect 561 563 577 581
rect 611 563 627 597
rect 285 477 301 511
rect 335 477 351 511
rect 285 423 351 477
rect 285 389 301 423
rect 335 389 351 423
rect 385 531 437 547
rect 385 497 387 531
rect 421 497 437 531
rect 385 413 437 497
rect 213 355 251 379
rect 385 379 387 413
rect 421 379 437 413
rect 385 355 437 379
rect 27 321 437 355
rect 475 531 527 547
rect 475 497 491 531
rect 525 497 527 531
rect 475 413 527 497
rect 475 379 491 413
rect 525 379 527 413
rect 561 521 627 563
rect 561 487 577 521
rect 611 487 627 521
rect 561 441 627 487
rect 561 407 577 441
rect 611 407 627 441
rect 661 599 699 615
rect 661 565 663 599
rect 697 565 699 599
rect 661 510 699 565
rect 661 476 663 510
rect 697 476 699 510
rect 661 413 699 476
rect 475 373 527 379
rect 661 379 663 413
rect 697 379 699 413
rect 733 607 875 649
rect 733 573 749 607
rect 783 573 825 607
rect 859 573 875 607
rect 733 526 875 573
rect 733 492 749 526
rect 783 492 825 526
rect 859 492 875 526
rect 733 441 875 492
rect 733 407 749 441
rect 783 407 825 441
rect 859 407 875 441
rect 909 599 947 615
rect 909 565 911 599
rect 945 565 947 599
rect 909 510 947 565
rect 909 476 911 510
rect 945 476 947 510
rect 909 413 947 476
rect 661 373 699 379
rect 909 379 911 413
rect 945 379 947 413
rect 981 607 1047 649
rect 981 573 997 607
rect 1031 573 1047 607
rect 981 526 1047 573
rect 981 492 997 526
rect 1031 492 1047 526
rect 981 445 1047 492
rect 981 411 997 445
rect 1031 411 1047 445
rect 1081 599 1133 615
rect 1081 565 1083 599
rect 1117 565 1133 599
rect 1081 510 1133 565
rect 1081 476 1083 510
rect 1117 476 1133 510
rect 1081 413 1133 476
rect 909 377 947 379
rect 1081 379 1083 413
rect 1117 379 1133 413
rect 1081 377 1133 379
rect 909 373 1133 377
rect 475 343 1133 373
rect 475 339 1025 343
rect 468 287 484 305
rect 31 253 71 287
rect 105 253 139 287
rect 173 253 189 287
rect 31 237 189 253
rect 223 253 262 287
rect 296 253 330 287
rect 364 253 380 287
rect 223 237 380 253
rect 414 271 484 287
rect 518 271 574 305
rect 608 271 641 305
rect 414 237 641 271
rect 694 287 857 303
rect 694 253 710 287
rect 744 253 778 287
rect 812 253 857 287
rect 694 237 857 253
rect 891 225 1025 339
rect 1059 275 1077 309
rect 1111 275 1135 309
rect 1059 242 1135 275
rect 27 169 43 203
rect 77 169 215 203
rect 249 169 390 203
rect 424 169 635 203
rect 669 169 857 203
rect 27 101 79 169
rect 27 67 43 101
rect 77 67 79 101
rect 27 51 79 67
rect 113 127 179 135
rect 113 93 129 127
rect 163 93 179 127
rect 113 17 179 93
rect 213 101 251 169
rect 213 67 215 101
rect 249 67 251 101
rect 213 51 251 67
rect 285 127 351 135
rect 285 93 301 127
rect 335 93 351 127
rect 285 17 351 93
rect 385 101 431 169
rect 385 67 390 101
rect 424 67 431 101
rect 385 51 431 67
rect 465 127 600 135
rect 465 93 481 127
rect 515 93 549 127
rect 583 93 600 127
rect 465 17 600 93
rect 634 101 671 169
rect 805 135 807 169
rect 841 135 857 169
rect 634 67 635 101
rect 669 67 671 101
rect 634 51 671 67
rect 705 127 771 135
rect 705 93 721 127
rect 755 93 771 127
rect 805 119 857 135
rect 891 191 911 225
rect 945 208 1025 225
rect 945 191 1083 208
rect 891 174 1083 191
rect 1117 174 1133 208
rect 891 153 961 174
rect 891 119 911 153
rect 945 119 961 153
rect 995 124 1045 140
rect 705 85 771 93
rect 995 90 997 124
rect 1031 90 1045 124
rect 995 85 1045 90
rect 705 51 1045 85
rect 1079 117 1133 174
rect 1079 83 1083 117
rect 1117 83 1133 117
rect 1079 67 1133 83
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o311ai_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1416736
string GDS_START 1405770
<< end >>
