magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 199 210 758 248
rect 1 49 758 210
rect 0 0 768 49
<< scpmos >>
rect 81 424 117 592
rect 276 368 312 592
rect 366 368 402 592
rect 561 368 597 592
rect 651 368 687 592
<< nmoslvt >>
rect 84 74 114 184
rect 282 74 312 222
rect 396 74 426 222
rect 474 74 504 222
rect 645 74 675 222
<< ndiff >>
rect 225 210 282 222
rect 27 146 84 184
rect 27 112 39 146
rect 73 112 84 146
rect 27 74 84 112
rect 114 146 171 184
rect 114 112 125 146
rect 159 112 171 146
rect 114 74 171 112
rect 225 176 237 210
rect 271 176 282 210
rect 225 120 282 176
rect 225 86 237 120
rect 271 86 282 120
rect 225 74 282 86
rect 312 152 396 222
rect 312 118 337 152
rect 371 118 396 152
rect 312 74 396 118
rect 426 74 474 222
rect 504 191 645 222
rect 504 157 515 191
rect 549 157 600 191
rect 634 157 645 191
rect 504 74 645 157
rect 675 186 732 222
rect 675 152 686 186
rect 720 152 732 186
rect 675 116 732 152
rect 675 82 686 116
rect 720 82 732 116
rect 675 74 732 82
<< pdiff >>
rect 27 580 81 592
rect 27 546 37 580
rect 71 546 81 580
rect 27 470 81 546
rect 27 436 37 470
rect 71 436 81 470
rect 27 424 81 436
rect 117 580 169 592
rect 117 546 127 580
rect 161 546 169 580
rect 117 470 169 546
rect 117 436 127 470
rect 161 436 169 470
rect 117 424 169 436
rect 223 580 276 592
rect 223 546 232 580
rect 266 546 276 580
rect 223 497 276 546
rect 223 463 232 497
rect 266 463 276 497
rect 223 414 276 463
rect 223 380 232 414
rect 266 380 276 414
rect 223 368 276 380
rect 312 580 366 592
rect 312 546 322 580
rect 356 546 366 580
rect 312 508 366 546
rect 312 474 322 508
rect 356 474 366 508
rect 312 368 366 474
rect 402 580 454 592
rect 402 546 412 580
rect 446 546 454 580
rect 402 508 454 546
rect 402 474 412 508
rect 446 474 454 508
rect 402 368 454 474
rect 508 531 561 592
rect 508 497 517 531
rect 551 497 561 531
rect 508 440 561 497
rect 508 406 517 440
rect 551 406 561 440
rect 508 368 561 406
rect 597 531 651 592
rect 597 497 607 531
rect 641 497 651 531
rect 597 414 651 497
rect 597 380 607 414
rect 641 380 651 414
rect 597 368 651 380
rect 687 580 741 592
rect 687 546 697 580
rect 731 546 741 580
rect 687 497 741 546
rect 687 463 697 497
rect 731 463 741 497
rect 687 414 741 463
rect 687 380 697 414
rect 731 380 741 414
rect 687 368 741 380
<< ndiffc >>
rect 39 112 73 146
rect 125 112 159 146
rect 237 176 271 210
rect 237 86 271 120
rect 337 118 371 152
rect 515 157 549 191
rect 600 157 634 191
rect 686 152 720 186
rect 686 82 720 116
<< pdiffc >>
rect 37 546 71 580
rect 37 436 71 470
rect 127 546 161 580
rect 127 436 161 470
rect 232 546 266 580
rect 232 463 266 497
rect 232 380 266 414
rect 322 546 356 580
rect 322 474 356 508
rect 412 546 446 580
rect 412 474 446 508
rect 517 497 551 531
rect 517 406 551 440
rect 607 497 641 531
rect 607 380 641 414
rect 697 546 731 580
rect 697 463 731 497
rect 697 380 731 414
<< poly >>
rect 81 592 117 618
rect 276 592 312 618
rect 366 592 402 618
rect 561 592 597 618
rect 651 592 687 618
rect 81 371 117 424
rect 44 355 114 371
rect 44 321 60 355
rect 94 321 114 355
rect 44 287 114 321
rect 44 253 60 287
rect 94 267 114 287
rect 276 267 312 368
rect 366 336 402 368
rect 561 336 597 368
rect 360 320 426 336
rect 360 286 376 320
rect 410 286 426 320
rect 507 320 591 336
rect 507 300 523 320
rect 360 270 426 286
rect 94 253 312 267
rect 44 237 312 253
rect 84 184 114 237
rect 282 222 312 237
rect 396 222 426 270
rect 474 286 523 300
rect 557 286 591 320
rect 651 310 687 368
rect 474 270 591 286
rect 645 294 745 310
rect 474 222 504 270
rect 645 260 695 294
rect 729 260 745 294
rect 645 244 745 260
rect 645 222 675 244
rect 84 48 114 74
rect 282 48 312 74
rect 396 48 426 74
rect 474 48 504 74
rect 645 48 675 74
<< polycont >>
rect 60 321 94 355
rect 60 253 94 287
rect 376 286 410 320
rect 523 286 557 320
rect 695 260 729 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 21 580 71 649
rect 21 546 37 580
rect 21 470 71 546
rect 21 436 37 470
rect 21 420 71 436
rect 111 580 178 596
rect 111 546 127 580
rect 161 546 178 580
rect 111 470 178 546
rect 111 436 127 470
rect 161 436 178 470
rect 111 420 178 436
rect 25 355 110 371
rect 25 321 60 355
rect 94 321 110 355
rect 25 287 110 321
rect 25 253 60 287
rect 94 253 110 287
rect 25 236 110 253
rect 144 304 178 420
rect 216 580 266 596
rect 216 546 232 580
rect 216 497 266 546
rect 216 463 232 497
rect 216 424 266 463
rect 306 580 372 649
rect 306 546 322 580
rect 356 546 372 580
rect 306 508 372 546
rect 306 474 322 508
rect 356 474 372 508
rect 306 458 372 474
rect 412 581 747 615
rect 412 580 462 581
rect 446 546 462 580
rect 681 580 747 581
rect 412 508 462 546
rect 446 474 462 508
rect 412 458 462 474
rect 501 531 567 547
rect 501 497 517 531
rect 551 497 567 531
rect 501 440 567 497
rect 501 424 517 440
rect 216 414 517 424
rect 216 380 232 414
rect 266 406 517 414
rect 551 406 567 440
rect 266 390 567 406
rect 607 531 645 547
rect 641 497 645 531
rect 607 414 645 497
rect 216 364 266 380
rect 641 380 645 414
rect 360 320 426 336
rect 360 304 376 320
rect 144 286 376 304
rect 410 286 426 320
rect 144 270 426 286
rect 505 320 573 356
rect 505 286 523 320
rect 557 286 573 320
rect 505 270 573 286
rect 144 181 178 270
rect 23 146 73 181
rect 23 112 39 146
rect 23 17 73 112
rect 109 146 178 181
rect 109 112 125 146
rect 159 112 178 146
rect 109 81 178 112
rect 221 210 455 236
rect 221 176 237 210
rect 271 202 455 210
rect 607 207 645 380
rect 681 546 697 580
rect 731 546 747 580
rect 681 497 747 546
rect 681 463 697 497
rect 731 463 747 497
rect 681 414 747 463
rect 681 380 697 414
rect 731 380 747 414
rect 681 364 747 380
rect 679 294 745 310
rect 679 260 695 294
rect 729 260 745 294
rect 679 236 745 260
rect 271 176 287 202
rect 221 120 287 176
rect 221 86 237 120
rect 271 86 287 120
rect 221 70 287 86
rect 321 152 387 168
rect 321 118 337 152
rect 371 118 387 152
rect 321 17 387 118
rect 421 104 455 202
rect 499 191 645 207
rect 499 157 515 191
rect 549 157 600 191
rect 634 157 645 191
rect 499 141 645 157
rect 679 186 736 202
rect 679 152 686 186
rect 720 152 736 186
rect 679 116 736 152
rect 679 104 686 116
rect 421 82 686 104
rect 720 82 736 116
rect 421 70 736 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2i_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 1712082
string GDS_START 1705246
<< end >>
