magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 332 1094 704
<< pwell >>
rect 103 248 570 256
rect 103 49 1035 248
rect 0 0 1056 49
<< scpmos >>
rect 176 392 212 592
rect 254 392 290 592
rect 476 368 512 592
rect 566 368 602 592
rect 656 368 692 592
rect 746 368 782 592
rect 836 368 872 592
rect 926 368 962 592
<< nmoslvt >>
rect 182 102 212 230
rect 277 102 307 230
rect 375 82 405 230
rect 461 82 491 230
rect 668 74 698 222
rect 754 74 784 222
rect 840 74 870 222
rect 926 74 956 222
<< ndiff >>
rect 129 218 182 230
rect 129 184 137 218
rect 171 184 182 218
rect 129 150 182 184
rect 129 116 137 150
rect 171 116 182 150
rect 129 102 182 116
rect 212 218 277 230
rect 212 184 227 218
rect 261 184 277 218
rect 212 148 277 184
rect 212 114 227 148
rect 261 114 277 148
rect 212 102 277 114
rect 307 166 375 230
rect 307 132 330 166
rect 364 132 375 166
rect 307 102 375 132
rect 322 82 375 102
rect 405 214 461 230
rect 405 180 416 214
rect 450 180 461 214
rect 405 128 461 180
rect 405 94 416 128
rect 450 94 461 128
rect 405 82 461 94
rect 491 146 544 230
rect 491 112 502 146
rect 536 112 544 146
rect 491 82 544 112
rect 615 120 668 222
rect 615 86 623 120
rect 657 86 668 120
rect 615 74 668 86
rect 698 207 754 222
rect 698 173 709 207
rect 743 173 754 207
rect 698 74 754 173
rect 784 210 840 222
rect 784 176 795 210
rect 829 176 840 210
rect 784 120 840 176
rect 784 86 795 120
rect 829 86 840 120
rect 784 74 840 86
rect 870 136 926 222
rect 870 102 881 136
rect 915 102 926 136
rect 870 74 926 102
rect 956 210 1009 222
rect 956 176 967 210
rect 1001 176 1009 210
rect 956 120 1009 176
rect 956 86 967 120
rect 1001 86 1009 120
rect 956 74 1009 86
<< pdiff >>
rect 124 580 176 592
rect 124 546 132 580
rect 166 546 176 580
rect 124 509 176 546
rect 124 475 132 509
rect 166 475 176 509
rect 124 438 176 475
rect 124 404 132 438
rect 166 404 176 438
rect 124 392 176 404
rect 212 392 254 592
rect 290 580 342 592
rect 290 546 300 580
rect 334 546 342 580
rect 290 510 342 546
rect 290 476 300 510
rect 334 476 342 510
rect 290 440 342 476
rect 290 406 300 440
rect 334 406 342 440
rect 290 392 342 406
rect 424 580 476 592
rect 424 546 432 580
rect 466 546 476 580
rect 424 497 476 546
rect 424 463 432 497
rect 466 463 476 497
rect 424 414 476 463
rect 424 380 432 414
rect 466 380 476 414
rect 424 368 476 380
rect 512 531 566 592
rect 512 497 522 531
rect 556 497 566 531
rect 512 414 566 497
rect 512 380 522 414
rect 556 380 566 414
rect 512 368 566 380
rect 602 580 656 592
rect 602 546 612 580
rect 646 546 656 580
rect 602 497 656 546
rect 602 463 612 497
rect 646 463 656 497
rect 602 414 656 463
rect 602 380 612 414
rect 646 380 656 414
rect 602 368 656 380
rect 692 580 746 592
rect 692 546 702 580
rect 736 546 746 580
rect 692 508 746 546
rect 692 474 702 508
rect 736 474 746 508
rect 692 368 746 474
rect 782 580 836 592
rect 782 546 792 580
rect 826 546 836 580
rect 782 510 836 546
rect 782 476 792 510
rect 826 476 836 510
rect 782 440 836 476
rect 782 406 792 440
rect 826 406 836 440
rect 782 368 836 406
rect 872 580 926 592
rect 872 546 882 580
rect 916 546 926 580
rect 872 508 926 546
rect 872 474 882 508
rect 916 474 926 508
rect 872 368 926 474
rect 962 580 1014 592
rect 962 546 972 580
rect 1006 546 1014 580
rect 962 497 1014 546
rect 962 463 972 497
rect 1006 463 1014 497
rect 962 414 1014 463
rect 962 380 972 414
rect 1006 380 1014 414
rect 962 368 1014 380
<< ndiffc >>
rect 137 184 171 218
rect 137 116 171 150
rect 227 184 261 218
rect 227 114 261 148
rect 330 132 364 166
rect 416 180 450 214
rect 416 94 450 128
rect 502 112 536 146
rect 623 86 657 120
rect 709 173 743 207
rect 795 176 829 210
rect 795 86 829 120
rect 881 102 915 136
rect 967 176 1001 210
rect 967 86 1001 120
<< pdiffc >>
rect 132 546 166 580
rect 132 475 166 509
rect 132 404 166 438
rect 300 546 334 580
rect 300 476 334 510
rect 300 406 334 440
rect 432 546 466 580
rect 432 463 466 497
rect 432 380 466 414
rect 522 497 556 531
rect 522 380 556 414
rect 612 546 646 580
rect 612 463 646 497
rect 612 380 646 414
rect 702 546 736 580
rect 702 474 736 508
rect 792 546 826 580
rect 792 476 826 510
rect 792 406 826 440
rect 882 546 916 580
rect 882 474 916 508
rect 972 546 1006 580
rect 972 463 1006 497
rect 972 380 1006 414
<< poly >>
rect 176 592 212 618
rect 254 592 290 618
rect 476 592 512 618
rect 566 592 602 618
rect 656 592 692 618
rect 746 592 782 618
rect 836 592 872 618
rect 926 592 962 618
rect 176 245 212 392
rect 254 356 290 392
rect 254 340 320 356
rect 254 306 270 340
rect 304 306 320 340
rect 476 330 512 368
rect 566 330 602 368
rect 254 290 320 306
rect 375 314 602 330
rect 182 230 212 245
rect 277 230 307 290
rect 375 280 391 314
rect 425 300 602 314
rect 656 330 692 368
rect 746 330 782 368
rect 656 314 782 330
rect 425 280 491 300
rect 375 264 491 280
rect 656 280 697 314
rect 731 294 782 314
rect 836 336 872 368
rect 926 336 962 368
rect 836 320 962 336
rect 731 280 784 294
rect 656 264 784 280
rect 836 286 852 320
rect 886 286 962 320
rect 836 270 962 286
rect 375 230 405 264
rect 461 230 491 264
rect 21 107 87 123
rect 21 73 37 107
rect 71 87 87 107
rect 182 87 212 102
rect 71 73 212 87
rect 277 76 307 102
rect 668 222 698 264
rect 754 222 784 264
rect 840 222 870 270
rect 926 222 956 270
rect 21 57 212 73
rect 375 56 405 82
rect 461 56 491 82
rect 668 48 698 74
rect 754 48 784 74
rect 840 48 870 74
rect 926 48 956 74
<< polycont >>
rect 270 306 304 340
rect 391 280 425 314
rect 697 280 731 314
rect 852 286 886 320
rect 37 73 71 107
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 116 580 182 649
rect 116 546 132 580
rect 166 546 182 580
rect 116 509 182 546
rect 116 475 132 509
rect 166 475 182 509
rect 116 438 182 475
rect 116 404 132 438
rect 166 404 182 438
rect 116 388 182 404
rect 284 580 382 596
rect 284 546 300 580
rect 334 546 382 580
rect 284 510 382 546
rect 284 476 300 510
rect 334 476 382 510
rect 284 440 382 476
rect 284 406 300 440
rect 334 406 382 440
rect 284 390 382 406
rect 217 340 314 356
rect 217 306 270 340
rect 304 306 314 340
rect 217 290 314 306
rect 348 330 382 390
rect 416 581 646 615
rect 416 580 466 581
rect 416 546 432 580
rect 596 580 646 581
rect 416 497 466 546
rect 416 463 432 497
rect 416 414 466 463
rect 416 380 432 414
rect 416 364 466 380
rect 505 531 556 547
rect 505 497 522 531
rect 505 414 556 497
rect 505 380 522 414
rect 348 314 441 330
rect 348 280 391 314
rect 425 280 441 314
rect 348 264 441 280
rect 505 282 556 380
rect 596 546 612 580
rect 596 497 646 546
rect 596 463 612 497
rect 596 424 646 463
rect 686 580 752 649
rect 686 546 702 580
rect 736 546 752 580
rect 686 508 752 546
rect 686 474 702 508
rect 736 474 752 508
rect 686 458 752 474
rect 792 580 826 596
rect 792 510 826 546
rect 792 440 826 476
rect 866 580 932 649
rect 866 546 882 580
rect 916 546 932 580
rect 866 508 932 546
rect 866 474 882 508
rect 916 474 932 508
rect 866 458 932 474
rect 972 580 1022 596
rect 1006 546 1022 580
rect 972 497 1022 546
rect 1006 463 1022 497
rect 596 414 792 424
rect 596 380 612 414
rect 646 406 792 414
rect 972 424 1022 463
rect 826 414 1022 424
rect 826 406 972 414
rect 646 390 972 406
rect 596 364 646 380
rect 1006 380 1022 414
rect 972 364 1022 380
rect 681 314 747 356
rect 348 256 382 264
rect 121 218 171 234
rect 121 184 137 218
rect 121 150 171 184
rect 21 107 87 134
rect 21 73 37 107
rect 71 73 87 107
rect 21 57 87 73
rect 121 116 137 150
rect 121 17 171 116
rect 207 222 382 256
rect 505 230 647 282
rect 681 280 697 314
rect 731 280 747 314
rect 681 264 747 280
rect 793 320 935 356
rect 793 286 852 320
rect 886 286 935 320
rect 793 270 935 286
rect 207 218 266 222
rect 207 184 227 218
rect 261 184 266 218
rect 416 214 759 230
rect 207 148 266 184
rect 207 114 227 148
rect 261 114 266 148
rect 207 98 266 114
rect 314 166 380 188
rect 314 132 330 166
rect 364 132 380 166
rect 314 17 380 132
rect 450 207 759 214
rect 450 196 709 207
rect 416 128 450 180
rect 693 173 709 196
rect 743 173 759 207
rect 416 78 450 94
rect 486 146 552 162
rect 693 154 759 173
rect 795 210 1017 236
rect 829 202 967 210
rect 486 112 502 146
rect 536 112 552 146
rect 795 120 829 176
rect 951 176 967 202
rect 1001 176 1017 210
rect 486 17 552 112
rect 607 86 623 120
rect 657 86 795 120
rect 607 70 829 86
rect 865 136 915 168
rect 865 102 881 136
rect 865 17 915 102
rect 951 120 1017 176
rect 951 86 967 120
rect 1001 86 1017 120
rect 951 70 1017 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2bb2oi_2
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 2008118
string GDS_START 1999424
<< end >>
