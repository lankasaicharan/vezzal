magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 1182 241 1628 259
rect 22 49 1628 241
rect 0 0 1632 49
<< scnmos >>
rect 101 47 131 215
rect 187 47 217 215
rect 273 47 303 215
rect 359 47 389 215
rect 481 47 511 215
rect 567 47 597 215
rect 813 47 843 215
rect 899 47 929 215
rect 985 47 1015 215
rect 1071 47 1101 215
rect 1261 65 1291 233
rect 1347 65 1377 233
rect 1433 65 1463 233
rect 1519 65 1549 233
<< scpmoshvt >>
rect 137 367 167 619
rect 223 367 253 619
rect 309 367 339 619
rect 395 367 425 619
rect 481 367 511 619
rect 567 367 597 619
rect 857 367 887 619
rect 943 367 973 619
rect 1029 367 1059 619
rect 1127 367 1157 619
rect 1213 367 1243 619
rect 1315 367 1345 619
rect 1431 367 1461 619
rect 1517 367 1547 619
<< ndiff >>
rect 48 173 101 215
rect 48 139 56 173
rect 90 139 101 173
rect 48 93 101 139
rect 48 59 56 93
rect 90 59 101 93
rect 48 47 101 59
rect 131 203 187 215
rect 131 169 142 203
rect 176 169 187 203
rect 131 101 187 169
rect 131 67 142 101
rect 176 67 187 101
rect 131 47 187 67
rect 217 173 273 215
rect 217 139 228 173
rect 262 139 273 173
rect 217 89 273 139
rect 217 55 228 89
rect 262 55 273 89
rect 217 47 273 55
rect 303 175 359 215
rect 303 141 314 175
rect 348 141 359 175
rect 303 101 359 141
rect 303 67 314 101
rect 348 67 359 101
rect 303 47 359 67
rect 389 177 481 215
rect 389 143 418 177
rect 452 143 481 177
rect 389 93 481 143
rect 389 59 418 93
rect 452 59 481 93
rect 389 47 481 59
rect 511 175 567 215
rect 511 141 522 175
rect 556 141 567 175
rect 511 89 567 141
rect 511 55 522 89
rect 556 55 567 89
rect 511 47 567 55
rect 597 97 650 215
rect 597 63 608 97
rect 642 63 650 97
rect 597 47 650 63
rect 760 175 813 215
rect 760 141 768 175
rect 802 141 813 175
rect 760 47 813 141
rect 843 92 899 215
rect 843 58 854 92
rect 888 58 899 92
rect 843 47 899 58
rect 929 169 985 215
rect 929 135 940 169
rect 974 135 985 169
rect 929 101 985 135
rect 929 67 940 101
rect 974 67 985 101
rect 929 47 985 67
rect 1015 173 1071 215
rect 1015 139 1026 173
rect 1060 139 1071 173
rect 1015 47 1071 139
rect 1101 165 1154 215
rect 1101 131 1112 165
rect 1146 131 1154 165
rect 1101 93 1154 131
rect 1101 59 1112 93
rect 1146 59 1154 93
rect 1208 151 1261 233
rect 1208 117 1216 151
rect 1250 117 1261 151
rect 1208 65 1261 117
rect 1291 225 1347 233
rect 1291 191 1302 225
rect 1336 191 1347 225
rect 1291 154 1347 191
rect 1291 120 1302 154
rect 1336 120 1347 154
rect 1291 65 1347 120
rect 1377 225 1433 233
rect 1377 191 1388 225
rect 1422 191 1433 225
rect 1377 111 1433 191
rect 1377 77 1388 111
rect 1422 77 1433 111
rect 1377 65 1433 77
rect 1463 179 1519 233
rect 1463 145 1474 179
rect 1508 145 1519 179
rect 1463 107 1519 145
rect 1463 73 1474 107
rect 1508 73 1519 107
rect 1463 65 1519 73
rect 1549 221 1602 233
rect 1549 187 1560 221
rect 1594 187 1602 221
rect 1549 111 1602 187
rect 1549 77 1560 111
rect 1594 77 1602 111
rect 1549 65 1602 77
rect 1101 47 1154 59
<< pdiff >>
rect 84 607 137 619
rect 84 573 92 607
rect 126 573 137 607
rect 84 533 137 573
rect 84 499 92 533
rect 126 499 137 533
rect 84 453 137 499
rect 84 419 92 453
rect 126 419 137 453
rect 84 367 137 419
rect 167 599 223 619
rect 167 565 178 599
rect 212 565 223 599
rect 167 508 223 565
rect 167 474 178 508
rect 212 474 223 508
rect 167 413 223 474
rect 167 379 178 413
rect 212 379 223 413
rect 167 367 223 379
rect 253 607 309 619
rect 253 573 264 607
rect 298 573 309 607
rect 253 533 309 573
rect 253 499 264 533
rect 298 499 309 533
rect 253 453 309 499
rect 253 419 264 453
rect 298 419 309 453
rect 253 367 309 419
rect 339 599 395 619
rect 339 565 350 599
rect 384 565 395 599
rect 339 508 395 565
rect 339 474 350 508
rect 384 474 395 508
rect 339 413 395 474
rect 339 379 350 413
rect 384 379 395 413
rect 339 367 395 379
rect 425 607 481 619
rect 425 573 436 607
rect 470 573 481 607
rect 425 508 481 573
rect 425 474 436 508
rect 470 474 481 508
rect 425 413 481 474
rect 425 379 436 413
rect 470 379 481 413
rect 425 367 481 379
rect 511 599 567 619
rect 511 565 522 599
rect 556 565 567 599
rect 511 515 567 565
rect 511 481 522 515
rect 556 481 567 515
rect 511 434 567 481
rect 511 400 522 434
rect 556 400 567 434
rect 511 367 567 400
rect 597 607 650 619
rect 597 573 608 607
rect 642 573 650 607
rect 597 492 650 573
rect 597 458 608 492
rect 642 458 650 492
rect 597 367 650 458
rect 804 599 857 619
rect 804 565 812 599
rect 846 565 857 599
rect 804 518 857 565
rect 804 484 812 518
rect 846 484 857 518
rect 804 434 857 484
rect 804 400 812 434
rect 846 400 857 434
rect 804 367 857 400
rect 887 607 943 619
rect 887 573 898 607
rect 932 573 943 607
rect 887 492 943 573
rect 887 458 898 492
rect 932 458 943 492
rect 887 367 943 458
rect 973 599 1029 619
rect 973 565 984 599
rect 1018 565 1029 599
rect 973 518 1029 565
rect 973 484 984 518
rect 1018 484 1029 518
rect 973 434 1029 484
rect 973 400 984 434
rect 1018 400 1029 434
rect 973 367 1029 400
rect 1059 607 1127 619
rect 1059 573 1070 607
rect 1104 573 1127 607
rect 1059 492 1127 573
rect 1059 458 1070 492
rect 1104 458 1127 492
rect 1059 367 1127 458
rect 1157 599 1213 619
rect 1157 565 1168 599
rect 1202 565 1213 599
rect 1157 516 1213 565
rect 1157 482 1168 516
rect 1202 482 1213 516
rect 1157 434 1213 482
rect 1157 400 1168 434
rect 1202 400 1213 434
rect 1157 367 1213 400
rect 1243 531 1315 619
rect 1243 497 1257 531
rect 1291 497 1315 531
rect 1243 436 1315 497
rect 1243 402 1257 436
rect 1291 402 1315 436
rect 1243 367 1315 402
rect 1345 599 1431 619
rect 1345 565 1371 599
rect 1405 565 1431 599
rect 1345 493 1431 565
rect 1345 459 1371 493
rect 1405 459 1431 493
rect 1345 367 1431 459
rect 1461 543 1517 619
rect 1461 509 1472 543
rect 1506 509 1517 543
rect 1461 424 1517 509
rect 1461 390 1472 424
rect 1506 390 1517 424
rect 1461 367 1517 390
rect 1547 599 1600 619
rect 1547 565 1558 599
rect 1592 565 1600 599
rect 1547 516 1600 565
rect 1547 482 1558 516
rect 1592 482 1600 516
rect 1547 434 1600 482
rect 1547 400 1558 434
rect 1592 400 1600 434
rect 1547 367 1600 400
<< ndiffc >>
rect 56 139 90 173
rect 56 59 90 93
rect 142 169 176 203
rect 142 67 176 101
rect 228 139 262 173
rect 228 55 262 89
rect 314 141 348 175
rect 314 67 348 101
rect 418 143 452 177
rect 418 59 452 93
rect 522 141 556 175
rect 522 55 556 89
rect 608 63 642 97
rect 768 141 802 175
rect 854 58 888 92
rect 940 135 974 169
rect 940 67 974 101
rect 1026 139 1060 173
rect 1112 131 1146 165
rect 1112 59 1146 93
rect 1216 117 1250 151
rect 1302 191 1336 225
rect 1302 120 1336 154
rect 1388 191 1422 225
rect 1388 77 1422 111
rect 1474 145 1508 179
rect 1474 73 1508 107
rect 1560 187 1594 221
rect 1560 77 1594 111
<< pdiffc >>
rect 92 573 126 607
rect 92 499 126 533
rect 92 419 126 453
rect 178 565 212 599
rect 178 474 212 508
rect 178 379 212 413
rect 264 573 298 607
rect 264 499 298 533
rect 264 419 298 453
rect 350 565 384 599
rect 350 474 384 508
rect 350 379 384 413
rect 436 573 470 607
rect 436 474 470 508
rect 436 379 470 413
rect 522 565 556 599
rect 522 481 556 515
rect 522 400 556 434
rect 608 573 642 607
rect 608 458 642 492
rect 812 565 846 599
rect 812 484 846 518
rect 812 400 846 434
rect 898 573 932 607
rect 898 458 932 492
rect 984 565 1018 599
rect 984 484 1018 518
rect 984 400 1018 434
rect 1070 573 1104 607
rect 1070 458 1104 492
rect 1168 565 1202 599
rect 1168 482 1202 516
rect 1168 400 1202 434
rect 1257 497 1291 531
rect 1257 402 1291 436
rect 1371 565 1405 599
rect 1371 459 1405 493
rect 1472 509 1506 543
rect 1472 390 1506 424
rect 1558 565 1592 599
rect 1558 482 1592 516
rect 1558 400 1592 434
<< poly >>
rect 137 619 167 645
rect 223 619 253 645
rect 309 619 339 645
rect 395 619 425 645
rect 481 619 511 645
rect 567 619 597 645
rect 857 619 887 645
rect 943 619 973 645
rect 1029 619 1059 645
rect 1127 619 1157 645
rect 1213 619 1243 645
rect 1315 619 1345 645
rect 1431 619 1461 645
rect 1517 619 1547 645
rect 137 329 167 367
rect 223 329 253 367
rect 309 329 339 367
rect 395 329 425 367
rect 481 335 511 367
rect 567 335 597 367
rect 857 345 887 367
rect 943 345 973 367
rect 101 313 439 329
rect 101 279 117 313
rect 151 279 185 313
rect 219 279 253 313
rect 287 279 321 313
rect 355 279 389 313
rect 423 279 439 313
rect 101 263 439 279
rect 481 319 597 335
rect 481 285 547 319
rect 581 285 597 319
rect 481 269 597 285
rect 700 319 973 345
rect 700 285 716 319
rect 750 285 784 319
rect 818 315 973 319
rect 1029 321 1059 367
rect 1127 321 1157 367
rect 1213 335 1243 367
rect 1315 335 1345 367
rect 1431 335 1461 367
rect 1517 335 1547 367
rect 818 285 929 315
rect 700 269 929 285
rect 101 215 131 263
rect 187 215 217 263
rect 273 215 303 263
rect 359 215 389 263
rect 481 215 511 269
rect 567 215 597 269
rect 813 215 843 269
rect 899 215 929 269
rect 1029 305 1167 321
rect 1029 271 1117 305
rect 1151 271 1167 305
rect 1029 267 1167 271
rect 1213 319 1389 335
rect 1213 285 1339 319
rect 1373 285 1389 319
rect 1431 319 1549 335
rect 1431 305 1487 319
rect 1213 269 1389 285
rect 1433 285 1487 305
rect 1521 285 1549 319
rect 1433 269 1549 285
rect 985 237 1167 267
rect 985 215 1015 237
rect 1071 215 1101 237
rect 1261 233 1291 269
rect 1347 233 1377 269
rect 1433 233 1463 269
rect 1519 233 1549 269
rect 101 21 131 47
rect 187 21 217 47
rect 273 21 303 47
rect 359 21 389 47
rect 481 21 511 47
rect 567 21 597 47
rect 813 21 843 47
rect 899 21 929 47
rect 985 21 1015 47
rect 1071 21 1101 47
rect 1261 39 1291 65
rect 1347 39 1377 65
rect 1433 39 1463 65
rect 1519 39 1549 65
<< polycont >>
rect 117 279 151 313
rect 185 279 219 313
rect 253 279 287 313
rect 321 279 355 313
rect 389 279 423 313
rect 547 285 581 319
rect 716 285 750 319
rect 784 285 818 319
rect 1117 271 1151 305
rect 1339 285 1373 319
rect 1487 285 1521 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 76 607 142 649
rect 76 573 92 607
rect 126 573 142 607
rect 76 533 142 573
rect 76 499 92 533
rect 126 499 142 533
rect 76 453 142 499
rect 76 419 92 453
rect 126 419 142 453
rect 176 599 214 615
rect 176 565 178 599
rect 212 565 214 599
rect 176 508 214 565
rect 176 474 178 508
rect 212 474 214 508
rect 176 413 214 474
rect 248 607 314 649
rect 248 573 264 607
rect 298 573 314 607
rect 248 533 314 573
rect 248 499 264 533
rect 298 499 314 533
rect 248 453 314 499
rect 248 419 264 453
rect 298 419 314 453
rect 348 599 394 615
rect 348 565 350 599
rect 384 565 394 599
rect 348 508 394 565
rect 348 474 350 508
rect 384 474 394 508
rect 176 385 178 413
rect 20 379 178 385
rect 212 385 214 413
rect 348 413 394 474
rect 348 385 350 413
rect 212 379 350 385
rect 384 379 394 413
rect 20 351 394 379
rect 428 607 474 649
rect 428 573 436 607
rect 470 573 474 607
rect 428 508 474 573
rect 428 474 436 508
rect 470 474 474 508
rect 428 413 474 474
rect 428 379 436 413
rect 470 379 474 413
rect 508 599 558 615
rect 508 565 522 599
rect 556 565 558 599
rect 508 515 558 565
rect 508 481 522 515
rect 556 481 558 515
rect 508 434 558 481
rect 592 607 658 649
rect 592 573 608 607
rect 642 573 658 607
rect 592 492 658 573
rect 592 458 608 492
rect 642 458 658 492
rect 592 452 658 458
rect 773 599 848 615
rect 773 565 812 599
rect 846 565 848 599
rect 773 518 848 565
rect 773 484 812 518
rect 846 484 848 518
rect 508 400 522 434
rect 556 418 558 434
rect 773 434 848 484
rect 882 607 948 649
rect 882 573 898 607
rect 932 573 948 607
rect 882 492 948 573
rect 882 458 898 492
rect 932 458 948 492
rect 882 452 948 458
rect 982 599 1020 615
rect 982 565 984 599
rect 1018 565 1020 599
rect 982 518 1020 565
rect 982 484 984 518
rect 1018 484 1020 518
rect 773 418 812 434
rect 556 400 812 418
rect 846 418 848 434
rect 982 434 1020 484
rect 1054 607 1120 649
rect 1054 573 1070 607
rect 1104 573 1120 607
rect 1054 492 1120 573
rect 1054 458 1070 492
rect 1104 458 1120 492
rect 1054 452 1120 458
rect 1154 599 1608 615
rect 1154 565 1168 599
rect 1202 581 1371 599
rect 1202 565 1217 581
rect 1154 516 1217 565
rect 1355 565 1371 581
rect 1405 581 1558 599
rect 1405 565 1421 581
rect 1154 482 1168 516
rect 1202 482 1217 516
rect 982 418 984 434
rect 846 400 984 418
rect 1018 418 1020 434
rect 1154 434 1217 482
rect 1154 418 1168 434
rect 1018 400 1168 418
rect 1202 400 1217 434
rect 508 384 1217 400
rect 1251 531 1307 547
rect 1251 497 1257 531
rect 1291 497 1307 531
rect 1251 436 1307 497
rect 1355 493 1421 565
rect 1556 565 1558 581
rect 1592 565 1608 599
rect 1355 459 1371 493
rect 1405 459 1421 493
rect 1355 454 1421 459
rect 1456 543 1522 547
rect 1456 509 1472 543
rect 1506 509 1522 543
rect 1251 402 1257 436
rect 1291 420 1307 436
rect 1456 424 1522 509
rect 1456 420 1472 424
rect 1291 402 1472 420
rect 1251 390 1472 402
rect 1506 390 1522 424
rect 1251 384 1522 390
rect 1556 516 1608 565
rect 1556 482 1558 516
rect 1592 482 1608 516
rect 1556 434 1608 482
rect 1556 400 1558 434
rect 1592 400 1608 434
rect 1556 384 1608 400
rect 428 363 474 379
rect 20 243 67 351
rect 508 319 649 350
rect 101 313 439 317
rect 101 279 117 313
rect 151 279 185 313
rect 219 279 253 313
rect 287 279 321 313
rect 355 279 389 313
rect 423 279 439 313
rect 508 285 547 319
rect 581 285 649 319
rect 691 319 841 350
rect 691 285 716 319
rect 750 285 784 319
rect 818 285 841 319
rect 1036 305 1217 350
rect 1036 287 1117 305
rect 691 283 841 285
rect 101 277 439 279
rect 405 249 439 277
rect 1085 271 1117 287
rect 1151 271 1217 305
rect 870 249 1051 253
rect 20 209 364 243
rect 405 235 1051 249
rect 1251 235 1287 384
rect 1323 319 1409 350
rect 1323 285 1339 319
rect 1373 285 1409 319
rect 1471 319 1601 350
rect 1471 285 1487 319
rect 1521 285 1601 319
rect 405 225 1352 235
rect 405 219 1302 225
rect 405 215 904 219
rect 140 203 178 209
rect 40 173 106 175
rect 40 139 56 173
rect 90 139 106 173
rect 40 93 106 139
rect 40 59 56 93
rect 90 59 106 93
rect 40 17 106 59
rect 140 169 142 203
rect 176 169 178 203
rect 312 175 364 209
rect 1013 201 1302 219
rect 140 101 178 169
rect 140 67 142 101
rect 176 67 178 101
rect 140 51 178 67
rect 212 173 278 175
rect 212 139 228 173
rect 262 139 278 173
rect 212 89 278 139
rect 212 55 228 89
rect 262 55 278 89
rect 212 17 278 55
rect 312 141 314 175
rect 348 141 364 175
rect 312 101 364 141
rect 312 67 314 101
rect 348 67 364 101
rect 312 51 364 67
rect 402 177 468 181
rect 402 143 418 177
rect 452 143 468 177
rect 402 93 468 143
rect 402 59 418 93
rect 452 59 468 93
rect 402 17 468 59
rect 506 175 716 181
rect 938 179 979 185
rect 506 141 522 175
rect 556 147 716 175
rect 556 141 572 147
rect 506 89 572 141
rect 506 55 522 89
rect 556 55 572 89
rect 506 51 572 55
rect 606 97 648 113
rect 606 63 608 97
rect 642 63 648 97
rect 606 17 648 63
rect 682 103 716 147
rect 752 175 979 179
rect 752 141 768 175
rect 802 169 979 175
rect 802 141 940 169
rect 752 137 940 141
rect 938 135 940 137
rect 974 135 979 169
rect 682 92 904 103
rect 682 58 854 92
rect 888 58 904 92
rect 682 51 904 58
rect 938 101 979 135
rect 1013 173 1062 201
rect 1013 139 1026 173
rect 1060 139 1062 173
rect 1286 191 1302 201
rect 1336 191 1352 225
rect 1013 123 1062 139
rect 1096 165 1162 167
rect 1096 131 1112 165
rect 1146 131 1162 165
rect 938 67 940 101
rect 974 89 979 101
rect 1096 93 1162 131
rect 1096 89 1112 93
rect 974 67 1112 89
rect 938 59 1112 67
rect 1146 59 1162 93
rect 938 51 1162 59
rect 1200 151 1252 167
rect 1200 117 1216 151
rect 1250 117 1252 151
rect 1286 154 1352 191
rect 1286 120 1302 154
rect 1336 120 1352 154
rect 1286 119 1352 120
rect 1386 225 1610 249
rect 1386 191 1388 225
rect 1422 221 1610 225
rect 1422 215 1560 221
rect 1422 191 1424 215
rect 1200 85 1252 117
rect 1386 111 1424 191
rect 1558 187 1560 215
rect 1594 187 1610 221
rect 1386 85 1388 111
rect 1200 77 1388 85
rect 1422 77 1424 111
rect 1200 51 1424 77
rect 1458 179 1524 181
rect 1458 145 1474 179
rect 1508 145 1524 179
rect 1458 107 1524 145
rect 1458 73 1474 107
rect 1508 73 1524 107
rect 1458 17 1524 73
rect 1558 111 1610 187
rect 1558 77 1560 111
rect 1594 77 1610 111
rect 1558 51 1610 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a32o_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2050362
string GDS_START 2036916
<< end >>
