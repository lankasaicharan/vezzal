magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 23 49 904 243
rect 0 0 960 49
<< scnmos >>
rect 106 133 136 217
rect 242 49 272 217
rect 328 49 358 217
rect 414 49 444 217
rect 500 49 530 217
rect 615 49 645 217
rect 687 49 717 217
rect 795 49 825 217
<< scpmoshvt >>
rect 106 367 136 451
rect 242 367 272 619
rect 328 367 358 619
rect 414 367 444 619
rect 500 367 530 619
rect 601 367 631 619
rect 687 367 717 619
rect 802 367 832 619
<< ndiff >>
rect 49 192 106 217
rect 49 158 57 192
rect 91 158 106 192
rect 49 133 106 158
rect 136 165 242 217
rect 136 133 197 165
rect 189 131 197 133
rect 231 131 242 165
rect 189 95 242 131
rect 189 61 197 95
rect 231 61 242 95
rect 189 49 242 61
rect 272 205 328 217
rect 272 171 283 205
rect 317 171 328 205
rect 272 101 328 171
rect 272 67 283 101
rect 317 67 328 101
rect 272 49 328 67
rect 358 174 414 217
rect 358 140 369 174
rect 403 140 414 174
rect 358 95 414 140
rect 358 61 369 95
rect 403 61 414 95
rect 358 49 414 61
rect 444 205 500 217
rect 444 171 455 205
rect 489 171 500 205
rect 444 101 500 171
rect 444 67 455 101
rect 489 67 500 101
rect 444 49 500 67
rect 530 161 615 217
rect 530 127 555 161
rect 589 127 615 161
rect 530 91 615 127
rect 530 57 555 91
rect 589 57 615 91
rect 530 49 615 57
rect 645 49 687 217
rect 717 49 795 217
rect 825 205 878 217
rect 825 171 836 205
rect 870 171 878 205
rect 825 101 878 171
rect 825 67 836 101
rect 870 67 878 101
rect 825 49 878 67
<< pdiff >>
rect 189 576 242 619
rect 189 542 197 576
rect 231 542 242 576
rect 189 451 242 542
rect 49 426 106 451
rect 49 392 57 426
rect 91 392 106 426
rect 49 367 106 392
rect 136 367 242 451
rect 272 413 328 619
rect 272 379 283 413
rect 317 379 328 413
rect 272 367 328 379
rect 358 576 414 619
rect 358 542 369 576
rect 403 542 414 576
rect 358 367 414 542
rect 444 413 500 619
rect 444 379 455 413
rect 489 379 500 413
rect 444 367 500 379
rect 530 598 601 619
rect 530 564 541 598
rect 575 564 601 598
rect 530 367 601 564
rect 631 436 687 619
rect 631 402 642 436
rect 676 402 687 436
rect 631 367 687 402
rect 717 598 802 619
rect 717 564 728 598
rect 762 564 802 598
rect 717 367 802 564
rect 832 599 885 619
rect 832 565 843 599
rect 877 565 885 599
rect 832 506 885 565
rect 832 472 843 506
rect 877 472 885 506
rect 832 413 885 472
rect 832 379 843 413
rect 877 379 885 413
rect 832 367 885 379
<< ndiffc >>
rect 57 158 91 192
rect 197 131 231 165
rect 197 61 231 95
rect 283 171 317 205
rect 283 67 317 101
rect 369 140 403 174
rect 369 61 403 95
rect 455 171 489 205
rect 455 67 489 101
rect 555 127 589 161
rect 555 57 589 91
rect 836 171 870 205
rect 836 67 870 101
<< pdiffc >>
rect 197 542 231 576
rect 57 392 91 426
rect 283 379 317 413
rect 369 542 403 576
rect 455 379 489 413
rect 541 564 575 598
rect 642 402 676 436
rect 728 564 762 598
rect 843 565 877 599
rect 843 472 877 506
rect 843 379 877 413
<< poly >>
rect 242 619 272 645
rect 328 619 358 645
rect 414 619 444 645
rect 500 619 530 645
rect 601 619 631 645
rect 687 619 717 645
rect 802 619 832 645
rect 106 451 136 477
rect 106 305 136 367
rect 242 335 272 367
rect 328 335 358 367
rect 414 335 444 367
rect 500 335 530 367
rect 601 335 631 367
rect 687 335 717 367
rect 802 335 832 367
rect 242 319 537 335
rect 106 289 177 305
rect 106 255 127 289
rect 161 255 177 289
rect 106 239 177 255
rect 242 285 283 319
rect 317 285 351 319
rect 385 285 419 319
rect 453 285 487 319
rect 521 285 537 319
rect 242 269 537 285
rect 579 319 645 335
rect 579 285 595 319
rect 629 285 645 319
rect 579 269 645 285
rect 106 217 136 239
rect 242 217 272 269
rect 328 217 358 269
rect 414 217 444 269
rect 500 217 530 269
rect 615 217 645 269
rect 687 319 753 335
rect 687 285 703 319
rect 737 285 753 319
rect 802 319 868 335
rect 802 299 818 319
rect 687 269 753 285
rect 795 285 818 299
rect 852 285 868 319
rect 795 269 868 285
rect 687 217 717 269
rect 795 217 825 269
rect 106 107 136 133
rect 242 23 272 49
rect 328 23 358 49
rect 414 23 444 49
rect 500 23 530 49
rect 615 23 645 49
rect 687 23 717 49
rect 795 23 825 49
<< polycont >>
rect 127 255 161 289
rect 283 285 317 319
rect 351 285 385 319
rect 419 285 453 319
rect 487 285 521 319
rect 595 285 629 319
rect 703 285 737 319
rect 818 285 852 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 181 576 247 649
rect 181 542 197 576
rect 231 542 247 576
rect 181 531 247 542
rect 353 576 419 649
rect 353 542 369 576
rect 403 542 419 576
rect 525 598 591 649
rect 525 564 541 598
rect 575 564 591 598
rect 525 556 591 564
rect 712 598 778 649
rect 712 564 728 598
rect 762 564 778 598
rect 712 556 778 564
rect 841 599 938 615
rect 841 565 843 599
rect 877 565 938 599
rect 353 531 419 542
rect 453 497 807 522
rect 41 486 807 497
rect 41 463 491 486
rect 41 426 91 463
rect 525 436 680 452
rect 41 392 57 426
rect 41 192 91 392
rect 41 158 57 192
rect 41 140 91 158
rect 125 289 161 424
rect 125 255 127 289
rect 125 94 161 255
rect 197 413 489 429
rect 197 379 283 413
rect 317 379 455 413
rect 197 363 489 379
rect 525 402 642 436
rect 676 402 680 436
rect 525 386 680 402
rect 197 249 231 363
rect 525 319 559 386
rect 267 285 283 319
rect 317 285 351 319
rect 385 285 419 319
rect 453 285 487 319
rect 521 285 559 319
rect 197 215 491 249
rect 273 205 319 215
rect 195 165 239 181
rect 195 131 197 165
rect 231 131 239 165
rect 195 95 239 131
rect 195 61 197 95
rect 231 61 239 95
rect 195 17 239 61
rect 273 171 283 205
rect 317 171 319 205
rect 453 205 491 215
rect 273 101 319 171
rect 273 67 283 101
rect 317 67 319 101
rect 273 51 319 67
rect 353 174 419 179
rect 353 140 369 174
rect 403 140 419 174
rect 353 95 419 140
rect 353 61 369 95
rect 403 61 419 95
rect 353 17 419 61
rect 453 171 455 205
rect 489 171 491 205
rect 525 233 559 285
rect 593 319 651 350
rect 593 285 595 319
rect 629 285 651 319
rect 593 269 651 285
rect 685 319 739 350
rect 685 285 703 319
rect 737 285 739 319
rect 685 269 739 285
rect 773 329 807 486
rect 841 506 938 565
rect 841 472 843 506
rect 877 472 938 506
rect 841 413 938 472
rect 841 379 843 413
rect 877 379 938 413
rect 841 363 938 379
rect 773 319 868 329
rect 773 285 818 319
rect 852 285 868 319
rect 773 267 868 285
rect 904 233 938 363
rect 525 205 938 233
rect 525 199 836 205
rect 453 101 491 171
rect 666 171 836 199
rect 870 171 938 205
rect 453 67 455 101
rect 489 67 491 101
rect 453 51 491 67
rect 539 161 605 165
rect 539 127 555 161
rect 589 127 605 161
rect 539 91 605 127
rect 539 57 555 91
rect 589 57 605 91
rect 539 17 605 57
rect 666 101 938 171
rect 666 67 836 101
rect 870 67 938 101
rect 666 51 938 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and3b_4
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6402480
string GDS_START 6394780
<< end >>
