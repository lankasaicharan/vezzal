magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 36 49 669 195
rect 0 0 672 49
<< scnmos >>
rect 115 85 145 169
rect 201 85 231 169
rect 287 85 317 169
rect 365 85 395 169
rect 560 85 590 169
<< scpmoshvt >>
rect 80 481 110 609
rect 158 481 188 609
rect 244 481 274 609
rect 330 481 360 609
rect 560 367 590 495
<< ndiff >>
rect 62 144 115 169
rect 62 110 70 144
rect 104 110 115 144
rect 62 85 115 110
rect 145 144 201 169
rect 145 110 156 144
rect 190 110 201 144
rect 145 85 201 110
rect 231 136 287 169
rect 231 102 242 136
rect 276 102 287 136
rect 231 85 287 102
rect 317 85 365 169
rect 395 135 560 169
rect 395 101 410 135
rect 444 101 513 135
rect 547 101 560 135
rect 395 85 560 101
rect 590 144 643 169
rect 590 110 601 144
rect 635 110 643 144
rect 590 85 643 110
<< pdiff >>
rect 27 597 80 609
rect 27 563 35 597
rect 69 563 80 597
rect 27 527 80 563
rect 27 493 35 527
rect 69 493 80 527
rect 27 481 80 493
rect 110 481 158 609
rect 188 597 244 609
rect 188 563 199 597
rect 233 563 244 597
rect 188 527 244 563
rect 188 493 199 527
rect 233 493 244 527
rect 188 481 244 493
rect 274 597 330 609
rect 274 563 285 597
rect 319 563 330 597
rect 274 527 330 563
rect 274 493 285 527
rect 319 493 330 527
rect 274 481 330 493
rect 360 591 413 609
rect 360 557 371 591
rect 405 557 413 591
rect 360 481 413 557
rect 507 483 560 495
rect 507 449 515 483
rect 549 449 560 483
rect 507 413 560 449
rect 507 379 515 413
rect 549 379 560 413
rect 507 367 560 379
rect 590 483 643 495
rect 590 449 601 483
rect 635 449 643 483
rect 590 413 643 449
rect 590 379 601 413
rect 635 379 643 413
rect 590 367 643 379
<< ndiffc >>
rect 70 110 104 144
rect 156 110 190 144
rect 242 102 276 136
rect 410 101 444 135
rect 513 101 547 135
rect 601 110 635 144
<< pdiffc >>
rect 35 563 69 597
rect 35 493 69 527
rect 199 563 233 597
rect 199 493 233 527
rect 285 563 319 597
rect 285 493 319 527
rect 371 557 405 591
rect 515 449 549 483
rect 515 379 549 413
rect 601 449 635 483
rect 601 379 635 413
<< poly >>
rect 80 609 110 635
rect 158 609 188 635
rect 244 609 274 635
rect 330 609 360 635
rect 560 495 590 521
rect 80 371 110 481
rect 158 449 188 481
rect 244 449 274 481
rect 158 419 274 449
rect 41 355 145 371
rect 41 321 57 355
rect 91 321 145 355
rect 41 287 145 321
rect 41 253 57 287
rect 91 253 145 287
rect 41 237 145 253
rect 115 169 145 237
rect 201 276 274 419
rect 330 370 360 481
rect 322 354 395 370
rect 322 320 338 354
rect 372 320 395 354
rect 322 304 395 320
rect 201 242 217 276
rect 251 256 274 276
rect 251 242 317 256
rect 201 226 317 242
rect 201 169 231 226
rect 287 169 317 226
rect 365 169 395 304
rect 443 309 509 325
rect 443 275 459 309
rect 493 275 509 309
rect 443 241 509 275
rect 443 207 459 241
rect 493 221 509 241
rect 560 221 590 367
rect 493 207 590 221
rect 443 191 590 207
rect 560 169 590 191
rect 115 59 145 85
rect 201 59 231 85
rect 287 59 317 85
rect 365 59 395 85
rect 560 59 590 85
<< polycont >>
rect 57 321 91 355
rect 57 253 91 287
rect 338 320 372 354
rect 217 242 251 276
rect 459 275 493 309
rect 459 207 493 241
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 19 597 85 613
rect 19 563 35 597
rect 69 563 85 597
rect 19 527 85 563
rect 19 493 35 527
rect 69 493 85 527
rect 19 439 85 493
rect 183 597 242 649
rect 183 563 199 597
rect 233 563 242 597
rect 183 527 242 563
rect 183 493 199 527
rect 233 493 242 527
rect 183 477 242 493
rect 276 597 328 613
rect 276 563 285 597
rect 319 563 328 597
rect 276 527 328 563
rect 362 591 407 649
rect 362 557 371 591
rect 405 557 407 591
rect 362 541 407 557
rect 276 493 285 527
rect 319 507 328 527
rect 441 533 651 567
rect 441 507 475 533
rect 319 493 475 507
rect 276 473 475 493
rect 509 483 563 499
rect 509 449 515 483
rect 549 449 563 483
rect 19 405 475 439
rect 41 355 388 371
rect 41 321 57 355
rect 91 354 388 355
rect 91 321 338 354
rect 41 320 338 321
rect 372 320 388 354
rect 41 313 388 320
rect 41 287 91 313
rect 41 253 57 287
rect 41 237 91 253
rect 125 276 270 279
rect 125 242 217 276
rect 251 242 270 276
rect 304 242 388 313
rect 441 325 475 405
rect 509 413 563 449
rect 509 379 515 413
rect 549 379 563 413
rect 509 363 563 379
rect 597 483 651 533
rect 597 449 601 483
rect 635 449 651 483
rect 597 413 651 449
rect 597 379 601 413
rect 635 379 651 413
rect 597 363 651 379
rect 441 309 495 325
rect 441 275 459 309
rect 493 275 495 309
rect 441 241 495 275
rect 441 208 459 241
rect 146 207 459 208
rect 493 207 495 241
rect 146 174 495 207
rect 54 144 112 160
rect 54 110 70 144
rect 104 110 112 144
rect 54 17 112 110
rect 146 144 192 174
rect 146 110 156 144
rect 190 110 192 144
rect 529 140 563 363
rect 146 79 192 110
rect 226 136 292 140
rect 226 102 242 136
rect 276 102 292 136
rect 226 17 292 102
rect 394 135 563 140
rect 394 101 410 135
rect 444 101 513 135
rect 547 101 563 135
rect 394 82 563 101
rect 597 144 651 160
rect 597 110 601 144
rect 635 110 651 144
rect 597 17 651 110
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xor2_0
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2201340
string GDS_START 2195104
<< end >>
