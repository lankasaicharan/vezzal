magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 749 165
rect 0 0 768 49
<< scnmos >>
rect 84 55 114 139
rect 156 55 186 139
rect 242 55 272 139
rect 320 55 350 139
rect 406 55 436 139
rect 478 55 508 139
rect 564 55 594 139
rect 636 55 666 139
<< scpmoshvt >>
rect 94 409 144 609
rect 202 409 252 609
rect 308 409 358 609
rect 526 419 576 619
rect 632 419 682 619
<< ndiff >>
rect 27 115 84 139
rect 27 81 39 115
rect 73 81 84 115
rect 27 55 84 81
rect 114 55 156 139
rect 186 114 242 139
rect 186 80 197 114
rect 231 80 242 114
rect 186 55 242 80
rect 272 55 320 139
rect 350 115 406 139
rect 350 81 361 115
rect 395 81 406 115
rect 350 55 406 81
rect 436 55 478 139
rect 508 101 564 139
rect 508 67 519 101
rect 553 67 564 101
rect 508 55 564 67
rect 594 55 636 139
rect 666 115 723 139
rect 666 81 677 115
rect 711 81 723 115
rect 666 55 723 81
<< pdiff >>
rect 37 597 94 609
rect 37 563 49 597
rect 83 563 94 597
rect 37 526 94 563
rect 37 492 49 526
rect 83 492 94 526
rect 37 455 94 492
rect 37 421 49 455
rect 83 421 94 455
rect 37 409 94 421
rect 144 597 202 609
rect 144 563 155 597
rect 189 563 202 597
rect 144 512 202 563
rect 144 478 155 512
rect 189 478 202 512
rect 144 409 202 478
rect 252 597 308 609
rect 252 563 263 597
rect 297 563 308 597
rect 252 512 308 563
rect 252 478 263 512
rect 297 478 308 512
rect 252 409 308 478
rect 358 527 415 609
rect 358 493 369 527
rect 403 493 415 527
rect 358 455 415 493
rect 358 421 369 455
rect 403 421 415 455
rect 358 409 415 421
rect 469 597 526 619
rect 469 563 481 597
rect 515 563 526 597
rect 469 473 526 563
rect 469 439 481 473
rect 515 439 526 473
rect 469 419 526 439
rect 576 607 632 619
rect 576 573 587 607
rect 621 573 632 607
rect 576 473 632 573
rect 576 439 587 473
rect 621 439 632 473
rect 576 419 632 439
rect 682 597 739 619
rect 682 563 693 597
rect 727 563 739 597
rect 682 465 739 563
rect 682 431 693 465
rect 727 431 739 465
rect 682 419 739 431
<< ndiffc >>
rect 39 81 73 115
rect 197 80 231 114
rect 361 81 395 115
rect 519 67 553 101
rect 677 81 711 115
<< pdiffc >>
rect 49 563 83 597
rect 49 492 83 526
rect 49 421 83 455
rect 155 563 189 597
rect 155 478 189 512
rect 263 563 297 597
rect 263 478 297 512
rect 369 493 403 527
rect 369 421 403 455
rect 481 563 515 597
rect 481 439 515 473
rect 587 573 621 607
rect 587 439 621 473
rect 693 563 727 597
rect 693 431 727 465
<< poly >>
rect 94 609 144 635
rect 202 609 252 635
rect 308 609 358 635
rect 526 619 576 645
rect 632 619 682 645
rect 94 313 144 409
rect 202 322 252 409
rect 308 394 358 409
rect 308 364 457 394
rect 526 387 576 419
rect 84 297 154 313
rect 84 263 104 297
rect 138 263 154 297
rect 84 229 154 263
rect 202 306 271 322
rect 202 272 221 306
rect 255 272 271 306
rect 202 256 271 272
rect 84 195 104 229
rect 138 208 154 229
rect 138 195 186 208
rect 84 178 186 195
rect 84 139 114 178
rect 156 139 186 178
rect 241 184 271 256
rect 319 300 385 316
rect 319 266 335 300
rect 369 266 385 300
rect 319 250 385 266
rect 241 154 272 184
rect 242 139 272 154
rect 320 139 350 250
rect 427 227 457 364
rect 499 371 576 387
rect 499 337 515 371
rect 549 337 576 371
rect 499 321 576 337
rect 632 285 682 419
rect 632 273 667 285
rect 601 257 667 273
rect 601 237 617 257
rect 427 211 516 227
rect 427 191 466 211
rect 406 177 466 191
rect 500 177 516 211
rect 406 161 516 177
rect 564 223 617 237
rect 651 223 667 257
rect 564 207 667 223
rect 406 139 436 161
rect 478 139 508 161
rect 564 139 594 207
rect 636 139 666 207
rect 84 29 114 55
rect 156 29 186 55
rect 242 29 272 55
rect 320 29 350 55
rect 406 29 436 55
rect 478 29 508 55
rect 564 29 594 55
rect 636 29 666 55
<< polycont >>
rect 104 263 138 297
rect 221 272 255 306
rect 104 195 138 229
rect 335 266 369 300
rect 515 337 549 371
rect 466 177 500 211
rect 617 223 651 257
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 18 597 99 613
rect 18 563 49 597
rect 83 563 99 597
rect 18 526 99 563
rect 18 492 49 526
rect 83 492 99 526
rect 18 455 99 492
rect 139 597 205 649
rect 139 563 155 597
rect 189 563 205 597
rect 139 512 205 563
rect 139 478 155 512
rect 189 478 205 512
rect 139 462 205 478
rect 247 597 531 613
rect 247 563 263 597
rect 297 579 481 597
rect 297 563 313 579
rect 247 512 313 563
rect 465 563 481 579
rect 515 563 531 597
rect 247 478 263 512
rect 297 478 313 512
rect 247 462 313 478
rect 353 527 419 543
rect 353 493 369 527
rect 403 493 419 527
rect 18 421 49 455
rect 83 421 99 455
rect 353 455 419 493
rect 353 426 369 455
rect 18 405 99 421
rect 135 421 369 426
rect 403 421 419 455
rect 465 473 531 563
rect 465 439 481 473
rect 515 439 531 473
rect 465 423 531 439
rect 571 607 637 649
rect 571 573 587 607
rect 621 573 637 607
rect 571 473 637 573
rect 571 439 587 473
rect 621 439 637 473
rect 571 423 637 439
rect 677 597 743 613
rect 677 563 693 597
rect 727 563 743 597
rect 677 465 743 563
rect 677 431 693 465
rect 727 431 743 465
rect 18 143 52 405
rect 135 392 419 421
rect 677 415 743 431
rect 135 313 169 392
rect 499 371 565 387
rect 88 297 169 313
rect 88 263 104 297
rect 138 263 169 297
rect 88 229 169 263
rect 205 306 271 356
rect 499 344 515 371
rect 205 272 221 306
rect 255 272 271 306
rect 205 256 271 272
rect 319 337 515 344
rect 549 337 565 371
rect 319 310 565 337
rect 319 300 385 310
rect 319 266 335 300
rect 369 266 385 300
rect 319 250 385 266
rect 601 257 667 356
rect 88 195 104 229
rect 138 213 169 229
rect 138 195 411 213
rect 88 179 411 195
rect 18 115 89 143
rect 18 81 39 115
rect 73 81 89 115
rect 18 53 89 81
rect 181 114 247 143
rect 181 80 197 114
rect 231 80 247 114
rect 181 17 247 80
rect 345 115 411 179
rect 450 211 516 227
rect 450 177 466 211
rect 500 177 516 211
rect 601 223 617 257
rect 651 223 667 257
rect 601 207 667 223
rect 450 171 516 177
rect 709 171 743 415
rect 450 137 743 171
rect 345 81 361 115
rect 395 81 411 115
rect 661 115 727 137
rect 345 53 411 81
rect 503 67 519 101
rect 553 67 569 101
rect 503 17 569 67
rect 661 81 677 115
rect 711 81 727 115
rect 661 53 727 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21bo_lp
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3736890
string GDS_START 3730242
<< end >>
