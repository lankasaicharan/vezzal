magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 4 49 1044 241
rect 0 0 1056 49
<< scnmos >>
rect 83 47 113 215
rect 169 47 199 215
rect 255 47 285 215
rect 341 47 371 215
rect 435 47 465 215
rect 521 47 551 215
rect 675 47 705 215
rect 761 47 791 215
rect 935 131 965 215
<< scpmoshvt >>
rect 83 367 113 619
rect 169 367 199 619
rect 255 367 285 619
rect 341 367 371 619
rect 449 367 479 619
rect 521 367 551 619
rect 629 367 659 619
rect 737 367 767 619
rect 946 525 976 609
<< ndiff >>
rect 30 167 83 215
rect 30 133 38 167
rect 72 133 83 167
rect 30 93 83 133
rect 30 59 38 93
rect 72 59 83 93
rect 30 47 83 59
rect 113 203 169 215
rect 113 169 124 203
rect 158 169 169 203
rect 113 101 169 169
rect 113 67 124 101
rect 158 67 169 101
rect 113 47 169 67
rect 199 89 255 215
rect 199 55 210 89
rect 244 55 255 89
rect 199 47 255 55
rect 285 147 341 215
rect 285 113 296 147
rect 330 113 341 147
rect 285 47 341 113
rect 371 165 435 215
rect 371 131 386 165
rect 420 131 435 165
rect 371 89 435 131
rect 371 55 386 89
rect 420 55 435 89
rect 371 47 435 55
rect 465 203 521 215
rect 465 169 476 203
rect 510 169 521 203
rect 465 101 521 169
rect 465 67 476 101
rect 510 67 521 101
rect 465 47 521 67
rect 551 165 675 215
rect 551 131 562 165
rect 596 131 630 165
rect 664 131 675 165
rect 551 89 675 131
rect 551 55 562 89
rect 596 55 630 89
rect 664 55 675 89
rect 551 47 675 55
rect 705 203 761 215
rect 705 169 716 203
rect 750 169 761 203
rect 705 101 761 169
rect 705 67 716 101
rect 750 67 761 101
rect 705 47 761 67
rect 791 198 935 215
rect 791 164 890 198
rect 924 164 935 198
rect 791 161 935 164
rect 791 127 802 161
rect 836 131 935 161
rect 965 190 1018 215
rect 965 156 976 190
rect 1010 156 1018 190
rect 965 131 1018 156
rect 836 127 844 131
rect 791 93 844 127
rect 791 59 802 93
rect 836 59 844 93
rect 791 47 844 59
<< pdiff >>
rect 30 607 83 619
rect 30 573 38 607
rect 72 573 83 607
rect 30 525 83 573
rect 30 491 38 525
rect 72 491 83 525
rect 30 441 83 491
rect 30 407 38 441
rect 72 407 83 441
rect 30 367 83 407
rect 113 599 169 619
rect 113 565 124 599
rect 158 565 169 599
rect 113 506 169 565
rect 113 472 124 506
rect 158 472 169 506
rect 113 413 169 472
rect 113 379 124 413
rect 158 379 169 413
rect 113 367 169 379
rect 199 607 255 619
rect 199 573 210 607
rect 244 573 255 607
rect 199 525 255 573
rect 199 491 210 525
rect 244 491 255 525
rect 199 441 255 491
rect 199 407 210 441
rect 244 407 255 441
rect 199 367 255 407
rect 285 599 341 619
rect 285 565 296 599
rect 330 565 341 599
rect 285 506 341 565
rect 285 472 296 506
rect 330 472 341 506
rect 285 413 341 472
rect 285 379 296 413
rect 330 379 341 413
rect 285 367 341 379
rect 371 607 449 619
rect 371 573 393 607
rect 427 573 449 607
rect 371 511 449 573
rect 371 477 393 511
rect 427 477 449 511
rect 371 418 449 477
rect 371 384 393 418
rect 427 384 449 418
rect 371 367 449 384
rect 479 367 521 619
rect 551 367 629 619
rect 659 367 737 619
rect 767 599 820 619
rect 767 565 778 599
rect 812 565 820 599
rect 767 506 820 565
rect 893 585 946 609
rect 893 551 901 585
rect 935 551 946 585
rect 893 525 946 551
rect 976 584 1029 609
rect 976 550 987 584
rect 1021 550 1029 584
rect 976 525 1029 550
rect 767 472 778 506
rect 812 472 820 506
rect 767 413 820 472
rect 767 379 778 413
rect 812 379 820 413
rect 767 367 820 379
<< ndiffc >>
rect 38 133 72 167
rect 38 59 72 93
rect 124 169 158 203
rect 124 67 158 101
rect 210 55 244 89
rect 296 113 330 147
rect 386 131 420 165
rect 386 55 420 89
rect 476 169 510 203
rect 476 67 510 101
rect 562 131 596 165
rect 630 131 664 165
rect 562 55 596 89
rect 630 55 664 89
rect 716 169 750 203
rect 716 67 750 101
rect 890 164 924 198
rect 802 127 836 161
rect 976 156 1010 190
rect 802 59 836 93
<< pdiffc >>
rect 38 573 72 607
rect 38 491 72 525
rect 38 407 72 441
rect 124 565 158 599
rect 124 472 158 506
rect 124 379 158 413
rect 210 573 244 607
rect 210 491 244 525
rect 210 407 244 441
rect 296 565 330 599
rect 296 472 330 506
rect 296 379 330 413
rect 393 573 427 607
rect 393 477 427 511
rect 393 384 427 418
rect 778 565 812 599
rect 901 551 935 585
rect 987 550 1021 584
rect 778 472 812 506
rect 778 379 812 413
<< poly >>
rect 83 619 113 645
rect 169 619 199 645
rect 255 619 285 645
rect 341 619 371 645
rect 449 619 479 645
rect 521 619 551 645
rect 629 619 659 645
rect 737 619 767 645
rect 946 609 976 635
rect 946 441 976 525
rect 946 425 1012 441
rect 946 391 962 425
rect 996 391 1012 425
rect 83 321 113 367
rect 169 321 199 367
rect 255 321 285 367
rect 341 321 371 367
rect 449 335 479 367
rect 83 305 371 321
rect 83 271 117 305
rect 151 271 185 305
rect 219 271 253 305
rect 287 271 321 305
rect 355 271 371 305
rect 83 255 371 271
rect 413 319 479 335
rect 413 285 429 319
rect 463 285 479 319
rect 413 269 479 285
rect 521 335 551 367
rect 521 319 587 335
rect 521 285 537 319
rect 571 285 587 319
rect 521 269 587 285
rect 629 319 659 367
rect 737 345 767 367
rect 946 357 1012 391
rect 629 303 695 319
rect 737 315 893 345
rect 946 337 962 357
rect 629 269 645 303
rect 679 269 695 303
rect 83 215 113 255
rect 169 215 199 255
rect 255 215 285 255
rect 341 215 371 255
rect 435 215 465 269
rect 521 215 551 269
rect 629 267 695 269
rect 761 287 893 315
rect 629 237 705 267
rect 675 215 705 237
rect 761 253 843 287
rect 877 253 893 287
rect 761 237 893 253
rect 935 323 962 337
rect 996 323 1012 357
rect 935 307 1012 323
rect 761 215 791 237
rect 935 215 965 307
rect 935 105 965 131
rect 83 21 113 47
rect 169 21 199 47
rect 255 21 285 47
rect 341 21 371 47
rect 435 21 465 47
rect 521 21 551 47
rect 675 21 705 47
rect 761 21 791 47
<< polycont >>
rect 962 391 996 425
rect 117 271 151 305
rect 185 271 219 305
rect 253 271 287 305
rect 321 271 355 305
rect 429 285 463 319
rect 537 285 571 319
rect 645 269 679 303
rect 843 253 877 287
rect 962 323 996 357
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 22 607 88 649
rect 22 573 38 607
rect 72 573 88 607
rect 22 525 88 573
rect 22 491 38 525
rect 72 491 88 525
rect 22 441 88 491
rect 22 407 38 441
rect 72 407 88 441
rect 122 599 160 615
rect 122 565 124 599
rect 158 565 160 599
rect 122 506 160 565
rect 122 472 124 506
rect 158 472 160 506
rect 122 413 160 472
rect 122 379 124 413
rect 158 379 160 413
rect 194 607 260 649
rect 194 573 210 607
rect 244 573 260 607
rect 194 525 260 573
rect 194 491 210 525
rect 244 491 260 525
rect 194 441 260 491
rect 194 407 210 441
rect 244 407 260 441
rect 294 599 343 615
rect 294 565 296 599
rect 330 565 343 599
rect 294 506 343 565
rect 294 472 296 506
rect 330 472 343 506
rect 294 413 343 472
rect 122 373 160 379
rect 294 379 296 413
rect 330 379 343 413
rect 377 607 443 649
rect 377 573 393 607
rect 427 573 443 607
rect 771 599 818 615
rect 377 511 443 573
rect 377 477 393 511
rect 427 477 443 511
rect 377 418 443 477
rect 377 384 393 418
rect 427 384 443 418
rect 477 384 571 588
rect 294 373 343 379
rect 18 339 343 373
rect 18 235 67 339
rect 415 319 463 350
rect 101 271 117 305
rect 151 271 185 305
rect 219 271 253 305
rect 287 271 321 305
rect 355 271 381 305
rect 347 235 381 271
rect 415 285 429 319
rect 415 269 463 285
rect 497 319 571 384
rect 497 285 537 319
rect 497 269 571 285
rect 605 303 737 588
rect 605 269 645 303
rect 679 269 737 303
rect 771 565 778 599
rect 812 565 818 599
rect 771 506 818 565
rect 885 585 951 649
rect 885 551 901 585
rect 935 551 951 585
rect 885 543 951 551
rect 985 584 1037 615
rect 985 550 987 584
rect 1021 550 1037 584
rect 985 509 1037 550
rect 771 472 778 506
rect 812 472 818 506
rect 771 413 818 472
rect 771 379 778 413
rect 812 379 818 413
rect 771 363 818 379
rect 852 475 1037 509
rect 771 235 807 363
rect 852 303 912 475
rect 946 425 1039 441
rect 946 391 962 425
rect 996 391 1039 425
rect 946 357 1039 391
rect 946 323 962 357
rect 996 323 1039 357
rect 946 307 1039 323
rect 843 287 912 303
rect 877 271 912 287
rect 877 253 1026 271
rect 843 237 1026 253
rect 18 203 158 235
rect 18 201 124 203
rect 122 169 124 201
rect 347 203 807 235
rect 347 199 476 203
rect 22 133 38 167
rect 72 133 88 167
rect 22 93 88 133
rect 22 59 38 93
rect 72 59 88 93
rect 22 17 88 59
rect 122 165 158 169
rect 470 169 476 199
rect 510 199 716 203
rect 510 169 512 199
rect 122 147 336 165
rect 122 131 296 147
rect 122 101 160 131
rect 122 67 124 101
rect 158 67 160 101
rect 294 113 296 131
rect 330 113 336 147
rect 294 97 336 113
rect 370 131 386 165
rect 420 131 436 165
rect 122 51 160 67
rect 194 89 260 97
rect 194 55 210 89
rect 244 55 260 89
rect 194 17 260 55
rect 370 89 436 131
rect 370 55 386 89
rect 420 55 436 89
rect 370 17 436 55
rect 470 101 512 169
rect 714 169 716 199
rect 750 201 807 203
rect 750 169 752 201
rect 470 67 476 101
rect 510 67 512 101
rect 470 51 512 67
rect 546 131 562 165
rect 596 131 630 165
rect 664 131 680 165
rect 546 89 680 131
rect 546 55 562 89
rect 596 55 630 89
rect 664 55 680 89
rect 546 17 680 55
rect 714 101 752 169
rect 841 198 940 203
rect 841 167 890 198
rect 714 67 716 101
rect 750 67 752 101
rect 714 51 752 67
rect 786 164 890 167
rect 924 164 940 198
rect 786 161 940 164
rect 786 127 802 161
rect 836 127 940 161
rect 974 190 1026 237
rect 974 156 976 190
rect 1010 156 1026 190
rect 974 140 1026 156
rect 786 93 940 127
rect 786 59 802 93
rect 836 59 940 93
rect 786 17 940 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or4b_4
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2943124
string GDS_START 2932838
<< end >>
