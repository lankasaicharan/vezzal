magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2678 1852
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 1 21 1337 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 747 47 777 177
rect 945 47 975 177
rect 1039 47 1069 177
rect 1133 47 1163 177
rect 1227 47 1257 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1125 297 1161 497
rect 1219 297 1255 497
<< ndiff >>
rect 27 165 89 177
rect 27 131 35 165
rect 69 131 89 165
rect 27 97 89 131
rect 27 63 35 97
rect 69 63 89 97
rect 27 47 89 63
rect 119 97 183 177
rect 119 63 129 97
rect 163 63 183 97
rect 119 47 183 63
rect 213 165 277 177
rect 213 131 223 165
rect 257 131 277 165
rect 213 97 277 131
rect 213 63 223 97
rect 257 63 277 97
rect 213 47 277 63
rect 307 97 371 177
rect 307 63 317 97
rect 351 63 371 97
rect 307 47 371 63
rect 401 165 455 177
rect 401 131 411 165
rect 445 131 455 165
rect 401 47 455 131
rect 485 97 549 177
rect 485 63 505 97
rect 539 63 549 97
rect 485 47 549 63
rect 579 165 643 177
rect 579 131 599 165
rect 633 131 643 165
rect 579 47 643 131
rect 673 97 747 177
rect 673 63 693 97
rect 727 63 747 97
rect 673 47 747 63
rect 777 165 829 177
rect 777 131 787 165
rect 821 131 829 165
rect 777 47 829 131
rect 883 97 945 177
rect 883 63 891 97
rect 925 63 945 97
rect 883 47 945 63
rect 975 165 1039 177
rect 975 131 985 165
rect 1019 131 1039 165
rect 975 47 1039 131
rect 1069 97 1133 177
rect 1069 63 1079 97
rect 1113 63 1133 97
rect 1069 47 1133 63
rect 1163 165 1227 177
rect 1163 131 1173 165
rect 1207 131 1227 165
rect 1163 47 1227 131
rect 1257 97 1311 177
rect 1257 63 1267 97
rect 1301 63 1311 97
rect 1257 47 1311 63
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 349 551 383
rect 493 315 505 349
rect 539 315 551 349
rect 493 297 551 315
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 417 645 451
rect 587 383 599 417
rect 633 383 645 417
rect 587 297 645 383
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 349 739 383
rect 681 315 693 349
rect 727 315 739 349
rect 681 297 739 315
rect 775 485 829 497
rect 775 451 787 485
rect 821 451 829 485
rect 775 417 829 451
rect 775 383 787 417
rect 821 383 829 417
rect 775 297 829 383
rect 883 485 937 497
rect 883 451 891 485
rect 925 451 937 485
rect 883 417 937 451
rect 883 383 891 417
rect 925 383 937 417
rect 883 297 937 383
rect 973 485 1031 497
rect 973 451 985 485
rect 1019 451 1031 485
rect 973 417 1031 451
rect 973 383 985 417
rect 1019 383 1031 417
rect 973 349 1031 383
rect 973 315 985 349
rect 1019 315 1031 349
rect 973 297 1031 315
rect 1067 485 1125 497
rect 1067 451 1079 485
rect 1113 451 1125 485
rect 1067 417 1125 451
rect 1067 383 1079 417
rect 1113 383 1125 417
rect 1067 297 1125 383
rect 1161 485 1219 497
rect 1161 451 1173 485
rect 1207 451 1219 485
rect 1161 417 1219 451
rect 1161 383 1173 417
rect 1207 383 1219 417
rect 1161 349 1219 383
rect 1161 315 1173 349
rect 1207 315 1219 349
rect 1161 297 1219 315
rect 1255 485 1311 497
rect 1255 451 1267 485
rect 1301 451 1311 485
rect 1255 417 1311 451
rect 1255 383 1267 417
rect 1301 383 1311 417
rect 1255 297 1311 383
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 129 63 163 97
rect 223 131 257 165
rect 223 63 257 97
rect 317 63 351 97
rect 411 131 445 165
rect 505 63 539 97
rect 599 131 633 165
rect 693 63 727 97
rect 787 131 821 165
rect 891 63 925 97
rect 985 131 1019 165
rect 1079 63 1113 97
rect 1173 131 1207 165
rect 1267 63 1301 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 505 451 539 485
rect 505 383 539 417
rect 505 315 539 349
rect 599 451 633 485
rect 599 383 633 417
rect 693 451 727 485
rect 693 383 727 417
rect 693 315 727 349
rect 787 451 821 485
rect 787 383 821 417
rect 891 451 925 485
rect 891 383 925 417
rect 985 451 1019 485
rect 985 383 1019 417
rect 985 315 1019 349
rect 1079 451 1113 485
rect 1079 383 1113 417
rect 1173 451 1207 485
rect 1173 383 1207 417
rect 1173 315 1207 349
rect 1267 451 1301 485
rect 1267 383 1301 417
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1125 497 1161 523
rect 1219 497 1255 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1125 282 1161 297
rect 1219 282 1255 297
rect 79 259 119 282
rect 173 259 213 282
rect 267 259 307 282
rect 361 259 401 282
rect 22 249 401 259
rect 22 215 38 249
rect 72 215 129 249
rect 163 215 223 249
rect 257 215 317 249
rect 351 215 401 249
rect 22 205 401 215
rect 89 177 119 205
rect 183 177 213 205
rect 277 177 307 205
rect 371 177 401 205
rect 455 259 495 282
rect 549 259 589 282
rect 643 259 683 282
rect 737 259 777 282
rect 935 259 975 282
rect 1029 259 1069 282
rect 1123 259 1163 282
rect 1217 259 1257 282
rect 455 249 777 259
rect 455 215 505 249
rect 539 215 599 249
rect 633 215 693 249
rect 727 215 777 249
rect 455 205 777 215
rect 869 249 1257 259
rect 869 215 885 249
rect 919 215 984 249
rect 1018 215 1079 249
rect 1113 215 1173 249
rect 1207 215 1257 249
rect 869 205 1257 215
rect 455 177 485 205
rect 549 177 579 205
rect 643 177 673 205
rect 747 177 777 205
rect 945 177 975 205
rect 1039 177 1069 205
rect 1133 177 1163 205
rect 1227 177 1257 205
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 747 21 777 47
rect 945 21 975 47
rect 1039 21 1069 47
rect 1133 21 1163 47
rect 1227 21 1257 47
<< polycont >>
rect 38 215 72 249
rect 129 215 163 249
rect 223 215 257 249
rect 317 215 351 249
rect 505 215 539 249
rect 599 215 633 249
rect 693 215 727 249
rect 885 215 919 249
rect 984 215 1018 249
rect 1079 215 1113 249
rect 1173 215 1207 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 289 69 315
rect 103 485 179 493
rect 103 451 129 485
rect 163 451 179 485
rect 103 417 179 451
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 223 485 257 527
rect 223 417 257 451
rect 223 367 257 383
rect 291 485 367 493
rect 291 451 317 485
rect 351 451 367 485
rect 291 417 367 451
rect 291 383 317 417
rect 351 383 367 417
rect 103 315 129 349
rect 163 333 179 349
rect 291 349 367 383
rect 411 485 445 527
rect 411 417 445 451
rect 411 367 445 383
rect 479 485 555 493
rect 479 451 505 485
rect 539 451 555 485
rect 479 417 555 451
rect 479 383 505 417
rect 539 383 555 417
rect 291 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 479 349 555 383
rect 599 485 633 527
rect 599 417 633 451
rect 599 367 633 383
rect 667 485 743 493
rect 667 451 693 485
rect 727 451 743 485
rect 667 417 743 451
rect 667 383 693 417
rect 727 383 743 417
rect 479 333 505 349
rect 351 315 505 333
rect 539 333 555 349
rect 667 349 743 383
rect 787 485 925 527
rect 821 451 891 485
rect 787 417 925 451
rect 821 383 891 417
rect 787 367 925 383
rect 959 485 1035 493
rect 959 451 985 485
rect 1019 451 1035 485
rect 959 417 1035 451
rect 959 383 985 417
rect 1019 383 1035 417
rect 667 333 693 349
rect 539 315 693 333
rect 727 333 743 349
rect 959 349 1035 383
rect 1079 485 1113 527
rect 1079 417 1113 451
rect 1079 367 1113 383
rect 1147 485 1223 493
rect 1147 451 1173 485
rect 1207 451 1223 485
rect 1147 417 1223 451
rect 1147 383 1173 417
rect 1207 383 1223 417
rect 959 333 985 349
rect 727 315 985 333
rect 1019 333 1035 349
rect 1147 349 1223 383
rect 1267 485 1320 527
rect 1301 451 1320 485
rect 1267 417 1320 451
rect 1301 383 1320 417
rect 1267 367 1320 383
rect 1147 333 1173 349
rect 1019 315 1173 333
rect 1207 333 1223 349
rect 1207 315 1357 333
rect 103 289 1357 315
rect 22 249 370 255
rect 22 215 38 249
rect 72 215 129 249
rect 163 215 223 249
rect 257 215 317 249
rect 351 215 370 249
rect 455 249 805 255
rect 455 215 505 249
rect 539 215 599 249
rect 633 215 693 249
rect 727 215 805 249
rect 850 249 1274 255
rect 850 215 885 249
rect 919 215 984 249
rect 1018 215 1079 249
rect 1113 215 1173 249
rect 1207 215 1274 249
rect 1311 181 1357 289
rect 18 165 837 181
rect 18 131 35 165
rect 69 147 223 165
rect 69 131 85 147
rect 18 97 85 131
rect 197 131 223 147
rect 257 147 411 165
rect 257 131 273 147
rect 385 131 411 147
rect 445 147 599 165
rect 445 131 461 147
rect 573 131 599 147
rect 633 147 787 165
rect 633 131 649 147
rect 761 131 787 147
rect 821 131 837 165
rect 959 165 1357 181
rect 959 131 985 165
rect 1019 131 1173 165
rect 1207 131 1357 165
rect 18 63 35 97
rect 69 63 85 97
rect 18 51 85 63
rect 129 97 163 113
rect 129 17 163 63
rect 197 97 273 131
rect 197 63 223 97
rect 257 63 273 97
rect 197 51 273 63
rect 317 97 351 113
rect 317 17 351 63
rect 479 63 505 97
rect 539 63 693 97
rect 727 63 891 97
rect 925 63 1079 97
rect 1113 63 1267 97
rect 1301 63 1320 97
rect 479 51 1320 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 1316 153 1350 187 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 1316 221 1350 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 1316 289 1350 323 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 1226 221 1260 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 950 221 984 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 765 221 799 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 675 221 709 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 580 221 614 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 307 221 341 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 215 221 249 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 1042 221 1076 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand3_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 640704
string GDS_START 629152
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
