magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 36 232 536 248
rect 15 228 536 232
rect 15 49 1631 228
rect 0 0 1632 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 273 368 309 592
rect 387 368 423 592
rect 501 388 537 588
rect 619 388 655 588
rect 709 388 745 588
rect 799 388 835 588
rect 1017 392 1053 592
rect 1111 392 1147 592
rect 1201 392 1237 592
rect 1329 392 1365 592
rect 1423 392 1459 592
rect 1513 392 1549 592
<< nmoslvt >>
rect 112 74 142 222
rect 198 74 228 222
rect 312 74 342 222
rect 423 74 453 222
rect 621 74 651 202
rect 707 74 737 202
rect 807 74 837 202
rect 907 74 937 202
rect 1013 74 1043 202
rect 1117 74 1147 202
rect 1207 74 1237 202
rect 1307 74 1337 202
rect 1393 74 1423 202
rect 1518 74 1548 202
<< ndiff >>
rect 62 206 112 222
rect 41 194 112 206
rect 41 160 53 194
rect 87 160 112 194
rect 41 120 112 160
rect 41 86 53 120
rect 87 86 112 120
rect 41 74 112 86
rect 142 210 198 222
rect 142 176 153 210
rect 187 176 198 210
rect 142 120 198 176
rect 142 86 153 120
rect 187 86 198 120
rect 142 74 198 86
rect 228 129 312 222
rect 228 95 253 129
rect 287 95 312 129
rect 228 74 312 95
rect 342 206 423 222
rect 342 172 353 206
rect 387 172 423 206
rect 342 120 423 172
rect 342 86 353 120
rect 387 86 423 120
rect 342 74 423 86
rect 453 188 510 222
rect 453 154 464 188
rect 498 154 510 188
rect 453 120 510 154
rect 453 86 464 120
rect 498 86 510 120
rect 453 74 510 86
rect 564 188 621 202
rect 564 154 576 188
rect 610 154 621 188
rect 564 120 621 154
rect 564 86 576 120
rect 610 86 621 120
rect 564 74 621 86
rect 651 179 707 202
rect 651 145 662 179
rect 696 145 707 179
rect 651 74 707 145
rect 737 136 807 202
rect 737 102 762 136
rect 796 102 807 136
rect 737 74 807 102
rect 837 179 907 202
rect 837 145 862 179
rect 896 145 907 179
rect 837 74 907 145
rect 937 194 1013 202
rect 937 160 962 194
rect 996 160 1013 194
rect 937 120 1013 160
rect 937 86 962 120
rect 996 86 1013 120
rect 937 74 1013 86
rect 1043 122 1117 202
rect 1043 88 1062 122
rect 1096 88 1117 122
rect 1043 74 1117 88
rect 1147 192 1207 202
rect 1147 158 1162 192
rect 1196 158 1207 192
rect 1147 120 1207 158
rect 1147 86 1162 120
rect 1196 86 1207 120
rect 1147 74 1207 86
rect 1237 121 1307 202
rect 1237 87 1262 121
rect 1296 87 1307 121
rect 1237 74 1307 87
rect 1337 190 1393 202
rect 1337 156 1348 190
rect 1382 156 1393 190
rect 1337 120 1393 156
rect 1337 86 1348 120
rect 1382 86 1393 120
rect 1337 74 1393 86
rect 1423 120 1518 202
rect 1423 86 1453 120
rect 1487 86 1518 120
rect 1423 74 1518 86
rect 1548 190 1605 202
rect 1548 156 1559 190
rect 1593 156 1605 190
rect 1548 120 1605 156
rect 1548 86 1559 120
rect 1593 86 1605 120
rect 1548 74 1605 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 497 173 546
rect 119 463 129 497
rect 163 463 173 497
rect 119 414 173 463
rect 119 380 129 414
rect 163 380 173 414
rect 119 368 173 380
rect 209 580 273 592
rect 209 546 229 580
rect 263 546 273 580
rect 209 474 273 546
rect 209 440 229 474
rect 263 440 273 474
rect 209 368 273 440
rect 309 580 387 592
rect 309 546 329 580
rect 363 546 387 580
rect 309 497 387 546
rect 309 463 329 497
rect 363 463 387 497
rect 309 414 387 463
rect 309 380 329 414
rect 363 380 387 414
rect 309 368 387 380
rect 423 588 479 592
rect 423 580 501 588
rect 423 546 433 580
rect 467 546 501 580
rect 423 510 501 546
rect 423 476 433 510
rect 467 476 501 510
rect 423 440 501 476
rect 423 406 433 440
rect 467 406 501 440
rect 423 388 501 406
rect 537 574 619 588
rect 537 540 561 574
rect 595 540 619 574
rect 537 388 619 540
rect 655 436 709 588
rect 655 402 665 436
rect 699 402 709 436
rect 655 388 709 402
rect 745 575 799 588
rect 745 541 755 575
rect 789 541 799 575
rect 745 388 799 541
rect 835 575 901 588
rect 835 541 855 575
rect 889 541 901 575
rect 835 388 901 541
rect 423 368 473 388
rect 961 577 1017 592
rect 961 543 973 577
rect 1007 543 1017 577
rect 961 392 1017 543
rect 1053 438 1111 592
rect 1053 404 1063 438
rect 1097 404 1111 438
rect 1053 392 1111 404
rect 1147 577 1201 592
rect 1147 543 1157 577
rect 1191 543 1201 577
rect 1147 392 1201 543
rect 1237 444 1329 592
rect 1237 410 1266 444
rect 1300 410 1329 444
rect 1237 392 1329 410
rect 1365 580 1423 592
rect 1365 546 1377 580
rect 1411 546 1423 580
rect 1365 392 1423 546
rect 1459 440 1513 592
rect 1459 406 1469 440
rect 1503 406 1513 440
rect 1459 392 1513 406
rect 1549 580 1605 592
rect 1549 546 1559 580
rect 1593 546 1605 580
rect 1549 511 1605 546
rect 1549 477 1559 511
rect 1593 477 1605 511
rect 1549 440 1605 477
rect 1549 406 1559 440
rect 1593 406 1605 440
rect 1549 392 1605 406
<< ndiffc >>
rect 53 160 87 194
rect 53 86 87 120
rect 153 176 187 210
rect 153 86 187 120
rect 253 95 287 129
rect 353 172 387 206
rect 353 86 387 120
rect 464 154 498 188
rect 464 86 498 120
rect 576 154 610 188
rect 576 86 610 120
rect 662 145 696 179
rect 762 102 796 136
rect 862 145 896 179
rect 962 160 996 194
rect 962 86 996 120
rect 1062 88 1096 122
rect 1162 158 1196 192
rect 1162 86 1196 120
rect 1262 87 1296 121
rect 1348 156 1382 190
rect 1348 86 1382 120
rect 1453 86 1487 120
rect 1559 156 1593 190
rect 1559 86 1593 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 229 546 263 580
rect 229 440 263 474
rect 329 546 363 580
rect 329 463 363 497
rect 329 380 363 414
rect 433 546 467 580
rect 433 476 467 510
rect 433 406 467 440
rect 561 540 595 574
rect 665 402 699 436
rect 755 541 789 575
rect 855 541 889 575
rect 973 543 1007 577
rect 1063 404 1097 438
rect 1157 543 1191 577
rect 1266 410 1300 444
rect 1377 546 1411 580
rect 1469 406 1503 440
rect 1559 546 1593 580
rect 1559 477 1593 511
rect 1559 406 1593 440
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 273 592 309 618
rect 387 592 423 618
rect 501 588 537 614
rect 619 588 655 614
rect 709 588 745 614
rect 799 603 946 633
rect 799 588 835 603
rect 83 286 119 368
rect 173 286 209 368
rect 273 322 309 368
rect 387 322 423 368
rect 501 356 537 388
rect 619 373 655 388
rect 709 373 745 388
rect 501 340 571 356
rect 619 343 745 373
rect 799 362 835 388
rect 916 356 946 603
rect 1017 592 1053 618
rect 1111 592 1147 618
rect 1201 592 1237 618
rect 1329 592 1365 618
rect 1423 592 1459 618
rect 1513 592 1549 618
rect 251 306 453 322
rect 251 286 267 306
rect 83 272 267 286
rect 301 272 335 306
rect 369 272 403 306
rect 437 272 453 306
rect 501 306 521 340
rect 555 306 571 340
rect 501 290 571 306
rect 715 320 745 343
rect 899 340 965 356
rect 715 304 851 320
rect 715 290 801 304
rect 83 256 453 272
rect 112 222 142 256
rect 198 222 228 256
rect 312 222 342 256
rect 423 222 453 256
rect 541 248 571 290
rect 785 270 801 290
rect 835 270 851 304
rect 899 306 915 340
rect 949 306 965 340
rect 899 290 965 306
rect 1017 302 1053 392
rect 1111 350 1147 392
rect 1117 302 1147 350
rect 785 248 851 270
rect 1013 286 1147 302
rect 1013 252 1029 286
rect 1063 252 1097 286
rect 1131 252 1147 286
rect 541 218 737 248
rect 785 218 937 248
rect 621 202 651 218
rect 707 202 737 218
rect 807 202 837 218
rect 907 202 937 218
rect 1013 236 1147 252
rect 1013 202 1043 236
rect 1117 202 1147 236
rect 1201 360 1237 392
rect 1329 377 1365 392
rect 1423 377 1459 392
rect 1201 344 1281 360
rect 1329 347 1459 377
rect 1201 310 1231 344
rect 1265 310 1281 344
rect 1201 276 1281 310
rect 1201 242 1231 276
rect 1265 247 1281 276
rect 1393 274 1459 347
rect 1513 356 1549 392
rect 1513 340 1579 356
rect 1513 306 1529 340
rect 1563 306 1579 340
rect 1513 290 1579 306
rect 1265 242 1337 247
rect 1201 226 1337 242
rect 1207 217 1337 226
rect 1207 202 1237 217
rect 1307 202 1337 217
rect 1393 240 1409 274
rect 1443 248 1459 274
rect 1443 240 1548 248
rect 1393 218 1548 240
rect 1393 202 1423 218
rect 1518 202 1548 218
rect 112 48 142 74
rect 198 48 228 74
rect 312 48 342 74
rect 423 48 453 74
rect 621 48 651 74
rect 707 48 737 74
rect 807 48 837 74
rect 907 48 937 74
rect 1013 48 1043 74
rect 1117 48 1147 74
rect 1207 48 1237 74
rect 1307 48 1337 74
rect 1393 48 1423 74
rect 1518 48 1548 74
<< polycont >>
rect 267 272 301 306
rect 335 272 369 306
rect 403 272 437 306
rect 521 306 555 340
rect 801 270 835 304
rect 915 306 949 340
rect 1029 252 1063 286
rect 1097 252 1131 286
rect 1231 310 1265 344
rect 1231 242 1265 276
rect 1529 306 1563 340
rect 1409 240 1443 274
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 497 179 546
rect 113 463 129 497
rect 163 463 179 497
rect 113 414 179 463
rect 213 580 279 649
rect 213 546 229 580
rect 263 546 279 580
rect 213 474 279 546
rect 213 440 229 474
rect 263 440 279 474
rect 213 424 279 440
rect 313 580 379 596
rect 313 546 329 580
rect 363 546 379 580
rect 313 497 379 546
rect 313 463 329 497
rect 363 463 379 497
rect 113 380 129 414
rect 163 390 179 414
rect 313 414 379 463
rect 313 390 329 414
rect 163 380 329 390
rect 363 380 379 414
rect 417 580 483 649
rect 417 546 433 580
rect 467 546 483 580
rect 417 510 483 546
rect 531 575 805 592
rect 531 574 755 575
rect 531 540 561 574
rect 595 541 755 574
rect 789 541 805 575
rect 595 540 805 541
rect 839 575 905 649
rect 839 541 855 575
rect 889 541 905 575
rect 839 540 905 541
rect 957 577 1249 596
rect 957 543 973 577
rect 1007 543 1157 577
rect 1191 543 1249 577
rect 1361 580 1427 649
rect 1361 546 1377 580
rect 1411 546 1427 580
rect 1543 580 1609 596
rect 1543 546 1559 580
rect 1593 546 1609 580
rect 957 540 1249 543
rect 417 476 433 510
rect 467 476 483 510
rect 1215 512 1249 540
rect 1543 512 1609 546
rect 1215 511 1609 512
rect 417 440 483 476
rect 417 406 433 440
rect 467 406 483 440
rect 417 390 483 406
rect 537 472 1181 506
rect 1215 478 1559 511
rect 113 356 379 380
rect 537 356 571 472
rect 113 330 179 356
rect 25 296 179 330
rect 505 340 571 356
rect 251 306 471 322
rect 25 262 71 296
rect 251 272 267 306
rect 301 272 335 306
rect 369 272 403 306
rect 437 272 471 306
rect 505 306 521 340
rect 555 306 571 340
rect 505 290 571 306
rect 646 436 1063 438
rect 646 402 665 436
rect 699 404 1063 436
rect 1097 404 1113 438
rect 699 402 715 404
rect 646 384 715 402
rect 25 228 203 262
rect 251 256 471 272
rect 646 256 712 384
rect 1147 370 1181 472
rect 1553 477 1559 478
rect 1593 477 1609 511
rect 1231 410 1266 444
rect 1300 440 1335 444
rect 1553 440 1609 477
rect 1300 410 1469 440
rect 1231 406 1469 410
rect 1503 406 1519 440
rect 1231 394 1519 406
rect 1453 390 1519 394
rect 1553 406 1559 440
rect 1593 406 1609 440
rect 1553 390 1609 406
rect 137 222 203 228
rect 437 222 712 256
rect 785 304 851 356
rect 785 270 801 304
rect 835 270 851 304
rect 899 340 1181 370
rect 899 306 915 340
rect 949 336 1181 340
rect 1215 356 1281 360
rect 1215 344 1607 356
rect 949 306 965 336
rect 899 290 965 306
rect 1215 310 1231 344
rect 1265 340 1607 344
rect 1265 316 1529 340
rect 1265 310 1281 316
rect 785 254 851 270
rect 1013 286 1147 302
rect 1013 252 1029 286
rect 1063 252 1097 286
rect 1131 252 1147 286
rect 1013 236 1147 252
rect 1215 276 1281 310
rect 1513 306 1529 316
rect 1563 306 1607 340
rect 1513 290 1607 306
rect 1215 242 1231 276
rect 1265 242 1281 276
rect 1215 226 1281 242
rect 1369 274 1459 282
rect 1369 240 1409 274
rect 1443 240 1459 274
rect 1369 224 1459 240
rect 137 210 403 222
rect 37 160 53 194
rect 87 160 103 194
rect 37 120 103 160
rect 37 86 53 120
rect 87 86 103 120
rect 37 17 103 86
rect 137 176 153 210
rect 187 206 403 210
rect 187 188 353 206
rect 187 176 203 188
rect 137 120 203 176
rect 337 172 353 188
rect 387 172 403 206
rect 660 220 712 222
rect 137 86 153 120
rect 187 86 203 120
rect 137 70 203 86
rect 237 129 303 154
rect 237 95 253 129
rect 287 95 303 129
rect 237 17 303 95
rect 337 120 403 172
rect 337 86 353 120
rect 387 86 403 120
rect 337 70 403 86
rect 448 154 464 188
rect 498 154 514 188
rect 448 120 514 154
rect 448 86 464 120
rect 498 86 514 120
rect 448 17 514 86
rect 560 154 576 188
rect 610 154 626 188
rect 560 120 626 154
rect 560 86 576 120
rect 610 86 626 120
rect 660 186 912 220
rect 660 179 712 186
rect 660 145 662 179
rect 696 145 712 179
rect 846 179 912 186
rect 660 119 712 145
rect 746 136 812 152
rect 560 85 626 86
rect 746 102 762 136
rect 796 102 812 136
rect 846 145 862 179
rect 896 145 912 179
rect 846 119 912 145
rect 946 194 1012 202
rect 946 160 962 194
rect 996 192 1012 194
rect 996 160 1162 192
rect 946 158 1162 160
rect 1196 190 1212 192
rect 1543 190 1609 206
rect 1196 158 1348 190
rect 946 120 1012 158
rect 1146 156 1348 158
rect 1382 156 1559 190
rect 1593 156 1609 190
rect 746 85 812 102
rect 946 86 962 120
rect 996 86 1012 120
rect 946 85 1012 86
rect 560 51 1012 85
rect 1046 122 1112 124
rect 1046 88 1062 122
rect 1096 88 1112 122
rect 1046 17 1112 88
rect 1146 120 1212 156
rect 1146 86 1162 120
rect 1196 86 1212 120
rect 1146 70 1212 86
rect 1246 121 1312 122
rect 1246 87 1262 121
rect 1296 87 1312 121
rect 1246 17 1312 87
rect 1348 120 1398 156
rect 1543 120 1609 156
rect 1382 86 1398 120
rect 1348 70 1398 86
rect 1432 86 1453 120
rect 1487 86 1509 120
rect 1432 17 1509 86
rect 1543 86 1559 120
rect 1593 86 1609 120
rect 1543 70 1609 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o32a_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 900420
string GDS_START 888010
<< end >>
