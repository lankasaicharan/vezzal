magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 1 49 549 157
rect 0 0 576 49
<< scnmos >>
rect 80 47 110 131
rect 177 47 207 131
rect 263 47 293 131
rect 349 47 379 131
rect 435 47 465 131
<< scpmoshvt >>
rect 80 367 110 619
rect 176 367 206 619
rect 262 367 292 619
rect 348 367 378 619
rect 434 367 464 619
<< ndiff >>
rect 27 105 80 131
rect 27 71 35 105
rect 69 71 80 105
rect 27 47 80 71
rect 110 105 177 131
rect 110 71 121 105
rect 155 71 177 105
rect 110 47 177 71
rect 207 105 263 131
rect 207 71 218 105
rect 252 71 263 105
rect 207 47 263 71
rect 293 105 349 131
rect 293 71 304 105
rect 338 71 349 105
rect 293 47 349 71
rect 379 105 435 131
rect 379 71 390 105
rect 424 71 435 105
rect 379 47 435 71
rect 465 105 523 131
rect 465 71 476 105
rect 510 71 523 105
rect 465 47 523 71
<< pdiff >>
rect 27 596 80 619
rect 27 562 35 596
rect 69 562 80 596
rect 27 511 80 562
rect 27 477 35 511
rect 69 477 80 511
rect 27 425 80 477
rect 27 391 35 425
rect 69 391 80 425
rect 27 367 80 391
rect 110 596 176 619
rect 110 562 121 596
rect 155 562 176 596
rect 110 511 176 562
rect 110 477 121 511
rect 155 477 176 511
rect 110 425 176 477
rect 110 391 121 425
rect 155 391 176 425
rect 110 367 176 391
rect 206 596 262 619
rect 206 562 217 596
rect 251 562 262 596
rect 206 511 262 562
rect 206 477 217 511
rect 251 477 262 511
rect 206 425 262 477
rect 206 391 217 425
rect 251 391 262 425
rect 206 367 262 391
rect 292 603 348 619
rect 292 569 303 603
rect 337 569 348 603
rect 292 531 348 569
rect 292 497 303 531
rect 337 497 348 531
rect 292 463 348 497
rect 292 429 303 463
rect 337 429 348 463
rect 292 367 348 429
rect 378 596 434 619
rect 378 562 389 596
rect 423 562 434 596
rect 378 511 434 562
rect 378 477 389 511
rect 423 477 434 511
rect 378 425 434 477
rect 378 391 389 425
rect 423 391 434 425
rect 378 367 434 391
rect 464 603 524 619
rect 464 569 475 603
rect 509 569 524 603
rect 464 531 524 569
rect 464 497 475 531
rect 509 497 524 531
rect 464 463 524 497
rect 464 429 475 463
rect 509 429 524 463
rect 464 367 524 429
<< ndiffc >>
rect 35 71 69 105
rect 121 71 155 105
rect 218 71 252 105
rect 304 71 338 105
rect 390 71 424 105
rect 476 71 510 105
<< pdiffc >>
rect 35 562 69 596
rect 35 477 69 511
rect 35 391 69 425
rect 121 562 155 596
rect 121 477 155 511
rect 121 391 155 425
rect 217 562 251 596
rect 217 477 251 511
rect 217 391 251 425
rect 303 569 337 603
rect 303 497 337 531
rect 303 429 337 463
rect 389 562 423 596
rect 389 477 423 511
rect 389 391 423 425
rect 475 569 509 603
rect 475 497 509 531
rect 475 429 509 463
<< poly >>
rect 80 619 110 645
rect 176 619 206 645
rect 262 619 292 645
rect 348 619 378 645
rect 434 619 464 645
rect 80 221 110 367
rect 176 307 206 367
rect 262 307 292 367
rect 348 307 378 367
rect 434 307 464 367
rect 176 291 465 307
rect 176 257 231 291
rect 265 257 299 291
rect 333 257 367 291
rect 401 257 465 291
rect 176 241 465 257
rect 69 205 135 221
rect 69 171 85 205
rect 119 171 135 205
rect 69 155 135 171
rect 80 131 110 155
rect 177 131 207 241
rect 263 131 293 241
rect 349 131 379 241
rect 435 131 465 241
rect 80 21 110 47
rect 177 21 207 47
rect 263 21 293 47
rect 349 21 379 47
rect 435 21 465 47
<< polycont >>
rect 231 257 265 291
rect 299 257 333 291
rect 367 257 401 291
rect 85 171 119 205
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 17 596 79 612
rect 17 562 35 596
rect 69 562 79 596
rect 17 511 79 562
rect 17 477 35 511
rect 69 477 79 511
rect 17 425 79 477
rect 17 391 35 425
rect 69 391 79 425
rect 17 307 79 391
rect 113 596 175 649
rect 113 562 121 596
rect 155 562 175 596
rect 113 511 175 562
rect 113 477 121 511
rect 155 477 175 511
rect 113 425 175 477
rect 113 391 121 425
rect 155 391 175 425
rect 113 375 175 391
rect 209 596 261 612
rect 209 562 217 596
rect 251 562 261 596
rect 209 511 261 562
rect 209 477 217 511
rect 251 477 261 511
rect 209 425 261 477
rect 209 391 217 425
rect 251 391 261 425
rect 295 603 346 649
rect 295 569 303 603
rect 337 569 346 603
rect 295 531 346 569
rect 295 497 303 531
rect 337 497 346 531
rect 295 463 346 497
rect 295 429 303 463
rect 337 429 346 463
rect 295 413 346 429
rect 381 596 433 612
rect 381 562 389 596
rect 423 562 433 596
rect 381 511 433 562
rect 381 477 389 511
rect 423 477 433 511
rect 381 425 433 477
rect 209 379 261 391
rect 381 391 389 425
rect 423 391 433 425
rect 467 603 524 649
rect 467 569 475 603
rect 509 569 524 603
rect 467 531 524 569
rect 467 497 475 531
rect 509 497 524 531
rect 467 463 524 497
rect 467 429 475 463
rect 509 429 524 463
rect 467 413 524 429
rect 381 379 433 391
rect 209 345 553 379
rect 17 291 417 307
rect 17 257 231 291
rect 265 257 299 291
rect 333 257 367 291
rect 401 257 417 291
rect 17 255 417 257
rect 17 121 51 255
rect 215 241 417 255
rect 85 205 161 221
rect 451 205 553 345
rect 119 171 161 205
rect 85 155 161 171
rect 209 155 553 205
rect 17 105 77 121
rect 17 71 35 105
rect 69 71 77 105
rect 17 55 77 71
rect 111 105 166 121
rect 111 71 121 105
rect 155 71 166 105
rect 111 17 166 71
rect 209 105 261 155
rect 209 71 218 105
rect 252 71 261 105
rect 209 55 261 71
rect 295 105 346 121
rect 295 71 304 105
rect 338 71 346 105
rect 295 17 346 71
rect 381 105 433 155
rect 381 71 390 105
rect 424 71 433 105
rect 381 55 433 71
rect 467 105 523 121
rect 467 71 476 105
rect 510 71 523 105
rect 467 17 523 71
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkbuf_4
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 687296
string GDS_START 681786
<< end >>
