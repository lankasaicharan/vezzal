* NGSPICE file created from sky130_fd_sc_hd__and2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR.t0 B.t0 a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X.t1 a_59_75# VPWR.t2 VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND.t0 B.t1 a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75# A.t0 VPWR.t1 VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X.t0 a_59_75# VGND.t1 VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A.t1 a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 B.n0 B.t0 261.886
R1 B.n0 B.t1 155.846
R2 B B.n0 12.136
R3 VPWR.n0 VPWR.t0 116.027
R4 VPWR.n1 VPWR.t1 115.039
R5 VPWR.n1 VPWR.n0 45.049
R6 VPWR.n0 VPWR.t2 28.735
R7 VPWR VPWR.n1 9.919
R8 X X.t0 91.583
R9 X.n0 X.t1 50.418
R10 X X.n2 10.736
R11 X X.n1 6.344
R12 X.n2 X 5.856
R13 X.n2 X 4.417
R14 X.n1 X 3.447
R15 X.n1 X.n0 3.29
R16 X.n0 X 1.823
R17 VGND.n0 VGND.t0 72.857
R18 VGND VGND.n0 50.612
R19 VGND.n0 VGND.t1 22.324
R20 A.n0 A.t0 256.068
R21 A.n0 A.t1 150.028
R22 A A.n1 8.792
R23 A.n1 A.n0 7.5
R24 A.n1 A 7.32
C0 VPWR VGND 0.01fF
C1 A X 0.01fF
C2 VPWR X 0.22fF
C3 VPWR A 0.03fF
C4 B a_59_75# 0.30fF
C5 VGND a_59_75# 0.20fF
C6 a_145_75# a_59_75# 0.02fF
C7 B VGND 0.01fF
C8 X a_59_75# 0.21fF
C9 A a_59_75# 0.19fF
C10 VPWR VPB 0.03fF
C11 B X 0.01fF
C12 VPWR a_59_75# 0.36fF
C13 B A 0.15fF
C14 X VGND 0.18fF
C15 A VGND 0.02fF
C16 VPWR B 0.01fF
.ends

