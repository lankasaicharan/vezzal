magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3322 1852
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 2022 157
rect 29 -17 63 21
<< scnmos >>
rect 90 47 120 131
rect 186 47 216 131
rect 282 47 312 131
rect 378 47 408 131
rect 464 47 494 131
rect 560 47 590 131
rect 656 47 686 131
rect 752 47 782 131
rect 848 47 878 131
rect 944 47 974 131
rect 1040 47 1070 131
rect 1136 47 1166 131
rect 1231 47 1261 131
rect 1327 47 1357 131
rect 1423 47 1453 131
rect 1519 47 1549 131
rect 1615 47 1645 131
rect 1711 47 1741 131
rect 1807 47 1837 131
rect 1913 47 1943 131
<< scpmoshvt >>
rect 82 297 118 497
rect 178 297 214 497
rect 274 297 310 497
rect 370 297 406 497
rect 466 297 502 497
rect 562 297 598 497
rect 658 297 694 497
rect 754 297 790 497
rect 850 297 886 497
rect 946 297 982 497
rect 1042 297 1078 497
rect 1138 297 1174 497
rect 1233 297 1269 497
rect 1329 297 1365 497
rect 1425 297 1461 497
rect 1521 297 1557 497
rect 1617 297 1653 497
rect 1713 297 1749 497
rect 1809 297 1845 497
rect 1905 297 1941 497
<< ndiff >>
rect 27 93 90 131
rect 27 59 35 93
rect 69 59 90 93
rect 27 47 90 59
rect 120 106 186 131
rect 120 72 131 106
rect 165 72 186 106
rect 120 47 186 72
rect 216 106 282 131
rect 216 72 227 106
rect 261 72 282 106
rect 216 47 282 72
rect 312 106 378 131
rect 312 72 323 106
rect 357 72 378 106
rect 312 47 378 72
rect 408 106 464 131
rect 408 72 419 106
rect 453 72 464 106
rect 408 47 464 72
rect 494 106 560 131
rect 494 72 515 106
rect 549 72 560 106
rect 494 47 560 72
rect 590 97 656 131
rect 590 63 611 97
rect 645 63 656 97
rect 590 47 656 63
rect 686 106 752 131
rect 686 72 707 106
rect 741 72 752 106
rect 686 47 752 72
rect 782 97 848 131
rect 782 63 803 97
rect 837 63 848 97
rect 782 47 848 63
rect 878 106 944 131
rect 878 72 899 106
rect 933 72 944 106
rect 878 47 944 72
rect 974 97 1040 131
rect 974 63 995 97
rect 1029 63 1040 97
rect 974 47 1040 63
rect 1070 106 1136 131
rect 1070 72 1091 106
rect 1125 72 1136 106
rect 1070 47 1136 72
rect 1166 97 1231 131
rect 1166 63 1187 97
rect 1221 63 1231 97
rect 1166 47 1231 63
rect 1261 106 1327 131
rect 1261 72 1282 106
rect 1316 72 1327 106
rect 1261 47 1327 72
rect 1357 97 1423 131
rect 1357 63 1378 97
rect 1412 63 1423 97
rect 1357 47 1423 63
rect 1453 106 1519 131
rect 1453 72 1474 106
rect 1508 72 1519 106
rect 1453 47 1519 72
rect 1549 97 1615 131
rect 1549 63 1570 97
rect 1604 63 1615 97
rect 1549 47 1615 63
rect 1645 106 1711 131
rect 1645 72 1666 106
rect 1700 72 1711 106
rect 1645 47 1711 72
rect 1741 97 1807 131
rect 1741 63 1762 97
rect 1796 63 1807 97
rect 1741 47 1807 63
rect 1837 106 1913 131
rect 1837 72 1858 106
rect 1892 72 1913 106
rect 1837 47 1913 72
rect 1943 97 1996 131
rect 1943 63 1954 97
rect 1988 63 1996 97
rect 1943 47 1996 63
<< pdiff >>
rect 27 485 82 497
rect 27 451 35 485
rect 69 451 82 485
rect 27 417 82 451
rect 27 383 35 417
rect 69 383 82 417
rect 27 297 82 383
rect 118 477 178 497
rect 118 443 131 477
rect 165 443 178 477
rect 118 409 178 443
rect 118 375 131 409
rect 165 375 178 409
rect 118 297 178 375
rect 214 485 274 497
rect 214 451 227 485
rect 261 451 274 485
rect 214 417 274 451
rect 214 383 227 417
rect 261 383 274 417
rect 214 297 274 383
rect 310 469 370 497
rect 310 435 323 469
rect 357 435 370 469
rect 310 401 370 435
rect 310 367 323 401
rect 357 367 370 401
rect 310 297 370 367
rect 406 485 466 497
rect 406 451 419 485
rect 453 451 466 485
rect 406 417 466 451
rect 406 383 419 417
rect 453 383 466 417
rect 406 297 466 383
rect 502 441 562 497
rect 502 407 515 441
rect 549 407 562 441
rect 502 355 562 407
rect 502 321 515 355
rect 549 321 562 355
rect 502 297 562 321
rect 598 461 658 497
rect 598 427 611 461
rect 645 427 658 461
rect 598 297 658 427
rect 694 441 754 497
rect 694 407 707 441
rect 741 407 754 441
rect 694 355 754 407
rect 694 321 707 355
rect 741 321 754 355
rect 694 297 754 321
rect 790 461 850 497
rect 790 427 803 461
rect 837 427 850 461
rect 790 297 850 427
rect 886 441 946 497
rect 886 407 899 441
rect 933 407 946 441
rect 886 355 946 407
rect 886 321 899 355
rect 933 321 946 355
rect 886 297 946 321
rect 982 461 1042 497
rect 982 427 995 461
rect 1029 427 1042 461
rect 982 297 1042 427
rect 1078 441 1138 497
rect 1078 407 1091 441
rect 1125 407 1138 441
rect 1078 355 1138 407
rect 1078 321 1091 355
rect 1125 321 1138 355
rect 1078 297 1138 321
rect 1174 461 1233 497
rect 1174 427 1187 461
rect 1221 427 1233 461
rect 1174 297 1233 427
rect 1269 441 1329 497
rect 1269 407 1282 441
rect 1316 407 1329 441
rect 1269 355 1329 407
rect 1269 321 1282 355
rect 1316 321 1329 355
rect 1269 297 1329 321
rect 1365 461 1425 497
rect 1365 427 1378 461
rect 1412 427 1425 461
rect 1365 297 1425 427
rect 1461 441 1521 497
rect 1461 407 1474 441
rect 1508 407 1521 441
rect 1461 355 1521 407
rect 1461 321 1474 355
rect 1508 321 1521 355
rect 1461 297 1521 321
rect 1557 461 1617 497
rect 1557 427 1570 461
rect 1604 427 1617 461
rect 1557 297 1617 427
rect 1653 441 1713 497
rect 1653 407 1666 441
rect 1700 407 1713 441
rect 1653 355 1713 407
rect 1653 321 1666 355
rect 1700 321 1713 355
rect 1653 297 1713 321
rect 1749 461 1809 497
rect 1749 427 1762 461
rect 1796 427 1809 461
rect 1749 297 1809 427
rect 1845 441 1905 497
rect 1845 407 1858 441
rect 1892 407 1905 441
rect 1845 355 1905 407
rect 1845 321 1858 355
rect 1892 321 1905 355
rect 1845 297 1905 321
rect 1941 461 1996 497
rect 1941 427 1954 461
rect 1988 427 1996 461
rect 1941 297 1996 427
<< ndiffc >>
rect 35 59 69 93
rect 131 72 165 106
rect 227 72 261 106
rect 323 72 357 106
rect 419 72 453 106
rect 515 72 549 106
rect 611 63 645 97
rect 707 72 741 106
rect 803 63 837 97
rect 899 72 933 106
rect 995 63 1029 97
rect 1091 72 1125 106
rect 1187 63 1221 97
rect 1282 72 1316 106
rect 1378 63 1412 97
rect 1474 72 1508 106
rect 1570 63 1604 97
rect 1666 72 1700 106
rect 1762 63 1796 97
rect 1858 72 1892 106
rect 1954 63 1988 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 131 443 165 477
rect 131 375 165 409
rect 227 451 261 485
rect 227 383 261 417
rect 323 435 357 469
rect 323 367 357 401
rect 419 451 453 485
rect 419 383 453 417
rect 515 407 549 441
rect 515 321 549 355
rect 611 427 645 461
rect 707 407 741 441
rect 707 321 741 355
rect 803 427 837 461
rect 899 407 933 441
rect 899 321 933 355
rect 995 427 1029 461
rect 1091 407 1125 441
rect 1091 321 1125 355
rect 1187 427 1221 461
rect 1282 407 1316 441
rect 1282 321 1316 355
rect 1378 427 1412 461
rect 1474 407 1508 441
rect 1474 321 1508 355
rect 1570 427 1604 461
rect 1666 407 1700 441
rect 1666 321 1700 355
rect 1762 427 1796 461
rect 1858 407 1892 441
rect 1858 321 1892 355
rect 1954 427 1988 461
<< poly >>
rect 82 497 118 523
rect 178 497 214 523
rect 274 497 310 523
rect 370 497 406 523
rect 466 497 502 523
rect 562 497 598 523
rect 658 497 694 523
rect 754 497 790 523
rect 850 497 886 523
rect 946 497 982 523
rect 1042 497 1078 523
rect 1138 497 1174 523
rect 1233 497 1269 523
rect 1329 497 1365 523
rect 1425 497 1461 523
rect 1521 497 1557 523
rect 1617 497 1653 523
rect 1713 497 1749 523
rect 1809 497 1845 523
rect 1905 497 1941 523
rect 82 282 118 297
rect 178 282 214 297
rect 274 282 310 297
rect 370 282 406 297
rect 466 282 502 297
rect 562 282 598 297
rect 658 282 694 297
rect 754 282 790 297
rect 850 282 886 297
rect 946 282 982 297
rect 1042 282 1078 297
rect 1138 282 1174 297
rect 1233 282 1269 297
rect 1329 282 1365 297
rect 1425 282 1461 297
rect 1521 282 1557 297
rect 1617 282 1653 297
rect 1713 282 1749 297
rect 1809 282 1845 297
rect 1905 282 1941 297
rect 21 249 408 282
rect 21 215 37 249
rect 71 215 408 249
rect 21 180 408 215
rect 90 131 120 180
rect 186 131 216 180
rect 282 131 312 180
rect 378 131 408 180
rect 464 265 504 282
rect 560 265 600 282
rect 656 265 696 282
rect 752 265 792 282
rect 848 265 888 282
rect 944 265 984 282
rect 1040 265 1080 282
rect 1136 265 1176 282
rect 1231 265 1271 282
rect 1327 265 1367 282
rect 1423 265 1463 282
rect 1519 265 1559 282
rect 1615 265 1655 282
rect 1711 265 1751 282
rect 1807 265 1847 282
rect 1903 265 1943 282
rect 464 249 1943 265
rect 464 215 514 249
rect 548 215 582 249
rect 616 215 660 249
rect 694 215 738 249
rect 772 215 816 249
rect 850 215 894 249
rect 928 215 962 249
rect 996 215 1040 249
rect 1074 215 1118 249
rect 1152 215 1196 249
rect 1230 215 1274 249
rect 1308 215 1342 249
rect 1376 215 1420 249
rect 1454 215 1498 249
rect 1532 215 1576 249
rect 1610 215 1644 249
rect 1678 215 1943 249
rect 464 190 1943 215
rect 464 131 494 190
rect 560 131 590 190
rect 656 131 686 190
rect 752 131 782 190
rect 848 131 878 190
rect 944 131 974 190
rect 1040 131 1070 190
rect 1136 131 1166 190
rect 1231 131 1261 190
rect 1327 131 1357 190
rect 1423 131 1453 190
rect 1519 131 1549 190
rect 1615 131 1645 190
rect 1711 131 1741 190
rect 1807 131 1837 190
rect 1913 131 1943 190
rect 90 21 120 47
rect 186 21 216 47
rect 282 21 312 47
rect 378 21 408 47
rect 464 21 494 47
rect 560 21 590 47
rect 656 21 686 47
rect 752 21 782 47
rect 848 21 878 47
rect 944 21 974 47
rect 1040 21 1070 47
rect 1136 21 1166 47
rect 1231 21 1261 47
rect 1327 21 1357 47
rect 1423 21 1453 47
rect 1519 21 1549 47
rect 1615 21 1645 47
rect 1711 21 1741 47
rect 1807 21 1837 47
rect 1913 21 1943 47
<< polycont >>
rect 37 215 71 249
rect 514 215 548 249
rect 582 215 616 249
rect 660 215 694 249
rect 738 215 772 249
rect 816 215 850 249
rect 894 215 928 249
rect 962 215 996 249
rect 1040 215 1074 249
rect 1118 215 1152 249
rect 1196 215 1230 249
rect 1274 215 1308 249
rect 1342 215 1376 249
rect 1420 215 1454 249
rect 1498 215 1532 249
rect 1576 215 1610 249
rect 1644 215 1678 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 19 485 78 527
rect 19 451 35 485
rect 69 451 78 485
rect 19 417 78 451
rect 19 383 35 417
rect 69 383 78 417
rect 19 365 78 383
rect 124 477 173 493
rect 124 443 131 477
rect 165 443 173 477
rect 124 409 173 443
rect 124 375 131 409
rect 165 375 173 409
rect 124 265 173 375
rect 218 485 270 527
rect 410 526 1805 527
rect 218 451 227 485
rect 261 451 270 485
rect 218 417 270 451
rect 218 383 227 417
rect 261 383 270 417
rect 218 365 270 383
rect 316 469 366 492
rect 316 435 323 469
rect 357 435 366 469
rect 316 401 366 435
rect 316 367 323 401
rect 357 367 366 401
rect 410 485 462 526
rect 410 451 419 485
rect 453 451 462 485
rect 410 417 462 451
rect 410 383 419 417
rect 453 383 462 417
rect 410 367 462 383
rect 506 441 558 492
rect 506 407 515 441
rect 549 407 558 441
rect 316 265 366 367
rect 506 355 558 407
rect 602 461 654 526
rect 602 427 611 461
rect 645 427 654 461
rect 602 381 654 427
rect 698 441 750 492
rect 698 407 707 441
rect 741 407 750 441
rect 506 321 515 355
rect 549 347 558 355
rect 698 355 750 407
rect 794 461 846 526
rect 794 427 803 461
rect 837 427 846 461
rect 794 381 846 427
rect 890 441 942 492
rect 890 407 899 441
rect 933 407 942 441
rect 698 347 707 355
rect 549 321 707 347
rect 741 347 750 355
rect 890 355 942 407
rect 986 461 1038 526
rect 986 427 995 461
rect 1029 427 1038 461
rect 986 381 1038 427
rect 1082 441 1134 492
rect 1082 407 1091 441
rect 1125 407 1134 441
rect 890 347 899 355
rect 741 321 899 347
rect 933 347 942 355
rect 1082 355 1134 407
rect 1178 461 1227 526
rect 1178 427 1187 461
rect 1221 427 1227 461
rect 1178 381 1227 427
rect 1271 441 1323 492
rect 1271 407 1282 441
rect 1316 407 1323 441
rect 1082 347 1091 355
rect 933 321 1091 347
rect 1125 347 1134 355
rect 1271 355 1323 407
rect 1370 461 1419 526
rect 1370 427 1378 461
rect 1412 427 1419 461
rect 1370 381 1419 427
rect 1463 441 1515 492
rect 1463 407 1474 441
rect 1508 407 1515 441
rect 1271 347 1282 355
rect 1125 321 1282 347
rect 1316 347 1323 355
rect 1463 355 1515 407
rect 1562 461 1611 526
rect 1562 427 1570 461
rect 1604 427 1611 461
rect 1562 381 1611 427
rect 1655 441 1707 492
rect 1655 407 1666 441
rect 1700 407 1707 441
rect 1463 347 1474 355
rect 1316 321 1474 347
rect 1508 347 1515 355
rect 1655 355 1707 407
rect 1754 461 1805 526
rect 1754 427 1762 461
rect 1796 427 1805 461
rect 1754 381 1805 427
rect 1849 441 1907 492
rect 1849 407 1858 441
rect 1892 407 1907 441
rect 1655 347 1666 355
rect 1508 321 1666 347
rect 1700 344 1707 355
rect 1849 355 1907 407
rect 1951 461 2005 527
rect 1951 427 1954 461
rect 1988 427 2005 461
rect 1951 378 2005 427
rect 1849 344 1858 355
rect 1700 321 1858 344
rect 1892 344 1907 355
rect 1892 321 2005 344
rect 506 299 2005 321
rect 17 249 80 265
rect 17 215 37 249
rect 71 215 80 249
rect 17 153 80 215
rect 124 249 1708 265
rect 124 215 514 249
rect 548 215 582 249
rect 616 215 660 249
rect 694 215 738 249
rect 772 215 816 249
rect 850 215 894 249
rect 928 215 962 249
rect 996 215 1040 249
rect 1074 215 1118 249
rect 1152 215 1196 249
rect 1230 215 1274 249
rect 1308 215 1342 249
rect 1376 215 1420 249
rect 1454 215 1498 249
rect 1532 215 1576 249
rect 1610 215 1644 249
rect 1678 215 1708 249
rect 17 93 78 119
rect 17 59 35 93
rect 69 59 78 93
rect 17 17 78 59
rect 124 106 174 215
rect 124 72 131 106
rect 165 72 174 106
rect 124 53 174 72
rect 218 106 270 122
rect 218 72 227 106
rect 261 72 270 106
rect 218 17 270 72
rect 316 106 366 215
rect 1752 181 2005 299
rect 506 147 2005 181
rect 316 72 323 106
rect 357 72 366 106
rect 316 53 366 72
rect 410 106 462 129
rect 410 72 419 106
rect 453 72 462 106
rect 410 17 462 72
rect 506 106 558 147
rect 506 72 515 106
rect 549 72 558 106
rect 506 56 558 72
rect 602 97 654 113
rect 602 63 611 97
rect 645 63 654 97
rect 602 17 654 63
rect 698 106 750 147
rect 698 72 707 106
rect 741 72 750 106
rect 698 56 750 72
rect 794 97 846 113
rect 794 63 803 97
rect 837 63 846 97
rect 794 17 846 63
rect 890 106 942 147
rect 890 72 899 106
rect 933 72 942 106
rect 890 56 942 72
rect 986 97 1035 113
rect 986 63 995 97
rect 1029 63 1035 97
rect 986 17 1035 63
rect 1069 106 1134 147
rect 1069 72 1091 106
rect 1125 72 1134 106
rect 1069 56 1134 72
rect 1178 97 1227 113
rect 1178 63 1187 97
rect 1221 63 1227 97
rect 1178 17 1227 63
rect 1271 106 1323 147
rect 1271 72 1282 106
rect 1316 72 1323 106
rect 1271 56 1323 72
rect 1369 97 1419 113
rect 1369 63 1378 97
rect 1412 63 1419 97
rect 1369 17 1419 63
rect 1463 106 1515 147
rect 1463 72 1474 106
rect 1508 72 1515 106
rect 1463 56 1515 72
rect 1561 97 1611 113
rect 1561 63 1570 97
rect 1604 63 1611 97
rect 1561 17 1611 63
rect 1655 106 1707 147
rect 1655 72 1666 106
rect 1700 72 1707 106
rect 1655 56 1707 72
rect 1753 97 1805 113
rect 1753 63 1762 97
rect 1796 63 1805 97
rect 1753 17 1805 63
rect 1849 106 1901 147
rect 1849 72 1858 106
rect 1892 72 1901 106
rect 1849 56 1901 72
rect 1945 97 2005 113
rect 1945 63 1954 97
rect 1988 63 2005 97
rect 1945 17 2005 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 1773 289 1807 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 1875 289 1909 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 1875 221 1909 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 1773 221 1807 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 1773 153 1807 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 1875 153 1909 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkbuf_16
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 890192
string GDS_START 876736
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
