magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 492 228 767 248
rect 1 49 767 228
rect 0 0 768 49
<< scnmos >>
rect 113 74 143 202
rect 199 74 229 202
rect 347 74 377 202
rect 433 74 463 202
rect 568 74 598 222
rect 654 74 684 222
<< scpmoshvt >>
rect 144 392 174 592
rect 228 392 258 592
rect 312 392 342 592
rect 428 392 458 592
rect 545 368 575 592
rect 635 368 665 592
<< ndiff >>
rect 518 202 568 222
rect 27 115 113 202
rect 27 81 45 115
rect 79 81 113 115
rect 27 74 113 81
rect 143 188 199 202
rect 143 154 154 188
rect 188 154 199 188
rect 143 120 199 154
rect 143 86 154 120
rect 188 86 199 120
rect 143 74 199 86
rect 229 115 347 202
rect 229 81 271 115
rect 305 81 347 115
rect 229 74 347 81
rect 377 190 433 202
rect 377 156 388 190
rect 422 156 433 190
rect 377 120 433 156
rect 377 86 388 120
rect 422 86 433 120
rect 377 74 433 86
rect 463 146 568 202
rect 463 112 500 146
rect 534 112 568 146
rect 463 74 568 112
rect 598 210 654 222
rect 598 176 609 210
rect 643 176 654 210
rect 598 120 654 176
rect 598 86 609 120
rect 643 86 654 120
rect 598 74 654 86
rect 684 139 741 222
rect 684 105 695 139
rect 729 105 741 139
rect 684 74 741 105
rect 27 69 98 74
rect 244 69 332 74
<< pdiff >>
rect 85 580 144 592
rect 85 546 97 580
rect 131 546 144 580
rect 85 509 144 546
rect 85 475 97 509
rect 131 475 144 509
rect 85 438 144 475
rect 85 404 97 438
rect 131 404 144 438
rect 85 392 144 404
rect 174 392 228 592
rect 258 392 312 592
rect 342 392 428 592
rect 458 580 545 592
rect 458 546 488 580
rect 522 546 545 580
rect 458 510 545 546
rect 458 476 488 510
rect 522 476 545 510
rect 458 440 545 476
rect 458 406 488 440
rect 522 406 545 440
rect 458 392 545 406
rect 476 368 545 392
rect 575 580 635 592
rect 575 546 588 580
rect 622 546 635 580
rect 575 497 635 546
rect 575 463 588 497
rect 622 463 635 497
rect 575 414 635 463
rect 575 380 588 414
rect 622 380 635 414
rect 575 368 635 380
rect 665 580 734 592
rect 665 546 688 580
rect 722 546 734 580
rect 665 462 734 546
rect 665 428 688 462
rect 722 428 734 462
rect 665 368 734 428
<< ndiffc >>
rect 45 81 79 115
rect 154 154 188 188
rect 154 86 188 120
rect 271 81 305 115
rect 388 156 422 190
rect 388 86 422 120
rect 500 112 534 146
rect 609 176 643 210
rect 609 86 643 120
rect 695 105 729 139
<< pdiffc >>
rect 97 546 131 580
rect 97 475 131 509
rect 97 404 131 438
rect 488 546 522 580
rect 488 476 522 510
rect 488 406 522 440
rect 588 546 622 580
rect 588 463 622 497
rect 588 380 622 414
rect 688 546 722 580
rect 688 428 722 462
<< poly >>
rect 144 592 174 618
rect 228 592 258 618
rect 312 592 342 618
rect 428 592 458 618
rect 545 592 575 618
rect 635 592 665 618
rect 144 377 174 392
rect 228 377 258 392
rect 312 377 342 392
rect 428 377 458 392
rect 85 347 177 377
rect 85 338 151 347
rect 85 304 101 338
rect 135 304 151 338
rect 85 288 151 304
rect 225 299 261 377
rect 309 336 345 377
rect 425 336 461 377
rect 545 353 575 368
rect 635 353 665 368
rect 309 320 377 336
rect 113 202 143 288
rect 199 283 267 299
rect 199 249 217 283
rect 251 249 267 283
rect 309 286 325 320
rect 359 286 377 320
rect 309 270 377 286
rect 425 320 491 336
rect 425 286 441 320
rect 475 286 491 320
rect 425 270 491 286
rect 542 326 578 353
rect 632 326 668 353
rect 542 310 668 326
rect 542 276 558 310
rect 592 290 668 310
rect 592 276 684 290
rect 199 233 267 249
rect 199 202 229 233
rect 347 202 377 270
rect 433 202 463 270
rect 542 260 684 276
rect 568 222 598 260
rect 654 222 684 260
rect 113 48 143 74
rect 199 48 229 74
rect 347 48 377 74
rect 433 48 463 74
rect 568 48 598 74
rect 654 48 684 74
<< polycont >>
rect 101 304 135 338
rect 217 249 251 283
rect 325 286 359 320
rect 441 286 475 320
rect 558 276 592 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 81 580 147 596
rect 81 546 97 580
rect 131 546 147 580
rect 472 580 538 649
rect 81 509 147 546
rect 81 475 97 509
rect 131 475 147 509
rect 81 438 147 475
rect 81 422 97 438
rect 17 404 97 422
rect 131 404 147 438
rect 17 388 147 404
rect 17 199 51 388
rect 85 338 167 354
rect 85 304 101 338
rect 135 304 167 338
rect 85 236 167 304
rect 201 283 267 578
rect 201 249 217 283
rect 251 249 267 283
rect 309 320 375 578
rect 472 546 488 580
rect 522 546 538 580
rect 472 510 538 546
rect 472 476 488 510
rect 522 476 538 510
rect 472 440 538 476
rect 472 406 488 440
rect 522 406 538 440
rect 472 390 538 406
rect 572 580 638 596
rect 572 546 588 580
rect 622 546 638 580
rect 572 497 638 546
rect 572 463 588 497
rect 622 463 638 497
rect 572 414 638 463
rect 672 580 738 649
rect 672 546 688 580
rect 722 546 738 580
rect 672 462 738 546
rect 672 428 688 462
rect 722 428 738 462
rect 572 380 588 414
rect 622 394 638 414
rect 622 380 743 394
rect 572 360 743 380
rect 309 286 325 320
rect 359 286 375 320
rect 309 270 375 286
rect 409 320 491 356
rect 409 286 441 320
rect 475 286 491 320
rect 409 270 491 286
rect 525 310 608 326
rect 525 276 558 310
rect 592 276 608 310
rect 201 233 267 249
rect 525 260 608 276
rect 525 236 559 260
rect 372 202 559 236
rect 697 226 743 360
rect 593 210 743 226
rect 372 199 438 202
rect 17 190 438 199
rect 17 188 388 190
rect 17 165 154 188
rect 138 154 154 165
rect 188 165 388 188
rect 188 154 204 165
rect 23 115 102 131
rect 23 81 45 115
rect 79 81 102 115
rect 23 17 102 81
rect 138 120 204 154
rect 372 156 388 165
rect 422 156 438 190
rect 593 176 609 210
rect 643 192 743 210
rect 138 86 154 120
rect 188 86 204 120
rect 138 70 204 86
rect 240 115 336 131
rect 240 81 271 115
rect 305 81 336 115
rect 240 17 336 81
rect 372 120 438 156
rect 372 86 388 120
rect 422 86 438 120
rect 372 70 438 86
rect 472 146 559 165
rect 472 112 500 146
rect 534 112 559 146
rect 472 17 559 112
rect 593 120 643 176
rect 593 86 609 120
rect 593 70 643 86
rect 679 139 745 155
rect 679 105 695 139
rect 729 105 745 139
rect 679 17 745 105
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or4_2
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 218144
string GDS_START 210716
<< end >>
