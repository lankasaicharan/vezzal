magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 50 49 548 157
rect 0 0 576 49
<< scnmos >>
rect 129 47 159 131
rect 207 47 237 131
rect 321 47 351 131
rect 435 47 465 131
<< scpmoshvt >>
rect 157 462 187 590
rect 243 462 273 590
rect 329 462 359 590
rect 415 462 445 590
<< ndiff >>
rect 76 106 129 131
rect 76 72 84 106
rect 118 72 129 106
rect 76 47 129 72
rect 159 47 207 131
rect 237 47 321 131
rect 351 47 435 131
rect 465 106 522 131
rect 465 72 480 106
rect 514 72 522 106
rect 465 47 522 72
<< pdiff >>
rect 104 578 157 590
rect 104 544 112 578
rect 146 544 157 578
rect 104 508 157 544
rect 104 474 112 508
rect 146 474 157 508
rect 104 462 157 474
rect 187 576 243 590
rect 187 542 198 576
rect 232 542 243 576
rect 187 508 243 542
rect 187 474 198 508
rect 232 474 243 508
rect 187 462 243 474
rect 273 578 329 590
rect 273 544 284 578
rect 318 544 329 578
rect 273 510 329 544
rect 273 476 284 510
rect 318 476 329 510
rect 273 462 329 476
rect 359 576 415 590
rect 359 542 370 576
rect 404 542 415 576
rect 359 508 415 542
rect 359 474 370 508
rect 404 474 415 508
rect 359 462 415 474
rect 445 578 498 590
rect 445 544 456 578
rect 490 544 498 578
rect 445 510 498 544
rect 445 476 456 510
rect 490 476 498 510
rect 445 462 498 476
<< ndiffc >>
rect 84 72 118 106
rect 480 72 514 106
<< pdiffc >>
rect 112 544 146 578
rect 112 474 146 508
rect 198 542 232 576
rect 198 474 232 508
rect 284 544 318 578
rect 284 476 318 510
rect 370 542 404 576
rect 370 474 404 508
rect 456 544 490 578
rect 456 476 490 510
<< poly >>
rect 157 590 187 616
rect 243 590 273 616
rect 329 590 359 616
rect 415 590 445 616
rect 157 365 187 462
rect 93 349 187 365
rect 93 315 109 349
rect 143 335 187 349
rect 143 315 159 335
rect 93 281 159 315
rect 243 287 273 462
rect 329 287 359 462
rect 415 365 445 462
rect 415 335 465 365
rect 435 302 465 335
rect 93 247 109 281
rect 143 247 159 281
rect 93 231 159 247
rect 129 131 159 231
rect 207 271 273 287
rect 207 237 223 271
rect 257 237 273 271
rect 207 203 273 237
rect 207 169 223 203
rect 257 169 273 203
rect 207 153 273 169
rect 321 271 387 287
rect 321 237 337 271
rect 371 237 387 271
rect 321 203 387 237
rect 321 169 337 203
rect 371 169 387 203
rect 321 153 387 169
rect 435 286 501 302
rect 435 252 451 286
rect 485 252 501 286
rect 435 218 501 252
rect 435 184 451 218
rect 485 184 501 218
rect 435 168 501 184
rect 207 131 237 153
rect 321 131 351 153
rect 435 131 465 168
rect 129 21 159 47
rect 207 21 237 47
rect 321 21 351 47
rect 435 21 465 47
<< polycont >>
rect 109 315 143 349
rect 109 247 143 281
rect 223 237 257 271
rect 223 169 257 203
rect 337 237 371 271
rect 337 169 371 203
rect 451 252 485 286
rect 451 184 485 218
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 96 578 155 649
rect 96 544 112 578
rect 146 544 155 578
rect 96 508 155 544
rect 96 474 112 508
rect 146 474 155 508
rect 96 458 155 474
rect 189 576 241 592
rect 189 542 198 576
rect 232 542 241 576
rect 189 508 241 542
rect 189 474 198 508
rect 232 474 241 508
rect 189 426 241 474
rect 275 578 327 649
rect 275 544 284 578
rect 318 544 327 578
rect 275 510 327 544
rect 275 476 284 510
rect 318 476 327 510
rect 275 460 327 476
rect 361 576 413 592
rect 361 542 370 576
rect 404 542 413 576
rect 361 508 413 542
rect 361 474 370 508
rect 404 474 413 508
rect 361 426 413 474
rect 447 578 506 649
rect 447 544 456 578
rect 490 544 506 578
rect 447 510 506 544
rect 447 476 456 510
rect 490 476 506 510
rect 447 460 506 476
rect 17 349 143 424
rect 189 384 559 426
rect 17 315 109 349
rect 17 281 143 315
rect 17 247 109 281
rect 17 168 143 247
rect 207 271 270 350
rect 207 237 223 271
rect 257 237 270 271
rect 207 203 270 237
rect 207 169 223 203
rect 257 169 270 203
rect 68 106 134 122
rect 68 72 84 106
rect 118 72 134 106
rect 207 75 270 169
rect 304 271 371 350
rect 304 237 337 271
rect 304 203 371 237
rect 304 169 337 203
rect 304 75 371 169
rect 405 286 485 350
rect 405 252 451 286
rect 405 218 485 252
rect 405 184 451 218
rect 405 156 485 184
rect 519 122 559 384
rect 456 106 559 122
rect 68 17 134 72
rect 456 72 480 106
rect 514 72 559 106
rect 456 56 559 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4_0
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4607888
string GDS_START 4601030
<< end >>
