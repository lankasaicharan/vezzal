magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 51 49 792 243
rect 0 0 864 49
<< scnmos >>
rect 130 49 160 217
rect 232 49 262 217
rect 318 49 348 217
rect 425 49 455 217
rect 511 49 541 217
rect 597 49 627 217
rect 683 49 713 217
<< scpmoshvt >>
rect 130 367 160 619
rect 202 367 232 619
rect 310 367 340 619
rect 425 367 455 619
rect 511 367 541 619
rect 597 367 627 619
rect 683 367 713 619
<< ndiff >>
rect 77 205 130 217
rect 77 171 85 205
rect 119 171 130 205
rect 77 101 130 171
rect 77 67 85 101
rect 119 67 130 101
rect 77 49 130 67
rect 160 165 232 217
rect 160 131 178 165
rect 212 131 232 165
rect 160 91 232 131
rect 160 57 178 91
rect 212 57 232 91
rect 160 49 232 57
rect 262 205 318 217
rect 262 171 273 205
rect 307 171 318 205
rect 262 101 318 171
rect 262 67 273 101
rect 307 67 318 101
rect 262 49 318 67
rect 348 165 425 217
rect 348 131 369 165
rect 403 131 425 165
rect 348 91 425 131
rect 348 57 369 91
rect 403 57 425 91
rect 348 49 425 57
rect 455 205 511 217
rect 455 171 466 205
rect 500 171 511 205
rect 455 101 511 171
rect 455 67 466 101
rect 500 67 511 101
rect 455 49 511 67
rect 541 181 597 217
rect 541 147 552 181
rect 586 147 597 181
rect 541 95 597 147
rect 541 61 552 95
rect 586 61 597 95
rect 541 49 597 61
rect 627 205 683 217
rect 627 171 638 205
rect 672 171 683 205
rect 627 101 683 171
rect 627 67 638 101
rect 672 67 683 101
rect 627 49 683 67
rect 713 165 766 217
rect 713 131 724 165
rect 758 131 766 165
rect 713 95 766 131
rect 713 61 724 95
rect 758 61 766 95
rect 713 49 766 61
<< pdiff >>
rect 77 607 130 619
rect 77 573 85 607
rect 119 573 130 607
rect 77 516 130 573
rect 77 482 85 516
rect 119 482 130 516
rect 77 426 130 482
rect 77 392 85 426
rect 119 392 130 426
rect 77 367 130 392
rect 160 367 202 619
rect 232 367 310 619
rect 340 607 425 619
rect 340 573 365 607
rect 399 573 425 607
rect 340 499 425 573
rect 340 465 365 499
rect 399 465 425 499
rect 340 367 425 465
rect 455 599 511 619
rect 455 565 466 599
rect 500 565 511 599
rect 455 507 511 565
rect 455 473 466 507
rect 500 473 511 507
rect 455 413 511 473
rect 455 379 466 413
rect 500 379 511 413
rect 455 367 511 379
rect 541 611 597 619
rect 541 577 552 611
rect 586 577 597 611
rect 541 536 597 577
rect 541 502 552 536
rect 586 502 597 536
rect 541 457 597 502
rect 541 423 552 457
rect 586 423 597 457
rect 541 367 597 423
rect 627 599 683 619
rect 627 565 638 599
rect 672 565 683 599
rect 627 507 683 565
rect 627 473 638 507
rect 672 473 683 507
rect 627 413 683 473
rect 627 379 638 413
rect 672 379 683 413
rect 627 367 683 379
rect 713 607 766 619
rect 713 573 724 607
rect 758 573 766 607
rect 713 536 766 573
rect 713 502 724 536
rect 758 502 766 536
rect 713 457 766 502
rect 713 423 724 457
rect 758 423 766 457
rect 713 367 766 423
<< ndiffc >>
rect 85 171 119 205
rect 85 67 119 101
rect 178 131 212 165
rect 178 57 212 91
rect 273 171 307 205
rect 273 67 307 101
rect 369 131 403 165
rect 369 57 403 91
rect 466 171 500 205
rect 466 67 500 101
rect 552 147 586 181
rect 552 61 586 95
rect 638 171 672 205
rect 638 67 672 101
rect 724 131 758 165
rect 724 61 758 95
<< pdiffc >>
rect 85 573 119 607
rect 85 482 119 516
rect 85 392 119 426
rect 365 573 399 607
rect 365 465 399 499
rect 466 565 500 599
rect 466 473 500 507
rect 466 379 500 413
rect 552 577 586 611
rect 552 502 586 536
rect 552 423 586 457
rect 638 565 672 599
rect 638 473 672 507
rect 638 379 672 413
rect 724 573 758 607
rect 724 502 758 536
rect 724 423 758 457
<< poly >>
rect 130 619 160 645
rect 202 619 232 645
rect 310 619 340 645
rect 425 619 455 645
rect 511 619 541 645
rect 597 619 627 645
rect 683 619 713 645
rect 130 325 160 367
rect 94 309 160 325
rect 94 275 110 309
rect 144 275 160 309
rect 94 259 160 275
rect 202 335 232 367
rect 310 335 340 367
rect 425 335 455 367
rect 511 335 541 367
rect 597 335 627 367
rect 683 335 713 367
rect 202 319 268 335
rect 202 285 218 319
rect 252 285 268 319
rect 202 269 268 285
rect 310 319 376 335
rect 310 285 326 319
rect 360 285 376 319
rect 310 269 376 285
rect 425 319 763 335
rect 425 285 441 319
rect 475 285 509 319
rect 543 285 577 319
rect 611 285 645 319
rect 679 285 713 319
rect 747 285 763 319
rect 425 269 763 285
rect 130 217 160 259
rect 232 217 262 269
rect 318 217 348 269
rect 425 217 455 269
rect 511 217 541 269
rect 597 217 627 269
rect 683 217 713 269
rect 130 23 160 49
rect 232 23 262 49
rect 318 23 348 49
rect 425 23 455 49
rect 511 23 541 49
rect 597 23 627 49
rect 683 23 713 49
<< polycont >>
rect 110 275 144 309
rect 218 285 252 319
rect 326 285 360 319
rect 441 285 475 319
rect 509 285 543 319
rect 577 285 611 319
rect 645 285 679 319
rect 713 285 747 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 69 607 135 615
rect 69 573 85 607
rect 119 573 135 607
rect 69 516 135 573
rect 69 482 85 516
rect 119 482 135 516
rect 69 426 135 482
rect 349 607 420 649
rect 349 573 365 607
rect 399 573 420 607
rect 349 499 420 573
rect 349 465 365 499
rect 399 465 420 499
rect 349 454 420 465
rect 464 599 502 615
rect 464 565 466 599
rect 500 565 502 599
rect 464 507 502 565
rect 464 473 466 507
rect 500 473 502 507
rect 69 392 85 426
rect 119 420 135 426
rect 119 392 430 420
rect 69 384 430 392
rect 17 309 171 350
rect 17 275 110 309
rect 144 275 171 309
rect 205 319 271 350
rect 205 285 218 319
rect 252 285 271 319
rect 205 269 271 285
rect 305 319 362 350
rect 305 285 326 319
rect 360 285 362 319
rect 305 269 362 285
rect 396 319 430 384
rect 464 413 502 473
rect 536 611 602 649
rect 536 577 552 611
rect 586 577 602 611
rect 536 536 602 577
rect 536 502 552 536
rect 586 502 602 536
rect 536 457 602 502
rect 536 423 552 457
rect 586 423 602 457
rect 636 599 674 615
rect 636 565 638 599
rect 672 565 674 599
rect 636 507 674 565
rect 636 473 638 507
rect 672 473 674 507
rect 464 379 466 413
rect 500 389 502 413
rect 636 413 674 473
rect 708 607 774 649
rect 708 573 724 607
rect 758 573 774 607
rect 708 536 774 573
rect 708 502 724 536
rect 758 502 774 536
rect 708 457 774 502
rect 708 423 724 457
rect 758 423 774 457
rect 636 389 638 413
rect 500 379 638 389
rect 672 389 674 413
rect 672 379 833 389
rect 464 355 833 379
rect 396 285 441 319
rect 475 285 509 319
rect 543 285 577 319
rect 611 285 645 319
rect 679 285 713 319
rect 747 285 763 319
rect 396 233 430 285
rect 797 249 833 355
rect 69 205 430 233
rect 69 171 85 205
rect 119 199 273 205
rect 119 171 128 199
rect 69 101 128 171
rect 262 171 273 199
rect 307 199 430 205
rect 464 215 833 249
rect 464 205 502 215
rect 307 171 319 199
rect 69 67 85 101
rect 119 67 128 101
rect 69 51 128 67
rect 162 131 178 165
rect 212 131 228 165
rect 162 91 228 131
rect 162 57 178 91
rect 212 57 228 91
rect 162 17 228 57
rect 262 101 319 171
rect 464 171 466 205
rect 500 171 502 205
rect 636 205 681 215
rect 262 67 273 101
rect 307 67 319 101
rect 262 51 319 67
rect 353 131 369 165
rect 403 131 426 165
rect 353 91 426 131
rect 353 57 369 91
rect 403 57 426 91
rect 353 17 426 57
rect 464 101 502 171
rect 464 67 466 101
rect 500 67 502 101
rect 464 51 502 67
rect 536 147 552 181
rect 586 147 602 181
rect 536 95 602 147
rect 536 61 552 95
rect 586 61 602 95
rect 536 17 602 61
rect 636 171 638 205
rect 672 171 681 205
rect 636 101 681 171
rect 636 67 638 101
rect 672 67 681 101
rect 636 51 681 67
rect 715 165 762 181
rect 715 131 724 165
rect 758 131 762 165
rect 715 95 762 131
rect 715 61 724 95
rect 758 61 762 95
rect 796 71 833 215
rect 715 17 762 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or3_4
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3189618
string GDS_START 3181942
<< end >>
