magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
rect 483 329 953 331
<< pwell >>
rect 13 49 1137 259
rect 0 0 1248 49
<< scnmos >>
rect 92 65 122 233
rect 178 65 208 233
rect 280 65 310 233
rect 382 65 412 233
rect 484 65 514 233
rect 676 65 706 233
rect 764 65 794 233
rect 856 65 886 233
rect 942 65 972 233
rect 1028 65 1058 233
<< scpmoshvt >>
rect 92 367 122 619
rect 178 367 208 619
rect 264 367 294 619
rect 350 367 380 619
rect 576 365 606 617
rect 662 365 692 617
rect 748 365 778 617
rect 834 365 864 617
rect 1024 367 1054 619
rect 1110 367 1140 619
<< ndiff >>
rect 39 221 92 233
rect 39 187 47 221
rect 81 187 92 221
rect 39 111 92 187
rect 39 77 47 111
rect 81 77 92 111
rect 39 65 92 77
rect 122 225 178 233
rect 122 191 133 225
rect 167 191 178 225
rect 122 153 178 191
rect 122 119 133 153
rect 167 119 178 153
rect 122 65 178 119
rect 208 181 280 233
rect 208 147 235 181
rect 269 147 280 181
rect 208 107 280 147
rect 208 73 235 107
rect 269 73 280 107
rect 208 65 280 73
rect 310 225 382 233
rect 310 191 337 225
rect 371 191 382 225
rect 310 153 382 191
rect 310 119 337 153
rect 371 119 382 153
rect 310 65 382 119
rect 412 181 484 233
rect 412 147 439 181
rect 473 147 484 181
rect 412 107 484 147
rect 412 73 439 107
rect 473 73 484 107
rect 412 65 484 73
rect 514 111 676 233
rect 514 77 539 111
rect 573 77 631 111
rect 665 77 676 111
rect 514 65 676 77
rect 706 208 764 233
rect 706 174 717 208
rect 751 174 764 208
rect 706 113 764 174
rect 706 79 717 113
rect 751 79 764 113
rect 706 65 764 79
rect 794 132 856 233
rect 794 98 805 132
rect 839 98 856 132
rect 794 65 856 98
rect 886 208 942 233
rect 886 174 897 208
rect 931 174 942 208
rect 886 113 942 174
rect 886 79 897 113
rect 931 79 942 113
rect 886 65 942 79
rect 972 132 1028 233
rect 972 98 983 132
rect 1017 98 1028 132
rect 972 65 1028 98
rect 1058 208 1111 233
rect 1058 174 1069 208
rect 1103 174 1111 208
rect 1058 113 1111 174
rect 1058 79 1069 113
rect 1103 79 1111 113
rect 1058 65 1111 79
<< pdiff >>
rect 39 599 92 619
rect 39 565 47 599
rect 81 565 92 599
rect 39 520 92 565
rect 39 486 47 520
rect 81 486 92 520
rect 39 434 92 486
rect 39 400 47 434
rect 81 400 92 434
rect 39 367 92 400
rect 122 543 178 619
rect 122 509 133 543
rect 167 509 178 543
rect 122 420 178 509
rect 122 386 133 420
rect 167 386 178 420
rect 122 367 178 386
rect 208 599 264 619
rect 208 565 219 599
rect 253 565 264 599
rect 208 502 264 565
rect 208 468 219 502
rect 253 468 264 502
rect 208 367 264 468
rect 294 566 350 619
rect 294 532 305 566
rect 339 532 350 566
rect 294 367 350 532
rect 380 599 433 619
rect 380 565 391 599
rect 425 565 433 599
rect 380 486 433 565
rect 380 452 391 486
rect 425 452 433 486
rect 380 367 433 452
rect 519 599 576 617
rect 519 565 527 599
rect 561 565 576 599
rect 519 502 576 565
rect 519 468 527 502
rect 561 468 576 502
rect 519 365 576 468
rect 606 547 662 617
rect 606 513 617 547
rect 651 513 662 547
rect 606 475 662 513
rect 606 441 617 475
rect 651 441 662 475
rect 606 407 662 441
rect 606 373 617 407
rect 651 373 662 407
rect 606 365 662 373
rect 692 599 748 617
rect 692 565 703 599
rect 737 565 748 599
rect 692 499 748 565
rect 692 465 703 499
rect 737 465 748 499
rect 692 413 748 465
rect 692 379 703 413
rect 737 379 748 413
rect 692 365 748 379
rect 778 547 834 617
rect 778 513 789 547
rect 823 513 834 547
rect 778 475 834 513
rect 778 441 789 475
rect 823 441 834 475
rect 778 407 834 441
rect 778 373 789 407
rect 823 373 834 407
rect 778 365 834 373
rect 864 599 917 617
rect 864 565 875 599
rect 909 565 917 599
rect 864 529 917 565
rect 864 495 875 529
rect 909 495 917 529
rect 864 459 917 495
rect 864 425 875 459
rect 909 425 917 459
rect 864 365 917 425
rect 971 607 1024 619
rect 971 573 979 607
rect 1013 573 1024 607
rect 971 526 1024 573
rect 971 492 979 526
rect 1013 492 1024 526
rect 971 443 1024 492
rect 971 409 979 443
rect 1013 409 1024 443
rect 971 367 1024 409
rect 1054 599 1110 619
rect 1054 565 1065 599
rect 1099 565 1110 599
rect 1054 504 1110 565
rect 1054 470 1065 504
rect 1099 470 1110 504
rect 1054 413 1110 470
rect 1054 379 1065 413
rect 1099 379 1110 413
rect 1054 367 1110 379
rect 1140 607 1193 619
rect 1140 573 1151 607
rect 1185 573 1193 607
rect 1140 505 1193 573
rect 1140 471 1151 505
rect 1185 471 1193 505
rect 1140 413 1193 471
rect 1140 379 1151 413
rect 1185 379 1193 413
rect 1140 367 1193 379
<< ndiffc >>
rect 47 187 81 221
rect 47 77 81 111
rect 133 191 167 225
rect 133 119 167 153
rect 235 147 269 181
rect 235 73 269 107
rect 337 191 371 225
rect 337 119 371 153
rect 439 147 473 181
rect 439 73 473 107
rect 539 77 573 111
rect 631 77 665 111
rect 717 174 751 208
rect 717 79 751 113
rect 805 98 839 132
rect 897 174 931 208
rect 897 79 931 113
rect 983 98 1017 132
rect 1069 174 1103 208
rect 1069 79 1103 113
<< pdiffc >>
rect 47 565 81 599
rect 47 486 81 520
rect 47 400 81 434
rect 133 509 167 543
rect 133 386 167 420
rect 219 565 253 599
rect 219 468 253 502
rect 305 532 339 566
rect 391 565 425 599
rect 391 452 425 486
rect 527 565 561 599
rect 527 468 561 502
rect 617 513 651 547
rect 617 441 651 475
rect 617 373 651 407
rect 703 565 737 599
rect 703 465 737 499
rect 703 379 737 413
rect 789 513 823 547
rect 789 441 823 475
rect 789 373 823 407
rect 875 565 909 599
rect 875 495 909 529
rect 875 425 909 459
rect 979 573 1013 607
rect 979 492 1013 526
rect 979 409 1013 443
rect 1065 565 1099 599
rect 1065 470 1099 504
rect 1065 379 1099 413
rect 1151 573 1185 607
rect 1151 471 1185 505
rect 1151 379 1185 413
<< poly >>
rect 92 619 122 645
rect 178 619 208 645
rect 264 619 294 645
rect 350 619 380 645
rect 576 617 606 643
rect 662 617 692 643
rect 748 617 778 643
rect 834 617 864 643
rect 1024 619 1054 645
rect 1110 619 1140 645
rect 92 335 122 367
rect 178 335 208 367
rect 92 319 208 335
rect 92 285 108 319
rect 142 285 208 319
rect 92 269 208 285
rect 264 335 294 367
rect 350 336 380 367
rect 350 335 412 336
rect 264 319 412 335
rect 576 333 606 365
rect 662 333 692 365
rect 264 285 309 319
rect 343 285 412 319
rect 264 269 412 285
rect 92 233 122 269
rect 178 233 208 269
rect 280 233 310 269
rect 382 233 412 269
rect 484 317 706 333
rect 484 283 500 317
rect 534 283 706 317
rect 484 267 706 283
rect 484 233 514 267
rect 676 233 706 267
rect 748 321 778 365
rect 834 321 864 365
rect 1024 321 1054 367
rect 1110 321 1140 367
rect 748 305 900 321
rect 748 271 764 305
rect 798 271 850 305
rect 884 271 900 305
rect 748 255 900 271
rect 942 305 1140 321
rect 942 271 979 305
rect 1013 271 1090 305
rect 1124 271 1140 305
rect 942 255 1140 271
rect 764 233 794 255
rect 856 233 886 255
rect 942 233 972 255
rect 1028 233 1058 255
rect 92 39 122 65
rect 178 39 208 65
rect 280 39 310 65
rect 382 39 412 65
rect 484 39 514 65
rect 676 39 706 65
rect 764 39 794 65
rect 856 39 886 65
rect 942 39 972 65
rect 1028 39 1058 65
<< polycont >>
rect 108 285 142 319
rect 309 285 343 319
rect 500 283 534 317
rect 764 271 798 305
rect 850 271 884 305
rect 979 271 1013 305
rect 1090 271 1124 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 31 599 255 615
rect 31 565 47 599
rect 81 581 219 599
rect 81 565 83 581
rect 31 520 83 565
rect 217 565 219 581
rect 253 565 255 599
rect 31 486 47 520
rect 81 486 83 520
rect 31 434 83 486
rect 31 400 47 434
rect 81 400 83 434
rect 31 384 83 400
rect 117 543 183 547
rect 117 509 133 543
rect 167 509 183 543
rect 117 420 183 509
rect 217 502 255 565
rect 289 566 355 649
rect 289 532 305 566
rect 339 532 355 566
rect 289 524 355 532
rect 389 599 441 615
rect 389 565 391 599
rect 425 565 441 599
rect 217 468 219 502
rect 253 490 255 502
rect 389 490 441 565
rect 253 486 441 490
rect 253 468 391 486
rect 217 452 391 468
rect 425 452 441 486
rect 511 599 925 615
rect 511 565 527 599
rect 561 581 703 599
rect 561 565 565 581
rect 511 502 565 565
rect 701 565 703 581
rect 737 581 875 599
rect 737 565 739 581
rect 511 468 527 502
rect 561 468 565 502
rect 511 452 565 468
rect 601 513 617 547
rect 651 513 667 547
rect 601 475 667 513
rect 117 386 133 420
rect 167 418 183 420
rect 601 441 617 475
rect 651 441 667 475
rect 601 418 667 441
rect 167 407 667 418
rect 167 386 617 407
rect 117 384 617 386
rect 601 373 617 384
rect 651 373 667 407
rect 17 319 259 350
rect 17 285 108 319
rect 142 285 259 319
rect 293 319 366 350
rect 293 285 309 319
rect 343 285 366 319
rect 400 317 567 350
rect 400 283 500 317
rect 534 283 567 317
rect 601 249 667 373
rect 701 499 739 565
rect 873 565 875 581
rect 909 565 925 599
rect 701 465 703 499
rect 737 465 739 499
rect 701 413 739 465
rect 701 379 703 413
rect 737 379 739 413
rect 701 363 739 379
rect 773 513 789 547
rect 823 513 839 547
rect 773 475 839 513
rect 773 441 789 475
rect 823 441 839 475
rect 773 407 839 441
rect 873 529 925 565
rect 873 495 875 529
rect 909 495 925 529
rect 873 459 925 495
rect 873 425 875 459
rect 909 425 925 459
rect 873 409 925 425
rect 963 607 1029 649
rect 963 573 979 607
rect 1013 573 1029 607
rect 963 526 1029 573
rect 963 492 979 526
rect 1013 492 1029 526
rect 963 443 1029 492
rect 963 409 979 443
rect 1013 409 1029 443
rect 1063 599 1108 615
rect 1063 565 1065 599
rect 1099 565 1108 599
rect 1063 504 1108 565
rect 1063 470 1065 504
rect 1099 470 1108 504
rect 1063 413 1108 470
rect 773 373 789 407
rect 823 375 839 407
rect 1063 379 1065 413
rect 1099 379 1108 413
rect 1063 375 1108 379
rect 823 373 1108 375
rect 773 341 1108 373
rect 1142 607 1201 649
rect 1142 573 1151 607
rect 1185 573 1201 607
rect 1142 505 1201 573
rect 1142 471 1151 505
rect 1185 471 1201 505
rect 1142 413 1201 471
rect 1142 379 1151 413
rect 1185 379 1201 413
rect 1142 363 1201 379
rect 31 221 83 237
rect 31 187 47 221
rect 81 187 83 221
rect 31 111 83 187
rect 117 225 667 249
rect 701 271 764 305
rect 798 271 850 305
rect 884 271 929 305
rect 701 242 929 271
rect 963 271 979 305
rect 1013 271 1090 305
rect 1124 271 1231 305
rect 963 242 1231 271
rect 117 191 133 225
rect 167 215 337 225
rect 167 191 183 215
rect 117 153 183 191
rect 321 191 337 215
rect 371 215 667 225
rect 371 191 387 215
rect 117 119 133 153
rect 167 119 183 153
rect 219 147 235 181
rect 269 147 285 181
rect 31 77 47 111
rect 81 85 83 111
rect 219 107 285 147
rect 321 153 387 191
rect 701 181 717 208
rect 321 119 337 153
rect 371 119 387 153
rect 423 147 439 181
rect 473 174 717 181
rect 751 174 897 208
rect 931 174 1069 208
rect 1103 174 1119 208
rect 473 147 755 174
rect 219 85 235 107
rect 81 77 235 85
rect 31 73 235 77
rect 269 85 285 107
rect 423 107 489 147
rect 715 113 755 147
rect 423 85 439 107
rect 269 73 439 85
rect 473 73 489 107
rect 31 51 489 73
rect 523 111 681 113
rect 523 77 539 111
rect 573 77 631 111
rect 665 77 681 111
rect 523 17 681 77
rect 715 79 717 113
rect 751 79 755 113
rect 715 63 755 79
rect 789 132 855 140
rect 789 98 805 132
rect 839 98 855 132
rect 789 17 855 98
rect 893 113 933 174
rect 893 79 897 113
rect 931 79 933 113
rect 893 63 933 79
rect 967 132 1033 140
rect 967 98 983 132
rect 1017 98 1033 132
rect 967 17 1033 98
rect 1067 113 1119 174
rect 1067 79 1069 113
rect 1103 79 1119 113
rect 1067 63 1119 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o32ai_2
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1784468
string GDS_START 1773078
<< end >>
