magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 756 243
rect 0 0 768 49
<< scnmos >>
rect 80 49 110 217
rect 166 49 196 217
rect 356 49 386 217
rect 446 49 476 217
rect 541 49 571 217
rect 647 49 677 217
<< scpmoshvt >>
rect 101 367 131 619
rect 187 367 217 619
rect 356 367 386 619
rect 428 367 458 619
rect 536 367 566 619
rect 647 367 677 619
<< ndiff >>
rect 27 205 80 217
rect 27 171 35 205
rect 69 171 80 205
rect 27 95 80 171
rect 27 61 35 95
rect 69 61 80 95
rect 27 49 80 61
rect 110 205 166 217
rect 110 171 121 205
rect 155 171 166 205
rect 110 101 166 171
rect 110 67 121 101
rect 155 67 166 101
rect 110 49 166 67
rect 196 181 249 217
rect 196 147 207 181
rect 241 147 249 181
rect 196 95 249 147
rect 196 61 207 95
rect 241 61 249 95
rect 196 49 249 61
rect 303 179 356 217
rect 303 145 311 179
rect 345 145 356 179
rect 303 95 356 145
rect 303 61 311 95
rect 345 61 356 95
rect 303 49 356 61
rect 386 169 446 217
rect 386 135 401 169
rect 435 135 446 169
rect 386 49 446 135
rect 476 205 541 217
rect 476 171 491 205
rect 525 171 541 205
rect 476 101 541 171
rect 476 67 491 101
rect 525 67 541 101
rect 476 49 541 67
rect 571 165 647 217
rect 571 131 591 165
rect 625 131 647 165
rect 571 91 647 131
rect 571 57 591 91
rect 625 57 647 91
rect 571 49 647 57
rect 677 205 730 217
rect 677 171 688 205
rect 722 171 730 205
rect 677 101 730 171
rect 677 67 688 101
rect 722 67 730 101
rect 677 49 730 67
<< pdiff >>
rect 43 607 101 619
rect 43 573 56 607
rect 90 573 101 607
rect 43 532 101 573
rect 43 498 56 532
rect 90 498 101 532
rect 43 449 101 498
rect 43 415 56 449
rect 90 415 101 449
rect 43 367 101 415
rect 131 599 187 619
rect 131 565 142 599
rect 176 565 187 599
rect 131 504 187 565
rect 131 470 142 504
rect 176 470 187 504
rect 131 413 187 470
rect 131 379 142 413
rect 176 379 187 413
rect 131 367 187 379
rect 217 607 356 619
rect 217 573 228 607
rect 262 573 311 607
rect 345 573 356 607
rect 217 492 356 573
rect 217 458 228 492
rect 262 458 311 492
rect 345 458 356 492
rect 217 367 356 458
rect 386 367 428 619
rect 458 599 536 619
rect 458 565 479 599
rect 513 565 536 599
rect 458 519 536 565
rect 458 485 479 519
rect 513 485 536 519
rect 458 436 536 485
rect 458 402 479 436
rect 513 402 536 436
rect 458 367 536 402
rect 566 367 647 619
rect 677 607 730 619
rect 677 573 688 607
rect 722 573 730 607
rect 677 518 730 573
rect 677 484 688 518
rect 722 484 730 518
rect 677 434 730 484
rect 677 400 688 434
rect 722 400 730 434
rect 677 367 730 400
<< ndiffc >>
rect 35 171 69 205
rect 35 61 69 95
rect 121 171 155 205
rect 121 67 155 101
rect 207 147 241 181
rect 207 61 241 95
rect 311 145 345 179
rect 311 61 345 95
rect 401 135 435 169
rect 491 171 525 205
rect 491 67 525 101
rect 591 131 625 165
rect 591 57 625 91
rect 688 171 722 205
rect 688 67 722 101
<< pdiffc >>
rect 56 573 90 607
rect 56 498 90 532
rect 56 415 90 449
rect 142 565 176 599
rect 142 470 176 504
rect 142 379 176 413
rect 228 573 262 607
rect 311 573 345 607
rect 228 458 262 492
rect 311 458 345 492
rect 479 565 513 599
rect 479 485 513 519
rect 479 402 513 436
rect 688 573 722 607
rect 688 484 722 518
rect 688 400 722 434
<< poly >>
rect 101 619 131 645
rect 187 619 217 645
rect 356 619 386 645
rect 428 619 458 645
rect 536 619 566 645
rect 647 619 677 645
rect 101 315 131 367
rect 187 315 217 367
rect 356 335 386 367
rect 313 319 386 335
rect 101 299 262 315
rect 101 279 212 299
rect 80 265 212 279
rect 246 265 262 299
rect 313 285 329 319
rect 363 285 386 319
rect 313 269 386 285
rect 428 335 458 367
rect 536 335 566 367
rect 428 319 494 335
rect 428 285 444 319
rect 478 285 494 319
rect 428 269 494 285
rect 536 319 602 335
rect 536 285 552 319
rect 586 285 602 319
rect 536 269 602 285
rect 647 325 677 367
rect 647 309 743 325
rect 647 275 693 309
rect 727 275 743 309
rect 80 249 262 265
rect 80 217 110 249
rect 166 217 196 249
rect 356 217 386 269
rect 446 217 476 269
rect 541 217 571 269
rect 647 259 743 275
rect 647 217 677 259
rect 80 23 110 49
rect 166 23 196 49
rect 356 23 386 49
rect 446 23 476 49
rect 541 23 571 49
rect 647 23 677 49
<< polycont >>
rect 212 265 246 299
rect 329 285 363 319
rect 444 285 478 319
rect 552 285 586 319
rect 693 275 727 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 40 607 90 649
rect 40 573 56 607
rect 40 532 90 573
rect 40 498 56 532
rect 40 449 90 498
rect 40 415 56 449
rect 40 399 90 415
rect 124 599 176 615
rect 124 565 142 599
rect 124 504 176 565
rect 124 470 142 504
rect 124 413 176 470
rect 212 607 361 649
rect 212 573 228 607
rect 262 573 311 607
rect 345 573 361 607
rect 212 492 361 573
rect 212 458 228 492
rect 262 458 311 492
rect 345 458 361 492
rect 212 454 361 458
rect 449 599 518 615
rect 449 565 479 599
rect 513 565 518 599
rect 675 607 738 649
rect 449 519 518 565
rect 449 485 479 519
rect 513 485 518 519
rect 449 436 518 485
rect 449 420 479 436
rect 124 379 142 413
rect 124 365 176 379
rect 19 205 73 221
rect 19 171 35 205
rect 69 171 73 205
rect 19 95 73 171
rect 19 61 35 95
rect 69 61 73 95
rect 19 17 73 61
rect 107 215 176 365
rect 210 402 479 420
rect 513 402 518 436
rect 210 386 518 402
rect 210 299 262 386
rect 210 265 212 299
rect 246 265 262 299
rect 296 319 379 350
rect 296 285 329 319
rect 363 285 379 319
rect 415 319 494 350
rect 415 285 444 319
rect 478 285 494 319
rect 552 319 641 588
rect 675 573 688 607
rect 722 573 738 607
rect 675 518 738 573
rect 675 484 688 518
rect 722 484 738 518
rect 675 434 738 484
rect 675 400 688 434
rect 722 400 738 434
rect 675 384 738 400
rect 586 285 641 319
rect 552 269 641 285
rect 677 309 751 350
rect 677 275 693 309
rect 727 275 751 309
rect 210 249 262 265
rect 210 215 441 249
rect 107 205 155 215
rect 107 171 121 205
rect 107 101 155 171
rect 107 67 121 101
rect 107 51 155 67
rect 191 147 207 181
rect 241 147 257 181
rect 191 95 257 147
rect 191 61 207 95
rect 241 61 257 95
rect 191 17 257 61
rect 295 145 311 179
rect 345 145 361 179
rect 295 95 361 145
rect 395 169 441 215
rect 395 135 401 169
rect 435 135 441 169
rect 395 119 441 135
rect 475 205 738 233
rect 475 171 491 205
rect 525 199 688 205
rect 525 171 541 199
rect 295 61 311 95
rect 345 85 361 95
rect 475 101 541 171
rect 675 171 688 199
rect 722 171 738 205
rect 475 85 491 101
rect 345 67 491 85
rect 525 67 541 101
rect 345 61 541 67
rect 295 51 541 61
rect 575 131 591 165
rect 625 131 641 165
rect 575 91 641 131
rect 575 57 591 91
rect 625 57 641 91
rect 575 17 641 57
rect 675 101 738 171
rect 675 67 688 101
rect 722 67 738 101
rect 675 51 738 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o22a_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 975574
string GDS_START 967794
<< end >>
