magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 4 49 758 167
rect 0 0 768 49
<< scnmos >>
rect 87 57 117 141
rect 159 57 189 141
rect 245 57 275 141
rect 323 57 353 141
rect 409 57 439 141
rect 481 57 511 141
rect 567 57 597 141
rect 645 57 675 141
<< scpmoshvt >>
rect 87 409 137 609
rect 347 409 397 609
rect 445 409 495 609
rect 608 409 658 609
<< ndiff >>
rect 30 116 87 141
rect 30 82 42 116
rect 76 82 87 116
rect 30 57 87 82
rect 117 57 159 141
rect 189 108 245 141
rect 189 74 200 108
rect 234 74 245 108
rect 189 57 245 74
rect 275 57 323 141
rect 353 116 409 141
rect 353 82 364 116
rect 398 82 409 116
rect 353 57 409 82
rect 439 57 481 141
rect 511 112 567 141
rect 511 78 522 112
rect 556 78 567 112
rect 511 57 567 78
rect 597 57 645 141
rect 675 116 732 141
rect 675 82 686 116
rect 720 82 732 116
rect 675 57 732 82
<< pdiff >>
rect 30 597 87 609
rect 30 563 42 597
rect 76 563 87 597
rect 30 526 87 563
rect 30 492 42 526
rect 76 492 87 526
rect 30 455 87 492
rect 30 421 42 455
rect 76 421 87 455
rect 30 409 87 421
rect 137 597 194 609
rect 137 563 148 597
rect 182 563 194 597
rect 137 526 194 563
rect 137 492 148 526
rect 182 492 194 526
rect 137 455 194 492
rect 137 421 148 455
rect 182 421 194 455
rect 137 409 194 421
rect 290 597 347 609
rect 290 563 302 597
rect 336 563 347 597
rect 290 526 347 563
rect 290 492 302 526
rect 336 492 347 526
rect 290 455 347 492
rect 290 421 302 455
rect 336 421 347 455
rect 290 409 347 421
rect 397 409 445 609
rect 495 597 608 609
rect 495 563 563 597
rect 597 563 608 597
rect 495 526 608 563
rect 495 492 563 526
rect 597 492 608 526
rect 495 455 608 492
rect 495 421 563 455
rect 597 421 608 455
rect 495 409 608 421
rect 658 597 715 609
rect 658 563 669 597
rect 703 563 715 597
rect 658 526 715 563
rect 658 492 669 526
rect 703 492 715 526
rect 658 455 715 492
rect 658 421 669 455
rect 703 421 715 455
rect 658 409 715 421
<< ndiffc >>
rect 42 82 76 116
rect 200 74 234 108
rect 364 82 398 116
rect 522 78 556 112
rect 686 82 720 116
<< pdiffc >>
rect 42 563 76 597
rect 42 492 76 526
rect 42 421 76 455
rect 148 563 182 597
rect 148 492 182 526
rect 148 421 182 455
rect 302 563 336 597
rect 302 492 336 526
rect 302 421 336 455
rect 563 563 597 597
rect 563 492 597 526
rect 563 421 597 455
rect 669 563 703 597
rect 669 492 703 526
rect 669 421 703 455
<< poly >>
rect 87 609 137 635
rect 347 609 397 635
rect 445 609 495 635
rect 608 609 658 635
rect 87 369 137 409
rect 87 353 178 369
rect 87 319 128 353
rect 162 319 178 353
rect 87 285 178 319
rect 347 299 397 409
rect 87 251 128 285
rect 162 265 178 285
rect 237 283 397 299
rect 162 251 189 265
rect 87 235 189 251
rect 87 141 117 235
rect 159 141 189 235
rect 237 249 253 283
rect 287 269 397 283
rect 445 377 495 409
rect 445 361 511 377
rect 445 327 461 361
rect 495 327 511 361
rect 445 293 511 327
rect 608 307 658 409
rect 287 249 353 269
rect 237 215 353 249
rect 445 259 461 293
rect 495 259 511 293
rect 445 243 511 259
rect 237 181 253 215
rect 287 181 353 215
rect 481 186 511 243
rect 237 165 353 181
rect 245 141 275 165
rect 323 141 353 165
rect 409 156 511 186
rect 409 141 439 156
rect 481 141 511 156
rect 567 291 638 307
rect 567 257 583 291
rect 617 257 638 291
rect 567 223 638 257
rect 567 189 583 223
rect 617 203 638 223
rect 617 189 675 203
rect 567 173 675 189
rect 567 141 597 173
rect 645 141 675 173
rect 87 31 117 57
rect 159 31 189 57
rect 245 31 275 57
rect 323 31 353 57
rect 409 31 439 57
rect 481 31 511 57
rect 567 31 597 57
rect 645 31 675 57
<< polycont >>
rect 128 319 162 353
rect 128 251 162 285
rect 253 249 287 283
rect 461 327 495 361
rect 461 259 495 293
rect 253 181 287 215
rect 583 257 617 291
rect 583 189 617 223
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 26 597 76 613
rect 26 563 42 597
rect 26 526 76 563
rect 26 492 42 526
rect 26 455 76 492
rect 26 421 42 455
rect 26 199 76 421
rect 132 597 198 649
rect 132 563 148 597
rect 182 563 198 597
rect 132 526 198 563
rect 132 492 148 526
rect 182 492 198 526
rect 132 455 198 492
rect 132 421 148 455
rect 182 421 198 455
rect 132 405 198 421
rect 286 597 373 613
rect 286 563 302 597
rect 336 563 373 597
rect 547 597 613 649
rect 286 526 373 563
rect 286 492 302 526
rect 336 492 373 526
rect 286 455 373 492
rect 286 421 302 455
rect 336 421 373 455
rect 286 405 373 421
rect 112 353 178 369
rect 112 319 128 353
rect 162 319 178 353
rect 112 285 178 319
rect 112 251 128 285
rect 162 251 178 285
rect 112 235 178 251
rect 237 283 303 299
rect 237 249 253 283
rect 287 249 303 283
rect 237 215 303 249
rect 237 199 253 215
rect 26 181 253 199
rect 287 181 303 215
rect 26 165 303 181
rect 339 207 373 405
rect 409 361 511 578
rect 547 563 563 597
rect 597 563 613 597
rect 547 526 613 563
rect 547 492 563 526
rect 597 492 613 526
rect 547 455 613 492
rect 547 421 563 455
rect 597 421 613 455
rect 547 405 613 421
rect 653 597 743 613
rect 653 563 669 597
rect 703 563 743 597
rect 653 526 743 563
rect 653 492 669 526
rect 703 492 743 526
rect 653 455 743 492
rect 653 421 669 455
rect 703 421 743 455
rect 653 405 743 421
rect 409 327 461 361
rect 495 327 511 361
rect 409 293 511 327
rect 409 259 461 293
rect 495 259 511 293
rect 409 243 511 259
rect 567 291 633 307
rect 567 257 583 291
rect 617 257 633 291
rect 567 223 633 257
rect 567 207 583 223
rect 339 189 583 207
rect 617 189 633 223
rect 339 173 633 189
rect 26 116 92 165
rect 26 82 42 116
rect 76 82 92 116
rect 26 53 92 82
rect 184 108 250 129
rect 184 74 200 108
rect 234 74 250 108
rect 184 17 250 74
rect 339 116 414 173
rect 339 82 364 116
rect 398 82 414 116
rect 339 53 414 82
rect 506 112 572 137
rect 506 78 522 112
rect 556 78 572 112
rect 506 17 572 78
rect 670 116 743 405
rect 670 82 686 116
rect 720 82 743 116
rect 670 53 743 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or2b_lp
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2244936
string GDS_START 2237600
<< end >>
