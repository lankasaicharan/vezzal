magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 479 158 863 252
rect 3 49 863 158
rect 0 0 864 49
<< scnmos >>
rect 86 48 116 132
rect 158 48 188 132
rect 244 48 274 132
rect 322 48 352 132
rect 574 142 604 226
rect 664 142 694 226
rect 750 142 780 226
<< scpmoshvt >>
rect 86 416 136 616
rect 248 416 298 616
rect 360 416 410 616
rect 518 416 568 616
rect 624 416 674 616
rect 730 416 780 616
<< ndiff >>
rect 29 111 86 132
rect 29 77 41 111
rect 75 77 86 111
rect 29 48 86 77
rect 116 48 158 132
rect 188 107 244 132
rect 188 73 199 107
rect 233 73 244 107
rect 188 48 244 73
rect 274 48 322 132
rect 352 111 409 132
rect 352 77 363 111
rect 397 77 409 111
rect 505 209 574 226
rect 505 175 517 209
rect 551 175 574 209
rect 505 142 574 175
rect 604 201 664 226
rect 604 167 619 201
rect 653 167 664 201
rect 604 142 664 167
rect 694 188 750 226
rect 694 154 705 188
rect 739 154 750 188
rect 694 142 750 154
rect 780 209 837 226
rect 780 175 791 209
rect 825 175 837 209
rect 780 142 837 175
rect 352 48 409 77
<< pdiff >>
rect 29 597 86 616
rect 29 563 41 597
rect 75 563 86 597
rect 29 462 86 563
rect 29 428 41 462
rect 75 428 86 462
rect 29 416 86 428
rect 136 603 248 616
rect 136 569 147 603
rect 181 569 248 603
rect 136 416 248 569
rect 298 462 360 616
rect 298 428 315 462
rect 349 428 360 462
rect 298 416 360 428
rect 410 603 518 616
rect 410 569 421 603
rect 455 569 518 603
rect 410 416 518 569
rect 568 597 624 616
rect 568 563 579 597
rect 613 563 624 597
rect 568 462 624 563
rect 568 428 579 462
rect 613 428 624 462
rect 568 416 624 428
rect 674 416 730 616
rect 780 604 837 616
rect 780 570 791 604
rect 825 570 837 604
rect 780 533 837 570
rect 780 499 791 533
rect 825 499 837 533
rect 780 462 837 499
rect 780 428 791 462
rect 825 428 837 462
rect 780 416 837 428
<< ndiffc >>
rect 41 77 75 111
rect 199 73 233 107
rect 363 77 397 111
rect 517 175 551 209
rect 619 167 653 201
rect 705 154 739 188
rect 791 175 825 209
<< pdiffc >>
rect 41 563 75 597
rect 41 428 75 462
rect 147 569 181 603
rect 315 428 349 462
rect 421 569 455 603
rect 579 563 613 597
rect 579 428 613 462
rect 791 570 825 604
rect 791 499 825 533
rect 791 428 825 462
<< poly >>
rect 86 616 136 642
rect 248 616 298 642
rect 360 616 410 642
rect 518 616 568 642
rect 624 616 674 642
rect 730 616 780 642
rect 86 286 136 416
rect 248 376 298 416
rect 360 376 410 416
rect 197 360 298 376
rect 197 326 213 360
rect 247 326 298 360
rect 197 310 298 326
rect 346 360 412 376
rect 518 366 568 416
rect 624 376 674 416
rect 730 376 780 416
rect 346 326 362 360
rect 396 326 412 360
rect 86 238 116 286
rect 86 222 193 238
rect 86 188 143 222
rect 177 188 193 222
rect 86 172 193 188
rect 86 132 116 172
rect 158 132 188 172
rect 244 132 274 310
rect 346 292 412 326
rect 346 258 362 292
rect 396 258 412 292
rect 346 242 412 258
rect 460 350 568 366
rect 460 316 507 350
rect 541 316 568 350
rect 460 300 568 316
rect 616 360 682 376
rect 616 326 632 360
rect 666 326 682 360
rect 616 310 682 326
rect 730 360 796 376
rect 730 326 746 360
rect 780 326 796 360
rect 730 310 796 326
rect 346 177 376 242
rect 322 147 376 177
rect 322 132 352 147
rect 460 119 490 300
rect 652 271 682 310
rect 574 226 604 252
rect 652 241 694 271
rect 664 226 694 241
rect 750 226 780 310
rect 574 119 604 142
rect 460 103 604 119
rect 664 116 694 142
rect 750 116 780 142
rect 460 89 517 103
rect 501 69 517 89
rect 551 69 604 103
rect 501 53 604 69
rect 86 22 116 48
rect 158 22 188 48
rect 244 22 274 48
rect 322 22 352 48
<< polycont >>
rect 213 326 247 360
rect 362 326 396 360
rect 143 188 177 222
rect 362 258 396 292
rect 507 316 541 350
rect 632 326 666 360
rect 746 326 780 360
rect 517 69 551 103
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 25 597 91 613
rect 25 563 41 597
rect 75 563 91 597
rect 131 603 197 649
rect 131 569 147 603
rect 181 569 197 603
rect 131 568 197 569
rect 405 603 471 649
rect 405 569 421 603
rect 455 569 471 603
rect 405 568 471 569
rect 563 597 629 613
rect 25 462 91 563
rect 563 563 579 597
rect 613 563 629 597
rect 563 532 629 563
rect 25 428 41 462
rect 75 428 91 462
rect 25 111 91 428
rect 127 498 629 532
rect 127 238 161 498
rect 563 462 629 498
rect 197 360 263 430
rect 299 428 315 462
rect 349 428 525 462
rect 299 412 525 428
rect 563 428 579 462
rect 613 428 629 462
rect 563 412 629 428
rect 775 604 841 649
rect 775 570 791 604
rect 825 570 841 604
rect 775 533 841 570
rect 775 499 791 533
rect 825 499 841 533
rect 775 462 841 499
rect 775 428 791 462
rect 825 428 841 462
rect 775 412 841 428
rect 197 326 213 360
rect 247 326 263 360
rect 197 310 263 326
rect 313 360 455 376
rect 313 326 362 360
rect 396 326 455 360
rect 313 292 455 326
rect 491 366 525 412
rect 491 350 557 366
rect 491 316 507 350
rect 541 316 557 350
rect 491 300 557 316
rect 601 360 682 376
rect 601 326 632 360
rect 666 326 682 360
rect 601 310 682 326
rect 730 360 844 376
rect 730 326 746 360
rect 780 326 844 360
rect 730 310 844 326
rect 313 258 362 292
rect 396 258 455 292
rect 313 242 455 258
rect 603 240 841 274
rect 127 222 193 238
rect 127 188 143 222
rect 177 206 193 222
rect 501 209 567 230
rect 501 206 517 209
rect 177 188 517 206
rect 127 175 517 188
rect 551 175 567 209
rect 127 172 567 175
rect 501 155 567 172
rect 603 201 653 240
rect 775 209 841 240
rect 603 167 619 201
rect 603 138 653 167
rect 689 188 739 204
rect 689 154 705 188
rect 775 175 791 209
rect 825 175 841 209
rect 775 170 841 175
rect 25 77 41 111
rect 75 77 91 111
rect 25 53 91 77
rect 183 107 249 136
rect 183 73 199 107
rect 233 73 249 107
rect 183 17 249 73
rect 347 119 413 136
rect 347 111 567 119
rect 347 77 363 111
rect 397 103 567 111
rect 397 77 517 103
rect 347 69 517 77
rect 551 69 567 103
rect 347 53 567 69
rect 689 17 739 154
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2bb2a_lp
flabel comment s 536 103 536 103 0 FreeSans 200 180 0 0 no_jumper_check
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3650056
string GDS_START 3642460
<< end >>
