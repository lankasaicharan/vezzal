magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
<< pwell >>
rect 23 239 1038 241
rect 23 49 1247 239
rect 0 0 1248 49
<< scnmos >>
rect 106 131 136 215
rect 254 47 284 215
rect 340 47 370 215
rect 426 47 456 215
rect 512 47 542 215
rect 641 47 671 215
rect 713 47 743 215
rect 821 47 851 215
rect 929 47 959 215
rect 1138 129 1168 213
<< scpmoshvt >>
rect 106 367 136 451
rect 254 367 284 619
rect 340 367 370 619
rect 426 367 456 619
rect 512 367 542 619
rect 627 367 657 619
rect 713 367 743 619
rect 821 367 851 619
rect 929 367 959 619
rect 1037 367 1067 451
<< ndiff >>
rect 49 190 106 215
rect 49 156 57 190
rect 91 156 106 190
rect 49 131 106 156
rect 136 165 254 215
rect 136 131 209 165
rect 243 131 254 165
rect 201 93 254 131
rect 201 59 209 93
rect 243 59 254 93
rect 201 47 254 59
rect 284 203 340 215
rect 284 169 295 203
rect 329 169 340 203
rect 284 101 340 169
rect 284 67 295 101
rect 329 67 340 101
rect 284 47 340 67
rect 370 179 426 215
rect 370 145 381 179
rect 415 145 426 179
rect 370 93 426 145
rect 370 59 381 93
rect 415 59 426 93
rect 370 47 426 59
rect 456 203 512 215
rect 456 169 467 203
rect 501 169 512 203
rect 456 101 512 169
rect 456 67 467 101
rect 501 67 512 101
rect 456 47 512 67
rect 542 124 641 215
rect 542 90 574 124
rect 608 90 641 124
rect 542 47 641 90
rect 671 47 713 215
rect 743 47 821 215
rect 851 47 929 215
rect 959 175 1012 215
rect 959 141 970 175
rect 1004 141 1012 175
rect 959 101 1012 141
rect 1085 177 1138 213
rect 1085 143 1093 177
rect 1127 143 1138 177
rect 1085 129 1138 143
rect 1168 189 1221 213
rect 1168 155 1179 189
rect 1213 155 1221 189
rect 1168 129 1221 155
rect 959 67 970 101
rect 1004 67 1012 101
rect 959 47 1012 67
<< pdiff >>
rect 201 607 254 619
rect 201 573 209 607
rect 243 573 254 607
rect 201 451 254 573
rect 49 426 106 451
rect 49 392 57 426
rect 91 392 106 426
rect 49 367 106 392
rect 136 367 254 451
rect 284 413 340 619
rect 284 379 295 413
rect 329 379 340 413
rect 284 367 340 379
rect 370 607 426 619
rect 370 573 381 607
rect 415 573 426 607
rect 370 367 426 573
rect 456 413 512 619
rect 456 379 467 413
rect 501 379 512 413
rect 456 367 512 379
rect 542 607 627 619
rect 542 573 569 607
rect 603 573 627 607
rect 542 367 627 573
rect 657 443 713 619
rect 657 409 668 443
rect 702 409 713 443
rect 657 367 713 409
rect 743 607 821 619
rect 743 573 766 607
rect 800 573 821 607
rect 743 367 821 573
rect 851 443 929 619
rect 851 409 873 443
rect 907 409 929 443
rect 851 367 929 409
rect 959 607 1012 619
rect 959 573 970 607
rect 1004 573 1012 607
rect 959 451 1012 573
rect 959 367 1037 451
rect 1067 436 1120 451
rect 1067 402 1078 436
rect 1112 402 1120 436
rect 1067 367 1120 402
<< ndiffc >>
rect 57 156 91 190
rect 209 131 243 165
rect 209 59 243 93
rect 295 169 329 203
rect 295 67 329 101
rect 381 145 415 179
rect 381 59 415 93
rect 467 169 501 203
rect 467 67 501 101
rect 574 90 608 124
rect 970 141 1004 175
rect 1093 143 1127 177
rect 1179 155 1213 189
rect 970 67 1004 101
<< pdiffc >>
rect 209 573 243 607
rect 57 392 91 426
rect 295 379 329 413
rect 381 573 415 607
rect 467 379 501 413
rect 569 573 603 607
rect 668 409 702 443
rect 766 573 800 607
rect 873 409 907 443
rect 970 573 1004 607
rect 1078 402 1112 436
<< poly >>
rect 254 619 284 645
rect 340 619 370 645
rect 426 619 456 645
rect 512 619 542 645
rect 627 619 657 645
rect 713 619 743 645
rect 821 619 851 645
rect 929 619 959 645
rect 106 451 136 477
rect 1037 451 1067 477
rect 106 303 136 367
rect 254 333 284 367
rect 340 333 370 367
rect 426 333 456 367
rect 512 333 542 367
rect 254 317 563 333
rect 106 287 177 303
rect 106 253 127 287
rect 161 253 177 287
rect 106 237 177 253
rect 254 283 309 317
rect 343 283 377 317
rect 411 283 445 317
rect 479 283 513 317
rect 547 283 563 317
rect 627 308 657 367
rect 713 308 743 367
rect 821 335 851 367
rect 821 319 887 335
rect 254 267 563 283
rect 605 292 671 308
rect 106 215 136 237
rect 254 215 284 267
rect 340 215 370 267
rect 426 215 456 267
rect 512 215 542 267
rect 605 258 621 292
rect 655 258 671 292
rect 605 242 671 258
rect 641 215 671 242
rect 713 292 779 308
rect 713 258 729 292
rect 763 258 779 292
rect 713 242 779 258
rect 821 285 837 319
rect 871 285 887 319
rect 821 269 887 285
rect 929 303 959 367
rect 1037 335 1067 367
rect 1037 319 1204 335
rect 1037 305 1154 319
rect 929 287 995 303
rect 713 215 743 242
rect 821 215 851 269
rect 929 253 945 287
rect 979 253 995 287
rect 929 237 995 253
rect 1138 285 1154 305
rect 1188 285 1204 319
rect 1138 269 1204 285
rect 929 215 959 237
rect 106 105 136 131
rect 1138 213 1168 269
rect 1138 103 1168 129
rect 254 21 284 47
rect 340 21 370 47
rect 426 21 456 47
rect 512 21 542 47
rect 641 21 671 47
rect 713 21 743 47
rect 821 21 851 47
rect 929 21 959 47
<< polycont >>
rect 127 253 161 287
rect 309 283 343 317
rect 377 283 411 317
rect 445 283 479 317
rect 513 283 547 317
rect 621 258 655 292
rect 729 258 763 292
rect 837 285 871 319
rect 945 253 979 287
rect 1154 285 1188 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 193 607 259 649
rect 193 573 209 607
rect 243 573 259 607
rect 193 563 259 573
rect 365 607 431 649
rect 365 573 381 607
rect 415 573 431 607
rect 365 563 431 573
rect 553 607 619 649
rect 553 573 569 607
rect 603 573 619 607
rect 553 563 619 573
rect 750 607 816 649
rect 750 573 766 607
rect 800 573 816 607
rect 750 563 816 573
rect 954 607 1020 649
rect 954 573 970 607
rect 1004 573 1020 607
rect 954 563 1020 573
rect 41 493 992 529
rect 41 426 91 493
rect 537 443 922 459
rect 41 392 57 426
rect 41 190 91 392
rect 41 156 57 190
rect 41 140 91 156
rect 125 287 171 424
rect 125 253 127 287
rect 161 253 171 287
rect 125 94 171 253
rect 223 413 501 429
rect 223 379 295 413
rect 329 379 467 413
rect 223 363 501 379
rect 537 409 668 443
rect 702 409 873 443
rect 907 409 922 443
rect 537 393 922 409
rect 223 249 259 363
rect 537 329 571 393
rect 293 317 571 329
rect 293 283 309 317
rect 343 283 377 317
rect 411 283 445 317
rect 479 283 513 317
rect 547 283 571 317
rect 223 215 503 249
rect 285 203 331 215
rect 205 165 251 181
rect 205 131 209 165
rect 243 131 251 165
rect 205 93 251 131
rect 205 59 209 93
rect 243 59 251 93
rect 205 17 251 59
rect 285 169 295 203
rect 329 169 331 203
rect 465 203 503 215
rect 285 101 331 169
rect 285 67 295 101
rect 329 67 331 101
rect 285 51 331 67
rect 365 179 431 181
rect 365 145 381 179
rect 415 145 431 179
rect 365 93 431 145
rect 365 59 381 93
rect 415 59 431 93
rect 365 17 431 59
rect 465 169 467 203
rect 501 169 503 203
rect 537 208 571 283
rect 607 292 662 359
rect 607 258 621 292
rect 655 258 662 292
rect 607 242 662 258
rect 696 292 780 358
rect 958 357 992 493
rect 696 258 729 292
rect 763 258 780 292
rect 821 323 992 357
rect 1068 436 1128 452
rect 1068 402 1078 436
rect 1112 402 1128 436
rect 1068 386 1128 402
rect 821 319 889 323
rect 821 285 837 319
rect 871 285 889 319
rect 821 269 889 285
rect 929 287 995 289
rect 696 242 780 258
rect 929 253 945 287
rect 979 253 995 287
rect 929 249 995 253
rect 1068 249 1102 386
rect 1138 319 1228 352
rect 1138 285 1154 319
rect 1188 285 1228 319
rect 929 215 1229 249
rect 537 181 881 208
rect 1177 189 1229 215
rect 537 175 1020 181
rect 537 174 970 175
rect 465 101 503 169
rect 692 141 970 174
rect 1004 141 1020 175
rect 465 67 467 101
rect 501 67 503 101
rect 465 51 503 67
rect 558 124 624 140
rect 558 90 574 124
rect 608 90 624 124
rect 558 17 624 90
rect 692 101 1020 141
rect 692 67 970 101
rect 1004 67 1020 101
rect 692 51 1020 67
rect 1077 177 1143 181
rect 1077 143 1093 177
rect 1127 143 1143 177
rect 1077 17 1143 143
rect 1177 155 1179 189
rect 1213 155 1229 189
rect 1177 139 1229 155
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4bb_4
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5243728
string GDS_START 5234652
<< end >>
