magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4562 1975
<< nwell >>
rect -38 331 3302 704
rect 1341 305 2358 331
<< pwell >>
rect 208 198 318 211
rect 490 198 1740 229
rect 12 176 1740 198
rect 12 157 1881 176
rect 2837 157 3263 200
rect 12 49 3263 157
rect 0 0 3264 49
<< scnmos >>
rect 111 88 141 172
rect 189 88 219 172
rect 307 88 337 172
rect 385 88 415 172
rect 471 88 501 172
rect 667 119 697 203
rect 739 119 769 203
rect 929 119 959 203
rect 1001 119 1031 203
rect 1119 119 1149 203
rect 1191 119 1221 203
rect 1402 119 1432 203
rect 1531 119 1561 203
rect 1605 119 1635 203
rect 1729 66 1759 150
rect 1870 47 1900 131
rect 1948 47 1978 131
rect 2062 47 2092 131
rect 2369 47 2399 131
rect 2477 47 2507 131
rect 2631 47 2661 131
rect 2709 47 2739 131
rect 2920 90 2950 174
rect 2992 90 3022 174
rect 3078 90 3108 174
rect 3150 90 3180 174
<< scpmoshvt >>
rect 173 419 223 619
rect 271 419 321 619
rect 389 419 439 619
rect 493 419 543 619
rect 599 419 649 619
rect 722 419 772 619
rect 945 408 995 608
rect 1097 408 1147 608
rect 1447 347 1497 547
rect 1583 347 1633 547
rect 1675 347 1725 547
rect 1781 347 1831 547
rect 2077 341 2127 541
rect 2199 341 2249 541
rect 2337 419 2387 619
rect 2435 419 2485 619
rect 2654 419 2704 619
rect 2760 419 2810 619
rect 2978 388 3028 588
rect 3084 388 3134 588
<< ndiff >>
rect 234 173 292 185
rect 234 172 246 173
rect 38 88 111 172
rect 141 88 189 172
rect 219 139 246 172
rect 280 172 292 173
rect 516 172 667 203
rect 280 139 307 172
rect 219 88 307 139
rect 337 88 385 172
rect 415 147 471 172
rect 415 113 426 147
rect 460 113 471 147
rect 415 88 471 113
rect 501 147 667 172
rect 501 113 528 147
rect 562 119 667 147
rect 697 119 739 203
rect 769 169 822 203
rect 769 135 780 169
rect 814 135 822 169
rect 769 119 822 135
rect 876 178 929 203
rect 876 144 884 178
rect 918 144 929 178
rect 876 119 929 144
rect 959 119 1001 203
rect 1031 141 1119 203
rect 1031 119 1058 141
rect 562 113 652 119
rect 501 88 652 113
rect 1046 107 1058 119
rect 1092 119 1119 141
rect 1149 119 1191 203
rect 1221 175 1278 203
rect 1221 141 1232 175
rect 1266 141 1278 175
rect 1221 119 1278 141
rect 1345 175 1402 203
rect 1345 141 1357 175
rect 1391 141 1402 175
rect 1345 119 1402 141
rect 1432 175 1531 203
rect 1432 141 1443 175
rect 1477 141 1531 175
rect 1432 119 1531 141
rect 1561 119 1605 203
rect 1635 150 1714 203
rect 1635 119 1729 150
rect 1092 107 1104 119
rect 1046 91 1104 107
rect 38 87 96 88
rect 38 53 50 87
rect 84 53 96 87
rect 38 41 96 53
rect 1650 66 1729 119
rect 1759 131 1855 150
rect 2863 149 2920 174
rect 1759 73 1870 131
rect 1759 66 1786 73
rect 1774 39 1786 66
rect 1820 47 1870 73
rect 1900 47 1948 131
rect 1978 89 2062 131
rect 1978 55 2017 89
rect 2051 55 2062 89
rect 1978 47 2062 55
rect 2092 111 2369 131
rect 2092 77 2318 111
rect 2352 77 2369 111
rect 2092 47 2369 77
rect 2399 47 2477 131
rect 2507 97 2631 131
rect 2507 63 2543 97
rect 2577 63 2631 97
rect 2507 47 2631 63
rect 2661 47 2709 131
rect 2739 97 2796 131
rect 2739 63 2750 97
rect 2784 63 2796 97
rect 2863 115 2875 149
rect 2909 115 2920 149
rect 2863 90 2920 115
rect 2950 90 2992 174
rect 3022 149 3078 174
rect 3022 115 3033 149
rect 3067 115 3078 149
rect 3022 90 3078 115
rect 3108 90 3150 174
rect 3180 149 3237 174
rect 3180 115 3191 149
rect 3225 115 3237 149
rect 3180 90 3237 115
rect 2739 47 2796 63
rect 1820 39 1832 47
rect 1774 27 1832 39
<< pdiff >>
rect 116 597 173 619
rect 116 563 128 597
rect 162 563 173 597
rect 116 465 173 563
rect 116 431 128 465
rect 162 431 173 465
rect 116 419 173 431
rect 223 419 271 619
rect 321 594 389 619
rect 321 560 332 594
rect 366 560 389 594
rect 321 419 389 560
rect 439 419 493 619
rect 543 597 599 619
rect 543 563 554 597
rect 588 563 599 597
rect 543 512 599 563
rect 543 478 554 512
rect 588 478 599 512
rect 543 419 599 478
rect 649 606 722 619
rect 649 572 660 606
rect 694 572 722 606
rect 649 419 722 572
rect 772 465 829 619
rect 772 431 783 465
rect 817 431 829 465
rect 772 419 829 431
rect 888 527 945 608
rect 888 493 900 527
rect 934 493 945 527
rect 888 454 945 493
rect 888 420 900 454
rect 934 420 945 454
rect 888 408 945 420
rect 995 596 1097 608
rect 995 562 1052 596
rect 1086 562 1097 596
rect 995 408 1097 562
rect 1147 456 1200 608
rect 1147 422 1158 456
rect 1192 422 1200 456
rect 1147 408 1200 422
rect 1365 535 1447 547
rect 1365 501 1373 535
rect 1407 501 1447 535
rect 1365 434 1447 501
rect 1365 400 1373 434
rect 1407 400 1447 434
rect 1365 388 1447 400
rect 1385 347 1447 388
rect 1497 535 1583 547
rect 1497 501 1508 535
rect 1542 501 1583 535
rect 1497 464 1583 501
rect 1497 430 1508 464
rect 1542 430 1583 464
rect 1497 393 1583 430
rect 1497 359 1508 393
rect 1542 359 1583 393
rect 1497 347 1583 359
rect 1633 347 1675 547
rect 1725 523 1781 547
rect 1725 489 1736 523
rect 1770 489 1781 523
rect 1725 347 1781 489
rect 1831 535 1917 547
rect 2264 597 2337 619
rect 2264 563 2276 597
rect 2310 563 2337 597
rect 2264 541 2337 563
rect 1831 501 1871 535
rect 1905 501 1917 535
rect 1831 464 1917 501
rect 1831 430 1871 464
rect 1905 430 1917 464
rect 1831 393 1917 430
rect 1831 359 1871 393
rect 1905 359 1917 393
rect 1831 347 1917 359
rect 2020 529 2077 541
rect 2020 495 2032 529
rect 2066 495 2077 529
rect 2020 458 2077 495
rect 2020 424 2032 458
rect 2066 424 2077 458
rect 2020 387 2077 424
rect 2020 353 2032 387
rect 2066 353 2077 387
rect 2020 341 2077 353
rect 2127 529 2199 541
rect 2127 495 2154 529
rect 2188 495 2199 529
rect 2127 458 2199 495
rect 2127 424 2154 458
rect 2188 424 2199 458
rect 2127 387 2199 424
rect 2127 353 2154 387
rect 2188 353 2199 387
rect 2127 341 2199 353
rect 2249 527 2337 541
rect 2249 493 2276 527
rect 2310 493 2337 527
rect 2249 457 2337 493
rect 2249 423 2276 457
rect 2310 423 2337 457
rect 2249 419 2337 423
rect 2387 419 2435 619
rect 2485 607 2654 619
rect 2485 573 2496 607
rect 2530 573 2654 607
rect 2485 536 2654 573
rect 2485 502 2496 536
rect 2530 502 2654 536
rect 2485 465 2654 502
rect 2485 431 2496 465
rect 2530 431 2654 465
rect 2485 419 2654 431
rect 2704 597 2760 619
rect 2704 563 2715 597
rect 2749 563 2760 597
rect 2704 473 2760 563
rect 2704 439 2715 473
rect 2749 439 2760 473
rect 2704 419 2760 439
rect 2810 607 2867 619
rect 2810 573 2821 607
rect 2855 573 2867 607
rect 2810 536 2867 573
rect 2810 502 2821 536
rect 2855 502 2867 536
rect 2810 465 2867 502
rect 2810 431 2821 465
rect 2855 431 2867 465
rect 2810 419 2867 431
rect 2921 576 2978 588
rect 2921 542 2933 576
rect 2967 542 2978 576
rect 2921 505 2978 542
rect 2921 471 2933 505
rect 2967 471 2978 505
rect 2921 434 2978 471
rect 2249 387 2322 419
rect 2249 353 2276 387
rect 2310 353 2322 387
rect 2249 341 2322 353
rect 2921 400 2933 434
rect 2967 400 2978 434
rect 2921 388 2978 400
rect 3028 576 3084 588
rect 3028 542 3039 576
rect 3073 542 3084 576
rect 3028 505 3084 542
rect 3028 471 3039 505
rect 3073 471 3084 505
rect 3028 434 3084 471
rect 3028 400 3039 434
rect 3073 400 3084 434
rect 3028 388 3084 400
rect 3134 576 3191 588
rect 3134 542 3145 576
rect 3179 542 3191 576
rect 3134 505 3191 542
rect 3134 471 3145 505
rect 3179 471 3191 505
rect 3134 434 3191 471
rect 3134 400 3145 434
rect 3179 400 3191 434
rect 3134 388 3191 400
<< ndiffc >>
rect 246 139 280 173
rect 426 113 460 147
rect 528 113 562 147
rect 780 135 814 169
rect 884 144 918 178
rect 1058 107 1092 141
rect 1232 141 1266 175
rect 1357 141 1391 175
rect 1443 141 1477 175
rect 50 53 84 87
rect 1786 39 1820 73
rect 2017 55 2051 89
rect 2318 77 2352 111
rect 2543 63 2577 97
rect 2750 63 2784 97
rect 2875 115 2909 149
rect 3033 115 3067 149
rect 3191 115 3225 149
<< pdiffc >>
rect 128 563 162 597
rect 128 431 162 465
rect 332 560 366 594
rect 554 563 588 597
rect 554 478 588 512
rect 660 572 694 606
rect 783 431 817 465
rect 900 493 934 527
rect 900 420 934 454
rect 1052 562 1086 596
rect 1158 422 1192 456
rect 1373 501 1407 535
rect 1373 400 1407 434
rect 1508 501 1542 535
rect 1508 430 1542 464
rect 1508 359 1542 393
rect 1736 489 1770 523
rect 2276 563 2310 597
rect 1871 501 1905 535
rect 1871 430 1905 464
rect 1871 359 1905 393
rect 2032 495 2066 529
rect 2032 424 2066 458
rect 2032 353 2066 387
rect 2154 495 2188 529
rect 2154 424 2188 458
rect 2154 353 2188 387
rect 2276 493 2310 527
rect 2276 423 2310 457
rect 2496 573 2530 607
rect 2496 502 2530 536
rect 2496 431 2530 465
rect 2715 563 2749 597
rect 2715 439 2749 473
rect 2821 573 2855 607
rect 2821 502 2855 536
rect 2821 431 2855 465
rect 2933 542 2967 576
rect 2933 471 2967 505
rect 2276 353 2310 387
rect 2933 400 2967 434
rect 3039 542 3073 576
rect 3039 471 3073 505
rect 3039 400 3073 434
rect 3145 542 3179 576
rect 3145 471 3179 505
rect 3145 400 3179 434
<< poly >>
rect 173 619 223 645
rect 271 619 321 645
rect 389 619 439 645
rect 493 619 543 645
rect 599 619 649 645
rect 722 619 772 645
rect 945 608 995 634
rect 1097 608 1147 634
rect 1215 615 2249 645
rect 2337 619 2387 645
rect 2435 619 2485 645
rect 2654 619 2704 645
rect 2760 619 2810 645
rect 173 380 223 419
rect 271 404 321 419
rect 173 368 203 380
rect 115 352 203 368
rect 115 318 131 352
rect 165 332 203 352
rect 271 371 337 404
rect 271 337 287 371
rect 321 337 337 371
rect 389 356 439 419
rect 493 356 543 419
rect 599 356 649 419
rect 722 377 772 419
rect 709 361 775 377
rect 165 318 219 332
rect 271 321 337 337
rect 115 302 219 318
rect 81 244 147 260
rect 81 210 97 244
rect 131 210 147 244
rect 81 194 147 210
rect 111 172 141 194
rect 189 172 219 302
rect 307 172 337 321
rect 379 340 445 356
rect 379 306 395 340
rect 429 306 445 340
rect 379 290 445 306
rect 487 340 553 356
rect 487 306 503 340
rect 537 306 553 340
rect 487 290 553 306
rect 595 340 661 356
rect 595 306 611 340
rect 645 306 661 340
rect 595 290 661 306
rect 709 327 725 361
rect 759 327 775 361
rect 709 311 775 327
rect 385 172 415 290
rect 595 248 625 290
rect 709 248 739 311
rect 945 300 995 408
rect 1097 370 1147 408
rect 1215 370 1245 615
rect 1447 547 1497 573
rect 1583 547 1633 615
rect 1675 547 1725 573
rect 1781 547 1831 573
rect 1095 354 1245 370
rect 1095 320 1111 354
rect 1145 320 1245 354
rect 945 284 1031 300
rect 945 264 981 284
rect 929 250 981 264
rect 1015 250 1031 284
rect 471 218 625 248
rect 667 218 769 248
rect 471 172 501 218
rect 667 203 697 218
rect 739 203 769 218
rect 929 234 1031 250
rect 1095 286 1245 320
rect 1287 340 1353 356
rect 2077 541 2127 567
rect 2199 541 2249 615
rect 1287 306 1303 340
rect 1337 332 1353 340
rect 1447 332 1497 347
rect 1337 306 1541 332
rect 1583 321 1633 347
rect 1675 321 1725 347
rect 1287 291 1541 306
rect 1675 291 1721 321
rect 1781 315 1831 347
rect 2978 588 3028 614
rect 3084 588 3134 614
rect 2337 374 2387 419
rect 2077 315 2127 341
rect 1770 311 1832 315
rect 1287 290 1553 291
rect 1095 252 1111 286
rect 1145 252 1245 286
rect 1095 248 1245 252
rect 1474 289 1553 290
rect 1663 289 1721 291
rect 1474 288 1555 289
rect 1661 288 1721 289
rect 1474 287 1556 288
rect 1660 287 1721 288
rect 1474 286 1557 287
rect 1659 286 1721 287
rect 1474 285 1558 286
rect 1658 285 1721 286
rect 1474 283 1559 285
rect 1657 283 1721 285
rect 1474 275 1561 283
rect 1655 279 1721 283
rect 1095 236 1432 248
rect 929 203 959 234
rect 1001 203 1031 234
rect 1119 203 1149 236
rect 1191 218 1432 236
rect 1474 241 1511 275
rect 1545 241 1561 275
rect 1474 225 1561 241
rect 1191 203 1221 218
rect 1402 203 1432 218
rect 1531 203 1561 225
rect 1605 275 1721 279
rect 1605 241 1671 275
rect 1705 241 1721 275
rect 1605 229 1721 241
rect 1766 299 1832 311
rect 1766 265 1782 299
rect 1816 265 1832 299
rect 1766 241 1832 265
rect 1874 299 2127 315
rect 1874 265 1890 299
rect 1924 285 2127 299
rect 2199 290 2249 341
rect 2357 326 2387 374
rect 1924 265 1978 285
rect 1605 227 1716 229
rect 1605 226 1713 227
rect 1605 225 1711 226
rect 1605 203 1635 225
rect 667 93 697 119
rect 739 93 769 119
rect 929 93 959 119
rect 1001 93 1031 119
rect 1766 195 1828 241
rect 1748 193 1828 195
rect 1744 191 1828 193
rect 1741 189 1828 191
rect 1737 187 1828 189
rect 1729 165 1828 187
rect 1874 185 1978 265
rect 2183 274 2249 290
rect 2183 240 2199 274
rect 2233 240 2249 274
rect 2183 224 2249 240
rect 2291 296 2387 326
rect 2435 326 2485 419
rect 2654 387 2704 419
rect 2631 371 2704 387
rect 2631 337 2647 371
rect 2681 337 2704 371
rect 2435 296 2507 326
rect 1729 150 1759 165
rect 1119 93 1149 119
rect 1191 93 1221 119
rect 1402 93 1432 119
rect 1531 93 1561 119
rect 1605 93 1635 119
rect 111 62 141 88
rect 189 62 219 88
rect 307 62 337 88
rect 385 62 415 88
rect 471 51 501 88
rect 1870 146 1978 185
rect 2026 203 2092 219
rect 2026 169 2042 203
rect 2076 176 2092 203
rect 2291 176 2321 296
rect 2477 274 2507 296
rect 2631 321 2704 337
rect 2477 258 2589 274
rect 2363 232 2429 248
rect 2363 198 2379 232
rect 2413 198 2429 232
rect 2363 182 2429 198
rect 2477 224 2539 258
rect 2573 224 2589 258
rect 2477 208 2589 224
rect 2076 169 2321 176
rect 2026 146 2321 169
rect 1870 131 1900 146
rect 1948 131 1978 146
rect 2062 131 2092 146
rect 2369 131 2399 182
rect 2477 131 2507 208
rect 2631 131 2661 321
rect 2760 219 2810 419
rect 2978 219 3028 388
rect 3084 348 3134 388
rect 2703 216 3028 219
rect 3070 332 3136 348
rect 3070 298 3086 332
rect 3120 298 3136 332
rect 3070 264 3136 298
rect 3070 230 3086 264
rect 3120 244 3136 264
rect 3120 230 3180 244
rect 2703 203 3022 216
rect 3070 214 3180 230
rect 2703 169 2719 203
rect 2753 189 3022 203
rect 2753 169 2790 189
rect 2920 174 2950 189
rect 2992 174 3022 189
rect 3078 174 3108 214
rect 3150 174 3180 214
rect 2703 153 2790 169
rect 2709 131 2739 153
rect 1729 51 1759 66
rect 471 21 1759 51
rect 2920 64 2950 90
rect 2992 64 3022 90
rect 3078 64 3108 90
rect 3150 64 3180 90
rect 1870 21 1900 47
rect 1948 21 1978 47
rect 2062 21 2092 47
rect 2369 21 2399 47
rect 2477 21 2507 47
rect 2631 21 2661 47
rect 2709 21 2739 47
<< polycont >>
rect 131 318 165 352
rect 287 337 321 371
rect 97 210 131 244
rect 395 306 429 340
rect 503 306 537 340
rect 611 306 645 340
rect 725 327 759 361
rect 1111 320 1145 354
rect 981 250 1015 284
rect 1303 306 1337 340
rect 1111 252 1145 286
rect 1511 241 1545 275
rect 1671 241 1705 275
rect 1782 265 1816 299
rect 1890 265 1924 299
rect 2199 240 2233 274
rect 2647 337 2681 371
rect 2042 169 2076 203
rect 2379 198 2413 232
rect 2539 224 2573 258
rect 3086 298 3120 332
rect 3086 230 3120 264
rect 2719 169 2753 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 18 597 178 613
rect 18 563 128 597
rect 162 563 178 597
rect 18 496 178 563
rect 316 594 382 649
rect 316 560 332 594
rect 366 560 382 594
rect 316 532 382 560
rect 538 597 604 613
rect 538 563 554 597
rect 588 563 604 597
rect 644 606 710 649
rect 644 572 660 606
rect 694 572 710 606
rect 644 571 710 572
rect 746 579 1002 613
rect 538 535 604 563
rect 746 535 780 579
rect 538 512 780 535
rect 538 496 554 512
rect 18 478 554 496
rect 588 501 780 512
rect 884 527 934 543
rect 588 478 604 501
rect 18 465 604 478
rect 884 493 900 527
rect 18 431 128 465
rect 162 462 604 465
rect 162 431 178 462
rect 18 415 178 431
rect 767 431 783 465
rect 817 431 845 465
rect 18 158 52 415
rect 217 392 731 426
rect 767 415 845 431
rect 217 371 337 392
rect 115 352 181 368
rect 115 318 131 352
rect 165 318 181 352
rect 115 302 181 318
rect 217 337 287 371
rect 321 337 337 371
rect 697 377 731 392
rect 697 361 775 377
rect 217 310 337 337
rect 379 340 451 356
rect 379 306 395 340
rect 429 306 451 340
rect 379 290 451 306
rect 487 340 553 356
rect 487 306 503 340
rect 537 306 553 340
rect 88 254 147 260
rect 487 254 553 306
rect 595 350 661 356
rect 595 316 607 350
rect 641 340 661 350
rect 595 306 611 316
rect 645 306 661 340
rect 697 327 725 361
rect 759 327 775 361
rect 697 311 775 327
rect 595 290 661 306
rect 811 254 845 415
rect 88 244 845 254
rect 88 210 97 244
rect 131 220 845 244
rect 131 210 147 220
rect 88 194 147 210
rect 230 158 246 173
rect 18 139 246 158
rect 280 139 296 173
rect 18 124 296 139
rect 230 123 296 124
rect 410 147 476 176
rect 410 113 426 147
rect 460 113 476 147
rect 34 87 100 88
rect 410 87 476 113
rect 34 53 50 87
rect 84 53 476 87
rect 512 147 578 176
rect 512 113 528 147
rect 562 113 578 147
rect 764 169 845 220
rect 764 135 780 169
rect 814 135 845 169
rect 764 119 845 135
rect 884 454 934 493
rect 968 526 1002 579
rect 1036 596 1102 649
rect 1036 562 1052 596
rect 1086 562 1102 596
rect 1373 535 1407 551
rect 968 501 1373 526
rect 968 492 1407 501
rect 884 420 900 454
rect 884 370 934 420
rect 1142 422 1158 456
rect 1192 422 1258 456
rect 1142 406 1258 422
rect 884 354 1161 370
rect 884 336 1111 354
rect 884 178 918 336
rect 1095 320 1111 336
rect 1145 320 1161 354
rect 965 284 1031 300
rect 965 250 981 284
rect 1015 250 1031 284
rect 965 234 1031 250
rect 1095 286 1161 320
rect 1195 356 1258 406
rect 1373 434 1407 492
rect 1195 340 1337 356
rect 1195 306 1303 340
rect 1195 290 1337 306
rect 1095 252 1111 286
rect 1145 252 1161 286
rect 1095 236 1161 252
rect 1214 175 1291 290
rect 1373 229 1407 400
rect 884 127 918 144
rect 1042 141 1108 145
rect 512 17 578 113
rect 1042 107 1058 141
rect 1092 107 1108 141
rect 1214 141 1232 175
rect 1266 141 1291 175
rect 1214 119 1291 141
rect 1341 175 1407 229
rect 1341 141 1357 175
rect 1391 141 1407 175
rect 1341 119 1407 141
rect 1443 535 1558 551
rect 1443 501 1508 535
rect 1542 501 1558 535
rect 1443 464 1558 501
rect 1443 430 1508 464
rect 1542 430 1558 464
rect 1717 523 1783 649
rect 1717 489 1736 523
rect 1770 489 1783 523
rect 1717 462 1783 489
rect 1855 535 1940 551
rect 1855 501 1871 535
rect 1905 501 1940 535
rect 1855 464 1940 501
rect 1443 426 1558 430
rect 1855 430 1871 464
rect 1905 430 1940 464
rect 1855 426 1940 430
rect 1443 393 1940 426
rect 1443 359 1508 393
rect 1542 392 1871 393
rect 1542 359 1558 392
rect 1443 358 1558 359
rect 1905 359 1940 393
rect 1443 175 1477 358
rect 1753 350 1837 356
rect 1753 316 1759 350
rect 1793 329 1837 350
rect 1871 343 1940 359
rect 1793 316 1840 329
rect 1443 125 1477 141
rect 1511 275 1545 305
rect 1511 159 1545 241
rect 1645 275 1711 305
rect 1645 241 1671 275
rect 1705 241 1711 275
rect 1753 299 1840 316
rect 1753 265 1782 299
rect 1816 265 1840 299
rect 1874 299 1940 343
rect 2016 529 2082 649
rect 2260 597 2326 613
rect 2260 563 2276 597
rect 2310 563 2326 597
rect 2016 495 2032 529
rect 2066 495 2082 529
rect 2016 458 2082 495
rect 2016 424 2032 458
rect 2066 424 2082 458
rect 2016 387 2082 424
rect 2016 353 2032 387
rect 2066 353 2082 387
rect 2016 337 2082 353
rect 2121 529 2204 545
rect 2121 495 2154 529
rect 2188 495 2204 529
rect 2121 458 2204 495
rect 2121 424 2154 458
rect 2188 424 2204 458
rect 2121 387 2204 424
rect 2121 353 2154 387
rect 2188 353 2204 387
rect 2121 337 2204 353
rect 2260 527 2326 563
rect 2260 493 2276 527
rect 2310 493 2326 527
rect 2260 457 2326 493
rect 2260 423 2276 457
rect 2310 423 2326 457
rect 2260 387 2326 423
rect 2480 607 2530 649
rect 2480 573 2496 607
rect 2699 597 2767 613
rect 2480 536 2530 573
rect 2480 502 2496 536
rect 2480 465 2530 502
rect 2480 431 2496 465
rect 2480 415 2530 431
rect 2260 353 2276 387
rect 2310 371 2326 387
rect 2617 387 2663 578
rect 2699 563 2715 597
rect 2749 563 2767 597
rect 2699 473 2767 563
rect 2699 439 2715 473
rect 2749 439 2767 473
rect 2699 423 2767 439
rect 2617 371 2697 387
rect 2310 353 2491 371
rect 2617 357 2647 371
rect 2260 337 2491 353
rect 1874 265 1890 299
rect 1924 265 1940 299
rect 2121 289 2155 337
rect 1645 229 1711 241
rect 1974 255 2155 289
rect 1974 229 2008 255
rect 1645 195 2008 229
rect 2042 203 2085 219
rect 2076 169 2085 203
rect 2042 159 2085 169
rect 1511 125 2085 159
rect 1042 17 1108 107
rect 2121 89 2155 255
rect 2191 274 2421 290
rect 2191 240 2199 274
rect 2233 240 2421 274
rect 2191 232 2421 240
rect 2191 224 2379 232
rect 2363 198 2379 224
rect 2413 198 2421 232
rect 2363 182 2421 198
rect 2457 172 2491 337
rect 2527 350 2647 357
rect 2561 337 2647 350
rect 2681 337 2697 371
rect 2561 323 2697 337
rect 2561 316 2567 323
rect 2527 310 2567 316
rect 2733 287 2767 423
rect 2805 607 2871 649
rect 2805 573 2821 607
rect 2855 573 2871 607
rect 2805 536 2871 573
rect 2805 502 2821 536
rect 2855 502 2871 536
rect 2805 465 2871 502
rect 2805 431 2821 465
rect 2855 431 2871 465
rect 2805 415 2871 431
rect 2907 576 2983 592
rect 2907 542 2933 576
rect 2967 542 2983 576
rect 2907 505 2983 542
rect 2907 471 2933 505
rect 2967 471 2983 505
rect 2907 434 2983 471
rect 2907 400 2933 434
rect 2967 400 2983 434
rect 2907 348 2983 400
rect 3023 576 3089 649
rect 3023 542 3039 576
rect 3073 542 3089 576
rect 3023 505 3089 542
rect 3023 471 3039 505
rect 3073 471 3089 505
rect 3023 434 3089 471
rect 3023 400 3039 434
rect 3073 400 3089 434
rect 3023 384 3089 400
rect 3129 576 3241 592
rect 3129 542 3145 576
rect 3179 542 3241 576
rect 3129 505 3241 542
rect 3129 471 3145 505
rect 3179 471 3241 505
rect 3129 434 3241 471
rect 3129 400 3145 434
rect 3179 400 3241 434
rect 3129 384 3241 400
rect 2907 332 3136 348
rect 2907 314 3086 332
rect 2603 274 2839 287
rect 2527 258 2839 274
rect 2527 224 2539 258
rect 2573 253 2839 258
rect 2573 224 2637 253
rect 2527 208 2637 224
rect 2703 203 2769 217
rect 2703 172 2719 203
rect 2457 169 2719 172
rect 2753 169 2769 203
rect 2457 138 2769 169
rect 2457 135 2491 138
rect 1770 73 1836 89
rect 1770 39 1786 73
rect 1820 39 1836 73
rect 2001 55 2017 89
rect 2051 55 2155 89
rect 2302 111 2491 135
rect 2302 77 2318 111
rect 2352 101 2491 111
rect 2805 102 2839 253
rect 2907 178 2941 314
rect 3070 298 3086 314
rect 3120 298 3136 332
rect 3070 264 3136 298
rect 3070 230 3086 264
rect 3120 230 3136 264
rect 3070 214 3136 230
rect 2352 77 2368 101
rect 2302 53 2368 77
rect 2527 97 2593 102
rect 2527 63 2543 97
rect 2577 63 2593 97
rect 1770 17 1836 39
rect 2527 17 2593 63
rect 2734 97 2839 102
rect 2734 63 2750 97
rect 2784 63 2839 97
rect 2875 149 2941 178
rect 2909 115 2941 149
rect 2875 86 2941 115
rect 3017 149 3083 178
rect 3017 115 3033 149
rect 3067 115 3083 149
rect 2734 59 2839 63
rect 3017 17 3083 115
rect 3175 149 3241 384
rect 3175 115 3191 149
rect 3225 115 3241 149
rect 3175 86 3241 115
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 607 340 641 350
rect 607 316 611 340
rect 611 316 641 340
rect 1759 316 1793 350
rect 2527 316 2561 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
<< metal1 >>
rect 0 683 3264 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3264 683
rect 0 617 3264 649
rect 595 350 653 356
rect 595 316 607 350
rect 641 347 653 350
rect 1747 350 1805 356
rect 1747 347 1759 350
rect 641 319 1759 347
rect 641 316 653 319
rect 595 310 653 316
rect 1747 316 1759 319
rect 1793 347 1805 350
rect 2515 350 2573 356
rect 2515 347 2527 350
rect 1793 319 2527 347
rect 1793 316 1805 319
rect 1747 310 1805 316
rect 2515 316 2527 319
rect 2561 316 2573 350
rect 2515 310 2573 316
rect 0 17 3264 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3264 17
rect 0 -49 3264 -17
<< labels >>
flabel pwell s 0 0 3264 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 3264 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfrtp_lp2
flabel comment s 1111 36 1111 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1739 630 1739 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1181 289 1181 289 0 FreeSans 200 180 0 0 no_jumper_check
flabel comment s 1363 310 1363 310 0 FreeSans 200 180 0 0 no_jumper_check
flabel metal1 s 2527 316 2561 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 3264 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 3264 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 3199 94 3233 128 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3199 168 3233 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3199 242 3233 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3199 316 3233 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3199 390 3233 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3199 464 3233 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3199 538 3233 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3264 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry R90
string GDS_END 3310868
string GDS_START 3289480
<< end >>
