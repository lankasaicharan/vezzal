magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 228 241 836 243
rect 1 49 836 241
rect 0 0 864 49
<< scnmos >>
rect 80 47 110 215
rect 307 49 337 217
rect 379 49 409 217
rect 487 49 517 217
rect 641 49 671 217
rect 727 49 757 217
<< scpmoshvt >>
rect 80 367 110 619
rect 293 367 323 619
rect 379 367 409 619
rect 547 367 577 619
rect 655 367 685 619
rect 727 367 757 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 101 80 169
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 187 163 215
rect 110 153 121 187
rect 155 153 163 187
rect 110 93 163 153
rect 110 59 121 93
rect 155 59 163 93
rect 110 47 163 59
rect 254 205 307 217
rect 254 171 262 205
rect 296 171 307 205
rect 254 101 307 171
rect 254 67 262 101
rect 296 67 307 101
rect 254 49 307 67
rect 337 49 379 217
rect 409 49 487 217
rect 517 205 641 217
rect 517 171 528 205
rect 562 171 596 205
rect 630 171 641 205
rect 517 101 641 171
rect 517 67 528 101
rect 562 67 596 101
rect 630 67 641 101
rect 517 49 641 67
rect 671 165 727 217
rect 671 131 682 165
rect 716 131 727 165
rect 671 91 727 131
rect 671 57 682 91
rect 716 57 727 91
rect 671 49 727 57
rect 757 205 810 217
rect 757 171 768 205
rect 802 171 810 205
rect 757 101 810 171
rect 757 67 768 101
rect 802 67 810 101
rect 757 49 810 67
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 506 80 565
rect 27 472 35 506
rect 69 472 80 506
rect 27 413 80 472
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 607 293 619
rect 110 573 121 607
rect 155 573 248 607
rect 282 573 293 607
rect 110 548 293 573
rect 110 514 185 548
rect 219 514 293 548
rect 110 488 293 514
rect 110 454 121 488
rect 155 454 248 488
rect 282 454 293 488
rect 110 413 293 454
rect 110 379 121 413
rect 155 379 293 413
rect 110 367 293 379
rect 323 599 379 619
rect 323 565 334 599
rect 368 565 379 599
rect 323 511 379 565
rect 323 477 334 511
rect 368 477 379 511
rect 323 420 379 477
rect 323 386 334 420
rect 368 386 379 420
rect 323 367 379 386
rect 409 607 547 619
rect 409 573 420 607
rect 454 573 502 607
rect 536 573 547 607
rect 409 493 547 573
rect 409 459 420 493
rect 454 459 502 493
rect 536 459 547 493
rect 409 367 547 459
rect 577 607 655 619
rect 577 573 602 607
rect 636 573 655 607
rect 577 517 655 573
rect 577 483 602 517
rect 636 483 655 517
rect 577 420 655 483
rect 577 386 602 420
rect 636 386 655 420
rect 577 367 655 386
rect 685 367 727 619
rect 757 607 810 619
rect 757 573 768 607
rect 802 573 810 607
rect 757 517 810 573
rect 757 483 768 517
rect 802 483 810 517
rect 757 420 810 483
rect 757 386 768 420
rect 802 386 810 420
rect 757 367 810 386
<< ndiffc >>
rect 35 169 69 203
rect 35 67 69 101
rect 121 153 155 187
rect 121 59 155 93
rect 262 171 296 205
rect 262 67 296 101
rect 528 171 562 205
rect 596 171 630 205
rect 528 67 562 101
rect 596 67 630 101
rect 682 131 716 165
rect 682 57 716 91
rect 768 171 802 205
rect 768 67 802 101
<< pdiffc >>
rect 35 565 69 599
rect 35 472 69 506
rect 35 379 69 413
rect 121 573 155 607
rect 248 573 282 607
rect 185 514 219 548
rect 121 454 155 488
rect 248 454 282 488
rect 121 379 155 413
rect 334 565 368 599
rect 334 477 368 511
rect 334 386 368 420
rect 420 573 454 607
rect 502 573 536 607
rect 420 459 454 493
rect 502 459 536 493
rect 602 573 636 607
rect 602 483 636 517
rect 602 386 636 420
rect 768 573 802 607
rect 768 483 802 517
rect 768 386 802 420
<< poly >>
rect 80 619 110 645
rect 293 619 323 645
rect 379 619 409 645
rect 547 619 577 645
rect 655 619 685 645
rect 727 619 757 645
rect 80 303 110 367
rect 293 335 323 367
rect 265 319 337 335
rect 80 287 159 303
rect 80 253 109 287
rect 143 253 159 287
rect 265 285 281 319
rect 315 285 337 319
rect 265 269 337 285
rect 80 237 159 253
rect 80 215 110 237
rect 307 217 337 269
rect 379 305 409 367
rect 547 335 577 367
rect 655 335 685 367
rect 487 319 577 335
rect 379 289 445 305
rect 379 255 395 289
rect 429 255 445 289
rect 379 239 445 255
rect 487 285 511 319
rect 545 285 577 319
rect 487 269 577 285
rect 619 319 685 335
rect 619 285 635 319
rect 669 285 685 319
rect 619 269 685 285
rect 727 325 757 367
rect 727 309 839 325
rect 727 275 789 309
rect 823 275 839 309
rect 379 217 409 239
rect 487 217 517 269
rect 641 217 671 269
rect 727 259 839 275
rect 727 217 757 259
rect 80 21 110 47
rect 307 23 337 49
rect 379 23 409 49
rect 487 23 517 49
rect 641 23 671 49
rect 727 23 757 49
<< polycont >>
rect 109 253 143 287
rect 281 285 315 319
rect 395 255 429 289
rect 511 285 545 319
rect 635 285 669 319
rect 789 275 823 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 19 599 73 615
rect 19 565 35 599
rect 69 565 73 599
rect 19 506 73 565
rect 19 472 35 506
rect 69 472 73 506
rect 19 413 73 472
rect 19 379 35 413
rect 69 379 73 413
rect 19 203 73 379
rect 107 607 298 649
rect 107 573 121 607
rect 155 573 248 607
rect 282 573 298 607
rect 107 548 298 573
rect 107 514 185 548
rect 219 514 298 548
rect 107 488 298 514
rect 107 454 121 488
rect 155 454 248 488
rect 282 454 298 488
rect 332 599 370 615
rect 332 565 334 599
rect 368 565 370 599
rect 332 511 370 565
rect 332 477 334 511
rect 368 477 370 511
rect 107 413 161 454
rect 332 420 370 477
rect 404 607 552 649
rect 404 573 420 607
rect 454 573 502 607
rect 536 573 552 607
rect 404 493 552 573
rect 404 459 420 493
rect 454 459 502 493
rect 536 459 552 493
rect 404 454 552 459
rect 586 607 652 615
rect 586 573 602 607
rect 636 573 652 607
rect 586 517 652 573
rect 586 483 602 517
rect 636 483 652 517
rect 586 420 652 483
rect 107 379 121 413
rect 155 379 161 413
rect 107 363 161 379
rect 195 386 334 420
rect 368 386 602 420
rect 636 386 652 420
rect 746 607 818 649
rect 746 573 768 607
rect 802 573 818 607
rect 746 517 818 573
rect 746 483 768 517
rect 802 483 818 517
rect 746 420 818 483
rect 746 386 768 420
rect 802 386 818 420
rect 195 303 229 386
rect 107 287 229 303
rect 107 253 109 287
rect 143 253 229 287
rect 265 319 361 352
rect 265 285 281 319
rect 315 285 361 319
rect 265 283 361 285
rect 395 289 461 352
rect 107 249 229 253
rect 429 255 461 289
rect 495 319 560 352
rect 495 285 511 319
rect 545 285 560 319
rect 495 269 560 285
rect 594 319 739 352
rect 594 285 635 319
rect 669 285 739 319
rect 594 267 739 285
rect 773 309 847 352
rect 773 275 789 309
rect 823 275 847 309
rect 773 267 847 275
rect 107 237 312 249
rect 195 215 312 237
rect 246 205 312 215
rect 19 169 35 203
rect 69 169 73 203
rect 19 101 73 169
rect 19 67 35 101
rect 69 67 73 101
rect 19 51 73 67
rect 107 187 161 203
rect 107 153 121 187
rect 155 181 161 187
rect 155 153 171 181
rect 107 93 171 153
rect 107 59 121 93
rect 155 59 171 93
rect 107 17 171 59
rect 246 171 262 205
rect 296 171 312 205
rect 246 101 312 171
rect 246 67 262 101
rect 296 67 312 101
rect 395 78 461 255
rect 512 205 818 233
rect 512 171 528 205
rect 562 171 596 205
rect 630 199 768 205
rect 630 171 632 199
rect 512 101 632 171
rect 766 171 768 199
rect 802 171 818 205
rect 246 51 312 67
rect 512 67 528 101
rect 562 67 596 101
rect 630 67 632 101
rect 512 51 632 67
rect 666 131 682 165
rect 716 131 732 165
rect 666 91 732 131
rect 666 57 682 91
rect 716 57 732 91
rect 666 17 732 57
rect 766 101 818 171
rect 766 67 768 101
rect 802 67 818 101
rect 766 51 818 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2111a_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4249668
string GDS_START 4240726
<< end >>
