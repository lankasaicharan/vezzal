magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 23 49 1012 243
rect 0 0 1056 49
<< scnmos >>
rect 106 133 136 217
rect 242 49 272 217
rect 328 49 358 217
rect 414 49 444 217
rect 500 49 530 217
rect 615 49 645 217
rect 687 49 717 217
rect 795 49 825 217
rect 903 49 933 217
<< scpmoshvt >>
rect 106 367 136 451
rect 242 367 272 619
rect 328 367 358 619
rect 414 367 444 619
rect 500 367 530 619
rect 601 367 631 619
rect 687 367 717 619
rect 817 367 847 619
rect 903 367 933 619
<< ndiff >>
rect 49 191 106 217
rect 49 157 57 191
rect 91 157 106 191
rect 49 133 106 157
rect 136 163 242 217
rect 136 133 197 163
rect 189 129 197 133
rect 231 129 242 163
rect 189 95 242 129
rect 189 61 197 95
rect 231 61 242 95
rect 189 49 242 61
rect 272 205 328 217
rect 272 171 283 205
rect 317 171 328 205
rect 272 101 328 171
rect 272 67 283 101
rect 317 67 328 101
rect 272 49 328 67
rect 358 181 414 217
rect 358 147 369 181
rect 403 147 414 181
rect 358 95 414 147
rect 358 61 369 95
rect 403 61 414 95
rect 358 49 414 61
rect 444 205 500 217
rect 444 171 455 205
rect 489 171 500 205
rect 444 101 500 171
rect 444 67 455 101
rect 489 67 500 101
rect 444 49 500 67
rect 530 165 615 217
rect 530 131 556 165
rect 590 131 615 165
rect 530 91 615 131
rect 530 57 556 91
rect 590 57 615 91
rect 530 49 615 57
rect 645 49 687 217
rect 717 49 795 217
rect 825 49 903 217
rect 933 205 986 217
rect 933 171 944 205
rect 978 171 986 205
rect 933 101 986 171
rect 933 67 944 101
rect 978 67 986 101
rect 933 49 986 67
<< pdiff >>
rect 189 597 242 619
rect 189 563 197 597
rect 231 563 242 597
rect 189 451 242 563
rect 49 425 106 451
rect 49 391 57 425
rect 91 391 106 425
rect 49 367 106 391
rect 136 367 242 451
rect 272 436 328 619
rect 272 402 283 436
rect 317 402 328 436
rect 272 367 328 402
rect 358 597 414 619
rect 358 563 369 597
rect 403 563 414 597
rect 358 367 414 563
rect 444 436 500 619
rect 444 402 455 436
rect 489 402 500 436
rect 444 367 500 402
rect 530 597 601 619
rect 530 563 541 597
rect 575 563 601 597
rect 530 367 601 563
rect 631 436 687 619
rect 631 402 642 436
rect 676 402 687 436
rect 631 367 687 402
rect 717 597 817 619
rect 717 563 728 597
rect 762 563 817 597
rect 717 367 817 563
rect 847 436 903 619
rect 847 402 858 436
rect 892 402 903 436
rect 847 367 903 402
rect 933 597 986 619
rect 933 563 944 597
rect 978 563 986 597
rect 933 367 986 563
<< ndiffc >>
rect 57 157 91 191
rect 197 129 231 163
rect 197 61 231 95
rect 283 171 317 205
rect 283 67 317 101
rect 369 147 403 181
rect 369 61 403 95
rect 455 171 489 205
rect 455 67 489 101
rect 556 131 590 165
rect 556 57 590 91
rect 944 171 978 205
rect 944 67 978 101
<< pdiffc >>
rect 197 563 231 597
rect 57 391 91 425
rect 283 402 317 436
rect 369 563 403 597
rect 455 402 489 436
rect 541 563 575 597
rect 642 402 676 436
rect 728 563 762 597
rect 858 402 892 436
rect 944 563 978 597
<< poly >>
rect 242 619 272 645
rect 328 619 358 645
rect 414 619 444 645
rect 500 619 530 645
rect 601 619 631 645
rect 687 619 717 645
rect 817 619 847 645
rect 903 619 933 645
rect 106 451 136 477
rect 106 305 136 367
rect 242 335 272 367
rect 328 335 358 367
rect 414 335 444 367
rect 500 335 530 367
rect 601 335 631 367
rect 687 335 717 367
rect 817 335 847 367
rect 242 319 537 335
rect 106 289 177 305
rect 106 255 127 289
rect 161 255 177 289
rect 106 239 177 255
rect 242 285 283 319
rect 317 285 351 319
rect 385 285 419 319
rect 453 285 487 319
rect 521 285 537 319
rect 242 269 537 285
rect 579 319 645 335
rect 579 285 595 319
rect 629 285 645 319
rect 579 269 645 285
rect 106 217 136 239
rect 242 217 272 269
rect 328 217 358 269
rect 414 217 444 269
rect 500 217 530 269
rect 615 217 645 269
rect 687 319 753 335
rect 687 285 703 319
rect 737 285 753 319
rect 687 269 753 285
rect 795 319 861 335
rect 795 285 811 319
rect 845 285 861 319
rect 795 269 861 285
rect 903 325 933 367
rect 903 309 1031 325
rect 903 275 981 309
rect 1015 275 1031 309
rect 687 217 717 269
rect 795 217 825 269
rect 903 259 1031 275
rect 903 217 933 259
rect 106 107 136 133
rect 242 23 272 49
rect 328 23 358 49
rect 414 23 444 49
rect 500 23 530 49
rect 615 23 645 49
rect 687 23 717 49
rect 795 23 825 49
rect 903 23 933 49
<< polycont >>
rect 127 255 161 289
rect 283 285 317 319
rect 351 285 385 319
rect 419 285 453 319
rect 487 285 521 319
rect 595 285 629 319
rect 703 285 737 319
rect 811 285 845 319
rect 981 275 1015 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 181 597 247 649
rect 181 563 197 597
rect 231 563 247 597
rect 181 556 247 563
rect 353 597 419 649
rect 353 563 369 597
rect 403 563 419 597
rect 353 556 419 563
rect 525 597 591 649
rect 525 563 541 597
rect 575 563 591 597
rect 525 556 591 563
rect 712 597 778 649
rect 712 563 728 597
rect 762 563 778 597
rect 712 556 778 563
rect 928 597 994 649
rect 928 563 944 597
rect 978 563 994 597
rect 928 556 994 563
rect 41 486 1031 522
rect 41 425 91 486
rect 41 391 57 425
rect 41 191 91 391
rect 41 157 57 191
rect 41 139 91 157
rect 127 289 163 438
rect 161 255 163 289
rect 127 76 163 255
rect 197 436 491 452
rect 197 402 283 436
rect 317 402 455 436
rect 489 402 491 436
rect 197 371 491 402
rect 525 436 896 452
rect 525 402 642 436
rect 676 402 858 436
rect 892 402 896 436
rect 525 386 896 402
rect 197 249 233 371
rect 525 335 559 386
rect 267 319 559 335
rect 267 285 283 319
rect 317 285 351 319
rect 385 285 419 319
rect 453 285 487 319
rect 521 285 559 319
rect 267 283 559 285
rect 197 215 491 249
rect 273 205 319 215
rect 197 163 239 179
rect 231 129 239 163
rect 197 95 239 129
rect 231 61 239 95
rect 197 17 239 61
rect 273 171 283 205
rect 317 171 319 205
rect 453 205 491 215
rect 273 101 319 171
rect 273 67 283 101
rect 317 67 319 101
rect 273 51 319 67
rect 353 147 369 181
rect 403 147 419 181
rect 353 95 419 147
rect 353 61 369 95
rect 403 61 419 95
rect 353 17 419 61
rect 453 171 455 205
rect 489 171 491 205
rect 525 233 559 283
rect 593 319 653 350
rect 593 285 595 319
rect 629 285 653 319
rect 593 269 653 285
rect 687 319 754 350
rect 687 285 703 319
rect 737 285 754 319
rect 687 269 754 285
rect 788 319 929 350
rect 788 285 811 319
rect 845 285 929 319
rect 788 267 929 285
rect 965 309 1031 486
rect 965 275 981 309
rect 1015 275 1031 309
rect 965 267 1031 275
rect 525 205 994 233
rect 525 199 944 205
rect 453 101 491 171
rect 659 171 944 199
rect 978 171 994 205
rect 453 67 455 101
rect 489 67 491 101
rect 453 51 491 67
rect 540 131 556 165
rect 590 131 606 165
rect 540 91 606 131
rect 540 57 556 91
rect 590 57 606 91
rect 540 17 606 57
rect 659 101 994 171
rect 659 67 944 101
rect 978 67 994 101
rect 659 51 994 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4b_4
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5337754
string GDS_START 5329562
<< end >>
