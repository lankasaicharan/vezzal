magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
<< pwell >>
rect 529 241 1247 259
rect 1 49 1247 241
rect 0 0 1248 49
<< scnmos >>
rect 80 47 110 215
rect 226 47 256 215
rect 312 47 342 215
rect 398 47 428 215
rect 608 65 638 233
rect 694 65 724 233
rect 780 65 810 233
rect 952 65 982 233
rect 1038 65 1068 233
rect 1124 65 1154 233
<< scpmoshvt >>
rect 132 367 162 619
rect 218 367 248 619
rect 312 367 342 619
rect 398 367 428 619
rect 515 367 545 619
rect 601 367 631 619
rect 880 367 910 619
rect 966 367 996 619
rect 1052 367 1082 619
rect 1138 367 1168 619
<< ndiff >>
rect 555 221 608 233
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 101 80 169
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 97 226 215
rect 110 63 127 97
rect 161 63 226 97
rect 110 47 226 63
rect 256 89 312 215
rect 256 55 267 89
rect 301 55 312 89
rect 256 47 312 55
rect 342 159 398 215
rect 342 125 353 159
rect 387 125 398 159
rect 342 47 398 125
rect 428 167 495 215
rect 428 133 453 167
rect 487 133 495 167
rect 428 93 495 133
rect 428 59 453 93
rect 487 59 495 93
rect 555 187 563 221
rect 597 187 608 221
rect 555 111 608 187
rect 555 77 563 111
rect 597 77 608 111
rect 555 65 608 77
rect 638 179 694 233
rect 638 145 649 179
rect 683 145 694 179
rect 638 107 694 145
rect 638 73 649 107
rect 683 73 694 107
rect 638 65 694 73
rect 724 221 780 233
rect 724 187 735 221
rect 769 187 780 221
rect 724 111 780 187
rect 724 77 735 111
rect 769 77 780 111
rect 724 65 780 77
rect 810 179 952 233
rect 810 145 821 179
rect 855 145 907 179
rect 941 145 952 179
rect 810 107 952 145
rect 810 73 821 107
rect 855 73 907 107
rect 941 73 952 107
rect 810 65 952 73
rect 982 225 1038 233
rect 982 191 993 225
rect 1027 191 1038 225
rect 982 111 1038 191
rect 982 77 993 111
rect 1027 77 1038 111
rect 982 65 1038 77
rect 1068 225 1124 233
rect 1068 191 1079 225
rect 1113 191 1124 225
rect 1068 153 1124 191
rect 1068 119 1079 153
rect 1113 119 1124 153
rect 1068 65 1124 119
rect 1154 179 1221 233
rect 1154 145 1179 179
rect 1213 145 1221 179
rect 1154 111 1221 145
rect 1154 77 1179 111
rect 1213 77 1221 111
rect 1154 65 1221 77
rect 428 47 495 59
<< pdiff >>
rect 56 607 132 619
rect 56 573 87 607
rect 121 573 132 607
rect 56 510 132 573
rect 56 476 87 510
rect 121 476 132 510
rect 56 413 132 476
rect 56 379 68 413
rect 102 379 132 413
rect 56 367 132 379
rect 162 599 218 619
rect 162 565 173 599
rect 207 565 218 599
rect 162 512 218 565
rect 162 478 173 512
rect 207 478 218 512
rect 162 420 218 478
rect 162 386 173 420
rect 207 386 218 420
rect 162 367 218 386
rect 248 607 312 619
rect 248 573 263 607
rect 297 573 312 607
rect 248 494 312 573
rect 248 460 263 494
rect 297 460 312 494
rect 248 367 312 460
rect 342 599 398 619
rect 342 565 353 599
rect 387 565 398 599
rect 342 516 398 565
rect 342 482 353 516
rect 387 482 398 516
rect 342 434 398 482
rect 342 400 353 434
rect 387 400 398 434
rect 342 367 398 400
rect 428 611 515 619
rect 428 577 455 611
rect 489 577 515 611
rect 428 525 515 577
rect 428 491 455 525
rect 489 491 515 525
rect 428 367 515 491
rect 545 607 601 619
rect 545 573 556 607
rect 590 573 601 607
rect 545 525 601 573
rect 545 491 556 525
rect 590 491 601 525
rect 545 367 601 491
rect 631 605 688 619
rect 631 571 642 605
rect 676 571 688 605
rect 631 367 688 571
rect 827 502 880 619
rect 827 468 835 502
rect 869 468 880 502
rect 827 367 880 468
rect 910 562 966 619
rect 910 528 921 562
rect 955 528 966 562
rect 910 367 966 528
rect 996 599 1052 619
rect 996 565 1007 599
rect 1041 565 1052 599
rect 996 508 1052 565
rect 996 474 1007 508
rect 1041 474 1052 508
rect 996 413 1052 474
rect 996 379 1007 413
rect 1041 379 1052 413
rect 996 367 1052 379
rect 1082 611 1138 619
rect 1082 577 1093 611
rect 1127 577 1138 611
rect 1082 536 1138 577
rect 1082 502 1093 536
rect 1127 502 1138 536
rect 1082 457 1138 502
rect 1082 423 1093 457
rect 1127 423 1138 457
rect 1082 367 1138 423
rect 1168 599 1221 619
rect 1168 565 1179 599
rect 1213 565 1221 599
rect 1168 508 1221 565
rect 1168 474 1179 508
rect 1213 474 1221 508
rect 1168 413 1221 474
rect 1168 379 1179 413
rect 1213 379 1221 413
rect 1168 367 1221 379
<< ndiffc >>
rect 35 169 69 203
rect 35 67 69 101
rect 127 63 161 97
rect 267 55 301 89
rect 353 125 387 159
rect 453 133 487 167
rect 453 59 487 93
rect 563 187 597 221
rect 563 77 597 111
rect 649 145 683 179
rect 649 73 683 107
rect 735 187 769 221
rect 735 77 769 111
rect 821 145 855 179
rect 907 145 941 179
rect 821 73 855 107
rect 907 73 941 107
rect 993 191 1027 225
rect 993 77 1027 111
rect 1079 191 1113 225
rect 1079 119 1113 153
rect 1179 145 1213 179
rect 1179 77 1213 111
<< pdiffc >>
rect 87 573 121 607
rect 87 476 121 510
rect 68 379 102 413
rect 173 565 207 599
rect 173 478 207 512
rect 173 386 207 420
rect 263 573 297 607
rect 263 460 297 494
rect 353 565 387 599
rect 353 482 387 516
rect 353 400 387 434
rect 455 577 489 611
rect 455 491 489 525
rect 556 573 590 607
rect 556 491 590 525
rect 642 571 676 605
rect 835 468 869 502
rect 921 528 955 562
rect 1007 565 1041 599
rect 1007 474 1041 508
rect 1007 379 1041 413
rect 1093 577 1127 611
rect 1093 502 1127 536
rect 1093 423 1127 457
rect 1179 565 1213 599
rect 1179 474 1213 508
rect 1179 379 1213 413
<< poly >>
rect 132 619 162 645
rect 218 619 248 645
rect 312 619 342 645
rect 398 619 428 645
rect 515 619 545 645
rect 601 619 631 645
rect 880 619 910 645
rect 966 619 996 645
rect 1052 619 1082 645
rect 1138 619 1168 645
rect 132 335 162 367
rect 218 335 248 367
rect 312 335 342 367
rect 398 335 428 367
rect 132 319 270 335
rect 132 299 220 319
rect 80 285 220 299
rect 254 285 270 319
rect 80 269 270 285
rect 312 319 451 335
rect 515 331 545 367
rect 601 331 631 367
rect 880 335 910 367
rect 966 335 996 367
rect 1052 335 1082 367
rect 1138 335 1168 367
rect 312 285 401 319
rect 435 285 451 319
rect 312 269 451 285
rect 493 315 724 331
rect 493 281 509 315
rect 543 281 577 315
rect 611 281 724 315
rect 80 215 110 269
rect 226 215 256 269
rect 312 215 342 269
rect 398 215 428 269
rect 493 265 724 281
rect 766 319 996 335
rect 766 285 782 319
rect 816 285 850 319
rect 884 285 996 319
rect 766 269 996 285
rect 1038 319 1168 335
rect 1038 285 1093 319
rect 1127 285 1168 319
rect 1038 269 1168 285
rect 608 233 638 265
rect 694 233 724 265
rect 780 233 810 269
rect 952 233 982 269
rect 1038 233 1068 269
rect 1124 233 1154 269
rect 80 21 110 47
rect 226 21 256 47
rect 312 21 342 47
rect 398 21 428 47
rect 608 39 638 65
rect 694 39 724 65
rect 780 39 810 65
rect 952 39 982 65
rect 1038 39 1068 65
rect 1124 39 1154 65
<< polycont >>
rect 220 285 254 319
rect 401 285 435 319
rect 509 281 543 315
rect 577 281 611 315
rect 782 285 816 319
rect 850 285 884 319
rect 1093 285 1127 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 60 607 129 649
rect 60 573 87 607
rect 121 573 129 607
rect 60 510 129 573
rect 60 476 87 510
rect 121 476 129 510
rect 60 454 129 476
rect 163 599 213 615
rect 163 565 173 599
rect 207 565 213 599
rect 163 512 213 565
rect 163 478 173 512
rect 207 478 213 512
rect 60 413 102 454
rect 163 420 213 478
rect 247 607 313 649
rect 247 573 263 607
rect 297 573 313 607
rect 247 494 313 573
rect 247 460 263 494
rect 297 460 313 494
rect 247 452 313 460
rect 349 599 403 615
rect 349 565 353 599
rect 387 565 403 599
rect 349 516 403 565
rect 349 482 353 516
rect 387 482 403 516
rect 439 611 505 649
rect 439 577 455 611
rect 489 577 505 611
rect 439 525 505 577
rect 439 491 455 525
rect 489 491 505 525
rect 439 487 505 491
rect 540 607 606 615
rect 540 573 556 607
rect 590 573 606 607
rect 540 525 606 573
rect 640 605 692 649
rect 640 571 642 605
rect 676 571 692 605
rect 640 555 692 571
rect 726 579 971 613
rect 540 491 556 525
rect 590 521 606 525
rect 726 521 771 579
rect 905 562 971 579
rect 905 528 921 562
rect 955 528 971 562
rect 590 491 771 521
rect 540 487 771 491
rect 819 502 871 527
rect 905 520 971 528
rect 1005 599 1043 615
rect 1005 565 1007 599
rect 1041 565 1043 599
rect 60 379 68 413
rect 60 363 102 379
rect 136 386 173 420
rect 207 418 213 420
rect 349 451 403 482
rect 819 468 835 502
rect 869 486 871 502
rect 1005 508 1043 565
rect 1005 486 1007 508
rect 869 474 1007 486
rect 1041 474 1043 508
rect 869 468 1043 474
rect 819 452 1043 468
rect 349 434 771 451
rect 349 418 353 434
rect 207 400 353 418
rect 387 418 771 434
rect 387 417 971 418
rect 387 400 389 417
rect 207 386 389 400
rect 136 384 389 386
rect 729 384 971 417
rect 136 249 170 384
rect 423 350 695 383
rect 204 319 365 350
rect 423 349 900 350
rect 423 335 457 349
rect 204 285 220 319
rect 254 285 365 319
rect 19 203 85 219
rect 136 215 297 249
rect 19 169 35 203
rect 69 181 85 203
rect 69 169 229 181
rect 19 147 229 169
rect 19 101 83 147
rect 19 67 35 101
rect 69 67 83 101
rect 19 51 83 67
rect 117 97 161 113
rect 117 63 127 97
rect 117 17 161 63
rect 195 89 229 147
rect 263 163 297 215
rect 331 235 365 285
rect 399 319 457 335
rect 399 285 401 319
rect 435 285 457 319
rect 661 319 900 349
rect 399 269 457 285
rect 493 281 509 315
rect 543 281 577 315
rect 611 281 627 315
rect 661 285 782 319
rect 816 285 850 319
rect 884 285 900 319
rect 661 281 900 285
rect 937 321 971 384
rect 1005 413 1043 452
rect 1077 611 1143 649
rect 1077 577 1093 611
rect 1127 577 1143 611
rect 1077 536 1143 577
rect 1077 502 1093 536
rect 1127 502 1143 536
rect 1077 457 1143 502
rect 1077 423 1093 457
rect 1127 423 1143 457
rect 1177 599 1231 615
rect 1177 565 1179 599
rect 1213 565 1231 599
rect 1177 508 1231 565
rect 1177 474 1179 508
rect 1213 474 1231 508
rect 1005 379 1007 413
rect 1041 389 1043 413
rect 1177 413 1231 474
rect 1177 389 1179 413
rect 1041 379 1179 389
rect 1213 379 1231 413
rect 1005 355 1231 379
rect 937 319 1143 321
rect 937 285 1093 319
rect 1127 285 1143 319
rect 937 281 1143 285
rect 493 235 527 281
rect 1177 247 1231 355
rect 331 201 527 235
rect 561 225 1029 247
rect 561 221 993 225
rect 561 187 563 221
rect 597 213 735 221
rect 597 187 599 213
rect 263 159 403 163
rect 263 125 353 159
rect 387 125 403 159
rect 263 123 403 125
rect 437 133 453 167
rect 487 133 503 167
rect 437 93 503 133
rect 437 89 453 93
rect 195 55 267 89
rect 301 59 453 89
rect 487 59 503 93
rect 561 111 599 187
rect 733 187 735 213
rect 769 213 993 221
rect 769 187 771 213
rect 561 77 563 111
rect 597 77 599 111
rect 561 60 599 77
rect 633 145 649 179
rect 683 145 699 179
rect 633 107 699 145
rect 633 73 649 107
rect 683 73 699 107
rect 301 55 503 59
rect 195 51 503 55
rect 633 17 699 73
rect 733 111 771 187
rect 991 191 993 213
rect 1027 191 1029 225
rect 733 77 735 111
rect 769 77 771 111
rect 733 60 771 77
rect 805 145 821 179
rect 855 145 907 179
rect 941 145 957 179
rect 805 107 957 145
rect 805 73 821 107
rect 855 73 907 107
rect 941 73 957 107
rect 805 17 957 73
rect 991 111 1029 191
rect 1063 225 1231 247
rect 1063 191 1079 225
rect 1113 213 1231 225
rect 1113 191 1129 213
rect 1063 153 1129 191
rect 1063 119 1079 153
rect 1113 119 1129 153
rect 1163 145 1179 179
rect 1213 145 1229 179
rect 991 77 993 111
rect 1027 85 1029 111
rect 1163 111 1229 145
rect 1163 85 1179 111
rect 1027 77 1179 85
rect 1213 77 1229 111
rect 991 51 1229 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xnor2_2
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1183 538 1217 572 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 1183 464 1217 498 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 1183 390 1217 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4370572
string GDS_START 4360050
<< end >>
