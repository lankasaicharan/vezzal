magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1778 1975
<< nwell >>
rect -38 331 518 704
<< pwell >>
rect 163 157 435 241
rect 58 49 435 157
rect 0 0 480 49
<< scnmos >>
rect 137 47 167 131
rect 239 47 269 215
rect 311 47 341 215
<< scpmoshvt >>
rect 93 367 123 451
rect 198 367 228 619
rect 284 367 314 619
<< ndiff >>
rect 189 131 239 215
rect 84 106 137 131
rect 84 72 92 106
rect 126 72 137 106
rect 84 47 137 72
rect 167 93 239 131
rect 167 59 178 93
rect 212 59 239 93
rect 167 47 239 59
rect 269 47 311 215
rect 341 203 409 215
rect 341 169 359 203
rect 393 169 409 203
rect 341 101 409 169
rect 341 67 359 101
rect 393 67 409 101
rect 341 47 409 67
<< pdiff >>
rect 145 607 198 619
rect 145 573 153 607
rect 187 573 198 607
rect 145 535 198 573
rect 145 501 153 535
rect 187 501 198 535
rect 145 457 198 501
rect 145 451 153 457
rect 40 426 93 451
rect 40 392 48 426
rect 82 392 93 426
rect 40 367 93 392
rect 123 423 153 451
rect 187 423 198 457
rect 123 367 198 423
rect 228 599 284 619
rect 228 565 239 599
rect 273 565 284 599
rect 228 512 284 565
rect 228 478 239 512
rect 273 478 284 512
rect 228 423 284 478
rect 228 389 239 423
rect 273 389 284 423
rect 228 367 284 389
rect 314 607 367 619
rect 314 573 325 607
rect 359 573 367 607
rect 314 500 367 573
rect 314 466 325 500
rect 359 466 367 500
rect 314 367 367 466
<< ndiffc >>
rect 92 72 126 106
rect 178 59 212 93
rect 359 169 393 203
rect 359 67 393 101
<< pdiffc >>
rect 153 573 187 607
rect 153 501 187 535
rect 48 392 82 426
rect 153 423 187 457
rect 239 565 273 599
rect 239 478 273 512
rect 239 389 273 423
rect 325 573 359 607
rect 325 466 359 500
<< poly >>
rect 198 619 228 645
rect 284 619 314 645
rect 93 451 123 477
rect 93 321 123 367
rect 25 305 123 321
rect 25 271 41 305
rect 75 271 123 305
rect 198 303 228 367
rect 284 345 314 367
rect 284 315 380 345
rect 311 305 380 315
rect 25 237 123 271
rect 176 287 242 303
rect 176 253 192 287
rect 226 267 242 287
rect 311 271 330 305
rect 364 271 380 305
rect 226 253 269 267
rect 176 237 269 253
rect 25 203 41 237
rect 75 203 123 237
rect 239 215 269 237
rect 311 237 380 271
rect 311 215 341 237
rect 25 189 123 203
rect 25 159 167 189
rect 137 131 167 159
rect 137 21 167 47
rect 239 21 269 47
rect 311 21 341 47
<< polycont >>
rect 41 271 75 305
rect 192 253 226 287
rect 330 271 364 305
rect 41 203 75 237
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 137 607 189 649
rect 137 573 153 607
rect 187 573 189 607
rect 137 535 189 573
rect 137 501 153 535
rect 187 501 189 535
rect 137 457 189 501
rect 32 426 98 442
rect 32 392 48 426
rect 82 392 98 426
rect 137 423 153 457
rect 187 423 189 457
rect 137 407 189 423
rect 223 599 275 615
rect 223 565 239 599
rect 273 565 275 599
rect 223 512 275 565
rect 223 478 239 512
rect 273 478 275 512
rect 223 423 275 478
rect 309 607 375 649
rect 309 573 325 607
rect 359 573 375 607
rect 309 500 375 573
rect 309 466 325 500
rect 359 466 375 500
rect 309 457 375 466
rect 32 373 98 392
rect 223 389 239 423
rect 273 389 463 423
rect 32 355 156 373
rect 32 339 327 355
rect 122 321 327 339
rect 291 305 380 321
rect 17 271 41 305
rect 75 271 91 305
rect 17 237 91 271
rect 17 203 41 237
rect 75 203 91 237
rect 125 253 192 287
rect 226 253 257 287
rect 125 203 257 253
rect 291 271 330 305
rect 364 271 380 305
rect 291 255 380 271
rect 291 169 325 255
rect 414 219 463 389
rect 76 135 325 169
rect 359 203 463 219
rect 393 169 463 203
rect 76 106 128 135
rect 76 72 92 106
rect 126 72 128 106
rect 359 101 463 169
rect 76 56 128 72
rect 162 93 228 101
rect 162 59 178 93
rect 212 59 228 93
rect 162 17 228 59
rect 393 67 463 101
rect 359 51 463 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2b_1
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4465538
string GDS_START 4460780
<< end >>
