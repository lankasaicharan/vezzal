magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 231 248 849 290
rect 1 49 849 248
rect 0 0 864 49
<< scnmos >>
rect 84 74 114 222
rect 323 136 353 264
rect 455 136 485 264
rect 632 136 662 264
rect 727 136 757 264
<< scpmoshvt >>
rect 86 368 116 592
rect 368 392 398 592
rect 452 392 482 592
rect 542 392 572 592
rect 748 392 778 592
<< ndiff >>
rect 257 253 323 264
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 210 185 222
rect 114 176 139 210
rect 173 176 185 210
rect 114 120 185 176
rect 257 219 269 253
rect 303 219 323 253
rect 257 182 323 219
rect 257 148 278 182
rect 312 148 323 182
rect 257 136 323 148
rect 353 185 455 264
rect 353 151 375 185
rect 409 151 455 185
rect 353 136 455 151
rect 485 196 632 264
rect 485 162 496 196
rect 530 162 587 196
rect 621 162 632 196
rect 485 136 632 162
rect 662 136 727 264
rect 757 256 823 264
rect 757 222 768 256
rect 802 222 823 256
rect 757 188 823 222
rect 757 154 777 188
rect 811 154 823 188
rect 757 136 823 154
rect 114 86 139 120
rect 173 86 185 120
rect 114 74 185 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 368 592
rect 116 546 139 580
rect 173 546 230 580
rect 264 546 321 580
rect 355 546 368 580
rect 116 496 368 546
rect 116 462 139 496
rect 173 462 230 496
rect 264 462 321 496
rect 355 462 368 496
rect 116 392 368 462
rect 398 392 452 592
rect 482 580 542 592
rect 482 546 495 580
rect 529 546 542 580
rect 482 509 542 546
rect 482 475 495 509
rect 529 475 542 509
rect 482 438 542 475
rect 482 404 495 438
rect 529 404 542 438
rect 482 392 542 404
rect 572 580 748 592
rect 572 546 595 580
rect 629 546 691 580
rect 725 546 748 580
rect 572 496 748 546
rect 572 462 595 496
rect 629 462 691 496
rect 725 462 748 496
rect 572 392 748 462
rect 778 580 837 592
rect 778 546 791 580
rect 825 546 837 580
rect 778 512 837 546
rect 778 478 791 512
rect 825 478 837 512
rect 778 444 837 478
rect 778 410 791 444
rect 825 410 837 444
rect 778 392 837 410
rect 116 368 169 392
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 176 173 210
rect 269 219 303 253
rect 278 148 312 182
rect 375 151 409 185
rect 496 162 530 196
rect 587 162 621 196
rect 768 222 802 256
rect 777 154 811 188
rect 139 86 173 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 546 173 580
rect 230 546 264 580
rect 321 546 355 580
rect 139 462 173 496
rect 230 462 264 496
rect 321 462 355 496
rect 495 546 529 580
rect 495 475 529 509
rect 495 404 529 438
rect 595 546 629 580
rect 691 546 725 580
rect 595 462 629 496
rect 691 462 725 496
rect 791 546 825 580
rect 791 478 825 512
rect 791 410 825 444
<< poly >>
rect 86 592 116 618
rect 368 592 398 618
rect 452 592 482 618
rect 542 592 572 618
rect 748 592 778 618
rect 368 377 398 392
rect 452 377 482 392
rect 542 377 572 392
rect 748 377 778 392
rect 86 353 116 368
rect 365 360 401 377
rect 83 330 119 353
rect 267 344 401 360
rect 83 314 219 330
rect 83 280 101 314
rect 135 280 169 314
rect 203 280 219 314
rect 267 310 283 344
rect 317 310 351 344
rect 385 310 401 344
rect 267 294 401 310
rect 83 264 219 280
rect 323 264 353 294
rect 449 282 485 377
rect 539 360 575 377
rect 745 360 781 377
rect 539 344 667 360
rect 539 310 617 344
rect 651 310 667 344
rect 539 294 667 310
rect 727 344 793 360
rect 727 310 743 344
rect 777 310 793 344
rect 727 294 793 310
rect 455 264 485 282
rect 632 264 662 294
rect 727 264 757 294
rect 84 222 114 264
rect 323 110 353 136
rect 455 114 485 136
rect 455 98 531 114
rect 632 110 662 136
rect 727 110 757 136
rect 84 48 114 74
rect 455 64 481 98
rect 515 64 531 98
rect 455 48 531 64
<< polycont >>
rect 101 280 135 314
rect 169 280 203 314
rect 283 310 317 344
rect 351 310 385 344
rect 617 310 651 344
rect 743 310 777 344
rect 481 64 515 98
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 17 580 89 596
rect 17 546 39 580
rect 73 546 89 580
rect 17 497 89 546
rect 17 463 39 497
rect 73 463 89 497
rect 17 414 89 463
rect 123 580 371 649
rect 123 546 139 580
rect 173 546 230 580
rect 264 546 321 580
rect 355 546 371 580
rect 123 496 371 546
rect 123 462 139 496
rect 173 462 230 496
rect 264 462 321 496
rect 355 462 371 496
rect 479 580 545 596
rect 479 546 495 580
rect 529 546 545 580
rect 479 509 545 546
rect 479 475 495 509
rect 529 475 545 509
rect 479 438 545 475
rect 579 580 741 649
rect 579 546 595 580
rect 629 546 691 580
rect 725 546 741 580
rect 579 496 741 546
rect 579 462 595 496
rect 629 462 691 496
rect 725 462 741 496
rect 775 580 841 596
rect 775 546 791 580
rect 825 546 841 580
rect 775 512 841 546
rect 775 478 791 512
rect 825 478 841 512
rect 479 428 495 438
rect 17 380 39 414
rect 73 380 89 414
rect 17 364 89 380
rect 185 404 495 428
rect 529 428 545 438
rect 775 444 841 478
rect 775 428 791 444
rect 529 410 791 428
rect 825 410 841 444
rect 529 404 841 410
rect 185 394 841 404
rect 17 226 51 364
rect 185 330 219 394
rect 479 388 567 394
rect 85 314 219 330
rect 85 280 101 314
rect 135 280 169 314
rect 203 280 219 314
rect 267 344 401 360
rect 267 310 283 344
rect 317 310 351 344
rect 385 310 401 344
rect 267 294 401 310
rect 85 264 219 280
rect 533 264 567 388
rect 601 344 667 360
rect 601 310 617 344
rect 651 310 667 344
rect 601 298 667 310
rect 727 344 839 360
rect 727 310 743 344
rect 777 310 839 344
rect 727 298 839 310
rect 253 253 499 260
rect 17 210 89 226
rect 17 176 39 210
rect 73 176 89 210
rect 17 120 89 176
rect 17 86 39 120
rect 73 86 89 120
rect 17 70 89 86
rect 123 210 189 226
rect 123 176 139 210
rect 173 176 189 210
rect 123 120 189 176
rect 253 219 269 253
rect 303 226 499 253
rect 533 256 827 264
rect 533 230 768 256
rect 303 219 319 226
rect 253 182 319 219
rect 465 196 499 226
rect 752 222 768 230
rect 802 222 827 256
rect 253 148 278 182
rect 312 148 319 182
rect 253 132 319 148
rect 353 151 375 185
rect 409 151 431 185
rect 465 162 496 196
rect 530 162 587 196
rect 621 162 637 196
rect 752 188 827 222
rect 752 167 777 188
rect 123 86 139 120
rect 173 86 189 120
rect 123 17 189 86
rect 353 17 431 151
rect 811 154 827 188
rect 777 132 827 154
rect 465 98 743 128
rect 465 64 481 98
rect 515 64 743 98
rect 465 51 743 64
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o211a_1
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 1063330
string GDS_START 1055350
<< end >>
