magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 331 1958 704
<< pwell >>
rect 11 49 1918 241
rect 0 0 1920 49
<< scnmos >>
rect 90 131 120 215
rect 192 131 222 215
rect 298 131 328 215
rect 384 131 414 215
rect 456 131 486 215
rect 574 131 604 215
rect 660 131 690 215
rect 768 131 798 215
rect 854 131 884 215
rect 948 131 978 215
rect 1020 131 1050 215
rect 1092 131 1122 215
rect 1207 47 1237 215
rect 1293 47 1323 215
rect 1379 47 1409 215
rect 1465 47 1495 215
rect 1551 47 1581 215
rect 1637 47 1667 215
rect 1723 47 1753 215
rect 1809 47 1839 215
<< scpmoshvt >>
rect 80 440 110 568
rect 166 440 196 568
rect 298 419 328 547
rect 415 419 445 547
rect 487 419 517 547
rect 574 419 604 547
rect 660 419 690 547
rect 768 419 798 547
rect 854 419 884 547
rect 948 419 978 547
rect 1020 419 1050 547
rect 1092 419 1122 547
rect 1207 367 1237 619
rect 1293 367 1323 619
rect 1379 367 1409 619
rect 1465 367 1495 619
rect 1551 367 1581 619
rect 1637 367 1667 619
rect 1723 367 1753 619
rect 1809 367 1839 619
<< ndiff >>
rect 37 191 90 215
rect 37 157 45 191
rect 79 157 90 191
rect 37 131 90 157
rect 120 173 192 215
rect 120 139 131 173
rect 165 139 192 173
rect 120 131 192 139
rect 222 203 298 215
rect 222 169 233 203
rect 267 169 298 203
rect 222 131 298 169
rect 328 203 384 215
rect 328 169 339 203
rect 373 169 384 203
rect 328 131 384 169
rect 414 131 456 215
rect 486 192 574 215
rect 486 158 501 192
rect 535 158 574 192
rect 486 131 574 158
rect 604 203 660 215
rect 604 169 615 203
rect 649 169 660 203
rect 604 131 660 169
rect 690 173 768 215
rect 690 139 705 173
rect 739 139 768 173
rect 690 131 768 139
rect 798 203 854 215
rect 798 169 809 203
rect 843 169 854 203
rect 798 131 854 169
rect 884 190 948 215
rect 884 156 903 190
rect 937 156 948 190
rect 884 131 948 156
rect 978 131 1020 215
rect 1050 131 1092 215
rect 1122 131 1207 215
rect 1150 100 1207 131
rect 1150 66 1158 100
rect 1192 66 1207 100
rect 1150 47 1207 66
rect 1237 203 1293 215
rect 1237 169 1248 203
rect 1282 169 1293 203
rect 1237 101 1293 169
rect 1237 67 1248 101
rect 1282 67 1293 101
rect 1237 47 1293 67
rect 1323 175 1379 215
rect 1323 141 1334 175
rect 1368 141 1379 175
rect 1323 89 1379 141
rect 1323 55 1334 89
rect 1368 55 1379 89
rect 1323 47 1379 55
rect 1409 203 1465 215
rect 1409 169 1420 203
rect 1454 169 1465 203
rect 1409 101 1465 169
rect 1409 67 1420 101
rect 1454 67 1465 101
rect 1409 47 1465 67
rect 1495 175 1551 215
rect 1495 141 1506 175
rect 1540 141 1551 175
rect 1495 89 1551 141
rect 1495 55 1506 89
rect 1540 55 1551 89
rect 1495 47 1551 55
rect 1581 186 1637 215
rect 1581 152 1592 186
rect 1626 152 1637 186
rect 1581 101 1637 152
rect 1581 67 1592 101
rect 1626 67 1637 101
rect 1581 47 1637 67
rect 1667 123 1723 215
rect 1667 89 1678 123
rect 1712 89 1723 123
rect 1667 47 1723 89
rect 1753 186 1809 215
rect 1753 152 1764 186
rect 1798 152 1809 186
rect 1753 101 1809 152
rect 1753 67 1764 101
rect 1798 67 1809 101
rect 1753 47 1809 67
rect 1839 123 1892 215
rect 1839 89 1850 123
rect 1884 89 1892 123
rect 1839 47 1892 89
<< pdiff >>
rect 27 554 80 568
rect 27 520 35 554
rect 69 520 80 554
rect 27 486 80 520
rect 27 452 35 486
rect 69 452 80 486
rect 27 440 80 452
rect 110 560 166 568
rect 110 526 121 560
rect 155 526 166 560
rect 110 440 166 526
rect 196 547 268 568
rect 1154 607 1207 619
rect 1154 573 1162 607
rect 1196 573 1207 607
rect 1154 547 1207 573
rect 196 506 298 547
rect 196 472 226 506
rect 260 472 298 506
rect 196 440 298 472
rect 218 419 298 440
rect 328 529 415 547
rect 328 495 370 529
rect 404 495 415 529
rect 328 461 415 495
rect 328 427 370 461
rect 404 427 415 461
rect 328 419 415 427
rect 445 419 487 547
rect 517 539 574 547
rect 517 505 529 539
rect 563 505 574 539
rect 517 471 574 505
rect 517 437 529 471
rect 563 437 574 471
rect 517 419 574 437
rect 604 537 660 547
rect 604 503 615 537
rect 649 503 660 537
rect 604 469 660 503
rect 604 435 615 469
rect 649 435 660 469
rect 604 419 660 435
rect 690 529 768 547
rect 690 495 712 529
rect 746 495 768 529
rect 690 419 768 495
rect 798 537 854 547
rect 798 503 809 537
rect 843 503 854 537
rect 798 469 854 503
rect 798 435 809 469
rect 843 435 854 469
rect 798 419 854 435
rect 884 537 948 547
rect 884 503 899 537
rect 933 503 948 537
rect 884 469 948 503
rect 884 435 899 469
rect 933 435 948 469
rect 884 419 948 435
rect 978 419 1020 547
rect 1050 419 1092 547
rect 1122 524 1207 547
rect 1122 490 1162 524
rect 1196 490 1207 524
rect 1122 419 1207 490
rect 1154 367 1207 419
rect 1237 599 1293 619
rect 1237 565 1248 599
rect 1282 565 1293 599
rect 1237 508 1293 565
rect 1237 474 1248 508
rect 1282 474 1293 508
rect 1237 413 1293 474
rect 1237 379 1248 413
rect 1282 379 1293 413
rect 1237 367 1293 379
rect 1323 607 1379 619
rect 1323 573 1334 607
rect 1368 573 1379 607
rect 1323 528 1379 573
rect 1323 494 1334 528
rect 1368 494 1379 528
rect 1323 455 1379 494
rect 1323 421 1334 455
rect 1368 421 1379 455
rect 1323 367 1379 421
rect 1409 599 1465 619
rect 1409 565 1420 599
rect 1454 565 1465 599
rect 1409 508 1465 565
rect 1409 474 1420 508
rect 1454 474 1465 508
rect 1409 413 1465 474
rect 1409 379 1420 413
rect 1454 379 1465 413
rect 1409 367 1465 379
rect 1495 607 1551 619
rect 1495 573 1506 607
rect 1540 573 1551 607
rect 1495 528 1551 573
rect 1495 494 1506 528
rect 1540 494 1551 528
rect 1495 455 1551 494
rect 1495 421 1506 455
rect 1540 421 1551 455
rect 1495 367 1551 421
rect 1581 599 1637 619
rect 1581 565 1592 599
rect 1626 565 1637 599
rect 1581 508 1637 565
rect 1581 474 1592 508
rect 1626 474 1637 508
rect 1581 413 1637 474
rect 1581 379 1592 413
rect 1626 379 1637 413
rect 1581 367 1637 379
rect 1667 607 1723 619
rect 1667 573 1678 607
rect 1712 573 1723 607
rect 1667 528 1723 573
rect 1667 494 1678 528
rect 1712 494 1723 528
rect 1667 455 1723 494
rect 1667 421 1678 455
rect 1712 421 1723 455
rect 1667 367 1723 421
rect 1753 599 1809 619
rect 1753 565 1764 599
rect 1798 565 1809 599
rect 1753 508 1809 565
rect 1753 474 1764 508
rect 1798 474 1809 508
rect 1753 413 1809 474
rect 1753 379 1764 413
rect 1798 379 1809 413
rect 1753 367 1809 379
rect 1839 607 1892 619
rect 1839 573 1850 607
rect 1884 573 1892 607
rect 1839 528 1892 573
rect 1839 494 1850 528
rect 1884 494 1892 528
rect 1839 455 1892 494
rect 1839 421 1850 455
rect 1884 421 1892 455
rect 1839 367 1892 421
<< ndiffc >>
rect 45 157 79 191
rect 131 139 165 173
rect 233 169 267 203
rect 339 169 373 203
rect 501 158 535 192
rect 615 169 649 203
rect 705 139 739 173
rect 809 169 843 203
rect 903 156 937 190
rect 1158 66 1192 100
rect 1248 169 1282 203
rect 1248 67 1282 101
rect 1334 141 1368 175
rect 1334 55 1368 89
rect 1420 169 1454 203
rect 1420 67 1454 101
rect 1506 141 1540 175
rect 1506 55 1540 89
rect 1592 152 1626 186
rect 1592 67 1626 101
rect 1678 89 1712 123
rect 1764 152 1798 186
rect 1764 67 1798 101
rect 1850 89 1884 123
<< pdiffc >>
rect 35 520 69 554
rect 35 452 69 486
rect 121 526 155 560
rect 1162 573 1196 607
rect 226 472 260 506
rect 370 495 404 529
rect 370 427 404 461
rect 529 505 563 539
rect 529 437 563 471
rect 615 503 649 537
rect 615 435 649 469
rect 712 495 746 529
rect 809 503 843 537
rect 809 435 843 469
rect 899 503 933 537
rect 899 435 933 469
rect 1162 490 1196 524
rect 1248 565 1282 599
rect 1248 474 1282 508
rect 1248 379 1282 413
rect 1334 573 1368 607
rect 1334 494 1368 528
rect 1334 421 1368 455
rect 1420 565 1454 599
rect 1420 474 1454 508
rect 1420 379 1454 413
rect 1506 573 1540 607
rect 1506 494 1540 528
rect 1506 421 1540 455
rect 1592 565 1626 599
rect 1592 474 1626 508
rect 1592 379 1626 413
rect 1678 573 1712 607
rect 1678 494 1712 528
rect 1678 421 1712 455
rect 1764 565 1798 599
rect 1764 474 1798 508
rect 1764 379 1798 413
rect 1850 573 1884 607
rect 1850 494 1884 528
rect 1850 421 1884 455
<< poly >>
rect 166 615 1050 645
rect 1207 619 1237 645
rect 1293 619 1323 645
rect 1379 619 1409 645
rect 1465 619 1495 645
rect 1551 619 1581 645
rect 1637 619 1667 645
rect 1723 619 1753 645
rect 1809 619 1839 645
rect 80 568 110 594
rect 166 568 196 615
rect 298 547 328 573
rect 415 547 445 615
rect 487 547 517 573
rect 574 547 604 573
rect 660 547 690 615
rect 768 547 798 573
rect 854 547 884 573
rect 948 547 978 573
rect 1020 547 1050 615
rect 1092 547 1122 573
rect 80 408 110 440
rect 52 392 120 408
rect 52 358 68 392
rect 102 358 120 392
rect 52 324 120 358
rect 52 290 68 324
rect 102 290 120 324
rect 166 366 196 440
rect 166 350 241 366
rect 166 316 191 350
rect 225 316 241 350
rect 166 300 241 316
rect 52 274 120 290
rect 90 215 120 274
rect 192 215 222 300
rect 298 215 328 419
rect 415 397 445 419
rect 378 367 445 397
rect 384 215 414 367
rect 487 319 517 419
rect 456 303 522 319
rect 456 269 472 303
rect 506 269 522 303
rect 456 253 522 269
rect 456 215 486 253
rect 574 215 604 419
rect 660 215 690 419
rect 768 387 798 419
rect 732 371 798 387
rect 732 337 748 371
rect 782 337 798 371
rect 732 321 798 337
rect 854 329 884 419
rect 768 215 798 321
rect 840 313 906 329
rect 840 279 856 313
rect 890 279 906 313
rect 840 263 906 279
rect 854 215 884 263
rect 948 215 978 419
rect 1020 215 1050 419
rect 1092 335 1122 419
rect 1092 319 1158 335
rect 1092 285 1108 319
rect 1142 285 1158 319
rect 1092 269 1158 285
rect 1207 329 1237 367
rect 1293 329 1323 367
rect 1379 329 1409 367
rect 1465 329 1495 367
rect 1207 313 1495 329
rect 1207 279 1223 313
rect 1257 279 1291 313
rect 1325 279 1359 313
rect 1393 279 1495 313
rect 1551 303 1581 367
rect 1637 303 1667 367
rect 1723 303 1753 367
rect 1809 303 1839 367
rect 1092 215 1122 269
rect 1207 263 1495 279
rect 1207 215 1237 263
rect 1293 215 1323 263
rect 1379 215 1409 263
rect 1465 215 1495 263
rect 1549 287 1839 303
rect 1549 253 1565 287
rect 1599 253 1633 287
rect 1667 253 1701 287
rect 1735 253 1769 287
rect 1803 253 1839 287
rect 1549 237 1839 253
rect 1551 215 1581 237
rect 1637 215 1667 237
rect 1723 215 1753 237
rect 1809 215 1839 237
rect 90 105 120 131
rect 192 105 222 131
rect 298 103 328 131
rect 384 105 414 131
rect 456 105 486 131
rect 270 87 336 103
rect 270 53 286 87
rect 320 57 336 87
rect 574 57 604 131
rect 660 105 690 131
rect 768 105 798 131
rect 854 105 884 131
rect 948 57 978 131
rect 1020 105 1050 131
rect 1092 105 1122 131
rect 320 53 978 57
rect 270 27 978 53
rect 1207 21 1237 47
rect 1293 21 1323 47
rect 1379 21 1409 47
rect 1465 21 1495 47
rect 1551 21 1581 47
rect 1637 21 1667 47
rect 1723 21 1753 47
rect 1809 21 1839 47
<< polycont >>
rect 68 358 102 392
rect 68 290 102 324
rect 191 316 225 350
rect 472 269 506 303
rect 748 337 782 371
rect 856 279 890 313
rect 1108 285 1142 319
rect 1223 279 1257 313
rect 1291 279 1325 313
rect 1359 279 1393 313
rect 1565 253 1599 287
rect 1633 253 1667 287
rect 1701 253 1735 287
rect 1769 253 1803 287
rect 286 53 320 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 19 554 69 570
rect 19 520 35 554
rect 105 560 171 649
rect 105 526 121 560
rect 155 526 171 560
rect 105 524 171 526
rect 300 579 493 615
rect 19 490 69 520
rect 222 506 264 522
rect 222 490 226 506
rect 19 486 226 490
rect 19 452 35 486
rect 69 472 226 486
rect 260 472 264 506
rect 69 456 264 472
rect 69 452 71 456
rect 19 436 71 452
rect 300 420 334 579
rect 105 402 334 420
rect 368 529 423 545
rect 368 495 370 529
rect 404 495 423 529
rect 368 461 423 495
rect 368 427 370 461
rect 404 427 423 461
rect 368 411 423 427
rect 52 392 334 402
rect 52 358 68 392
rect 102 386 334 392
rect 102 358 139 386
rect 52 324 139 358
rect 52 290 68 324
rect 102 290 139 324
rect 175 350 355 351
rect 175 316 191 350
rect 225 316 355 350
rect 175 310 355 316
rect 52 281 139 290
rect 389 276 423 411
rect 41 213 283 247
rect 41 191 81 213
rect 41 157 45 191
rect 79 157 81 191
rect 217 203 283 213
rect 41 141 81 157
rect 115 173 181 177
rect 115 139 131 173
rect 165 139 181 173
rect 217 169 233 203
rect 267 169 283 203
rect 217 162 283 169
rect 353 242 423 276
rect 459 383 493 579
rect 527 539 571 649
rect 527 505 529 539
rect 563 505 571 539
rect 527 471 571 505
rect 527 437 529 471
rect 563 437 571 471
rect 527 421 571 437
rect 605 537 655 553
rect 605 503 615 537
rect 649 503 655 537
rect 605 469 655 503
rect 696 529 762 649
rect 1146 607 1212 649
rect 1146 573 1162 607
rect 1196 573 1212 607
rect 696 495 712 529
rect 746 495 762 529
rect 696 487 762 495
rect 796 537 852 553
rect 796 503 809 537
rect 843 503 852 537
rect 605 435 615 469
rect 649 453 655 469
rect 796 469 852 503
rect 796 453 809 469
rect 649 435 809 453
rect 843 435 852 469
rect 605 419 852 435
rect 886 537 949 553
rect 886 503 899 537
rect 933 503 949 537
rect 886 469 949 503
rect 1146 524 1212 573
rect 1146 490 1162 524
rect 1196 490 1212 524
rect 1146 487 1212 490
rect 1246 599 1284 615
rect 1246 565 1248 599
rect 1282 565 1284 599
rect 1246 508 1284 565
rect 886 435 899 469
rect 933 453 949 469
rect 1246 474 1248 508
rect 1282 474 1284 508
rect 933 435 1212 453
rect 886 419 1212 435
rect 459 371 999 383
rect 459 337 748 371
rect 782 349 999 371
rect 782 337 798 349
rect 459 303 798 337
rect 965 335 999 349
rect 965 319 1144 335
rect 459 269 472 303
rect 506 277 798 303
rect 840 313 931 315
rect 840 279 856 313
rect 890 279 931 313
rect 840 277 931 279
rect 459 253 506 269
rect 895 276 931 277
rect 319 203 389 242
rect 611 209 847 243
rect 929 242 931 276
rect 965 285 1108 319
rect 1142 285 1144 319
rect 965 269 1144 285
rect 1178 313 1212 419
rect 1246 413 1284 474
rect 1318 607 1384 649
rect 1318 573 1334 607
rect 1368 573 1384 607
rect 1318 528 1384 573
rect 1318 494 1334 528
rect 1368 494 1384 528
rect 1318 455 1384 494
rect 1318 421 1334 455
rect 1368 421 1384 455
rect 1418 599 1456 615
rect 1418 565 1420 599
rect 1454 565 1456 599
rect 1418 508 1456 565
rect 1418 474 1420 508
rect 1454 474 1456 508
rect 1246 379 1248 413
rect 1282 385 1284 413
rect 1418 413 1456 474
rect 1490 607 1556 649
rect 1490 573 1506 607
rect 1540 573 1556 607
rect 1490 528 1556 573
rect 1490 494 1506 528
rect 1540 494 1556 528
rect 1490 455 1556 494
rect 1490 421 1506 455
rect 1540 421 1556 455
rect 1590 599 1628 615
rect 1590 565 1592 599
rect 1626 565 1628 599
rect 1590 508 1628 565
rect 1590 474 1592 508
rect 1626 474 1628 508
rect 1418 385 1420 413
rect 1282 379 1420 385
rect 1454 385 1456 413
rect 1590 413 1628 474
rect 1662 607 1728 649
rect 1662 573 1678 607
rect 1712 573 1728 607
rect 1662 528 1728 573
rect 1662 494 1678 528
rect 1712 494 1728 528
rect 1662 455 1728 494
rect 1662 421 1678 455
rect 1712 421 1728 455
rect 1762 599 1800 615
rect 1762 565 1764 599
rect 1798 565 1800 599
rect 1762 508 1800 565
rect 1762 474 1764 508
rect 1798 474 1800 508
rect 1454 379 1515 385
rect 1246 347 1515 379
rect 1590 379 1592 413
rect 1626 385 1628 413
rect 1762 413 1800 474
rect 1834 607 1900 649
rect 1834 573 1850 607
rect 1884 573 1900 607
rect 1834 528 1900 573
rect 1834 494 1850 528
rect 1884 494 1900 528
rect 1834 455 1900 494
rect 1834 421 1850 455
rect 1884 421 1900 455
rect 1762 385 1764 413
rect 1626 379 1764 385
rect 1798 385 1800 413
rect 1798 379 1902 385
rect 1590 351 1902 379
rect 1178 279 1223 313
rect 1257 279 1291 313
rect 1325 279 1359 313
rect 1393 279 1409 313
rect 895 240 931 242
rect 319 169 339 203
rect 373 169 389 203
rect 319 162 389 169
rect 485 192 551 208
rect 115 17 181 139
rect 485 158 501 192
rect 535 158 551 192
rect 215 87 449 128
rect 215 53 286 87
rect 320 53 449 87
rect 485 17 551 158
rect 611 203 653 209
rect 611 169 615 203
rect 649 169 653 203
rect 805 203 847 209
rect 1178 206 1212 279
rect 1443 245 1515 347
rect 611 153 653 169
rect 689 139 705 173
rect 739 139 755 173
rect 805 169 809 203
rect 843 169 847 203
rect 805 153 847 169
rect 899 190 1212 206
rect 899 156 903 190
rect 937 156 1212 190
rect 899 140 1212 156
rect 1246 209 1515 245
rect 1549 287 1819 303
rect 1549 253 1565 287
rect 1599 276 1633 287
rect 1601 253 1633 276
rect 1667 253 1701 287
rect 1735 253 1769 287
rect 1803 253 1819 287
rect 1549 242 1567 253
rect 1601 242 1819 253
rect 1549 236 1819 242
rect 1246 203 1284 209
rect 1246 169 1248 203
rect 1282 169 1284 203
rect 1418 203 1456 209
rect 689 17 755 139
rect 1142 100 1208 106
rect 1142 66 1158 100
rect 1192 66 1208 100
rect 1142 17 1208 66
rect 1246 101 1284 169
rect 1246 67 1248 101
rect 1282 67 1284 101
rect 1246 51 1284 67
rect 1318 141 1334 175
rect 1368 141 1384 175
rect 1318 89 1384 141
rect 1318 55 1334 89
rect 1368 55 1384 89
rect 1318 17 1384 55
rect 1418 169 1420 203
rect 1454 169 1456 203
rect 1853 202 1902 351
rect 1590 186 1902 202
rect 1418 101 1456 169
rect 1418 67 1420 101
rect 1454 67 1456 101
rect 1418 51 1456 67
rect 1490 141 1506 175
rect 1540 141 1556 175
rect 1490 89 1556 141
rect 1490 55 1506 89
rect 1540 55 1556 89
rect 1490 17 1556 55
rect 1590 152 1592 186
rect 1626 168 1764 186
rect 1626 152 1628 168
rect 1590 101 1628 152
rect 1762 152 1764 168
rect 1798 168 1902 186
rect 1798 152 1800 168
rect 1590 67 1592 101
rect 1626 67 1628 101
rect 1590 51 1628 67
rect 1662 123 1728 134
rect 1662 89 1678 123
rect 1712 89 1728 123
rect 1662 17 1728 89
rect 1762 101 1800 152
rect 1762 67 1764 101
rect 1798 67 1800 101
rect 1762 51 1800 67
rect 1834 123 1900 134
rect 1834 89 1850 123
rect 1884 89 1900 123
rect 1834 17 1900 89
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 319 242 353 276
rect 895 242 929 276
rect 1567 253 1599 276
rect 1599 253 1601 276
rect 1567 242 1601 253
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 307 276 365 282
rect 307 242 319 276
rect 353 273 365 276
rect 883 276 941 282
rect 883 273 895 276
rect 353 245 895 273
rect 353 242 365 245
rect 307 236 365 242
rect 883 242 895 245
rect 929 273 941 276
rect 1555 276 1613 282
rect 1555 273 1567 276
rect 929 245 1567 273
rect 929 242 941 245
rect 883 236 941 242
rect 1555 242 1567 245
rect 1601 242 1613 276
rect 1555 236 1613 242
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fa_4
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1855 168 1889 202 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2472800
string GDS_START 2457840
<< end >>
