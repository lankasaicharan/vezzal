magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 4 49 1119 259
rect 0 0 1152 49
<< scnmos >>
rect 83 65 113 233
rect 169 65 199 233
rect 255 65 285 233
rect 357 65 387 233
rect 459 65 489 233
rect 545 65 575 233
rect 752 65 782 233
rect 838 65 868 233
rect 924 65 954 233
rect 1010 65 1040 233
<< scpmoshvt >>
rect 83 367 113 619
rect 169 367 199 619
rect 255 367 285 619
rect 373 367 403 619
rect 459 367 489 619
rect 545 367 575 619
rect 752 367 782 619
rect 838 367 868 619
rect 924 367 954 619
rect 1010 367 1040 619
<< ndiff >>
rect 30 221 83 233
rect 30 187 38 221
rect 72 187 83 221
rect 30 111 83 187
rect 30 77 38 111
rect 72 77 83 111
rect 30 65 83 77
rect 113 221 169 233
rect 113 187 124 221
rect 158 187 169 221
rect 113 111 169 187
rect 113 77 124 111
rect 158 77 169 111
rect 113 65 169 77
rect 199 225 255 233
rect 199 191 210 225
rect 244 191 255 225
rect 199 157 255 191
rect 199 123 210 157
rect 244 123 255 157
rect 199 65 255 123
rect 285 175 357 233
rect 285 141 312 175
rect 346 141 357 175
rect 285 107 357 141
rect 285 73 312 107
rect 346 73 357 107
rect 285 65 357 73
rect 387 175 459 233
rect 387 141 414 175
rect 448 141 459 175
rect 387 107 459 141
rect 387 73 414 107
rect 448 73 459 107
rect 387 65 459 73
rect 489 212 545 233
rect 489 178 500 212
rect 534 178 545 212
rect 489 107 545 178
rect 489 73 500 107
rect 534 73 545 107
rect 489 65 545 73
rect 575 175 752 233
rect 575 141 600 175
rect 634 141 707 175
rect 741 141 752 175
rect 575 107 752 141
rect 575 73 600 107
rect 634 73 707 107
rect 741 73 752 107
rect 575 65 752 73
rect 782 221 838 233
rect 782 187 793 221
rect 827 187 838 221
rect 782 111 838 187
rect 782 77 793 111
rect 827 77 838 111
rect 782 65 838 77
rect 868 175 924 233
rect 868 141 879 175
rect 913 141 924 175
rect 868 107 924 141
rect 868 73 879 107
rect 913 73 924 107
rect 868 65 924 73
rect 954 221 1010 233
rect 954 187 965 221
rect 999 187 1010 221
rect 954 111 1010 187
rect 954 77 965 111
rect 999 77 1010 111
rect 954 65 1010 77
rect 1040 208 1093 233
rect 1040 174 1051 208
rect 1085 174 1093 208
rect 1040 111 1093 174
rect 1040 77 1051 111
rect 1085 77 1093 111
rect 1040 65 1093 77
<< pdiff >>
rect 30 599 83 619
rect 30 565 38 599
rect 72 565 83 599
rect 30 511 83 565
rect 30 477 38 511
rect 72 477 83 511
rect 30 413 83 477
rect 30 379 38 413
rect 72 379 83 413
rect 30 367 83 379
rect 113 572 169 619
rect 113 538 124 572
rect 158 538 169 572
rect 113 367 169 538
rect 199 599 255 619
rect 199 565 210 599
rect 244 565 255 599
rect 199 508 255 565
rect 199 474 210 508
rect 244 474 255 508
rect 199 367 255 474
rect 285 572 373 619
rect 285 538 314 572
rect 348 538 373 572
rect 285 367 373 538
rect 403 599 459 619
rect 403 565 414 599
rect 448 565 459 599
rect 403 505 459 565
rect 403 471 414 505
rect 448 471 459 505
rect 403 415 459 471
rect 403 381 414 415
rect 448 381 459 415
rect 403 367 459 381
rect 489 547 545 619
rect 489 513 500 547
rect 534 513 545 547
rect 489 479 545 513
rect 489 445 500 479
rect 534 445 545 479
rect 489 411 545 445
rect 489 377 500 411
rect 534 377 545 411
rect 489 367 545 377
rect 575 599 628 619
rect 575 565 586 599
rect 620 565 628 599
rect 575 505 628 565
rect 575 471 586 505
rect 620 471 628 505
rect 575 415 628 471
rect 575 381 586 415
rect 620 381 628 415
rect 575 367 628 381
rect 699 599 752 619
rect 699 565 707 599
rect 741 565 752 599
rect 699 529 752 565
rect 699 495 707 529
rect 741 495 752 529
rect 699 459 752 495
rect 699 425 707 459
rect 741 425 752 459
rect 699 367 752 425
rect 782 607 838 619
rect 782 573 793 607
rect 827 573 838 607
rect 782 515 838 573
rect 782 481 793 515
rect 827 481 838 515
rect 782 367 838 481
rect 868 599 924 619
rect 868 565 879 599
rect 913 565 924 599
rect 868 529 924 565
rect 868 495 879 529
rect 913 495 924 529
rect 868 459 924 495
rect 868 425 879 459
rect 913 425 924 459
rect 868 367 924 425
rect 954 531 1010 619
rect 954 497 965 531
rect 999 497 1010 531
rect 954 413 1010 497
rect 954 379 965 413
rect 999 379 1010 413
rect 954 367 1010 379
rect 1040 599 1093 619
rect 1040 565 1051 599
rect 1085 565 1093 599
rect 1040 514 1093 565
rect 1040 480 1051 514
rect 1085 480 1093 514
rect 1040 434 1093 480
rect 1040 400 1051 434
rect 1085 400 1093 434
rect 1040 367 1093 400
<< ndiffc >>
rect 38 187 72 221
rect 38 77 72 111
rect 124 187 158 221
rect 124 77 158 111
rect 210 191 244 225
rect 210 123 244 157
rect 312 141 346 175
rect 312 73 346 107
rect 414 141 448 175
rect 414 73 448 107
rect 500 178 534 212
rect 500 73 534 107
rect 600 141 634 175
rect 707 141 741 175
rect 600 73 634 107
rect 707 73 741 107
rect 793 187 827 221
rect 793 77 827 111
rect 879 141 913 175
rect 879 73 913 107
rect 965 187 999 221
rect 965 77 999 111
rect 1051 174 1085 208
rect 1051 77 1085 111
<< pdiffc >>
rect 38 565 72 599
rect 38 477 72 511
rect 38 379 72 413
rect 124 538 158 572
rect 210 565 244 599
rect 210 474 244 508
rect 314 538 348 572
rect 414 565 448 599
rect 414 471 448 505
rect 414 381 448 415
rect 500 513 534 547
rect 500 445 534 479
rect 500 377 534 411
rect 586 565 620 599
rect 586 471 620 505
rect 586 381 620 415
rect 707 565 741 599
rect 707 495 741 529
rect 707 425 741 459
rect 793 573 827 607
rect 793 481 827 515
rect 879 565 913 599
rect 879 495 913 529
rect 879 425 913 459
rect 965 497 999 531
rect 965 379 999 413
rect 1051 565 1085 599
rect 1051 480 1085 514
rect 1051 400 1085 434
<< poly >>
rect 83 619 113 645
rect 169 619 199 645
rect 255 619 285 645
rect 373 619 403 645
rect 459 619 489 645
rect 545 619 575 645
rect 752 619 782 645
rect 838 619 868 645
rect 924 619 954 645
rect 1010 619 1040 645
rect 83 325 113 367
rect 47 309 113 325
rect 47 275 63 309
rect 97 275 113 309
rect 47 259 113 275
rect 83 233 113 259
rect 169 335 199 367
rect 255 335 285 367
rect 373 335 403 367
rect 169 319 285 335
rect 169 285 198 319
rect 232 285 285 319
rect 169 269 285 285
rect 337 319 403 335
rect 337 285 353 319
rect 387 285 403 319
rect 337 269 403 285
rect 459 315 489 367
rect 545 315 575 367
rect 752 335 782 367
rect 838 335 868 367
rect 459 285 575 315
rect 617 305 683 321
rect 617 285 633 305
rect 169 233 199 269
rect 255 233 285 269
rect 357 233 387 269
rect 459 233 489 285
rect 545 271 633 285
rect 667 271 683 305
rect 545 255 683 271
rect 725 319 868 335
rect 725 285 741 319
rect 775 285 868 319
rect 725 269 868 285
rect 545 233 575 255
rect 752 233 782 269
rect 838 233 868 269
rect 924 285 954 367
rect 1010 321 1040 367
rect 1010 305 1085 321
rect 1010 285 1035 305
rect 924 271 1035 285
rect 1069 271 1085 305
rect 924 255 1085 271
rect 924 233 954 255
rect 1010 233 1040 255
rect 83 39 113 65
rect 169 39 199 65
rect 255 39 285 65
rect 357 39 387 65
rect 459 39 489 65
rect 545 39 575 65
rect 752 39 782 65
rect 838 39 868 65
rect 924 39 954 65
rect 1010 39 1040 65
<< polycont >>
rect 63 275 97 309
rect 198 285 232 319
rect 353 285 387 319
rect 633 271 667 305
rect 741 285 775 319
rect 1035 271 1069 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 22 599 74 615
rect 22 565 38 599
rect 72 565 74 599
rect 22 511 74 565
rect 108 572 174 649
rect 108 538 124 572
rect 158 538 174 572
rect 108 526 174 538
rect 208 599 248 615
rect 208 565 210 599
rect 244 565 248 599
rect 22 477 38 511
rect 72 492 74 511
rect 208 508 248 565
rect 298 572 364 649
rect 298 538 314 572
rect 348 538 364 572
rect 298 526 364 538
rect 410 599 636 615
rect 410 565 414 599
rect 448 581 586 599
rect 448 565 450 581
rect 208 492 210 508
rect 72 477 210 492
rect 22 474 210 477
rect 244 492 248 508
rect 410 505 450 565
rect 584 565 586 581
rect 620 565 636 599
rect 410 492 414 505
rect 244 474 414 492
rect 22 471 414 474
rect 448 471 450 505
rect 22 458 450 471
rect 22 413 76 458
rect 22 379 38 413
rect 72 379 76 413
rect 22 363 76 379
rect 110 384 376 424
rect 110 325 146 384
rect 47 309 146 325
rect 47 275 63 309
rect 97 275 146 309
rect 182 319 285 350
rect 182 285 198 319
rect 232 285 285 319
rect 319 331 376 384
rect 410 415 450 458
rect 410 381 414 415
rect 448 381 450 415
rect 410 365 450 381
rect 484 513 500 547
rect 534 513 550 547
rect 484 479 550 513
rect 484 445 500 479
rect 534 445 550 479
rect 484 411 550 445
rect 484 377 500 411
rect 534 377 550 411
rect 484 361 550 377
rect 584 505 636 565
rect 584 471 586 505
rect 620 471 636 505
rect 584 415 636 471
rect 584 381 586 415
rect 620 381 636 415
rect 691 599 743 615
rect 691 565 707 599
rect 741 565 743 599
rect 691 529 743 565
rect 691 495 707 529
rect 741 495 743 529
rect 691 459 743 495
rect 777 607 843 649
rect 777 573 793 607
rect 827 573 843 607
rect 777 515 843 573
rect 777 481 793 515
rect 827 481 843 515
rect 777 477 843 481
rect 877 599 1101 615
rect 877 565 879 599
rect 913 581 1051 599
rect 913 565 923 581
rect 877 529 923 565
rect 1035 565 1051 581
rect 1085 565 1101 599
rect 877 495 879 529
rect 913 495 923 529
rect 691 425 707 459
rect 741 443 743 459
rect 877 459 923 495
rect 877 443 879 459
rect 741 425 879 443
rect 913 425 923 459
rect 691 409 923 425
rect 957 531 1001 547
rect 957 497 965 531
rect 999 497 1001 531
rect 957 413 1001 497
rect 584 365 636 381
rect 957 379 965 413
rect 999 379 1001 413
rect 1035 514 1101 565
rect 1035 480 1051 514
rect 1085 480 1101 514
rect 1035 434 1101 480
rect 1035 400 1051 434
rect 1085 400 1101 434
rect 1035 384 1101 400
rect 957 375 1001 379
rect 319 319 403 331
rect 319 285 353 319
rect 387 285 403 319
rect 500 249 550 361
rect 22 221 81 237
rect 22 187 38 221
rect 72 187 81 221
rect 22 111 81 187
rect 22 77 38 111
rect 72 77 81 111
rect 22 17 81 77
rect 115 221 160 237
rect 115 187 124 221
rect 158 187 160 221
rect 115 111 160 187
rect 194 225 550 249
rect 194 191 210 225
rect 244 215 550 225
rect 617 305 667 321
rect 617 271 633 305
rect 701 319 791 375
rect 701 285 741 319
rect 775 285 791 319
rect 701 283 791 285
rect 827 341 1001 375
rect 617 249 667 271
rect 827 249 861 341
rect 1035 305 1135 350
rect 1069 271 1135 305
rect 617 221 999 249
rect 1035 242 1135 271
rect 617 215 793 221
rect 244 191 260 215
rect 194 157 260 191
rect 498 212 550 215
rect 194 123 210 157
rect 244 123 260 157
rect 194 121 260 123
rect 294 175 364 181
rect 294 141 312 175
rect 346 141 364 175
rect 115 77 124 111
rect 158 87 160 111
rect 294 107 364 141
rect 294 87 312 107
rect 158 77 312 87
rect 115 73 312 77
rect 346 73 364 107
rect 115 53 364 73
rect 398 175 464 179
rect 398 141 414 175
rect 448 141 464 175
rect 398 107 464 141
rect 398 73 414 107
rect 448 73 464 107
rect 398 17 464 73
rect 498 178 500 212
rect 534 178 550 212
rect 791 187 793 215
rect 827 215 965 221
rect 827 187 829 215
rect 498 107 550 178
rect 498 73 500 107
rect 534 73 550 107
rect 498 57 550 73
rect 584 175 757 179
rect 584 141 600 175
rect 634 141 707 175
rect 741 141 757 175
rect 584 107 757 141
rect 584 73 600 107
rect 634 73 707 107
rect 741 73 757 107
rect 584 17 757 73
rect 791 111 829 187
rect 791 77 793 111
rect 827 77 829 111
rect 791 61 829 77
rect 863 175 929 179
rect 863 141 879 175
rect 913 141 929 175
rect 863 107 929 141
rect 863 73 879 107
rect 913 73 929 107
rect 863 17 929 73
rect 965 111 999 187
rect 965 61 999 77
rect 1035 174 1051 208
rect 1085 174 1101 208
rect 1035 111 1101 174
rect 1035 77 1051 111
rect 1085 77 1101 111
rect 1035 17 1101 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2bb2oi_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3088054
string GDS_START 3077874
<< end >>
