magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 45 49 629 241
rect 0 0 672 49
<< scnmos >>
rect 124 131 154 215
rect 232 47 262 215
rect 304 47 334 215
rect 412 47 442 215
rect 520 47 550 215
<< scpmoshvt >>
rect 124 367 154 451
rect 232 367 262 619
rect 318 367 348 619
rect 434 367 464 619
rect 520 367 550 619
<< ndiff >>
rect 71 187 124 215
rect 71 153 79 187
rect 113 153 124 187
rect 71 131 124 153
rect 154 196 232 215
rect 154 162 175 196
rect 209 162 232 196
rect 154 131 232 162
rect 176 93 232 131
rect 176 59 184 93
rect 218 59 232 93
rect 176 47 232 59
rect 262 47 304 215
rect 334 47 412 215
rect 442 47 520 215
rect 550 203 603 215
rect 550 169 561 203
rect 595 169 603 203
rect 550 101 603 169
rect 550 67 561 101
rect 595 67 603 101
rect 550 47 603 67
<< pdiff >>
rect 179 607 232 619
rect 179 573 187 607
rect 221 573 232 607
rect 179 526 232 573
rect 179 492 187 526
rect 221 492 232 526
rect 179 451 232 492
rect 71 424 124 451
rect 71 390 79 424
rect 113 390 124 424
rect 71 367 124 390
rect 154 441 232 451
rect 154 407 165 441
rect 199 407 232 441
rect 154 367 232 407
rect 262 599 318 619
rect 262 565 273 599
rect 307 565 318 599
rect 262 526 318 565
rect 262 492 273 526
rect 307 492 318 526
rect 262 457 318 492
rect 262 423 273 457
rect 307 423 318 457
rect 262 367 318 423
rect 348 607 434 619
rect 348 573 373 607
rect 407 573 434 607
rect 348 513 434 573
rect 348 479 373 513
rect 407 479 434 513
rect 348 367 434 479
rect 464 599 520 619
rect 464 565 475 599
rect 509 565 520 599
rect 464 525 520 565
rect 464 491 475 525
rect 509 491 520 525
rect 464 441 520 491
rect 464 407 475 441
rect 509 407 520 441
rect 464 367 520 407
rect 550 607 603 619
rect 550 573 561 607
rect 595 573 603 607
rect 550 514 603 573
rect 550 480 561 514
rect 595 480 603 514
rect 550 367 603 480
<< ndiffc >>
rect 79 153 113 187
rect 175 162 209 196
rect 184 59 218 93
rect 561 169 595 203
rect 561 67 595 101
<< pdiffc >>
rect 187 573 221 607
rect 187 492 221 526
rect 79 390 113 424
rect 165 407 199 441
rect 273 565 307 599
rect 273 492 307 526
rect 273 423 307 457
rect 373 573 407 607
rect 373 479 407 513
rect 475 565 509 599
rect 475 491 509 525
rect 475 407 509 441
rect 561 573 595 607
rect 561 480 595 514
<< poly >>
rect 232 619 262 645
rect 318 619 348 645
rect 434 619 464 645
rect 520 619 550 645
rect 124 451 154 477
rect 124 303 154 367
rect 232 303 262 367
rect 318 303 348 367
rect 434 303 464 367
rect 520 335 550 367
rect 520 319 586 335
rect 88 287 154 303
rect 88 253 104 287
rect 138 253 154 287
rect 88 237 154 253
rect 196 287 262 303
rect 196 253 212 287
rect 246 253 262 287
rect 196 237 262 253
rect 124 215 154 237
rect 232 215 262 237
rect 304 287 370 303
rect 304 253 320 287
rect 354 253 370 287
rect 304 237 370 253
rect 412 287 478 303
rect 412 253 428 287
rect 462 253 478 287
rect 412 237 478 253
rect 520 285 536 319
rect 570 285 586 319
rect 520 269 586 285
rect 304 215 334 237
rect 412 215 442 237
rect 520 215 550 269
rect 124 105 154 131
rect 232 21 262 47
rect 304 21 334 47
rect 412 21 442 47
rect 520 21 550 47
<< polycont >>
rect 104 253 138 287
rect 212 253 246 287
rect 320 253 354 287
rect 428 253 462 287
rect 536 285 570 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 149 607 232 649
rect 149 573 187 607
rect 221 573 232 607
rect 149 526 232 573
rect 149 492 187 526
rect 221 492 232 526
rect 149 441 232 492
rect 17 424 115 440
rect 17 390 79 424
rect 113 390 115 424
rect 149 407 165 441
rect 199 407 232 441
rect 266 599 323 615
rect 266 565 273 599
rect 307 565 323 599
rect 266 526 323 565
rect 266 492 273 526
rect 307 492 323 526
rect 266 457 323 492
rect 357 607 423 649
rect 357 573 373 607
rect 407 573 423 607
rect 357 513 423 573
rect 357 479 373 513
rect 407 479 423 513
rect 357 475 423 479
rect 459 599 511 615
rect 459 565 475 599
rect 509 565 511 599
rect 459 525 511 565
rect 459 491 475 525
rect 509 491 511 525
rect 266 423 273 457
rect 307 441 323 457
rect 459 441 511 491
rect 545 607 611 649
rect 545 573 561 607
rect 595 573 611 607
rect 545 514 611 573
rect 545 480 561 514
rect 595 480 611 514
rect 545 475 611 480
rect 307 423 475 441
rect 266 407 475 423
rect 509 407 655 441
rect 17 373 115 390
rect 17 339 570 373
rect 17 203 70 339
rect 520 319 570 339
rect 104 287 178 303
rect 138 253 178 287
rect 104 237 178 253
rect 212 287 272 303
rect 246 253 272 287
rect 212 237 272 253
rect 306 287 365 303
rect 306 253 320 287
rect 354 253 365 287
rect 17 187 125 203
rect 17 153 79 187
rect 113 153 125 187
rect 17 137 125 153
rect 159 196 225 203
rect 159 162 175 196
rect 209 162 225 196
rect 159 93 225 162
rect 159 59 184 93
rect 218 59 225 93
rect 306 74 365 253
rect 399 287 478 303
rect 399 253 428 287
rect 462 253 478 287
rect 520 285 536 319
rect 520 269 570 285
rect 399 74 478 253
rect 604 219 655 407
rect 545 203 655 219
rect 545 169 561 203
rect 595 169 655 203
rect 545 101 655 169
rect 159 17 225 59
rect 545 67 561 101
rect 595 67 655 101
rect 545 51 655 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4b_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 768656
string GDS_START 761898
<< end >>
