magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
<< pwell >>
rect 21 49 1243 259
rect 0 0 1248 49
<< scnmos >>
rect 119 65 149 233
rect 205 65 235 233
rect 323 65 353 233
rect 455 65 485 233
rect 580 65 610 233
rect 666 65 696 233
rect 784 65 814 233
rect 870 65 900 233
rect 961 65 991 233
rect 1120 65 1150 233
<< scpmoshvt >>
rect 119 367 149 619
rect 205 367 235 619
rect 291 367 321 619
rect 395 367 425 619
rect 585 367 615 619
rect 671 367 701 619
rect 757 367 787 619
rect 875 367 905 619
rect 961 367 991 619
rect 1079 367 1109 619
<< ndiff >>
rect 47 89 119 233
rect 47 55 55 89
rect 89 65 119 89
rect 149 225 205 233
rect 149 191 160 225
rect 194 191 205 225
rect 149 65 205 191
rect 235 89 323 233
rect 235 65 262 89
rect 89 55 97 65
rect 47 39 97 55
rect 250 55 262 65
rect 296 65 323 89
rect 353 225 455 233
rect 353 191 387 225
rect 421 191 455 225
rect 353 65 455 191
rect 485 89 580 233
rect 485 65 512 89
rect 296 55 308 65
rect 250 43 308 55
rect 500 55 512 65
rect 546 65 580 89
rect 610 225 666 233
rect 610 191 621 225
rect 655 191 666 225
rect 610 65 666 191
rect 696 89 784 233
rect 696 65 723 89
rect 546 55 558 65
rect 500 43 558 55
rect 711 55 723 65
rect 757 65 784 89
rect 814 221 870 233
rect 814 187 825 221
rect 859 187 870 221
rect 814 107 870 187
rect 814 73 825 107
rect 859 73 870 107
rect 814 65 870 73
rect 900 225 961 233
rect 900 191 911 225
rect 945 191 961 225
rect 900 153 961 191
rect 900 119 911 153
rect 945 119 961 153
rect 900 65 961 119
rect 991 181 1120 233
rect 991 147 1075 181
rect 1109 147 1120 181
rect 991 112 1120 147
rect 991 78 1002 112
rect 1036 78 1075 112
rect 1109 78 1120 112
rect 991 65 1120 78
rect 1150 181 1217 233
rect 1150 147 1175 181
rect 1209 147 1217 181
rect 1150 111 1217 147
rect 1150 77 1175 111
rect 1209 77 1217 111
rect 1150 65 1217 77
rect 757 55 769 65
rect 711 43 769 55
<< pdiff >>
rect 802 622 860 638
rect 802 619 814 622
rect 59 607 119 619
rect 59 573 74 607
rect 108 573 119 607
rect 59 508 119 573
rect 59 474 74 508
rect 108 474 119 508
rect 59 414 119 474
rect 59 380 67 414
rect 101 380 119 414
rect 59 367 119 380
rect 149 599 205 619
rect 149 565 160 599
rect 194 565 205 599
rect 149 508 205 565
rect 149 474 160 508
rect 194 474 205 508
rect 149 367 205 474
rect 235 510 291 619
rect 235 476 246 510
rect 280 476 291 510
rect 235 367 291 476
rect 321 568 395 619
rect 321 534 336 568
rect 370 534 395 568
rect 321 367 395 534
rect 425 568 478 619
rect 425 534 436 568
rect 470 534 478 568
rect 425 367 478 534
rect 532 576 585 619
rect 532 542 540 576
rect 574 542 585 576
rect 532 367 585 542
rect 615 486 671 619
rect 615 452 626 486
rect 660 452 671 486
rect 615 418 671 452
rect 615 384 626 418
rect 660 384 671 418
rect 615 367 671 384
rect 701 574 757 619
rect 701 540 712 574
rect 746 540 757 574
rect 701 367 757 540
rect 787 588 814 619
rect 848 619 860 622
rect 1006 622 1064 638
rect 1006 619 1018 622
rect 848 588 875 619
rect 787 367 875 588
rect 905 554 961 619
rect 905 520 916 554
rect 950 520 961 554
rect 905 367 961 520
rect 991 588 1018 619
rect 1052 619 1064 622
rect 1052 588 1079 619
rect 991 367 1079 588
rect 1109 554 1162 619
rect 1109 520 1120 554
rect 1154 520 1162 554
rect 1109 367 1162 520
<< ndiffc >>
rect 55 55 89 89
rect 160 191 194 225
rect 262 55 296 89
rect 387 191 421 225
rect 512 55 546 89
rect 621 191 655 225
rect 723 55 757 89
rect 825 187 859 221
rect 825 73 859 107
rect 911 191 945 225
rect 911 119 945 153
rect 1075 147 1109 181
rect 1002 78 1036 112
rect 1075 78 1109 112
rect 1175 147 1209 181
rect 1175 77 1209 111
<< pdiffc >>
rect 74 573 108 607
rect 74 474 108 508
rect 67 380 101 414
rect 160 565 194 599
rect 160 474 194 508
rect 246 476 280 510
rect 336 534 370 568
rect 436 534 470 568
rect 540 542 574 576
rect 626 452 660 486
rect 626 384 660 418
rect 712 540 746 574
rect 814 588 848 622
rect 916 520 950 554
rect 1018 588 1052 622
rect 1120 520 1154 554
<< poly >>
rect 119 619 149 645
rect 205 619 235 645
rect 291 619 321 645
rect 395 619 425 645
rect 585 619 615 645
rect 671 619 701 645
rect 757 619 787 645
rect 875 619 905 645
rect 961 619 991 645
rect 1079 619 1109 645
rect 119 321 149 367
rect 83 305 149 321
rect 83 271 99 305
rect 133 271 149 305
rect 83 255 149 271
rect 119 233 149 255
rect 205 335 235 367
rect 291 335 321 367
rect 395 335 425 367
rect 205 319 353 335
rect 205 285 249 319
rect 283 285 353 319
rect 205 269 353 285
rect 395 319 485 335
rect 585 321 615 367
rect 671 321 701 367
rect 757 321 787 367
rect 875 335 905 367
rect 961 335 991 367
rect 395 285 417 319
rect 451 285 485 319
rect 395 269 485 285
rect 205 233 235 269
rect 323 233 353 269
rect 455 233 485 269
rect 540 305 701 321
rect 540 271 556 305
rect 590 271 701 305
rect 540 255 701 271
rect 748 305 814 321
rect 748 271 764 305
rect 798 271 814 305
rect 748 255 814 271
rect 857 319 991 335
rect 857 285 873 319
rect 907 285 941 319
rect 975 285 991 319
rect 857 269 991 285
rect 1079 335 1109 367
rect 1079 319 1150 335
rect 1079 285 1095 319
rect 1129 285 1150 319
rect 1079 269 1150 285
rect 580 233 610 255
rect 666 233 696 255
rect 784 233 814 255
rect 870 233 900 269
rect 961 233 991 269
rect 1120 233 1150 269
rect 119 39 149 65
rect 205 39 235 65
rect 323 39 353 65
rect 455 39 485 65
rect 580 39 610 65
rect 666 39 696 65
rect 784 39 814 65
rect 870 39 900 65
rect 961 39 991 65
rect 1120 39 1150 65
<< polycont >>
rect 99 271 133 305
rect 249 285 283 319
rect 417 285 451 319
rect 556 271 590 305
rect 764 271 798 305
rect 873 285 907 319
rect 941 285 975 319
rect 1095 285 1129 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 51 607 124 649
rect 51 573 74 607
rect 108 573 124 607
rect 51 508 124 573
rect 51 474 74 508
rect 108 474 124 508
rect 51 458 124 474
rect 158 599 386 615
rect 158 565 160 599
rect 194 568 386 599
rect 194 565 336 568
rect 158 560 336 565
rect 158 508 204 560
rect 320 534 336 560
rect 370 534 386 568
rect 320 526 386 534
rect 420 568 486 649
rect 798 622 864 649
rect 420 534 436 568
rect 470 534 486 568
rect 420 526 486 534
rect 524 576 762 615
rect 798 588 814 622
rect 848 588 864 622
rect 1002 622 1068 649
rect 1002 588 1018 622
rect 1052 588 1068 622
rect 524 542 540 576
rect 574 574 762 576
rect 574 542 712 574
rect 524 540 712 542
rect 746 554 762 574
rect 746 540 916 554
rect 524 526 916 540
rect 158 474 160 508
rect 194 474 204 508
rect 158 458 204 474
rect 238 510 286 526
rect 593 520 916 526
rect 950 520 1120 554
rect 1154 520 1170 554
rect 238 476 246 510
rect 280 492 286 510
rect 280 476 540 492
rect 238 458 540 476
rect 51 414 101 458
rect 51 380 67 414
rect 51 364 101 380
rect 135 390 467 424
rect 135 321 169 390
rect 74 305 169 321
rect 74 271 99 305
rect 133 271 169 305
rect 74 269 169 271
rect 203 350 285 356
rect 203 316 223 350
rect 257 319 285 350
rect 203 285 249 316
rect 283 285 285 319
rect 203 269 285 285
rect 319 319 467 390
rect 319 285 417 319
rect 451 285 467 319
rect 319 269 467 285
rect 506 321 540 458
rect 610 452 626 486
rect 660 452 1231 486
rect 610 418 676 452
rect 610 384 626 418
rect 660 384 676 418
rect 610 368 676 384
rect 506 305 606 321
rect 506 271 556 305
rect 590 271 606 305
rect 74 157 108 269
rect 506 266 606 271
rect 506 235 540 266
rect 144 225 540 235
rect 642 232 676 368
rect 780 384 1145 418
rect 780 321 814 384
rect 144 191 160 225
rect 194 191 387 225
rect 421 191 540 225
rect 605 225 676 232
rect 605 191 621 225
rect 655 191 676 225
rect 748 305 814 321
rect 748 271 764 305
rect 798 271 814 305
rect 857 319 895 350
rect 929 319 991 350
rect 857 285 873 319
rect 929 316 941 319
rect 907 285 941 316
rect 975 285 991 319
rect 857 283 991 285
rect 1079 319 1145 384
rect 1079 285 1095 319
rect 1129 285 1145 319
rect 1079 283 1145 285
rect 748 157 784 271
rect 1179 249 1231 452
rect 74 123 784 157
rect 818 221 861 237
rect 818 187 825 221
rect 859 187 861 221
rect 818 107 861 187
rect 895 225 1231 249
rect 895 191 911 225
rect 945 215 1231 225
rect 945 191 1025 215
rect 895 162 1025 191
rect 895 153 961 162
rect 895 119 911 153
rect 945 119 961 153
rect 1059 147 1075 181
rect 1109 147 1125 181
rect 1059 128 1125 147
rect 39 55 55 89
rect 89 55 105 89
rect 39 17 105 55
rect 246 55 262 89
rect 296 55 312 89
rect 246 17 312 55
rect 496 55 512 89
rect 546 55 562 89
rect 496 17 562 55
rect 707 55 723 89
rect 757 55 773 89
rect 707 17 773 55
rect 818 73 825 107
rect 859 85 861 107
rect 995 112 1125 128
rect 995 85 1002 112
rect 859 78 1002 85
rect 1036 78 1075 112
rect 1109 78 1125 112
rect 859 73 1125 78
rect 818 51 1125 73
rect 1159 147 1175 181
rect 1209 147 1225 181
rect 1159 111 1225 147
rect 1159 77 1175 111
rect 1209 77 1225 111
rect 1159 17 1225 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 223 319 257 350
rect 223 316 249 319
rect 249 316 257 319
rect 895 319 929 350
rect 895 316 907 319
rect 907 316 929 319
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 211 350 269 356
rect 211 316 223 350
rect 257 347 269 350
rect 883 350 941 356
rect 883 347 895 350
rect 257 319 895 347
rect 257 316 269 319
rect 211 310 269 316
rect 883 316 895 319
rect 929 316 941 350
rect 883 310 941 316
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xor2_2
flabel metal1 s 895 316 929 350 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 991 168 1025 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1183 390 1217 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2195048
string GDS_START 2185628
<< end >>
