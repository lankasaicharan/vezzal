magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 6 49 722 243
rect 0 0 768 49
<< scnmos >>
rect 85 49 115 217
rect 171 49 201 217
rect 325 49 355 217
rect 397 49 427 217
rect 505 49 535 217
rect 613 49 643 217
<< scpmoshvt >>
rect 124 367 154 619
rect 210 367 240 619
rect 312 367 342 619
rect 398 367 428 619
rect 527 367 557 619
rect 613 367 643 619
<< ndiff >>
rect 32 204 85 217
rect 32 170 40 204
rect 74 170 85 204
rect 32 95 85 170
rect 32 61 40 95
rect 74 61 85 95
rect 32 49 85 61
rect 115 209 171 217
rect 115 175 126 209
rect 160 175 171 209
rect 115 101 171 175
rect 115 67 126 101
rect 160 67 171 101
rect 115 49 171 67
rect 201 128 325 217
rect 201 94 212 128
rect 246 94 280 128
rect 314 94 325 128
rect 201 49 325 94
rect 355 49 397 217
rect 427 49 505 217
rect 535 199 613 217
rect 535 165 554 199
rect 588 165 613 199
rect 535 96 613 165
rect 535 62 554 96
rect 588 62 613 96
rect 535 49 613 62
rect 643 205 696 217
rect 643 171 654 205
rect 688 171 696 205
rect 643 95 696 171
rect 643 61 654 95
rect 688 61 696 95
rect 643 49 696 61
<< pdiff >>
rect 49 607 124 619
rect 49 573 57 607
rect 91 573 124 607
rect 49 509 124 573
rect 49 475 57 509
rect 91 475 124 509
rect 49 415 124 475
rect 49 381 57 415
rect 91 381 124 415
rect 49 367 124 381
rect 154 597 210 619
rect 154 563 165 597
rect 199 563 210 597
rect 154 529 210 563
rect 154 495 165 529
rect 199 495 210 529
rect 154 459 210 495
rect 154 425 165 459
rect 199 425 210 459
rect 154 367 210 425
rect 240 607 312 619
rect 240 573 260 607
rect 294 573 312 607
rect 240 529 312 573
rect 240 495 260 529
rect 294 495 312 529
rect 240 443 312 495
rect 240 409 260 443
rect 294 409 312 443
rect 240 367 312 409
rect 342 599 398 619
rect 342 565 353 599
rect 387 565 398 599
rect 342 529 398 565
rect 342 495 353 529
rect 387 495 398 529
rect 342 459 398 495
rect 342 425 353 459
rect 387 425 398 459
rect 342 367 398 425
rect 428 607 527 619
rect 428 573 461 607
rect 495 573 527 607
rect 428 531 527 573
rect 428 497 461 531
rect 495 497 527 531
rect 428 367 527 497
rect 557 604 613 619
rect 557 570 568 604
rect 602 570 613 604
rect 557 525 613 570
rect 557 491 568 525
rect 602 491 613 525
rect 557 443 613 491
rect 557 409 568 443
rect 602 409 613 443
rect 557 367 613 409
rect 643 599 696 619
rect 643 565 654 599
rect 688 565 696 599
rect 643 510 696 565
rect 643 476 654 510
rect 688 476 696 510
rect 643 413 696 476
rect 643 379 654 413
rect 688 379 696 413
rect 643 367 696 379
<< ndiffc >>
rect 40 170 74 204
rect 40 61 74 95
rect 126 175 160 209
rect 126 67 160 101
rect 212 94 246 128
rect 280 94 314 128
rect 554 165 588 199
rect 554 62 588 96
rect 654 171 688 205
rect 654 61 688 95
<< pdiffc >>
rect 57 573 91 607
rect 57 475 91 509
rect 57 381 91 415
rect 165 563 199 597
rect 165 495 199 529
rect 165 425 199 459
rect 260 573 294 607
rect 260 495 294 529
rect 260 409 294 443
rect 353 565 387 599
rect 353 495 387 529
rect 353 425 387 459
rect 461 573 495 607
rect 461 497 495 531
rect 568 570 602 604
rect 568 491 602 525
rect 568 409 602 443
rect 654 565 688 599
rect 654 476 688 510
rect 654 379 688 413
<< poly >>
rect 124 619 154 645
rect 210 619 240 645
rect 312 619 342 645
rect 398 619 428 645
rect 527 619 557 645
rect 613 619 643 645
rect 124 305 154 367
rect 210 305 240 367
rect 312 305 342 367
rect 398 305 428 367
rect 527 305 557 367
rect 613 305 643 367
rect 85 289 247 305
rect 85 275 197 289
rect 85 217 115 275
rect 171 255 197 275
rect 231 255 247 289
rect 171 239 247 255
rect 289 289 355 305
rect 289 255 305 289
rect 339 255 355 289
rect 289 239 355 255
rect 171 217 201 239
rect 325 217 355 239
rect 397 289 463 305
rect 397 255 413 289
rect 447 255 463 289
rect 397 239 463 255
rect 505 289 571 305
rect 505 255 521 289
rect 555 255 571 289
rect 505 239 571 255
rect 613 289 727 305
rect 613 255 677 289
rect 711 255 727 289
rect 613 239 727 255
rect 397 217 427 239
rect 505 217 535 239
rect 613 217 643 239
rect 85 23 115 49
rect 171 23 201 49
rect 325 23 355 49
rect 397 23 427 49
rect 505 23 535 49
rect 613 23 643 49
<< polycont >>
rect 197 255 231 289
rect 305 255 339 289
rect 413 255 447 289
rect 521 255 555 289
rect 677 255 711 289
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 41 607 93 649
rect 41 573 57 607
rect 91 573 93 607
rect 41 509 93 573
rect 41 475 57 509
rect 91 475 93 509
rect 41 415 93 475
rect 41 381 57 415
rect 91 381 93 415
rect 41 365 93 381
rect 127 597 210 613
rect 127 563 165 597
rect 199 563 210 597
rect 127 529 210 563
rect 127 495 165 529
rect 199 495 210 529
rect 127 459 210 495
rect 127 425 165 459
rect 199 425 210 459
rect 127 409 210 425
rect 244 607 310 649
rect 244 573 260 607
rect 294 573 310 607
rect 244 529 310 573
rect 244 495 260 529
rect 294 495 310 529
rect 244 443 310 495
rect 244 409 260 443
rect 294 409 310 443
rect 344 599 403 615
rect 344 565 353 599
rect 387 565 403 599
rect 344 529 403 565
rect 344 495 353 529
rect 387 495 403 529
rect 344 459 403 495
rect 445 607 511 649
rect 445 573 461 607
rect 495 573 511 607
rect 445 531 511 573
rect 445 497 461 531
rect 495 497 511 531
rect 445 489 511 497
rect 552 604 618 613
rect 552 570 568 604
rect 602 570 618 604
rect 552 525 618 570
rect 552 491 568 525
rect 602 491 618 525
rect 344 425 353 459
rect 387 445 403 459
rect 552 445 618 491
rect 387 443 618 445
rect 387 425 568 443
rect 344 409 568 425
rect 602 409 618 443
rect 652 599 704 615
rect 652 565 654 599
rect 688 565 704 599
rect 652 510 704 565
rect 652 476 654 510
rect 688 476 704 510
rect 652 413 704 476
rect 127 225 162 409
rect 652 379 654 413
rect 688 379 704 413
rect 652 375 704 379
rect 197 341 704 375
rect 197 289 269 341
rect 231 255 269 289
rect 197 239 269 255
rect 303 289 363 305
rect 303 255 305 289
rect 339 255 363 289
rect 303 239 363 255
rect 397 289 463 305
rect 677 289 751 305
rect 397 255 413 289
rect 447 255 463 289
rect 397 239 463 255
rect 497 255 521 289
rect 555 255 643 289
rect 497 239 643 255
rect 711 255 751 289
rect 677 239 751 255
rect 24 204 90 220
rect 24 170 40 204
rect 74 170 90 204
rect 24 95 90 170
rect 24 61 40 95
rect 74 61 90 95
rect 24 17 90 61
rect 124 209 162 225
rect 124 175 126 209
rect 160 175 162 209
rect 124 101 162 175
rect 235 205 269 239
rect 235 199 604 205
rect 235 171 554 199
rect 538 165 554 171
rect 588 165 604 199
rect 124 67 126 101
rect 160 67 162 101
rect 124 51 162 67
rect 196 128 330 137
rect 196 94 212 128
rect 246 94 280 128
rect 314 94 330 128
rect 196 17 330 94
rect 538 96 604 165
rect 538 62 554 96
rect 588 62 604 96
rect 538 51 604 62
rect 638 171 654 205
rect 688 171 704 205
rect 638 95 704 171
rect 638 61 654 95
rect 688 61 704 95
rect 638 17 704 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a31o_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2780304
string GDS_START 2772700
<< end >>
