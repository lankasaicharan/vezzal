magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 36 49 718 167
rect 0 0 768 49
<< scnmos >>
rect 119 57 149 141
rect 197 57 227 141
rect 283 57 313 141
rect 361 57 391 141
rect 447 57 477 141
rect 519 57 549 141
rect 605 57 635 141
<< scpmoshvt >>
rect 85 431 115 515
rect 157 431 187 515
rect 289 431 319 515
rect 361 431 391 515
rect 447 431 477 515
rect 519 431 549 515
rect 629 387 659 515
<< ndiff >>
rect 62 116 119 141
rect 62 82 74 116
rect 108 82 119 116
rect 62 57 119 82
rect 149 57 197 141
rect 227 116 283 141
rect 227 82 238 116
rect 272 82 283 116
rect 227 57 283 82
rect 313 57 361 141
rect 391 116 447 141
rect 391 82 402 116
rect 436 82 447 116
rect 391 57 447 82
rect 477 57 519 141
rect 549 116 605 141
rect 549 82 560 116
rect 594 82 605 116
rect 549 57 605 82
rect 635 116 692 141
rect 635 82 646 116
rect 680 82 692 116
rect 635 57 692 82
<< pdiff >>
rect 28 490 85 515
rect 28 456 40 490
rect 74 456 85 490
rect 28 431 85 456
rect 115 431 157 515
rect 187 490 289 515
rect 187 456 221 490
rect 255 456 289 490
rect 187 431 289 456
rect 319 431 361 515
rect 391 490 447 515
rect 391 456 402 490
rect 436 456 447 490
rect 391 431 447 456
rect 477 431 519 515
rect 549 475 629 515
rect 549 441 584 475
rect 618 441 629 475
rect 549 431 629 441
rect 572 387 629 431
rect 659 503 739 515
rect 659 469 693 503
rect 727 469 739 503
rect 659 433 739 469
rect 659 399 693 433
rect 727 399 739 433
rect 659 387 739 399
<< ndiffc >>
rect 74 82 108 116
rect 238 82 272 116
rect 402 82 436 116
rect 560 82 594 116
rect 646 82 680 116
<< pdiffc >>
rect 40 456 74 490
rect 221 456 255 490
rect 402 456 436 490
rect 584 441 618 475
rect 693 469 727 503
rect 693 399 727 433
<< poly >>
rect 85 597 585 619
rect 85 589 535 597
rect 85 515 115 589
rect 519 563 535 589
rect 569 563 585 597
rect 519 547 585 563
rect 157 515 187 541
rect 289 515 319 541
rect 361 515 391 541
rect 447 515 477 541
rect 519 515 549 547
rect 629 515 659 541
rect 85 331 115 431
rect 157 409 187 431
rect 157 379 227 409
rect 85 301 149 331
rect 119 141 149 301
rect 197 315 227 379
rect 289 315 319 431
rect 197 299 319 315
rect 197 265 253 299
rect 287 285 319 299
rect 361 315 391 431
rect 447 315 477 431
rect 361 299 477 315
rect 287 265 313 285
rect 197 231 313 265
rect 197 197 253 231
rect 287 197 313 231
rect 197 181 313 197
rect 197 141 227 181
rect 283 141 313 181
rect 361 265 425 299
rect 459 265 477 299
rect 361 231 477 265
rect 361 197 425 231
rect 459 197 477 231
rect 361 181 477 197
rect 361 141 391 181
rect 447 141 477 181
rect 519 141 549 431
rect 629 355 659 387
rect 591 339 659 355
rect 591 305 607 339
rect 641 305 659 339
rect 591 271 659 305
rect 591 237 607 271
rect 641 237 659 271
rect 591 221 659 237
rect 605 141 635 221
rect 119 31 149 57
rect 197 31 227 57
rect 283 31 313 57
rect 361 31 391 57
rect 447 31 477 57
rect 519 31 549 57
rect 605 31 635 57
<< polycont >>
rect 535 563 569 597
rect 253 265 287 299
rect 253 197 287 231
rect 425 265 459 299
rect 425 197 459 231
rect 607 305 641 339
rect 607 237 641 271
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 24 490 90 519
rect 24 456 40 490
rect 74 456 90 490
rect 24 385 90 456
rect 205 490 271 649
rect 505 597 585 613
rect 505 563 535 597
rect 569 563 585 597
rect 505 532 585 563
rect 205 456 221 490
rect 255 456 271 490
rect 205 427 271 456
rect 386 490 452 519
rect 621 496 655 649
rect 386 456 402 490
rect 436 456 452 490
rect 386 385 452 456
rect 568 475 655 496
rect 568 441 584 475
rect 618 441 655 475
rect 568 421 655 441
rect 693 503 743 519
rect 727 469 743 503
rect 693 433 743 469
rect 727 399 743 433
rect 24 351 657 385
rect 24 145 58 351
rect 121 299 303 315
rect 121 265 253 299
rect 287 265 303 299
rect 121 231 303 265
rect 121 197 253 231
rect 287 197 303 231
rect 121 181 303 197
rect 339 145 373 351
rect 591 339 657 351
rect 409 299 551 315
rect 409 265 425 299
rect 459 265 551 299
rect 409 231 551 265
rect 409 197 425 231
rect 459 197 551 231
rect 591 305 607 339
rect 641 305 657 339
rect 591 271 657 305
rect 591 237 607 271
rect 641 237 657 271
rect 591 221 657 237
rect 409 181 551 197
rect 693 145 743 399
rect 24 116 124 145
rect 24 82 74 116
rect 108 82 124 116
rect 24 53 124 82
rect 222 116 288 145
rect 222 82 238 116
rect 272 82 288 116
rect 222 17 288 82
rect 339 116 452 145
rect 339 82 402 116
rect 436 82 452 116
rect 339 53 452 82
rect 544 116 594 145
rect 544 82 560 116
rect 544 17 594 82
rect 630 116 743 145
rect 630 82 646 116
rect 680 82 743 116
rect 630 53 743 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 maj3_0
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6737606
string GDS_START 6731530
<< end >>
