magic
tech sky130A
magscale 1 2
timestamp 1627201166
<< checkpaint >>
rect -1250 -1349 1722 1723
<< pwell >>
rect 10 10 462 392
<< nmoslvt >>
rect 92 36 122 366
rect 178 36 208 366
rect 264 36 294 366
rect 350 36 380 366
<< ndiff >>
rect 36 329 92 366
rect 36 295 47 329
rect 81 295 92 329
rect 36 257 92 295
rect 36 223 47 257
rect 81 223 92 257
rect 36 185 92 223
rect 36 151 47 185
rect 81 151 92 185
rect 36 113 92 151
rect 36 79 47 113
rect 81 79 92 113
rect 36 36 92 79
rect 122 329 178 366
rect 122 295 133 329
rect 167 295 178 329
rect 122 257 178 295
rect 122 223 133 257
rect 167 223 178 257
rect 122 185 178 223
rect 122 151 133 185
rect 167 151 178 185
rect 122 113 178 151
rect 122 79 133 113
rect 167 79 178 113
rect 122 36 178 79
rect 208 329 264 366
rect 208 295 219 329
rect 253 295 264 329
rect 208 257 264 295
rect 208 223 219 257
rect 253 223 264 257
rect 208 185 264 223
rect 208 151 219 185
rect 253 151 264 185
rect 208 113 264 151
rect 208 79 219 113
rect 253 79 264 113
rect 208 36 264 79
rect 294 329 350 366
rect 294 295 305 329
rect 339 295 350 329
rect 294 257 350 295
rect 294 223 305 257
rect 339 223 350 257
rect 294 185 350 223
rect 294 151 305 185
rect 339 151 350 185
rect 294 113 350 151
rect 294 79 305 113
rect 339 79 350 113
rect 294 36 350 79
rect 380 329 436 366
rect 380 295 391 329
rect 425 295 436 329
rect 380 257 436 295
rect 380 223 391 257
rect 425 223 436 257
rect 380 185 436 223
rect 380 151 391 185
rect 425 151 436 185
rect 380 113 436 151
rect 380 79 391 113
rect 425 79 436 113
rect 380 36 436 79
<< ndiffc >>
rect 47 295 81 329
rect 47 223 81 257
rect 47 151 81 185
rect 47 79 81 113
rect 133 295 167 329
rect 133 223 167 257
rect 133 151 167 185
rect 133 79 167 113
rect 219 295 253 329
rect 219 223 253 257
rect 219 151 253 185
rect 219 79 253 113
rect 305 295 339 329
rect 305 223 339 257
rect 305 151 339 185
rect 305 79 339 113
rect 391 295 425 329
rect 391 223 425 257
rect 391 151 425 185
rect 391 79 425 113
<< poly >>
rect 92 447 380 463
rect 92 413 117 447
rect 151 413 185 447
rect 219 413 253 447
rect 287 413 321 447
rect 355 413 380 447
rect 92 392 380 413
rect 92 366 122 392
rect 178 366 208 392
rect 264 366 294 392
rect 350 366 380 392
rect 92 10 122 36
rect 178 10 208 36
rect 264 10 294 36
rect 350 10 380 36
<< polycont >>
rect 117 413 151 447
rect 185 413 219 447
rect 253 413 287 447
rect 321 413 355 447
<< locali >>
rect 101 447 371 463
rect 101 413 111 447
rect 151 413 183 447
rect 219 413 253 447
rect 289 413 321 447
rect 361 413 371 447
rect 101 397 371 413
rect 47 329 81 357
rect 47 257 81 295
rect 47 185 81 223
rect 47 113 81 151
rect 47 51 81 79
rect 133 329 167 357
rect 133 257 167 295
rect 133 185 167 223
rect 133 113 167 151
rect 133 51 167 79
rect 219 329 253 357
rect 219 257 253 295
rect 219 185 253 223
rect 219 113 253 151
rect 219 51 253 79
rect 305 329 339 357
rect 305 257 339 295
rect 305 185 339 223
rect 305 113 339 151
rect 305 51 339 79
rect 391 329 425 357
rect 391 257 425 295
rect 391 185 425 223
rect 391 113 425 151
rect 391 51 425 79
<< viali >>
rect 111 413 117 447
rect 117 413 145 447
rect 183 413 185 447
rect 185 413 217 447
rect 255 413 287 447
rect 287 413 289 447
rect 327 413 355 447
rect 355 413 361 447
rect 47 295 81 329
rect 47 223 81 257
rect 47 151 81 185
rect 47 79 81 113
rect 133 295 167 329
rect 133 223 167 257
rect 133 151 167 185
rect 133 79 167 113
rect 219 295 253 329
rect 219 223 253 257
rect 219 151 253 185
rect 219 79 253 113
rect 305 295 339 329
rect 305 223 339 257
rect 305 151 339 185
rect 305 79 339 113
rect 391 295 425 329
rect 391 223 425 257
rect 391 151 425 185
rect 391 79 425 113
<< metal1 >>
rect 99 447 373 459
rect 99 413 111 447
rect 145 413 183 447
rect 217 413 255 447
rect 289 413 327 447
rect 361 413 373 447
rect 99 401 373 413
rect 41 329 87 357
rect 41 295 47 329
rect 81 295 87 329
rect 41 257 87 295
rect 41 223 47 257
rect 81 223 87 257
rect 41 185 87 223
rect 41 151 47 185
rect 81 151 87 185
rect 41 113 87 151
rect 41 79 47 113
rect 81 79 87 113
rect 41 -29 87 79
rect 124 338 176 357
rect 124 274 176 286
rect 124 185 176 222
rect 124 151 133 185
rect 167 151 176 185
rect 124 113 176 151
rect 124 79 133 113
rect 167 79 176 113
rect 124 51 176 79
rect 213 329 259 357
rect 213 295 219 329
rect 253 295 259 329
rect 213 257 259 295
rect 213 223 219 257
rect 253 223 259 257
rect 213 185 259 223
rect 213 151 219 185
rect 253 151 259 185
rect 213 113 259 151
rect 213 79 219 113
rect 253 79 259 113
rect 213 -29 259 79
rect 296 338 348 357
rect 296 274 348 286
rect 296 185 348 222
rect 296 151 305 185
rect 339 151 348 185
rect 296 113 348 151
rect 296 79 305 113
rect 339 79 348 113
rect 296 51 348 79
rect 385 329 431 357
rect 385 295 391 329
rect 425 295 431 329
rect 385 257 431 295
rect 385 223 391 257
rect 425 223 431 257
rect 385 185 431 223
rect 385 151 391 185
rect 425 151 431 185
rect 385 113 431 151
rect 385 79 391 113
rect 425 79 431 113
rect 385 -29 431 79
rect 41 -89 431 -29
<< via1 >>
rect 124 329 176 338
rect 124 295 133 329
rect 133 295 167 329
rect 167 295 176 329
rect 124 286 176 295
rect 124 257 176 274
rect 124 223 133 257
rect 133 223 167 257
rect 167 223 176 257
rect 124 222 176 223
rect 296 329 348 338
rect 296 295 305 329
rect 305 295 339 329
rect 339 295 348 329
rect 296 286 348 295
rect 296 257 348 274
rect 296 223 305 257
rect 305 223 339 257
rect 339 223 348 257
rect 296 222 348 223
<< metal2 >>
rect 117 348 183 357
rect 117 292 122 348
rect 178 292 183 348
rect 117 286 124 292
rect 176 286 183 292
rect 117 274 183 286
rect 117 268 124 274
rect 176 268 183 274
rect 117 212 122 268
rect 178 212 183 268
rect 117 203 183 212
rect 289 348 355 357
rect 289 292 294 348
rect 350 292 355 348
rect 289 286 296 292
rect 348 286 355 292
rect 289 274 355 286
rect 289 268 296 274
rect 348 268 355 274
rect 289 212 294 268
rect 350 212 355 268
rect 289 203 355 212
<< via2 >>
rect 122 338 178 348
rect 122 292 124 338
rect 124 292 176 338
rect 176 292 178 338
rect 122 222 124 268
rect 124 222 176 268
rect 176 222 178 268
rect 122 212 178 222
rect 294 338 350 348
rect 294 292 296 338
rect 296 292 348 338
rect 348 292 350 338
rect 294 222 296 268
rect 296 222 348 268
rect 348 222 350 268
rect 294 212 350 222
<< metal3 >>
rect 117 348 355 357
rect 117 292 122 348
rect 178 292 294 348
rect 350 292 355 348
rect 117 291 355 292
rect 117 268 183 291
rect 117 212 122 268
rect 178 212 183 268
rect 117 203 183 212
rect 289 268 355 291
rect 289 212 294 268
rect 350 212 355 268
rect 289 203 355 212
<< labels >>
flabel metal3 s 117 291 355 357 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 99 401 373 459 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 41 -89 431 -29 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel pwell s 74 370 90 389 0 FreeSans 200 0 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 5856414
string GDS_START 5848448
string path 10.200 8.925 10.200 -2.225 
<< end >>
