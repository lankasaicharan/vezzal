magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 157 210 648 248
rect 36 49 648 210
rect 0 0 672 49
<< scpmos >>
rect 113 368 149 536
rect 227 368 263 592
rect 311 368 347 592
rect 413 368 449 592
rect 527 368 563 592
<< nmoslvt >>
rect 119 74 149 184
rect 233 74 263 222
rect 319 74 349 222
rect 435 74 465 222
rect 521 74 551 222
<< ndiff >>
rect 183 184 233 222
rect 62 146 119 184
rect 62 112 74 146
rect 108 112 119 146
rect 62 74 119 112
rect 149 146 233 184
rect 149 112 174 146
rect 208 112 233 146
rect 149 74 233 112
rect 263 210 319 222
rect 263 176 274 210
rect 308 176 319 210
rect 263 120 319 176
rect 263 86 274 120
rect 308 86 319 120
rect 263 74 319 86
rect 349 136 435 222
rect 349 102 374 136
rect 408 102 435 136
rect 349 74 435 102
rect 465 210 521 222
rect 465 176 476 210
rect 510 176 521 210
rect 465 120 521 176
rect 465 86 476 120
rect 510 86 521 120
rect 465 74 521 86
rect 551 136 622 222
rect 551 102 576 136
rect 610 102 622 136
rect 551 74 622 102
<< pdiff >>
rect 171 580 227 592
rect 171 546 183 580
rect 217 546 227 580
rect 171 536 227 546
rect 57 524 113 536
rect 57 490 69 524
rect 103 490 113 524
rect 57 414 113 490
rect 57 380 69 414
rect 103 380 113 414
rect 57 368 113 380
rect 149 508 227 536
rect 149 474 183 508
rect 217 474 227 508
rect 149 368 227 474
rect 263 368 311 592
rect 347 368 413 592
rect 449 368 527 592
rect 563 580 643 592
rect 563 546 597 580
rect 631 546 643 580
rect 563 500 643 546
rect 563 466 597 500
rect 631 466 643 500
rect 563 420 643 466
rect 563 386 597 420
rect 631 386 643 420
rect 563 368 643 386
<< ndiffc >>
rect 74 112 108 146
rect 174 112 208 146
rect 274 176 308 210
rect 274 86 308 120
rect 374 102 408 136
rect 476 176 510 210
rect 476 86 510 120
rect 576 102 610 136
<< pdiffc >>
rect 183 546 217 580
rect 69 490 103 524
rect 69 380 103 414
rect 183 474 217 508
rect 597 546 631 580
rect 597 466 631 500
rect 597 386 631 420
<< poly >>
rect 227 592 263 618
rect 311 592 347 618
rect 413 592 449 618
rect 527 592 563 618
rect 113 536 149 562
rect 113 288 149 368
rect 227 336 263 368
rect 311 336 347 368
rect 413 336 449 368
rect 527 336 563 368
rect 197 320 263 336
rect 89 272 155 288
rect 89 238 105 272
rect 139 238 155 272
rect 197 286 213 320
rect 247 286 263 320
rect 197 270 263 286
rect 305 320 371 336
rect 305 286 321 320
rect 355 286 371 320
rect 305 270 371 286
rect 413 320 479 336
rect 413 286 429 320
rect 463 286 479 320
rect 413 270 479 286
rect 521 320 587 336
rect 521 286 537 320
rect 571 286 587 320
rect 521 270 587 286
rect 89 222 155 238
rect 233 222 263 270
rect 319 222 349 270
rect 435 222 465 270
rect 521 222 551 270
rect 119 184 149 222
rect 119 48 149 74
rect 233 48 263 74
rect 319 48 349 74
rect 435 48 465 74
rect 521 48 551 74
<< polycont >>
rect 105 238 139 272
rect 213 286 247 320
rect 321 286 355 320
rect 429 286 463 320
rect 537 286 571 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 167 580 233 649
rect 167 546 183 580
rect 217 546 233 580
rect 21 524 119 540
rect 21 490 69 524
rect 103 490 119 524
rect 21 424 119 490
rect 167 508 233 546
rect 167 474 183 508
rect 217 474 233 508
rect 167 458 233 474
rect 581 580 655 596
rect 581 546 597 580
rect 631 546 655 580
rect 581 500 655 546
rect 581 466 597 500
rect 631 466 655 500
rect 21 414 547 424
rect 21 380 69 414
rect 103 390 547 414
rect 103 380 119 390
rect 21 364 119 380
rect 21 188 55 364
rect 197 320 263 356
rect 89 272 163 288
rect 89 238 105 272
rect 139 238 163 272
rect 197 286 213 320
rect 247 286 263 320
rect 197 270 263 286
rect 305 320 371 356
rect 305 286 321 320
rect 355 286 371 320
rect 305 270 371 286
rect 409 320 479 356
rect 409 286 429 320
rect 463 286 479 320
rect 409 270 479 286
rect 513 336 547 390
rect 581 420 655 466
rect 581 386 597 420
rect 631 386 655 420
rect 581 370 655 386
rect 513 320 587 336
rect 513 286 537 320
rect 571 286 587 320
rect 513 270 587 286
rect 89 222 163 238
rect 621 236 655 370
rect 258 210 655 236
rect 21 146 124 188
rect 21 112 74 146
rect 108 112 124 146
rect 21 70 124 112
rect 158 146 224 188
rect 158 112 174 146
rect 208 112 224 146
rect 158 17 224 112
rect 258 176 274 210
rect 308 202 476 210
rect 308 176 324 202
rect 258 120 324 176
rect 460 176 476 202
rect 510 202 655 210
rect 510 176 526 202
rect 258 86 274 120
rect 308 86 324 120
rect 258 70 324 86
rect 358 136 424 168
rect 358 102 374 136
rect 408 102 424 136
rect 358 17 424 102
rect 460 120 526 176
rect 460 86 476 120
rect 510 86 526 120
rect 460 70 526 86
rect 560 136 626 168
rect 560 102 576 136
rect 610 102 626 136
rect 560 17 626 102
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4b_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 921770
string GDS_START 915928
<< end >>
