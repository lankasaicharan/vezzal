magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3026 1975
<< nwell >>
rect -38 331 1766 704
rect 176 321 1081 331
rect 176 317 344 321
<< pwell >>
rect 19 157 293 246
rect 831 157 1727 263
rect 19 49 1727 157
rect 0 0 1728 49
<< scnmos >>
rect 98 136 128 220
rect 184 136 214 220
rect 407 47 437 131
rect 517 47 547 131
rect 589 47 619 131
rect 707 47 737 131
rect 805 47 835 131
rect 937 69 967 237
rect 1195 153 1225 237
rect 1328 69 1358 237
rect 1414 69 1444 237
rect 1532 69 1562 237
rect 1618 69 1648 237
<< scpmoshvt >>
rect 112 415 142 543
rect 198 415 228 543
rect 415 491 445 619
rect 559 491 589 619
rect 631 491 661 619
rect 739 491 769 575
rect 811 491 841 575
rect 962 357 992 609
rect 1195 367 1225 495
rect 1328 367 1358 619
rect 1414 367 1444 619
rect 1516 367 1546 619
rect 1602 367 1632 619
<< ndiff >>
rect 45 192 98 220
rect 45 158 53 192
rect 87 158 98 192
rect 45 136 98 158
rect 128 192 184 220
rect 128 158 139 192
rect 173 158 184 192
rect 128 136 184 158
rect 214 202 267 220
rect 214 168 225 202
rect 259 168 267 202
rect 214 136 267 168
rect 857 177 937 237
rect 857 143 869 177
rect 903 143 937 177
rect 857 131 937 143
rect 354 106 407 131
rect 354 72 362 106
rect 396 72 407 106
rect 354 47 407 72
rect 437 87 517 131
rect 437 53 460 87
rect 494 53 517 87
rect 437 47 517 53
rect 547 47 589 131
rect 619 87 707 131
rect 619 53 646 87
rect 680 53 707 87
rect 619 47 707 53
rect 737 47 805 131
rect 835 89 937 131
rect 835 55 869 89
rect 903 69 937 89
rect 967 209 1024 237
rect 967 175 978 209
rect 1012 175 1024 209
rect 967 111 1024 175
rect 1138 229 1195 237
rect 1138 195 1150 229
rect 1184 195 1195 229
rect 1138 153 1195 195
rect 1225 153 1328 237
rect 967 77 978 111
rect 1012 77 1024 111
rect 967 69 1024 77
rect 903 55 915 69
rect 835 47 915 55
rect 452 41 502 47
rect 634 45 692 47
rect 1248 89 1328 153
rect 1248 55 1260 89
rect 1294 69 1328 89
rect 1358 229 1414 237
rect 1358 195 1369 229
rect 1403 195 1414 229
rect 1358 69 1414 195
rect 1444 89 1532 237
rect 1444 69 1471 89
rect 1294 55 1306 69
rect 1248 47 1306 55
rect 1459 55 1471 69
rect 1505 69 1532 89
rect 1562 229 1618 237
rect 1562 195 1573 229
rect 1607 195 1618 229
rect 1562 116 1618 195
rect 1562 82 1573 116
rect 1607 82 1618 116
rect 1562 69 1618 82
rect 1648 225 1701 237
rect 1648 191 1659 225
rect 1693 191 1701 225
rect 1648 115 1701 191
rect 1648 81 1659 115
rect 1693 81 1701 115
rect 1648 69 1701 81
rect 1505 55 1517 69
rect 1459 47 1517 55
<< pdiff >>
rect 362 607 415 619
rect 362 573 370 607
rect 404 573 415 607
rect 48 530 112 543
rect 48 496 56 530
rect 90 496 112 530
rect 48 462 112 496
rect 48 428 56 462
rect 90 428 112 462
rect 48 415 112 428
rect 142 535 198 543
rect 142 501 153 535
rect 187 501 198 535
rect 142 415 198 501
rect 228 415 308 543
rect 362 539 415 573
rect 362 505 370 539
rect 404 505 415 539
rect 362 491 415 505
rect 445 606 559 619
rect 445 572 484 606
rect 518 572 559 606
rect 445 491 559 572
rect 589 491 631 619
rect 661 605 714 619
rect 1267 611 1328 619
rect 661 571 672 605
rect 706 575 714 605
rect 905 601 962 609
rect 905 575 917 601
rect 706 571 739 575
rect 661 537 739 571
rect 661 503 672 537
rect 706 503 739 537
rect 661 491 739 503
rect 769 491 811 575
rect 841 567 917 575
rect 951 567 962 601
rect 841 533 962 567
rect 841 499 852 533
rect 886 499 962 533
rect 841 491 962 499
rect 250 395 308 415
rect 250 361 262 395
rect 296 361 308 395
rect 250 353 308 361
rect 909 481 962 491
rect 909 447 917 481
rect 951 447 962 481
rect 909 357 962 447
rect 992 597 1045 609
rect 992 563 1003 597
rect 1037 563 1045 597
rect 992 502 1045 563
rect 1267 577 1283 611
rect 1317 577 1328 611
rect 1267 543 1328 577
rect 992 468 1003 502
rect 1037 468 1045 502
rect 1267 509 1283 543
rect 1317 509 1328 543
rect 1267 495 1328 509
rect 992 403 1045 468
rect 992 369 1003 403
rect 1037 369 1045 403
rect 992 357 1045 369
rect 1142 481 1195 495
rect 1142 447 1150 481
rect 1184 447 1195 481
rect 1142 413 1195 447
rect 1142 379 1150 413
rect 1184 379 1195 413
rect 1142 367 1195 379
rect 1225 477 1328 495
rect 1225 443 1236 477
rect 1270 443 1328 477
rect 1225 409 1328 443
rect 1225 375 1236 409
rect 1270 375 1328 409
rect 1225 367 1328 375
rect 1358 599 1414 619
rect 1358 565 1369 599
rect 1403 565 1414 599
rect 1358 497 1414 565
rect 1358 463 1369 497
rect 1403 463 1414 497
rect 1358 420 1414 463
rect 1358 386 1369 420
rect 1403 386 1414 420
rect 1358 367 1414 386
rect 1444 571 1516 619
rect 1444 537 1469 571
rect 1503 537 1516 571
rect 1444 367 1516 537
rect 1546 419 1602 619
rect 1546 385 1557 419
rect 1591 385 1602 419
rect 1546 367 1602 385
rect 1632 571 1685 619
rect 1632 537 1643 571
rect 1677 537 1685 571
rect 1632 367 1685 537
<< ndiffc >>
rect 53 158 87 192
rect 139 158 173 192
rect 225 168 259 202
rect 869 143 903 177
rect 362 72 396 106
rect 460 53 494 87
rect 646 53 680 87
rect 869 55 903 89
rect 978 175 1012 209
rect 1150 195 1184 229
rect 978 77 1012 111
rect 1260 55 1294 89
rect 1369 195 1403 229
rect 1471 55 1505 89
rect 1573 195 1607 229
rect 1573 82 1607 116
rect 1659 191 1693 225
rect 1659 81 1693 115
<< pdiffc >>
rect 370 573 404 607
rect 56 496 90 530
rect 56 428 90 462
rect 153 501 187 535
rect 370 505 404 539
rect 484 572 518 606
rect 672 571 706 605
rect 672 503 706 537
rect 917 567 951 601
rect 852 499 886 533
rect 262 361 296 395
rect 917 447 951 481
rect 1003 563 1037 597
rect 1283 577 1317 611
rect 1003 468 1037 502
rect 1283 509 1317 543
rect 1003 369 1037 403
rect 1150 447 1184 481
rect 1150 379 1184 413
rect 1236 443 1270 477
rect 1236 375 1270 409
rect 1369 565 1403 599
rect 1369 463 1403 497
rect 1369 386 1403 420
rect 1469 537 1503 571
rect 1557 385 1591 419
rect 1643 537 1677 571
<< poly >>
rect 415 619 445 645
rect 559 619 589 645
rect 631 619 661 645
rect 112 543 142 569
rect 198 543 228 569
rect 962 609 992 635
rect 1328 619 1358 645
rect 1414 619 1444 645
rect 1516 619 1546 645
rect 1602 619 1632 645
rect 739 575 769 601
rect 811 575 841 601
rect 415 459 445 491
rect 559 459 589 491
rect 112 376 142 415
rect 76 360 142 376
rect 76 326 92 360
rect 126 326 142 360
rect 76 292 142 326
rect 76 258 92 292
rect 126 258 142 292
rect 198 272 228 415
rect 400 429 445 459
rect 487 443 589 459
rect 400 327 430 429
rect 487 409 503 443
rect 537 429 589 443
rect 631 459 661 491
rect 631 443 697 459
rect 537 409 553 429
rect 487 393 553 409
rect 631 409 647 443
rect 681 409 697 443
rect 631 393 697 409
rect 487 391 538 393
rect 364 311 430 327
rect 472 375 538 391
rect 472 341 488 375
rect 522 341 538 375
rect 739 351 769 491
rect 472 325 538 341
rect 587 335 769 351
rect 364 277 380 311
rect 414 277 430 311
rect 76 242 142 258
rect 184 242 322 272
rect 98 220 128 242
rect 184 220 214 242
rect 98 110 128 136
rect 184 110 214 136
rect 292 114 322 242
rect 364 243 430 277
rect 364 209 380 243
rect 414 209 430 243
rect 364 193 430 209
rect 400 176 430 193
rect 488 176 518 325
rect 587 301 603 335
rect 637 301 769 335
rect 587 285 769 301
rect 811 413 841 491
rect 811 397 877 413
rect 811 363 827 397
rect 861 363 877 397
rect 811 329 877 363
rect 1195 495 1225 521
rect 811 295 827 329
rect 861 295 877 329
rect 962 325 992 357
rect 587 283 632 285
rect 566 267 632 283
rect 566 233 582 267
rect 616 233 632 267
rect 811 279 877 295
rect 919 309 992 325
rect 566 217 632 233
rect 674 221 740 237
rect 400 146 437 176
rect 488 146 547 176
rect 407 131 437 146
rect 517 131 547 146
rect 589 131 619 217
rect 674 187 690 221
rect 724 187 740 221
rect 674 171 740 187
rect 811 183 841 279
rect 919 275 935 309
rect 969 275 992 309
rect 919 259 992 275
rect 937 237 967 259
rect 1195 237 1225 367
rect 1328 325 1358 367
rect 1267 309 1358 325
rect 1267 275 1283 309
rect 1317 289 1358 309
rect 1414 289 1444 367
rect 1317 275 1444 289
rect 1267 259 1444 275
rect 1516 289 1546 367
rect 1602 325 1632 367
rect 1602 309 1697 325
rect 1602 289 1647 309
rect 1516 275 1647 289
rect 1681 275 1697 309
rect 1516 259 1697 275
rect 1328 237 1358 259
rect 1414 237 1444 259
rect 1532 237 1562 259
rect 1618 237 1648 259
rect 707 131 737 171
rect 805 153 841 183
rect 805 131 835 153
rect 256 98 322 114
rect 256 64 272 98
rect 306 64 322 98
rect 256 48 322 64
rect 1195 105 1225 153
rect 1142 89 1225 105
rect 407 21 437 47
rect 517 21 547 47
rect 589 21 619 47
rect 707 21 737 47
rect 805 21 835 47
rect 937 43 967 69
rect 1142 55 1158 89
rect 1192 55 1225 89
rect 1142 39 1225 55
rect 1328 43 1358 69
rect 1414 43 1444 69
rect 1532 43 1562 69
rect 1618 43 1648 69
<< polycont >>
rect 92 326 126 360
rect 92 258 126 292
rect 503 409 537 443
rect 647 409 681 443
rect 488 341 522 375
rect 380 277 414 311
rect 380 209 414 243
rect 603 301 637 335
rect 827 363 861 397
rect 827 295 861 329
rect 582 233 616 267
rect 690 187 724 221
rect 935 275 969 309
rect 1283 275 1317 309
rect 1647 275 1681 309
rect 272 64 306 98
rect 1158 55 1192 89
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 22 530 103 546
rect 22 496 56 530
rect 90 496 103 530
rect 137 535 203 649
rect 137 501 153 535
rect 187 501 203 535
rect 137 499 203 501
rect 354 607 420 615
rect 354 573 370 607
rect 404 573 420 607
rect 354 539 420 573
rect 468 606 534 649
rect 468 572 484 606
rect 518 572 534 606
rect 468 567 534 572
rect 656 605 722 615
rect 656 571 672 605
rect 706 571 722 605
rect 354 505 370 539
rect 404 533 420 539
rect 656 537 722 571
rect 404 505 620 533
rect 354 499 620 505
rect 22 465 103 496
rect 22 462 552 465
rect 22 428 56 462
rect 90 443 552 462
rect 90 431 503 443
rect 90 428 106 431
rect 22 412 106 428
rect 22 208 56 412
rect 487 409 503 431
rect 537 409 552 443
rect 246 395 312 397
rect 90 360 182 376
rect 90 326 92 360
rect 126 326 182 360
rect 90 292 182 326
rect 90 258 92 292
rect 126 258 182 292
rect 90 242 182 258
rect 246 361 262 395
rect 296 391 312 395
rect 296 361 437 391
rect 246 311 437 361
rect 487 375 552 409
rect 586 444 620 499
rect 656 503 672 537
rect 706 512 722 537
rect 849 601 967 649
rect 849 567 917 601
rect 951 567 967 601
rect 849 533 967 567
rect 706 503 792 512
rect 656 478 792 503
rect 586 443 724 444
rect 586 409 647 443
rect 681 409 724 443
rect 586 393 724 409
rect 487 341 488 375
rect 522 341 552 375
rect 487 325 552 341
rect 587 335 642 351
rect 246 277 380 311
rect 414 277 437 311
rect 246 275 437 277
rect 587 301 603 335
rect 637 301 642 335
rect 587 275 642 301
rect 246 267 642 275
rect 246 243 582 267
rect 246 218 380 243
rect 209 209 380 218
rect 414 233 582 243
rect 616 233 642 267
rect 414 209 642 233
rect 22 192 97 208
rect 22 158 53 192
rect 87 158 97 192
rect 22 140 97 158
rect 131 192 175 208
rect 131 158 139 192
rect 173 158 175 192
rect 209 202 642 209
rect 209 168 225 202
rect 259 193 642 202
rect 676 221 724 393
rect 259 168 280 193
rect 209 164 280 168
rect 676 187 690 221
rect 676 159 724 187
rect 131 17 175 158
rect 223 98 322 130
rect 223 64 272 98
rect 306 64 322 98
rect 356 125 724 159
rect 758 245 792 478
rect 849 499 852 533
rect 886 499 967 533
rect 849 481 967 499
rect 849 447 917 481
rect 951 447 967 481
rect 1001 597 1053 615
rect 1001 563 1003 597
rect 1037 563 1053 597
rect 1001 502 1053 563
rect 1001 468 1003 502
rect 1037 468 1053 502
rect 1227 611 1317 649
rect 1227 577 1283 611
rect 1227 543 1317 577
rect 1227 509 1283 543
rect 1001 413 1053 468
rect 826 403 1053 413
rect 826 397 1003 403
rect 826 363 827 397
rect 861 369 1003 397
rect 1037 369 1053 403
rect 861 363 1053 369
rect 826 359 1053 363
rect 826 329 867 359
rect 826 295 827 329
rect 861 295 867 329
rect 826 279 867 295
rect 901 309 983 325
rect 901 275 935 309
rect 969 275 983 309
rect 901 259 983 275
rect 901 245 935 259
rect 758 211 935 245
rect 1017 225 1053 359
rect 356 106 410 125
rect 356 72 362 106
rect 396 72 410 106
rect 758 91 792 211
rect 969 209 1053 225
rect 356 56 410 72
rect 444 87 510 91
rect 444 53 460 87
rect 494 53 510 87
rect 444 17 510 53
rect 630 87 792 91
rect 630 53 646 87
rect 680 53 792 87
rect 630 51 792 53
rect 853 143 869 177
rect 903 143 919 177
rect 853 89 919 143
rect 853 55 869 89
rect 903 55 919 89
rect 853 17 919 55
rect 969 175 978 209
rect 1012 175 1053 209
rect 1134 481 1193 497
rect 1134 447 1150 481
rect 1184 447 1193 481
rect 1134 413 1193 447
rect 1134 379 1150 413
rect 1184 379 1193 413
rect 1134 325 1193 379
rect 1227 477 1317 509
rect 1227 443 1236 477
rect 1270 443 1317 477
rect 1227 409 1317 443
rect 1227 375 1236 409
rect 1270 375 1317 409
rect 1227 359 1317 375
rect 1353 599 1419 615
rect 1353 565 1369 599
rect 1403 565 1419 599
rect 1353 497 1419 565
rect 1453 571 1519 649
rect 1453 537 1469 571
rect 1503 537 1519 571
rect 1453 529 1519 537
rect 1627 571 1693 649
rect 1627 537 1643 571
rect 1677 537 1693 571
rect 1627 529 1693 537
rect 1353 463 1369 497
rect 1403 463 1419 497
rect 1353 420 1419 463
rect 1353 386 1369 420
rect 1403 386 1419 420
rect 1134 309 1317 325
rect 1134 275 1283 309
rect 1134 259 1317 275
rect 1134 229 1200 259
rect 1134 195 1150 229
rect 1184 195 1200 229
rect 1134 193 1200 195
rect 1353 229 1419 386
rect 1353 195 1369 229
rect 1403 195 1419 229
rect 1353 193 1419 195
rect 1455 461 1698 495
rect 969 111 1053 175
rect 1455 159 1489 461
rect 969 77 978 111
rect 1012 91 1053 111
rect 1142 125 1489 159
rect 1541 419 1609 427
rect 1541 385 1557 419
rect 1591 385 1609 419
rect 1541 229 1609 385
rect 1645 309 1698 461
rect 1645 275 1647 309
rect 1681 275 1698 309
rect 1645 259 1698 275
rect 1541 195 1573 229
rect 1607 195 1609 229
rect 1541 131 1609 195
rect 1142 91 1208 125
rect 1555 116 1609 131
rect 1012 89 1208 91
rect 1012 77 1158 89
rect 969 55 1158 77
rect 1192 55 1208 89
rect 969 51 1208 55
rect 1244 89 1310 91
rect 1244 55 1260 89
rect 1294 55 1310 89
rect 1244 17 1310 55
rect 1455 89 1521 91
rect 1455 55 1471 89
rect 1505 55 1521 89
rect 1555 82 1573 116
rect 1607 82 1609 116
rect 1555 66 1609 82
rect 1643 191 1659 225
rect 1693 191 1709 225
rect 1643 115 1709 191
rect 1643 81 1659 115
rect 1693 81 1709 115
rect 1455 17 1521 55
rect 1643 17 1709 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlxbn_2
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1375 390 1409 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1375 464 1409 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1375 538 1409 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5953208
string GDS_START 5939398
<< end >>
