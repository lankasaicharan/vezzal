magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2034 1852
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 687 203
rect 29 -17 63 21
<< scnmos >>
rect 83 47 113 177
rect 271 47 301 177
rect 355 47 385 177
rect 473 47 503 177
rect 569 47 599 177
<< scpmoshvt >>
rect 85 297 121 497
rect 263 297 299 497
rect 357 297 393 497
rect 475 297 511 497
rect 571 297 607 497
<< ndiff >>
rect 27 136 83 177
rect 27 102 35 136
rect 69 102 83 136
rect 27 47 83 102
rect 113 93 165 177
rect 113 59 123 93
rect 157 59 165 93
rect 113 47 165 59
rect 219 95 271 177
rect 219 61 227 95
rect 261 61 271 95
rect 219 47 271 61
rect 301 163 355 177
rect 301 129 311 163
rect 345 129 355 163
rect 301 47 355 129
rect 385 163 473 177
rect 385 129 429 163
rect 463 129 473 163
rect 385 95 473 129
rect 385 61 429 95
rect 463 61 473 95
rect 385 47 473 61
rect 503 89 569 177
rect 503 55 525 89
rect 559 55 569 89
rect 503 47 569 55
rect 599 163 661 177
rect 599 129 619 163
rect 653 129 661 163
rect 599 95 661 129
rect 599 61 619 95
rect 653 61 661 95
rect 599 47 661 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 263 497
rect 121 443 137 477
rect 171 443 208 477
rect 242 443 263 477
rect 121 409 263 443
rect 121 375 137 409
rect 171 375 208 409
rect 242 375 263 409
rect 121 297 263 375
rect 299 297 357 497
rect 393 477 475 497
rect 393 443 405 477
rect 439 443 475 477
rect 393 409 475 443
rect 393 375 405 409
rect 439 375 475 409
rect 393 341 475 375
rect 393 307 405 341
rect 439 307 475 341
rect 393 297 475 307
rect 511 297 571 497
rect 607 485 661 497
rect 607 451 619 485
rect 653 451 661 485
rect 607 417 661 451
rect 607 383 619 417
rect 653 383 661 417
rect 607 349 661 383
rect 607 315 619 349
rect 653 315 661 349
rect 607 297 661 315
<< ndiffc >>
rect 35 102 69 136
rect 123 59 157 93
rect 227 61 261 95
rect 311 129 345 163
rect 429 129 463 163
rect 429 61 463 95
rect 525 55 559 89
rect 619 129 653 163
rect 619 61 653 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 137 443 171 477
rect 208 443 242 477
rect 137 375 171 409
rect 208 375 242 409
rect 405 443 439 477
rect 405 375 439 409
rect 405 307 439 341
rect 619 451 653 485
rect 619 383 653 417
rect 619 315 653 349
<< poly >>
rect 85 497 121 523
rect 263 497 299 523
rect 357 497 393 523
rect 475 497 511 523
rect 571 497 607 523
rect 85 282 121 297
rect 263 282 299 297
rect 357 282 393 297
rect 475 282 511 297
rect 571 282 607 297
rect 83 265 123 282
rect 261 265 301 282
rect 83 249 151 265
rect 83 215 107 249
rect 141 215 151 249
rect 83 199 151 215
rect 247 249 301 265
rect 247 215 257 249
rect 291 215 301 249
rect 247 199 301 215
rect 83 177 113 199
rect 271 177 301 199
rect 355 265 395 282
rect 473 265 513 282
rect 569 265 609 282
rect 355 249 409 265
rect 355 215 365 249
rect 399 215 409 249
rect 355 199 409 215
rect 473 249 527 265
rect 473 215 483 249
rect 517 215 527 249
rect 473 199 527 215
rect 569 249 627 265
rect 569 215 583 249
rect 617 215 627 249
rect 569 199 627 215
rect 355 177 385 199
rect 473 177 503 199
rect 569 177 599 199
rect 83 21 113 47
rect 271 21 301 47
rect 355 21 385 47
rect 473 21 503 47
rect 569 21 599 47
<< polycont >>
rect 107 215 141 249
rect 257 215 291 249
rect 365 215 399 249
rect 483 215 517 249
rect 583 215 617 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 477 73 493
rect 17 443 39 477
rect 17 409 73 443
rect 17 375 39 409
rect 121 477 272 527
rect 121 443 137 477
rect 171 443 208 477
rect 242 443 272 477
rect 121 409 272 443
rect 121 375 137 409
rect 171 375 208 409
rect 242 375 272 409
rect 361 477 455 493
rect 597 485 708 527
rect 361 443 405 477
rect 439 443 455 477
rect 361 409 455 443
rect 361 375 405 409
rect 439 375 455 409
rect 17 341 73 375
rect 361 341 455 375
rect 17 307 39 341
rect 17 136 73 307
rect 107 307 405 341
rect 439 307 455 341
rect 107 299 455 307
rect 107 249 172 299
rect 489 265 533 481
rect 597 451 619 485
rect 653 451 708 485
rect 597 417 708 451
rect 597 383 619 417
rect 653 383 708 417
rect 597 349 708 383
rect 597 315 619 349
rect 653 315 708 349
rect 597 291 708 315
rect 141 215 172 249
rect 213 249 307 265
rect 213 215 257 249
rect 291 215 307 249
rect 346 249 431 265
rect 346 215 365 249
rect 399 215 431 249
rect 467 249 533 265
rect 467 215 483 249
rect 517 215 533 249
rect 567 249 662 255
rect 567 215 583 249
rect 617 215 662 249
rect 107 179 172 215
rect 107 163 361 179
rect 107 143 311 163
rect 17 102 35 136
rect 69 102 73 136
rect 288 129 311 143
rect 345 129 361 163
rect 413 163 671 173
rect 413 129 429 163
rect 463 139 619 163
rect 463 129 479 139
rect 17 73 73 102
rect 123 93 157 109
rect 413 95 479 129
rect 593 129 619 139
rect 653 129 671 163
rect 211 61 227 95
rect 261 61 429 95
rect 463 61 479 95
rect 211 59 479 61
rect 525 89 559 105
rect 123 17 157 59
rect 593 95 671 129
rect 593 61 619 95
rect 653 61 671 95
rect 593 56 671 61
rect 525 17 559 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 489 357 523 391 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 29 425 63 459 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 259 221 293 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 594 221 628 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 370 221 404 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o22a_1
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 948062
string GDS_START 941852
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
