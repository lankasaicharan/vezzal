magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 17 49 897 259
rect 0 0 960 49
<< scnmos >>
rect 96 65 126 233
rect 182 65 212 233
rect 284 65 314 233
rect 370 65 400 233
rect 530 65 560 233
rect 616 65 646 233
rect 702 65 732 233
rect 788 65 818 233
<< scpmoshvt >>
rect 96 367 126 619
rect 182 367 212 619
rect 268 367 298 619
rect 354 367 384 619
rect 544 367 574 619
rect 630 367 660 619
rect 716 367 746 619
rect 802 367 832 619
<< ndiff >>
rect 43 192 96 233
rect 43 158 51 192
rect 85 158 96 192
rect 43 111 96 158
rect 43 77 51 111
rect 85 77 96 111
rect 43 65 96 77
rect 126 225 182 233
rect 126 191 137 225
rect 171 191 182 225
rect 126 153 182 191
rect 126 119 137 153
rect 171 119 182 153
rect 126 65 182 119
rect 212 114 284 233
rect 212 80 227 114
rect 261 80 284 114
rect 212 65 284 80
rect 314 202 370 233
rect 314 168 325 202
rect 359 168 370 202
rect 314 65 370 168
rect 400 192 530 233
rect 400 158 485 192
rect 519 158 530 192
rect 400 122 530 158
rect 400 88 411 122
rect 445 111 530 122
rect 445 88 485 111
rect 400 77 485 88
rect 519 77 530 111
rect 400 65 530 77
rect 560 132 616 233
rect 560 98 571 132
rect 605 98 616 132
rect 560 65 616 98
rect 646 208 702 233
rect 646 174 657 208
rect 691 174 702 208
rect 646 113 702 174
rect 646 79 657 113
rect 691 79 702 113
rect 646 65 702 79
rect 732 132 788 233
rect 732 98 743 132
rect 777 98 788 132
rect 732 65 788 98
rect 818 208 871 233
rect 818 174 829 208
rect 863 174 871 208
rect 818 113 871 174
rect 818 79 829 113
rect 863 79 871 113
rect 818 65 871 79
<< pdiff >>
rect 43 599 96 619
rect 43 565 51 599
rect 85 565 96 599
rect 43 507 96 565
rect 43 473 51 507
rect 85 473 96 507
rect 43 413 96 473
rect 43 379 51 413
rect 85 379 96 413
rect 43 367 96 379
rect 126 607 182 619
rect 126 573 137 607
rect 171 573 182 607
rect 126 535 182 573
rect 126 501 137 535
rect 171 501 182 535
rect 126 457 182 501
rect 126 423 137 457
rect 171 423 182 457
rect 126 367 182 423
rect 212 599 268 619
rect 212 565 223 599
rect 257 565 268 599
rect 212 506 268 565
rect 212 472 223 506
rect 257 472 268 506
rect 212 413 268 472
rect 212 379 223 413
rect 257 379 268 413
rect 212 367 268 379
rect 298 543 354 619
rect 298 509 309 543
rect 343 509 354 543
rect 298 413 354 509
rect 298 379 309 413
rect 343 379 354 413
rect 298 367 354 379
rect 384 599 437 619
rect 384 565 395 599
rect 429 565 437 599
rect 384 529 437 565
rect 384 495 395 529
rect 429 495 437 529
rect 384 457 437 495
rect 384 423 395 457
rect 429 423 437 457
rect 384 367 437 423
rect 491 599 544 619
rect 491 565 499 599
rect 533 565 544 599
rect 491 529 544 565
rect 491 495 499 529
rect 533 495 544 529
rect 491 457 544 495
rect 491 423 499 457
rect 533 423 544 457
rect 491 367 544 423
rect 574 543 630 619
rect 574 509 585 543
rect 619 509 630 543
rect 574 413 630 509
rect 574 379 585 413
rect 619 379 630 413
rect 574 367 630 379
rect 660 599 716 619
rect 660 565 671 599
rect 705 565 716 599
rect 660 505 716 565
rect 660 471 671 505
rect 705 471 716 505
rect 660 413 716 471
rect 660 379 671 413
rect 705 379 716 413
rect 660 367 716 379
rect 746 611 802 619
rect 746 577 757 611
rect 791 577 802 611
rect 746 526 802 577
rect 746 492 757 526
rect 791 492 802 526
rect 746 441 802 492
rect 746 407 757 441
rect 791 407 802 441
rect 746 367 802 407
rect 832 599 885 619
rect 832 565 843 599
rect 877 565 885 599
rect 832 504 885 565
rect 832 470 843 504
rect 877 470 885 504
rect 832 413 885 470
rect 832 379 843 413
rect 877 379 885 413
rect 832 367 885 379
<< ndiffc >>
rect 51 158 85 192
rect 51 77 85 111
rect 137 191 171 225
rect 137 119 171 153
rect 227 80 261 114
rect 325 168 359 202
rect 485 158 519 192
rect 411 88 445 122
rect 485 77 519 111
rect 571 98 605 132
rect 657 174 691 208
rect 657 79 691 113
rect 743 98 777 132
rect 829 174 863 208
rect 829 79 863 113
<< pdiffc >>
rect 51 565 85 599
rect 51 473 85 507
rect 51 379 85 413
rect 137 573 171 607
rect 137 501 171 535
rect 137 423 171 457
rect 223 565 257 599
rect 223 472 257 506
rect 223 379 257 413
rect 309 509 343 543
rect 309 379 343 413
rect 395 565 429 599
rect 395 495 429 529
rect 395 423 429 457
rect 499 565 533 599
rect 499 495 533 529
rect 499 423 533 457
rect 585 509 619 543
rect 585 379 619 413
rect 671 565 705 599
rect 671 471 705 505
rect 671 379 705 413
rect 757 577 791 611
rect 757 492 791 526
rect 757 407 791 441
rect 843 565 877 599
rect 843 470 877 504
rect 843 379 877 413
<< poly >>
rect 96 619 126 645
rect 182 619 212 645
rect 268 619 298 645
rect 354 619 384 645
rect 544 619 574 645
rect 630 619 660 645
rect 716 619 746 645
rect 802 619 832 645
rect 96 321 126 367
rect 182 321 212 367
rect 35 305 212 321
rect 35 271 51 305
rect 85 271 137 305
rect 171 271 212 305
rect 35 255 212 271
rect 268 321 298 367
rect 354 321 384 367
rect 544 321 574 367
rect 630 321 660 367
rect 268 305 384 321
rect 268 271 284 305
rect 318 285 384 305
rect 508 305 660 321
rect 318 271 400 285
rect 268 255 400 271
rect 508 271 524 305
rect 558 271 610 305
rect 644 271 660 305
rect 716 321 746 367
rect 802 321 832 367
rect 716 305 854 321
rect 716 285 804 305
rect 508 255 660 271
rect 702 271 804 285
rect 838 271 854 305
rect 702 255 854 271
rect 96 233 126 255
rect 182 233 212 255
rect 284 233 314 255
rect 370 233 400 255
rect 530 233 560 255
rect 616 233 646 255
rect 702 233 732 255
rect 788 233 818 255
rect 96 39 126 65
rect 182 39 212 65
rect 284 39 314 65
rect 370 39 400 65
rect 530 39 560 65
rect 616 39 646 65
rect 702 39 732 65
rect 788 39 818 65
<< polycont >>
rect 51 271 85 305
rect 137 271 171 305
rect 284 271 318 305
rect 524 271 558 305
rect 610 271 644 305
rect 804 271 838 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 35 599 87 615
rect 35 565 51 599
rect 85 565 87 599
rect 35 507 87 565
rect 35 473 51 507
rect 85 473 87 507
rect 35 413 87 473
rect 121 607 187 649
rect 121 573 137 607
rect 171 573 187 607
rect 121 535 187 573
rect 121 501 137 535
rect 171 501 187 535
rect 121 457 187 501
rect 121 423 137 457
rect 171 423 187 457
rect 221 599 445 615
rect 221 565 223 599
rect 257 581 395 599
rect 257 565 259 581
rect 221 506 259 565
rect 393 565 395 581
rect 429 565 445 599
rect 221 472 223 506
rect 257 472 259 506
rect 35 379 51 413
rect 85 389 87 413
rect 221 413 259 472
rect 221 389 223 413
rect 85 379 223 389
rect 257 379 259 413
rect 35 355 259 379
rect 293 543 359 547
rect 293 509 309 543
rect 343 509 359 543
rect 293 413 359 509
rect 293 379 309 413
rect 343 379 359 413
rect 393 529 445 565
rect 393 495 395 529
rect 429 495 445 529
rect 393 457 445 495
rect 393 423 395 457
rect 429 423 445 457
rect 393 407 445 423
rect 483 599 707 615
rect 483 565 499 599
rect 533 581 671 599
rect 533 565 535 581
rect 483 529 535 565
rect 669 565 671 581
rect 705 565 707 599
rect 483 495 499 529
rect 533 495 535 529
rect 483 457 535 495
rect 483 423 499 457
rect 533 423 535 457
rect 483 407 535 423
rect 569 543 635 547
rect 569 509 585 543
rect 619 509 635 543
rect 569 413 635 509
rect 293 373 359 379
rect 569 379 585 413
rect 619 379 635 413
rect 569 373 635 379
rect 293 339 635 373
rect 669 505 707 565
rect 669 471 671 505
rect 705 471 707 505
rect 669 413 707 471
rect 669 379 671 413
rect 705 379 707 413
rect 741 611 807 649
rect 741 577 757 611
rect 791 577 807 611
rect 741 526 807 577
rect 741 492 757 526
rect 791 492 807 526
rect 741 441 807 492
rect 741 407 757 441
rect 791 407 807 441
rect 841 599 893 615
rect 841 565 843 599
rect 877 565 893 599
rect 841 504 893 565
rect 841 470 843 504
rect 877 470 893 504
rect 841 413 893 470
rect 669 373 707 379
rect 841 379 843 413
rect 877 379 893 413
rect 841 373 893 379
rect 669 339 893 373
rect 31 305 187 321
rect 31 271 51 305
rect 85 271 137 305
rect 171 271 187 305
rect 221 271 284 305
rect 318 271 366 305
rect 31 242 87 271
rect 221 242 366 271
rect 121 225 187 237
rect 35 192 87 208
rect 35 158 51 192
rect 85 158 87 192
rect 35 111 87 158
rect 121 191 137 225
rect 171 206 187 225
rect 400 206 451 339
rect 490 271 524 305
rect 558 271 610 305
rect 644 271 754 305
rect 490 242 754 271
rect 788 271 804 305
rect 838 271 943 305
rect 788 242 943 271
rect 171 202 451 206
rect 171 191 325 202
rect 121 168 325 191
rect 359 168 451 202
rect 121 164 451 168
rect 485 192 657 208
rect 121 153 187 164
rect 121 119 137 153
rect 171 119 187 153
rect 519 174 657 192
rect 691 174 829 208
rect 863 174 879 208
rect 519 158 521 174
rect 485 130 521 158
rect 221 122 521 130
rect 35 77 51 111
rect 85 85 87 111
rect 221 114 411 122
rect 221 85 227 114
rect 85 80 227 85
rect 261 88 411 114
rect 445 111 521 122
rect 445 88 485 111
rect 261 80 485 88
rect 85 77 485 80
rect 519 77 521 111
rect 35 51 521 77
rect 555 132 621 140
rect 555 98 571 132
rect 605 98 621 132
rect 555 17 621 98
rect 657 113 693 174
rect 691 79 693 113
rect 657 63 693 79
rect 727 132 793 140
rect 727 98 743 132
rect 777 98 793 132
rect 727 17 793 98
rect 827 113 879 174
rect 827 79 829 113
rect 863 79 879 113
rect 827 63 879 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o22ai_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1325670
string GDS_START 1316686
<< end >>
