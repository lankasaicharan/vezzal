magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 23 49 1517 241
rect 0 0 1536 49
<< scnmos >>
rect 102 47 132 215
rect 188 47 218 215
rect 274 47 304 215
rect 376 47 406 215
rect 462 47 492 215
rect 548 47 578 215
rect 738 47 768 215
rect 824 47 854 215
rect 910 47 940 215
rect 996 47 1026 215
rect 1150 47 1180 215
rect 1236 47 1266 215
rect 1322 47 1352 215
rect 1408 47 1438 215
<< scpmoshvt >>
rect 102 367 132 619
rect 188 367 218 619
rect 274 367 304 619
rect 360 367 390 619
rect 495 367 525 619
rect 581 367 611 619
rect 735 367 765 619
rect 821 367 851 619
rect 910 367 940 619
rect 996 367 1026 619
rect 1097 367 1127 619
rect 1183 367 1213 619
rect 1269 367 1299 619
rect 1355 367 1385 619
<< ndiff >>
rect 49 203 102 215
rect 49 169 57 203
rect 91 169 102 203
rect 49 101 102 169
rect 49 67 57 101
rect 91 67 102 101
rect 49 47 102 67
rect 132 175 188 215
rect 132 141 143 175
rect 177 141 188 175
rect 132 93 188 141
rect 132 59 143 93
rect 177 59 188 93
rect 132 47 188 59
rect 218 203 274 215
rect 218 169 229 203
rect 263 169 274 203
rect 218 101 274 169
rect 218 67 229 101
rect 263 67 274 101
rect 218 47 274 67
rect 304 92 376 215
rect 304 58 315 92
rect 349 58 376 92
rect 304 47 376 58
rect 406 162 462 215
rect 406 128 417 162
rect 451 128 462 162
rect 406 91 462 128
rect 406 57 417 91
rect 451 57 462 91
rect 406 47 462 57
rect 492 171 548 215
rect 492 137 503 171
rect 537 137 548 171
rect 492 47 548 137
rect 578 187 631 215
rect 578 153 589 187
rect 623 153 631 187
rect 578 101 631 153
rect 578 67 589 101
rect 623 67 631 101
rect 578 47 631 67
rect 685 95 738 215
rect 685 61 693 95
rect 727 61 738 95
rect 685 47 738 61
rect 768 93 824 215
rect 768 59 779 93
rect 813 59 824 93
rect 768 47 824 59
rect 854 175 910 215
rect 854 141 865 175
rect 899 141 910 175
rect 854 47 910 141
rect 940 167 996 215
rect 940 133 951 167
rect 985 133 996 167
rect 940 93 996 133
rect 940 59 951 93
rect 985 59 996 93
rect 940 47 996 59
rect 1026 167 1150 215
rect 1026 133 1037 167
rect 1071 133 1105 167
rect 1139 133 1150 167
rect 1026 93 1150 133
rect 1026 59 1037 93
rect 1071 59 1105 93
rect 1139 59 1150 93
rect 1026 47 1150 59
rect 1180 203 1236 215
rect 1180 169 1191 203
rect 1225 169 1236 203
rect 1180 101 1236 169
rect 1180 67 1191 101
rect 1225 67 1236 101
rect 1180 47 1236 67
rect 1266 172 1322 215
rect 1266 138 1277 172
rect 1311 138 1322 172
rect 1266 89 1322 138
rect 1266 55 1277 89
rect 1311 55 1322 89
rect 1266 47 1322 55
rect 1352 203 1408 215
rect 1352 169 1363 203
rect 1397 169 1408 203
rect 1352 101 1408 169
rect 1352 67 1363 101
rect 1397 67 1408 101
rect 1352 47 1408 67
rect 1438 172 1491 215
rect 1438 138 1449 172
rect 1483 138 1491 172
rect 1438 93 1491 138
rect 1438 59 1449 93
rect 1483 59 1491 93
rect 1438 47 1491 59
<< pdiff >>
rect 49 607 102 619
rect 49 573 57 607
rect 91 573 102 607
rect 49 502 102 573
rect 49 468 57 502
rect 91 468 102 502
rect 49 413 102 468
rect 49 379 57 413
rect 91 379 102 413
rect 49 367 102 379
rect 132 584 188 619
rect 132 550 143 584
rect 177 550 188 584
rect 132 367 188 550
rect 218 424 274 619
rect 218 390 229 424
rect 263 390 274 424
rect 218 367 274 390
rect 304 584 360 619
rect 304 550 315 584
rect 349 550 360 584
rect 304 367 360 550
rect 390 610 495 619
rect 390 576 401 610
rect 435 576 495 610
rect 390 545 495 576
rect 390 511 450 545
rect 484 511 495 545
rect 390 477 495 511
rect 390 443 450 477
rect 484 443 495 477
rect 390 409 495 443
rect 390 375 450 409
rect 484 375 495 409
rect 390 367 495 375
rect 525 599 581 619
rect 525 565 536 599
rect 570 565 581 599
rect 525 504 581 565
rect 525 470 536 504
rect 570 470 581 504
rect 525 413 581 470
rect 525 379 536 413
rect 570 379 581 413
rect 525 367 581 379
rect 611 595 735 619
rect 611 561 622 595
rect 656 561 690 595
rect 724 561 735 595
rect 611 367 735 561
rect 765 436 821 619
rect 765 402 776 436
rect 810 402 821 436
rect 765 367 821 402
rect 851 595 910 619
rect 851 561 862 595
rect 896 561 910 595
rect 851 367 910 561
rect 940 436 996 619
rect 940 402 951 436
rect 985 402 996 436
rect 940 367 996 402
rect 1026 595 1097 619
rect 1026 561 1037 595
rect 1071 561 1097 595
rect 1026 367 1097 561
rect 1127 599 1183 619
rect 1127 565 1138 599
rect 1172 565 1183 599
rect 1127 508 1183 565
rect 1127 474 1138 508
rect 1172 474 1183 508
rect 1127 413 1183 474
rect 1127 379 1138 413
rect 1172 379 1183 413
rect 1127 367 1183 379
rect 1213 607 1269 619
rect 1213 573 1224 607
rect 1258 573 1269 607
rect 1213 532 1269 573
rect 1213 498 1224 532
rect 1258 498 1269 532
rect 1213 453 1269 498
rect 1213 419 1224 453
rect 1258 419 1269 453
rect 1213 367 1269 419
rect 1299 599 1355 619
rect 1299 565 1310 599
rect 1344 565 1355 599
rect 1299 508 1355 565
rect 1299 474 1310 508
rect 1344 474 1355 508
rect 1299 413 1355 474
rect 1299 379 1310 413
rect 1344 379 1355 413
rect 1299 367 1355 379
rect 1385 607 1438 619
rect 1385 573 1396 607
rect 1430 573 1438 607
rect 1385 532 1438 573
rect 1385 498 1396 532
rect 1430 498 1438 532
rect 1385 453 1438 498
rect 1385 419 1396 453
rect 1430 419 1438 453
rect 1385 367 1438 419
<< ndiffc >>
rect 57 169 91 203
rect 57 67 91 101
rect 143 141 177 175
rect 143 59 177 93
rect 229 169 263 203
rect 229 67 263 101
rect 315 58 349 92
rect 417 128 451 162
rect 417 57 451 91
rect 503 137 537 171
rect 589 153 623 187
rect 589 67 623 101
rect 693 61 727 95
rect 779 59 813 93
rect 865 141 899 175
rect 951 133 985 167
rect 951 59 985 93
rect 1037 133 1071 167
rect 1105 133 1139 167
rect 1037 59 1071 93
rect 1105 59 1139 93
rect 1191 169 1225 203
rect 1191 67 1225 101
rect 1277 138 1311 172
rect 1277 55 1311 89
rect 1363 169 1397 203
rect 1363 67 1397 101
rect 1449 138 1483 172
rect 1449 59 1483 93
<< pdiffc >>
rect 57 573 91 607
rect 57 468 91 502
rect 57 379 91 413
rect 143 550 177 584
rect 229 390 263 424
rect 315 550 349 584
rect 401 576 435 610
rect 450 511 484 545
rect 450 443 484 477
rect 450 375 484 409
rect 536 565 570 599
rect 536 470 570 504
rect 536 379 570 413
rect 622 561 656 595
rect 690 561 724 595
rect 776 402 810 436
rect 862 561 896 595
rect 951 402 985 436
rect 1037 561 1071 595
rect 1138 565 1172 599
rect 1138 474 1172 508
rect 1138 379 1172 413
rect 1224 573 1258 607
rect 1224 498 1258 532
rect 1224 419 1258 453
rect 1310 565 1344 599
rect 1310 474 1344 508
rect 1310 379 1344 413
rect 1396 573 1430 607
rect 1396 498 1430 532
rect 1396 419 1430 453
<< poly >>
rect 102 619 132 645
rect 188 619 218 645
rect 274 619 304 645
rect 360 619 390 645
rect 495 619 525 645
rect 581 619 611 645
rect 735 619 765 645
rect 821 619 851 645
rect 910 619 940 645
rect 996 619 1026 645
rect 1097 619 1127 645
rect 1183 619 1213 645
rect 1269 619 1299 645
rect 1355 619 1385 645
rect 102 335 132 367
rect 66 319 132 335
rect 66 285 82 319
rect 116 285 132 319
rect 66 269 132 285
rect 102 215 132 269
rect 188 335 218 367
rect 274 335 304 367
rect 360 335 390 367
rect 188 319 304 335
rect 188 285 213 319
rect 247 285 304 319
rect 188 269 304 285
rect 353 319 419 335
rect 353 285 369 319
rect 403 285 419 319
rect 495 303 525 367
rect 581 303 611 367
rect 735 303 765 367
rect 821 345 851 367
rect 910 345 940 367
rect 821 319 940 345
rect 821 315 885 319
rect 353 269 419 285
rect 462 287 636 303
rect 188 215 218 269
rect 274 215 304 269
rect 376 215 406 269
rect 462 253 586 287
rect 620 253 636 287
rect 462 237 636 253
rect 713 287 779 303
rect 713 253 729 287
rect 763 253 779 287
rect 713 237 779 253
rect 824 285 885 315
rect 919 285 940 319
rect 996 303 1026 367
rect 1097 331 1127 367
rect 1183 331 1213 367
rect 1269 331 1299 367
rect 1355 331 1385 367
rect 1097 315 1438 331
rect 824 237 940 285
rect 982 287 1048 303
rect 982 253 998 287
rect 1032 253 1048 287
rect 1097 281 1113 315
rect 1147 281 1181 315
rect 1215 281 1249 315
rect 1283 281 1317 315
rect 1351 281 1385 315
rect 1419 281 1438 315
rect 1097 265 1438 281
rect 982 237 1048 253
rect 462 215 492 237
rect 548 215 578 237
rect 738 215 768 237
rect 824 215 854 237
rect 910 215 940 237
rect 996 215 1026 237
rect 1150 215 1180 265
rect 1236 215 1266 265
rect 1322 215 1352 265
rect 1408 215 1438 265
rect 102 21 132 47
rect 188 21 218 47
rect 274 21 304 47
rect 376 21 406 47
rect 462 21 492 47
rect 548 21 578 47
rect 738 21 768 47
rect 824 21 854 47
rect 910 21 940 47
rect 996 21 1026 47
rect 1150 21 1180 47
rect 1236 21 1266 47
rect 1322 21 1352 47
rect 1408 21 1438 47
<< polycont >>
rect 82 285 116 319
rect 213 285 247 319
rect 369 285 403 319
rect 586 253 620 287
rect 729 253 763 287
rect 885 285 919 319
rect 998 253 1032 287
rect 1113 281 1147 315
rect 1181 281 1215 315
rect 1249 281 1283 315
rect 1317 281 1351 315
rect 1385 281 1419 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 41 607 91 649
rect 41 573 57 607
rect 387 610 484 649
rect 41 502 91 573
rect 125 584 353 600
rect 125 550 143 584
rect 177 550 315 584
rect 349 550 353 584
rect 125 534 353 550
rect 387 576 401 610
rect 435 576 484 610
rect 387 545 484 576
rect 387 534 450 545
rect 41 468 57 502
rect 439 511 450 534
rect 41 413 91 468
rect 41 379 57 413
rect 41 363 91 379
rect 125 462 405 500
rect 125 329 163 462
rect 197 424 333 428
rect 197 390 229 424
rect 263 390 333 424
rect 197 386 333 390
rect 66 319 163 329
rect 66 285 82 319
rect 116 285 163 319
rect 66 281 163 285
rect 197 319 263 352
rect 197 285 213 319
rect 247 285 263 319
rect 197 281 263 285
rect 41 213 263 247
rect 41 203 93 213
rect 41 169 57 203
rect 91 169 93 203
rect 227 203 263 213
rect 41 101 93 169
rect 41 67 57 101
rect 91 67 93 101
rect 41 51 93 67
rect 127 175 193 179
rect 127 141 143 175
rect 177 141 193 175
rect 127 93 193 141
rect 127 59 143 93
rect 177 59 193 93
rect 127 17 193 59
rect 227 169 229 203
rect 297 235 333 386
rect 369 330 405 462
rect 439 477 484 511
rect 439 443 450 477
rect 439 409 484 443
rect 439 375 450 409
rect 439 359 484 375
rect 518 599 572 615
rect 518 565 536 599
rect 570 565 572 599
rect 518 522 572 565
rect 606 595 740 649
rect 606 561 622 595
rect 656 561 690 595
rect 724 561 740 595
rect 606 556 740 561
rect 846 595 912 649
rect 846 561 862 595
rect 896 561 912 595
rect 846 556 912 561
rect 1021 595 1087 649
rect 1021 561 1037 595
rect 1071 561 1087 595
rect 1021 556 1087 561
rect 1136 599 1174 615
rect 1136 565 1138 599
rect 1172 565 1174 599
rect 518 504 1102 522
rect 518 470 536 504
rect 570 486 1102 504
rect 570 470 586 486
rect 518 413 586 470
rect 518 379 536 413
rect 570 379 586 413
rect 518 346 586 379
rect 659 436 989 452
rect 659 402 776 436
rect 810 402 951 436
rect 985 402 989 436
rect 659 386 989 402
rect 369 319 419 330
rect 403 285 419 319
rect 369 269 419 285
rect 518 235 552 346
rect 659 303 695 386
rect 869 319 950 352
rect 586 287 695 303
rect 620 253 695 287
rect 586 237 695 253
rect 297 199 552 235
rect 227 165 263 169
rect 501 171 552 199
rect 227 162 467 165
rect 227 131 417 162
rect 227 101 265 131
rect 227 67 229 101
rect 263 67 265 101
rect 401 128 417 131
rect 451 128 467 162
rect 227 51 265 67
rect 299 92 365 97
rect 299 58 315 92
rect 349 58 365 92
rect 299 17 365 58
rect 401 91 467 128
rect 501 137 503 171
rect 537 137 552 171
rect 501 121 552 137
rect 586 187 625 203
rect 586 153 589 187
rect 623 153 625 187
rect 401 57 417 91
rect 451 87 467 91
rect 586 101 625 153
rect 659 183 695 237
rect 729 287 835 303
rect 763 253 835 287
rect 869 285 885 319
rect 919 285 950 319
rect 1068 315 1102 486
rect 1136 508 1174 565
rect 1136 474 1138 508
rect 1172 474 1174 508
rect 1136 413 1174 474
rect 1208 607 1274 649
rect 1208 573 1224 607
rect 1258 573 1274 607
rect 1208 532 1274 573
rect 1208 498 1224 532
rect 1258 498 1274 532
rect 1208 453 1274 498
rect 1208 419 1224 453
rect 1258 419 1274 453
rect 1308 599 1344 615
rect 1308 565 1310 599
rect 1308 508 1344 565
rect 1308 474 1310 508
rect 1136 379 1138 413
rect 1172 385 1174 413
rect 1308 413 1344 474
rect 1380 607 1446 649
rect 1380 573 1396 607
rect 1430 573 1446 607
rect 1380 532 1446 573
rect 1380 498 1396 532
rect 1430 498 1446 532
rect 1380 453 1446 498
rect 1380 419 1396 453
rect 1430 419 1446 453
rect 1308 385 1310 413
rect 1172 379 1310 385
rect 1344 379 1519 385
rect 1136 349 1519 379
rect 984 287 1034 303
rect 729 251 835 253
rect 984 253 998 287
rect 1032 253 1034 287
rect 1068 281 1113 315
rect 1147 281 1181 315
rect 1215 281 1249 315
rect 1283 281 1317 315
rect 1351 281 1385 315
rect 1419 281 1435 315
rect 984 251 1034 253
rect 729 217 1034 251
rect 1469 247 1519 349
rect 1175 209 1519 247
rect 1175 203 1227 209
rect 659 175 915 183
rect 659 145 865 175
rect 849 141 865 145
rect 899 141 915 175
rect 849 131 915 141
rect 949 167 1001 183
rect 949 133 951 167
rect 985 133 1001 167
rect 586 87 589 101
rect 451 67 589 87
rect 623 67 625 101
rect 451 57 625 67
rect 401 51 625 57
rect 677 95 729 111
rect 949 97 1001 133
rect 677 61 693 95
rect 727 61 729 95
rect 677 17 729 61
rect 763 93 1001 97
rect 763 59 779 93
rect 813 59 951 93
rect 985 59 1001 93
rect 763 51 1001 59
rect 1035 167 1141 183
rect 1035 133 1037 167
rect 1071 133 1105 167
rect 1139 133 1141 167
rect 1035 93 1141 133
rect 1035 59 1037 93
rect 1071 59 1105 93
rect 1139 59 1141 93
rect 1035 17 1141 59
rect 1175 169 1191 203
rect 1225 169 1227 203
rect 1361 203 1399 209
rect 1175 101 1227 169
rect 1175 67 1191 101
rect 1225 67 1227 101
rect 1175 51 1227 67
rect 1261 172 1327 175
rect 1261 138 1277 172
rect 1311 138 1327 172
rect 1261 89 1327 138
rect 1261 55 1277 89
rect 1311 55 1327 89
rect 1261 17 1327 55
rect 1361 169 1363 203
rect 1397 169 1399 203
rect 1361 101 1399 169
rect 1361 67 1363 101
rect 1397 67 1399 101
rect 1361 51 1399 67
rect 1433 172 1499 175
rect 1433 138 1449 172
rect 1483 138 1499 172
rect 1433 93 1499 138
rect 1433 59 1449 93
rect 1483 59 1499 93
rect 1433 17 1499 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2bb2a_4
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3617080
string GDS_START 3604870
<< end >>
