magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 4274 1975
<< nwell >>
rect -38 332 3014 704
<< pwell >>
rect 582 191 877 248
rect 582 184 1314 191
rect 1535 184 2117 228
rect 2585 184 2975 252
rect 1 49 2975 184
rect 0 0 2976 49
<< scpmos >>
rect 83 464 119 592
rect 173 464 209 592
rect 257 464 293 592
rect 383 464 419 592
rect 467 464 503 592
rect 679 368 715 592
rect 769 368 805 592
rect 977 457 1013 541
rect 1084 483 1120 567
rect 1188 463 1224 547
rect 1325 463 1361 547
rect 1424 463 1460 547
rect 1551 379 1587 547
rect 1641 379 1677 547
rect 1870 424 1906 592
rect 1960 424 1996 592
rect 2108 508 2144 592
rect 2186 508 2222 592
rect 2276 508 2312 592
rect 2472 508 2508 592
rect 2668 392 2704 592
rect 2769 368 2805 592
rect 2859 368 2895 592
<< nmoslvt >>
rect 84 74 114 158
rect 209 74 239 158
rect 287 74 317 158
rect 373 74 403 158
rect 467 74 497 158
rect 665 74 695 222
rect 765 74 795 222
rect 961 81 991 165
rect 1113 81 1143 165
rect 1185 81 1215 165
rect 1399 74 1429 158
rect 1477 74 1507 158
rect 1611 74 1641 202
rect 1697 74 1727 202
rect 1925 74 1955 202
rect 2011 74 2041 202
rect 2111 74 2141 158
rect 2189 74 2219 158
rect 2303 74 2333 158
rect 2470 74 2500 158
rect 2668 98 2698 226
rect 2773 78 2803 226
rect 2859 78 2889 226
<< ndiff >>
rect 608 202 665 222
rect 608 168 620 202
rect 654 168 665 202
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 120 209 158
rect 114 86 151 120
rect 185 86 209 120
rect 114 74 209 86
rect 239 74 287 158
rect 317 133 373 158
rect 317 99 328 133
rect 362 99 373 133
rect 317 74 373 99
rect 403 74 467 158
rect 497 126 554 158
rect 497 92 508 126
rect 542 92 554 126
rect 497 74 554 92
rect 608 120 665 168
rect 608 86 620 120
rect 654 86 665 120
rect 608 74 665 86
rect 695 202 765 222
rect 695 168 720 202
rect 754 168 765 202
rect 695 120 765 168
rect 695 86 720 120
rect 754 86 765 120
rect 695 74 765 86
rect 795 210 851 222
rect 795 176 806 210
rect 840 176 851 210
rect 795 120 851 176
rect 795 86 806 120
rect 840 86 851 120
rect 795 74 851 86
rect 905 153 961 165
rect 905 119 916 153
rect 950 119 961 153
rect 905 81 961 119
rect 991 140 1113 165
rect 991 106 1068 140
rect 1102 106 1113 140
rect 991 81 1113 106
rect 1143 81 1185 165
rect 1215 81 1288 165
rect 1561 158 1611 202
rect 1230 72 1288 81
rect 1342 122 1399 158
rect 1342 88 1354 122
rect 1388 88 1399 122
rect 1342 74 1399 88
rect 1429 74 1477 158
rect 1507 120 1611 158
rect 1507 86 1535 120
rect 1569 86 1611 120
rect 1507 74 1611 86
rect 1641 190 1697 202
rect 1641 156 1652 190
rect 1686 156 1697 190
rect 1641 120 1697 156
rect 1641 86 1652 120
rect 1686 86 1697 120
rect 1641 74 1697 86
rect 1727 123 1800 202
rect 1727 89 1754 123
rect 1788 89 1800 123
rect 1727 74 1800 89
rect 1854 123 1925 202
rect 1854 89 1866 123
rect 1900 89 1925 123
rect 1854 74 1925 89
rect 1955 179 2011 202
rect 1955 145 1966 179
rect 2000 145 2011 179
rect 1955 74 2011 145
rect 2041 158 2091 202
rect 2611 214 2668 226
rect 2611 180 2623 214
rect 2657 180 2668 214
rect 2041 133 2111 158
rect 2041 99 2066 133
rect 2100 99 2111 133
rect 2041 74 2111 99
rect 2141 74 2189 158
rect 2219 74 2303 158
rect 2333 120 2470 158
rect 2333 86 2344 120
rect 2378 86 2416 120
rect 2450 86 2470 120
rect 2333 74 2470 86
rect 2500 133 2557 158
rect 2500 99 2511 133
rect 2545 99 2557 133
rect 2500 74 2557 99
rect 2611 144 2668 180
rect 2611 110 2623 144
rect 2657 110 2668 144
rect 2611 98 2668 110
rect 2698 214 2773 226
rect 2698 180 2727 214
rect 2761 180 2773 214
rect 2698 124 2773 180
rect 2698 98 2727 124
rect 1230 38 1242 72
rect 1276 38 1288 72
rect 2715 90 2727 98
rect 2761 90 2773 124
rect 2715 78 2773 90
rect 2803 214 2859 226
rect 2803 180 2814 214
rect 2848 180 2859 214
rect 2803 124 2859 180
rect 2803 90 2814 124
rect 2848 90 2859 124
rect 2803 78 2859 90
rect 2889 214 2949 226
rect 2889 180 2903 214
rect 2937 180 2949 214
rect 2889 122 2949 180
rect 2889 88 2903 122
rect 2937 88 2949 122
rect 2889 78 2949 88
rect 1230 27 1288 38
<< pdiff >>
rect 518 616 571 628
rect 518 592 528 616
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 512 83 546
rect 27 478 39 512
rect 73 478 83 512
rect 27 464 83 478
rect 119 573 173 592
rect 119 539 129 573
rect 163 539 173 573
rect 119 464 173 539
rect 209 464 257 592
rect 293 566 383 592
rect 293 532 321 566
rect 355 532 383 566
rect 293 464 383 532
rect 419 464 467 592
rect 503 582 528 592
rect 562 582 571 616
rect 503 464 571 582
rect 625 414 679 592
rect 625 380 635 414
rect 669 380 679 414
rect 625 368 679 380
rect 715 573 769 592
rect 715 539 725 573
rect 759 539 769 573
rect 715 368 769 539
rect 805 573 861 592
rect 805 539 815 573
rect 849 539 861 573
rect 805 520 861 539
rect 805 368 855 520
rect 1804 580 1870 592
rect 1034 541 1084 567
rect 921 516 977 541
rect 921 482 933 516
rect 967 482 977 516
rect 921 457 977 482
rect 1013 516 1084 541
rect 1013 482 1023 516
rect 1057 483 1084 516
rect 1120 547 1170 567
rect 1120 483 1188 547
rect 1057 482 1069 483
rect 1013 457 1069 482
rect 1138 463 1188 483
rect 1224 535 1325 547
rect 1224 501 1235 535
rect 1269 501 1325 535
rect 1224 463 1325 501
rect 1361 520 1424 547
rect 1361 486 1371 520
rect 1405 486 1424 520
rect 1361 463 1424 486
rect 1460 531 1551 547
rect 1460 497 1507 531
rect 1541 497 1551 531
rect 1460 463 1551 497
rect 1495 429 1507 463
rect 1541 429 1551 463
rect 1495 379 1551 429
rect 1587 535 1641 547
rect 1587 501 1597 535
rect 1631 501 1641 535
rect 1587 463 1641 501
rect 1587 429 1597 463
rect 1631 429 1641 463
rect 1587 379 1641 429
rect 1677 533 1730 547
rect 1677 499 1687 533
rect 1721 499 1730 533
rect 1677 379 1730 499
rect 1804 546 1816 580
rect 1850 546 1870 580
rect 1804 497 1870 546
rect 1804 463 1816 497
rect 1850 463 1870 497
rect 1804 424 1870 463
rect 1906 547 1960 592
rect 1906 513 1916 547
rect 1950 513 1960 547
rect 1906 470 1960 513
rect 1906 436 1916 470
rect 1950 436 1960 470
rect 1906 424 1960 436
rect 1996 566 2108 592
rect 1996 532 2037 566
rect 2071 532 2108 566
rect 1996 508 2108 532
rect 2144 508 2186 592
rect 2222 579 2276 592
rect 2222 545 2232 579
rect 2266 545 2276 579
rect 2222 508 2276 545
rect 2312 567 2365 592
rect 2312 533 2322 567
rect 2356 533 2365 567
rect 2312 508 2365 533
rect 2419 567 2472 592
rect 2419 533 2428 567
rect 2462 533 2472 567
rect 2419 508 2472 533
rect 2508 580 2561 592
rect 2508 546 2518 580
rect 2552 546 2561 580
rect 2508 508 2561 546
rect 2615 580 2668 592
rect 2615 546 2624 580
rect 2658 546 2668 580
rect 2615 509 2668 546
rect 1996 424 2046 508
rect 2615 475 2624 509
rect 2658 475 2668 509
rect 2615 438 2668 475
rect 2615 404 2624 438
rect 2658 404 2668 438
rect 2615 392 2668 404
rect 2704 580 2769 592
rect 2704 546 2724 580
rect 2758 546 2769 580
rect 2704 505 2769 546
rect 2704 471 2724 505
rect 2758 471 2769 505
rect 2704 434 2769 471
rect 2704 400 2724 434
rect 2758 400 2769 434
rect 2704 392 2769 400
rect 2719 368 2769 392
rect 2805 580 2859 592
rect 2805 546 2815 580
rect 2849 546 2859 580
rect 2805 499 2859 546
rect 2805 465 2815 499
rect 2849 465 2859 499
rect 2805 414 2859 465
rect 2805 380 2815 414
rect 2849 380 2859 414
rect 2805 368 2859 380
rect 2895 580 2949 592
rect 2895 546 2905 580
rect 2939 546 2949 580
rect 2895 498 2949 546
rect 2895 464 2905 498
rect 2939 464 2949 498
rect 2895 368 2949 464
<< ndiffc >>
rect 620 168 654 202
rect 39 99 73 133
rect 151 86 185 120
rect 328 99 362 133
rect 508 92 542 126
rect 620 86 654 120
rect 720 168 754 202
rect 720 86 754 120
rect 806 176 840 210
rect 806 86 840 120
rect 916 119 950 153
rect 1068 106 1102 140
rect 1354 88 1388 122
rect 1535 86 1569 120
rect 1652 156 1686 190
rect 1652 86 1686 120
rect 1754 89 1788 123
rect 1866 89 1900 123
rect 1966 145 2000 179
rect 2623 180 2657 214
rect 2066 99 2100 133
rect 2344 86 2378 120
rect 2416 86 2450 120
rect 2511 99 2545 133
rect 2623 110 2657 144
rect 2727 180 2761 214
rect 1242 38 1276 72
rect 2727 90 2761 124
rect 2814 180 2848 214
rect 2814 90 2848 124
rect 2903 180 2937 214
rect 2903 88 2937 122
<< pdiffc >>
rect 39 546 73 580
rect 39 478 73 512
rect 129 539 163 573
rect 321 532 355 566
rect 528 582 562 616
rect 635 380 669 414
rect 725 539 759 573
rect 815 539 849 573
rect 933 482 967 516
rect 1023 482 1057 516
rect 1235 501 1269 535
rect 1371 486 1405 520
rect 1507 497 1541 531
rect 1507 429 1541 463
rect 1597 501 1631 535
rect 1597 429 1631 463
rect 1687 499 1721 533
rect 1816 546 1850 580
rect 1816 463 1850 497
rect 1916 513 1950 547
rect 1916 436 1950 470
rect 2037 532 2071 566
rect 2232 545 2266 579
rect 2322 533 2356 567
rect 2428 533 2462 567
rect 2518 546 2552 580
rect 2624 546 2658 580
rect 2624 475 2658 509
rect 2624 404 2658 438
rect 2724 546 2758 580
rect 2724 471 2758 505
rect 2724 400 2758 434
rect 2815 546 2849 580
rect 2815 465 2849 499
rect 2815 380 2849 414
rect 2905 546 2939 580
rect 2905 464 2939 498
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 257 592 293 618
rect 383 592 419 618
rect 467 592 503 618
rect 679 592 715 618
rect 769 592 805 618
rect 876 615 1996 645
rect 83 428 119 464
rect 173 428 209 464
rect 257 430 293 464
rect 383 432 419 464
rect 83 412 209 428
rect 83 378 111 412
rect 145 398 209 412
rect 251 414 317 430
rect 145 378 161 398
rect 83 344 161 378
rect 251 380 267 414
rect 301 380 317 414
rect 251 364 317 380
rect 359 416 425 432
rect 359 382 375 416
rect 409 382 425 416
rect 359 366 425 382
rect 467 430 503 464
rect 467 414 566 430
rect 467 380 516 414
rect 550 380 566 414
rect 83 310 111 344
rect 145 310 161 344
rect 83 294 161 310
rect 84 158 114 294
rect 179 230 245 246
rect 179 196 195 230
rect 229 196 245 230
rect 179 180 245 196
rect 209 158 239 180
rect 287 158 317 364
rect 467 346 566 380
rect 876 424 906 615
rect 1084 567 1120 615
rect 1870 592 1906 615
rect 1960 592 1996 615
rect 2108 592 2144 618
rect 2186 592 2222 618
rect 2276 592 2312 618
rect 2472 592 2508 618
rect 2668 592 2704 618
rect 2769 592 2805 618
rect 2859 592 2895 618
rect 977 541 1013 567
rect 1188 547 1224 573
rect 1325 547 1361 573
rect 1424 547 1460 573
rect 1551 547 1587 573
rect 1641 547 1677 573
rect 1084 457 1120 483
rect 870 394 906 424
rect 359 300 425 316
rect 359 266 375 300
rect 409 266 425 300
rect 359 250 425 266
rect 467 312 516 346
rect 550 312 566 346
rect 467 278 566 312
rect 679 310 715 368
rect 769 336 805 368
rect 870 336 900 394
rect 977 346 1013 457
rect 1080 393 1146 409
rect 1080 359 1096 393
rect 1130 359 1146 393
rect 1080 346 1146 359
rect 765 320 900 336
rect 373 158 403 250
rect 467 244 516 278
rect 550 244 566 278
rect 651 294 717 310
rect 651 260 667 294
rect 701 260 717 294
rect 651 244 717 260
rect 765 286 793 320
rect 827 286 900 320
rect 765 270 900 286
rect 942 330 1146 346
rect 1188 396 1224 463
rect 1188 380 1254 396
rect 1188 346 1204 380
rect 1238 346 1254 380
rect 1188 330 1254 346
rect 942 296 958 330
rect 992 316 1146 330
rect 992 296 1013 316
rect 942 280 1013 296
rect 467 228 566 244
rect 467 158 497 228
rect 665 222 695 244
rect 765 222 795 270
rect 870 238 900 270
rect 1107 252 1143 316
rect 870 208 991 238
rect 961 165 991 208
rect 1113 165 1143 252
rect 1196 253 1226 330
rect 1325 314 1361 463
rect 1310 298 1376 314
rect 1310 264 1326 298
rect 1360 264 1376 298
rect 1196 237 1262 253
rect 1196 217 1212 237
rect 1185 203 1212 217
rect 1246 203 1262 237
rect 1185 187 1262 203
rect 1310 230 1376 264
rect 1424 311 1460 463
rect 2108 427 2144 508
rect 1551 311 1587 379
rect 1641 311 1677 379
rect 1424 295 1507 311
rect 1424 261 1457 295
rect 1491 261 1507 295
rect 1424 245 1507 261
rect 1551 295 1677 311
rect 1762 345 1828 361
rect 1762 311 1778 345
rect 1812 311 1828 345
rect 1762 295 1828 311
rect 1551 261 1567 295
rect 1601 261 1677 295
rect 1551 247 1677 261
rect 1798 247 1828 295
rect 1870 319 1906 424
rect 1960 398 1996 424
rect 2078 411 2144 427
rect 2078 377 2094 411
rect 2128 377 2144 411
rect 2078 361 2144 377
rect 2186 367 2222 508
rect 1870 289 2141 319
rect 1551 245 1727 247
rect 1310 196 1326 230
rect 1360 203 1376 230
rect 1360 196 1429 203
rect 1185 165 1215 187
rect 1310 173 1429 196
rect 1399 158 1429 173
rect 1477 158 1507 245
rect 1611 217 1727 245
rect 1798 217 2041 247
rect 1611 202 1641 217
rect 1697 202 1727 217
rect 1925 202 1955 217
rect 2011 202 2041 217
rect 84 48 114 74
rect 209 48 239 74
rect 287 48 317 74
rect 373 48 403 74
rect 467 48 497 74
rect 665 48 695 74
rect 765 48 795 74
rect 961 55 991 81
rect 1113 55 1143 81
rect 1185 55 1215 81
rect 2111 158 2141 289
rect 2192 246 2222 367
rect 2276 360 2312 508
rect 2472 428 2508 508
rect 2427 412 2508 428
rect 2427 378 2443 412
rect 2477 398 2508 412
rect 2477 378 2502 398
rect 2276 344 2355 360
rect 2276 310 2305 344
rect 2339 310 2355 344
rect 2276 294 2355 310
rect 2427 344 2502 378
rect 2427 310 2443 344
rect 2477 310 2502 344
rect 2427 305 2502 310
rect 2668 305 2704 392
rect 2769 330 2805 368
rect 2859 330 2895 368
rect 2189 230 2255 246
rect 2189 196 2205 230
rect 2239 196 2255 230
rect 2189 180 2255 196
rect 2189 158 2219 180
rect 2303 158 2333 294
rect 2427 276 2704 305
rect 2427 242 2443 276
rect 2477 242 2704 276
rect 2746 314 2895 330
rect 2746 280 2762 314
rect 2796 280 2895 314
rect 2746 264 2895 280
rect 2427 241 2704 242
rect 2427 226 2502 241
rect 2668 226 2698 241
rect 2773 226 2803 264
rect 2859 241 2895 264
rect 2859 226 2889 241
rect 2470 158 2500 226
rect 1399 48 1429 74
rect 1477 48 1507 74
rect 1611 48 1641 74
rect 1697 48 1727 74
rect 1925 48 1955 74
rect 2011 48 2041 74
rect 2111 48 2141 74
rect 2189 48 2219 74
rect 2303 48 2333 74
rect 2470 48 2500 74
rect 2668 72 2698 98
rect 2773 52 2803 78
rect 2859 52 2889 78
<< polycont >>
rect 111 378 145 412
rect 267 380 301 414
rect 375 382 409 416
rect 516 380 550 414
rect 111 310 145 344
rect 195 196 229 230
rect 375 266 409 300
rect 516 312 550 346
rect 1096 359 1130 393
rect 516 244 550 278
rect 667 260 701 294
rect 793 286 827 320
rect 1204 346 1238 380
rect 958 296 992 330
rect 1326 264 1360 298
rect 1212 203 1246 237
rect 1457 261 1491 295
rect 1778 311 1812 345
rect 1567 261 1601 295
rect 2094 377 2128 411
rect 1326 196 1360 230
rect 2443 378 2477 412
rect 2305 310 2339 344
rect 2443 310 2477 344
rect 2205 196 2239 230
rect 2443 242 2477 276
rect 2762 280 2796 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 23 580 73 596
rect 23 546 39 580
rect 23 512 73 546
rect 113 573 179 649
rect 512 616 578 649
rect 512 582 528 616
rect 562 582 578 616
rect 113 539 129 573
rect 163 539 179 573
rect 113 532 179 539
rect 287 566 477 582
rect 512 566 578 582
rect 709 573 775 649
rect 287 532 321 566
rect 355 532 477 566
rect 709 539 725 573
rect 759 539 775 573
rect 23 478 39 512
rect 443 498 624 532
rect 709 516 775 539
rect 815 579 1146 613
rect 815 573 865 579
rect 849 539 865 573
rect 815 516 865 539
rect 917 516 983 545
rect 73 478 409 498
rect 23 464 409 478
rect 23 462 73 464
rect 23 246 57 462
rect 95 412 161 428
rect 95 378 111 412
rect 145 378 161 412
rect 95 344 161 378
rect 217 414 317 430
rect 217 380 267 414
rect 301 380 317 414
rect 217 364 317 380
rect 359 416 409 464
rect 359 382 375 416
rect 359 366 409 382
rect 95 310 111 344
rect 145 316 161 344
rect 145 310 409 316
rect 95 300 409 310
rect 95 282 375 300
rect 359 266 375 282
rect 359 250 409 266
rect 23 230 245 246
rect 23 196 195 230
rect 229 196 245 230
rect 443 216 477 498
rect 590 482 624 498
rect 917 482 933 516
rect 967 482 983 516
rect 590 448 983 482
rect 1023 516 1073 545
rect 1057 482 1073 516
rect 1023 453 1073 482
rect 511 414 556 430
rect 917 414 983 448
rect 511 380 516 414
rect 550 380 556 414
rect 511 346 556 380
rect 511 312 516 346
rect 550 312 556 346
rect 511 278 556 312
rect 511 244 516 278
rect 550 244 556 278
rect 511 228 556 244
rect 592 380 635 414
rect 669 380 843 414
rect 592 364 843 380
rect 23 180 245 196
rect 312 182 477 216
rect 592 202 626 364
rect 777 320 843 364
rect 660 294 743 310
rect 660 260 667 294
rect 701 260 743 294
rect 777 286 793 320
rect 827 286 843 320
rect 777 270 843 286
rect 884 380 983 414
rect 660 236 743 260
rect 806 210 840 226
rect 23 133 89 180
rect 23 99 39 133
rect 73 99 89 133
rect 23 70 89 99
rect 123 120 214 136
rect 123 86 151 120
rect 185 86 214 120
rect 123 17 214 86
rect 312 133 378 182
rect 592 168 620 202
rect 654 168 670 202
rect 312 99 328 133
rect 362 99 378 133
rect 312 70 378 99
rect 492 126 558 148
rect 492 92 508 126
rect 542 92 558 126
rect 492 17 558 92
rect 592 120 670 168
rect 592 86 620 120
rect 654 86 670 120
rect 592 70 670 86
rect 704 168 720 202
rect 754 168 770 202
rect 704 120 770 168
rect 704 86 720 120
rect 754 86 770 120
rect 704 17 770 86
rect 806 120 840 176
rect 884 169 918 380
rect 952 330 993 346
rect 952 296 958 330
rect 992 296 993 330
rect 952 237 993 296
rect 1027 309 1061 453
rect 1112 451 1146 579
rect 1219 535 1269 649
rect 1219 501 1235 535
rect 1219 485 1269 501
rect 1303 581 1473 615
rect 1303 451 1337 581
rect 1112 417 1337 451
rect 1371 520 1405 547
rect 1112 409 1146 417
rect 1095 393 1146 409
rect 1095 359 1096 393
rect 1130 359 1146 393
rect 1371 383 1405 486
rect 1095 343 1146 359
rect 1188 380 1405 383
rect 1188 346 1204 380
rect 1238 349 1405 380
rect 1439 379 1473 581
rect 1507 531 1541 649
rect 1507 463 1541 497
rect 1507 413 1541 429
rect 1581 535 1647 551
rect 1581 501 1597 535
rect 1631 501 1647 535
rect 1581 463 1647 501
rect 1687 533 1737 649
rect 1721 499 1737 533
rect 1687 481 1737 499
rect 1800 581 2087 615
rect 1800 580 1866 581
rect 1800 546 1816 580
rect 1850 546 1866 580
rect 2021 566 2087 581
rect 1800 497 1866 546
rect 1800 463 1816 497
rect 1850 463 1866 497
rect 1900 513 1916 547
rect 1950 513 1966 547
rect 1900 470 1966 513
rect 1581 429 1597 463
rect 1631 447 1647 463
rect 1631 429 1753 447
rect 1900 436 1916 470
rect 1950 436 1966 470
rect 2021 532 2037 566
rect 2071 532 2087 566
rect 2021 495 2087 532
rect 2216 579 2266 649
rect 2216 545 2232 579
rect 2216 529 2266 545
rect 2306 567 2372 596
rect 2306 533 2322 567
rect 2356 533 2372 567
rect 2306 495 2372 533
rect 2021 461 2372 495
rect 2412 567 2462 596
rect 2412 533 2428 567
rect 2412 496 2462 533
rect 2502 580 2568 649
rect 2502 546 2518 580
rect 2552 546 2568 580
rect 2502 530 2568 546
rect 2607 580 2674 596
rect 2607 546 2624 580
rect 2658 546 2674 580
rect 2607 509 2674 546
rect 2412 462 2561 496
rect 1900 429 1966 436
rect 1581 413 1966 429
rect 2178 428 2372 461
rect 1719 395 1966 413
rect 2000 411 2144 427
rect 1439 361 1685 379
rect 2000 377 2094 411
rect 2128 377 2144 411
rect 2000 361 2144 377
rect 2178 412 2493 428
rect 2178 394 2443 412
rect 1238 346 1254 349
rect 1188 343 1254 346
rect 1439 345 2034 361
rect 1310 309 1376 314
rect 1651 311 1778 345
rect 1812 311 2034 345
rect 2178 314 2212 394
rect 2427 378 2443 394
rect 2477 378 2493 412
rect 1027 298 1376 309
rect 1027 275 1326 298
rect 952 203 1034 237
rect 884 153 966 169
rect 884 119 916 153
rect 950 119 966 153
rect 806 85 840 86
rect 1000 85 1034 203
rect 806 51 1034 85
rect 1068 140 1118 275
rect 1310 264 1326 275
rect 1360 264 1376 298
rect 1102 106 1118 140
rect 1196 237 1262 241
rect 1196 203 1212 237
rect 1246 203 1262 237
rect 1196 140 1262 203
rect 1310 230 1376 264
rect 1441 295 1511 311
rect 1441 261 1457 295
rect 1491 276 1511 295
rect 1441 242 1471 261
rect 1505 242 1511 276
rect 1551 295 1617 311
rect 1651 295 2034 311
rect 1551 261 1567 295
rect 1601 261 1617 295
rect 1551 245 1617 261
rect 2082 280 2212 314
rect 2289 344 2375 360
rect 2289 310 2305 344
rect 2339 310 2375 344
rect 1310 196 1326 230
rect 1360 208 1376 230
rect 1551 208 1585 245
rect 1360 196 1585 208
rect 1310 174 1585 196
rect 1636 190 2016 211
rect 1636 156 1652 190
rect 1686 179 2016 190
rect 1686 177 1966 179
rect 1686 156 1702 177
rect 1196 122 1404 140
rect 1196 106 1354 122
rect 1068 77 1118 106
rect 1338 88 1354 106
rect 1388 88 1404 122
rect 1226 38 1242 72
rect 1276 38 1292 72
rect 1338 70 1404 88
rect 1502 120 1602 136
rect 1502 86 1535 120
rect 1569 86 1602 120
rect 1226 17 1292 38
rect 1502 17 1602 86
rect 1636 120 1702 156
rect 1950 145 1966 177
rect 2000 145 2016 179
rect 2082 162 2116 280
rect 2289 276 2375 310
rect 1636 86 1652 120
rect 1686 86 1702 120
rect 1636 70 1702 86
rect 1738 123 1804 143
rect 1738 89 1754 123
rect 1788 89 1804 123
rect 1738 17 1804 89
rect 1850 123 1916 143
rect 1850 89 1866 123
rect 1900 89 1916 123
rect 1950 119 2016 145
rect 2050 133 2116 162
rect 2189 230 2255 246
rect 2289 242 2335 276
rect 2369 242 2375 276
rect 2289 236 2375 242
rect 2427 344 2493 378
rect 2427 310 2443 344
rect 2477 310 2493 344
rect 2427 276 2493 310
rect 2427 242 2443 276
rect 2477 242 2493 276
rect 2189 196 2205 230
rect 2239 196 2255 230
rect 2427 226 2493 242
rect 2189 192 2255 196
rect 2527 192 2561 462
rect 2189 158 2561 192
rect 1850 85 1916 89
rect 2050 99 2066 133
rect 2100 99 2116 133
rect 2500 133 2561 158
rect 2050 85 2116 99
rect 1850 51 2116 85
rect 2328 86 2344 120
rect 2378 86 2416 120
rect 2450 86 2466 120
rect 2328 17 2466 86
rect 2500 99 2511 133
rect 2545 99 2561 133
rect 2500 70 2561 99
rect 2607 475 2624 509
rect 2658 475 2674 509
rect 2607 438 2674 475
rect 2607 404 2624 438
rect 2658 404 2674 438
rect 2607 330 2674 404
rect 2708 580 2765 649
rect 2708 546 2724 580
rect 2758 546 2765 580
rect 2708 505 2765 546
rect 2708 471 2724 505
rect 2758 471 2765 505
rect 2708 434 2765 471
rect 2708 400 2724 434
rect 2758 400 2765 434
rect 2708 364 2765 400
rect 2799 580 2855 596
rect 2799 546 2815 580
rect 2849 546 2855 580
rect 2799 499 2855 546
rect 2799 465 2815 499
rect 2849 465 2855 499
rect 2799 430 2855 465
rect 2889 580 2955 649
rect 2889 546 2905 580
rect 2939 546 2955 580
rect 2889 498 2955 546
rect 2889 464 2905 498
rect 2939 464 2955 498
rect 2799 414 2951 430
rect 2799 380 2815 414
rect 2849 380 2951 414
rect 2799 364 2951 380
rect 2607 314 2801 330
rect 2607 280 2762 314
rect 2796 280 2801 314
rect 2865 298 2951 364
rect 2607 264 2801 280
rect 2835 264 2951 298
rect 2607 214 2673 264
rect 2835 230 2869 264
rect 2607 180 2623 214
rect 2657 180 2673 214
rect 2607 144 2673 180
rect 2607 110 2623 144
rect 2657 110 2673 144
rect 2607 94 2673 110
rect 2711 214 2761 230
rect 2711 180 2727 214
rect 2711 124 2761 180
rect 2711 90 2727 124
rect 2711 17 2761 90
rect 2798 214 2869 230
rect 2798 180 2814 214
rect 2848 180 2869 214
rect 2798 124 2869 180
rect 2798 90 2814 124
rect 2848 90 2869 124
rect 2798 74 2869 90
rect 2903 214 2953 230
rect 2937 180 2953 214
rect 2903 122 2953 180
rect 2937 88 2953 122
rect 2903 17 2953 88
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 1471 261 1491 276
rect 1491 261 1505 276
rect 1471 242 1505 261
rect 2335 242 2369 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< metal1 >>
rect 0 683 2976 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 0 617 2976 649
rect 1459 276 1517 282
rect 1459 242 1471 276
rect 1505 273 1517 276
rect 2323 276 2381 282
rect 2323 273 2335 276
rect 1505 245 2335 273
rect 1505 242 1517 245
rect 1459 236 1517 242
rect 2323 242 2335 245
rect 2369 242 2381 276
rect 2323 236 2381 242
rect 0 17 2976 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
rect 0 -49 2976 -17
<< labels >>
flabel pwell s 0 0 2976 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2976 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfstp_2
flabel comment s 1209 268 1209 268 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 1021 323 1021 323 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 2335 242 2369 276 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel metal1 s 0 0 2976 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 0 617 2976 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 2911 316 2945 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2911 390 2945 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2976 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 182238
string GDS_START 161308
<< end >>
