magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1778 1975
<< nwell >>
rect -38 331 518 704
<< pwell >>
rect 11 49 479 157
rect 0 0 480 49
<< scnmos >>
rect 90 47 120 131
rect 221 47 251 131
rect 293 47 323 131
rect 365 47 395 131
<< scpmoshvt >>
rect 112 391 142 475
rect 198 391 228 475
rect 284 391 314 475
rect 370 391 400 475
<< ndiff >>
rect 37 119 90 131
rect 37 85 45 119
rect 79 85 90 119
rect 37 47 90 85
rect 120 93 221 131
rect 120 59 131 93
rect 165 59 221 93
rect 120 47 221 59
rect 251 47 293 131
rect 323 47 365 131
rect 395 119 453 131
rect 395 85 411 119
rect 445 85 453 119
rect 395 47 453 85
<< pdiff >>
rect 59 463 112 475
rect 59 429 67 463
rect 101 429 112 463
rect 59 391 112 429
rect 142 463 198 475
rect 142 429 153 463
rect 187 429 198 463
rect 142 391 198 429
rect 228 437 284 475
rect 228 403 239 437
rect 273 403 284 437
rect 228 391 284 403
rect 314 463 370 475
rect 314 429 325 463
rect 359 429 370 463
rect 314 391 370 429
rect 400 437 453 475
rect 400 403 411 437
rect 445 403 453 437
rect 400 391 453 403
<< ndiffc >>
rect 45 85 79 119
rect 131 59 165 93
rect 411 85 445 119
<< pdiffc >>
rect 67 429 101 463
rect 153 429 187 463
rect 239 403 273 437
rect 325 429 359 463
rect 411 403 445 437
<< poly >>
rect 82 593 400 609
rect 82 559 98 593
rect 132 579 400 593
rect 132 559 148 579
rect 82 543 148 559
rect 112 475 142 501
rect 198 475 228 501
rect 284 475 314 501
rect 370 475 400 579
rect 112 302 142 391
rect 76 286 142 302
rect 198 287 228 391
rect 284 365 314 391
rect 370 369 400 391
rect 284 335 323 365
rect 370 339 437 369
rect 293 291 323 335
rect 76 252 92 286
rect 126 252 142 286
rect 76 218 142 252
rect 76 184 92 218
rect 126 184 142 218
rect 76 168 142 184
rect 185 271 251 287
rect 185 237 201 271
rect 235 237 251 271
rect 185 203 251 237
rect 185 169 201 203
rect 235 169 251 203
rect 90 131 120 168
rect 185 153 251 169
rect 221 131 251 153
rect 293 275 359 291
rect 293 241 309 275
rect 343 241 359 275
rect 293 225 359 241
rect 293 131 323 225
rect 407 183 437 339
rect 365 153 437 183
rect 365 131 395 153
rect 90 21 120 47
rect 221 21 251 47
rect 293 21 323 47
rect 365 21 395 47
<< polycont >>
rect 98 559 132 593
rect 92 252 126 286
rect 92 184 126 218
rect 201 237 235 271
rect 201 169 235 203
rect 309 241 343 275
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 51 593 140 609
rect 51 559 98 593
rect 132 559 140 593
rect 51 543 140 559
rect 51 467 117 543
rect 174 509 208 649
rect 325 509 359 649
rect 22 463 117 467
rect 22 429 67 463
rect 101 429 117 463
rect 22 425 117 429
rect 153 475 359 509
rect 153 463 187 475
rect 325 463 359 475
rect 22 123 56 425
rect 153 413 187 429
rect 223 437 289 441
rect 223 403 239 437
rect 273 403 289 437
rect 325 413 359 429
rect 395 437 461 441
rect 223 377 289 403
rect 395 403 411 437
rect 445 403 461 437
rect 395 377 461 403
rect 92 286 161 350
rect 223 343 461 377
rect 319 316 461 343
rect 126 252 161 286
rect 92 218 161 252
rect 126 184 161 218
rect 92 168 161 184
rect 201 271 257 287
rect 235 237 257 271
rect 201 203 257 237
rect 235 169 257 203
rect 22 119 95 123
rect 22 85 45 119
rect 79 85 95 119
rect 22 81 95 85
rect 131 93 165 109
rect 201 94 257 169
rect 293 275 359 276
rect 293 241 309 275
rect 343 241 359 275
rect 293 94 359 241
rect 395 119 461 316
rect 395 85 411 119
rect 445 85 461 119
rect 395 81 461 85
rect 131 17 165 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand3b_m
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3642402
string GDS_START 3636708
<< end >>
