magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 1 157 189 196
rect 572 157 959 245
rect 1 49 959 157
rect 0 0 960 49
<< scnmos >>
rect 80 86 110 170
rect 277 47 307 131
rect 363 47 393 131
rect 449 47 479 131
rect 657 135 687 219
rect 729 135 759 219
rect 850 135 880 219
<< scpmoshvt >>
rect 99 491 129 619
rect 204 491 234 575
rect 363 491 393 575
rect 441 491 471 575
rect 631 491 661 575
rect 717 491 747 575
rect 826 491 856 619
<< ndiff >>
rect 27 145 80 170
rect 27 111 35 145
rect 69 111 80 145
rect 27 86 80 111
rect 110 145 163 170
rect 110 111 121 145
rect 155 111 163 145
rect 110 86 163 111
rect 220 106 277 131
rect 220 72 228 106
rect 262 72 277 106
rect 220 47 277 72
rect 307 106 363 131
rect 307 72 318 106
rect 352 72 363 106
rect 307 47 363 72
rect 393 106 449 131
rect 393 72 404 106
rect 438 72 449 106
rect 393 47 449 72
rect 479 106 532 131
rect 479 72 490 106
rect 524 72 532 106
rect 479 47 532 72
rect 598 194 657 219
rect 598 160 606 194
rect 640 160 657 194
rect 598 135 657 160
rect 687 135 729 219
rect 759 194 850 219
rect 759 160 787 194
rect 821 160 850 194
rect 759 135 850 160
rect 880 181 933 219
rect 880 147 891 181
rect 925 147 933 181
rect 880 135 933 147
<< pdiff >>
rect 42 607 99 619
rect 42 573 50 607
rect 84 573 99 607
rect 42 537 99 573
rect 42 503 50 537
rect 84 503 99 537
rect 42 491 99 503
rect 129 607 182 619
rect 129 573 140 607
rect 174 575 182 607
rect 769 607 826 619
rect 769 575 777 607
rect 174 573 204 575
rect 129 537 204 573
rect 129 503 159 537
rect 193 503 204 537
rect 129 491 204 503
rect 234 550 363 575
rect 234 516 245 550
rect 279 516 318 550
rect 352 516 363 550
rect 234 491 363 516
rect 393 491 441 575
rect 471 550 631 575
rect 471 516 482 550
rect 516 516 586 550
rect 620 516 631 550
rect 471 491 631 516
rect 661 550 717 575
rect 661 516 672 550
rect 706 516 717 550
rect 661 491 717 516
rect 747 573 777 575
rect 811 573 826 607
rect 747 537 826 573
rect 747 503 758 537
rect 792 503 826 537
rect 747 491 826 503
rect 856 605 909 619
rect 856 571 867 605
rect 901 571 909 605
rect 856 537 909 571
rect 856 503 867 537
rect 901 503 909 537
rect 856 491 909 503
<< ndiffc >>
rect 35 111 69 145
rect 121 111 155 145
rect 228 72 262 106
rect 318 72 352 106
rect 404 72 438 106
rect 490 72 524 106
rect 606 160 640 194
rect 787 160 821 194
rect 891 147 925 181
<< pdiffc >>
rect 50 573 84 607
rect 50 503 84 537
rect 140 573 174 607
rect 159 503 193 537
rect 245 516 279 550
rect 318 516 352 550
rect 482 516 516 550
rect 586 516 620 550
rect 672 516 706 550
rect 777 573 811 607
rect 758 503 792 537
rect 867 571 901 605
rect 867 503 901 537
<< poly >>
rect 99 619 129 645
rect 826 619 856 645
rect 204 575 234 601
rect 363 575 393 601
rect 441 575 471 601
rect 631 575 661 601
rect 717 575 747 601
rect 99 453 129 491
rect 80 437 151 453
rect 80 403 101 437
rect 135 403 151 437
rect 80 369 151 403
rect 80 335 101 369
rect 135 335 151 369
rect 80 319 151 335
rect 204 345 234 491
rect 363 459 393 491
rect 290 443 393 459
rect 290 409 335 443
rect 369 409 393 443
rect 290 393 393 409
rect 204 329 315 345
rect 80 170 110 319
rect 204 315 265 329
rect 249 295 265 315
rect 299 295 315 329
rect 249 261 315 295
rect 249 227 265 261
rect 299 227 315 261
rect 249 211 315 227
rect 277 131 307 211
rect 363 131 393 393
rect 441 277 471 491
rect 631 433 661 491
rect 575 417 661 433
rect 575 383 591 417
rect 625 383 661 417
rect 575 367 661 383
rect 441 261 577 277
rect 441 227 479 261
rect 513 227 577 261
rect 631 271 661 367
rect 717 343 747 491
rect 826 453 856 491
rect 801 437 880 453
rect 801 403 817 437
rect 851 403 880 437
rect 801 369 880 403
rect 717 313 759 343
rect 801 335 817 369
rect 851 335 880 369
rect 801 319 880 335
rect 631 241 687 271
rect 441 211 577 227
rect 657 219 687 241
rect 729 219 759 313
rect 850 219 880 319
rect 449 131 479 211
rect 80 60 110 86
rect 547 67 577 211
rect 657 109 687 135
rect 729 67 759 135
rect 850 109 880 135
rect 277 21 307 47
rect 363 21 393 47
rect 449 21 479 47
rect 547 37 759 67
<< polycont >>
rect 101 403 135 437
rect 101 335 135 369
rect 335 409 369 443
rect 265 295 299 329
rect 265 227 299 261
rect 591 383 625 417
rect 479 227 513 261
rect 817 403 851 437
rect 817 335 851 369
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 19 607 100 615
rect 19 573 50 607
rect 84 573 100 607
rect 19 537 100 573
rect 19 503 50 537
rect 84 503 100 537
rect 19 499 100 503
rect 134 607 200 649
rect 134 573 140 607
rect 174 573 200 607
rect 134 537 200 573
rect 134 503 159 537
rect 193 503 200 537
rect 19 285 65 499
rect 134 487 200 503
rect 234 550 368 566
rect 234 516 245 550
rect 279 516 318 550
rect 352 516 368 550
rect 234 500 368 516
rect 466 550 636 649
rect 756 607 817 649
rect 756 573 777 607
rect 811 573 817 607
rect 466 516 482 550
rect 516 516 586 550
rect 620 516 636 550
rect 466 500 636 516
rect 670 550 722 566
rect 670 516 672 550
rect 706 516 722 550
rect 670 500 722 516
rect 234 453 283 500
rect 101 437 283 453
rect 135 419 283 437
rect 317 443 654 459
rect 135 403 229 419
rect 101 369 229 403
rect 317 409 335 443
rect 369 417 654 443
rect 369 409 591 417
rect 317 383 591 409
rect 625 383 654 417
rect 688 453 722 500
rect 756 537 817 573
rect 756 503 758 537
rect 792 503 817 537
rect 756 487 817 503
rect 851 605 943 615
rect 851 571 867 605
rect 901 571 943 605
rect 851 537 943 571
rect 851 503 867 537
rect 901 503 943 537
rect 851 487 943 503
rect 688 437 853 453
rect 688 403 817 437
rect 851 403 853 437
rect 135 335 229 369
rect 688 369 853 403
rect 688 347 817 369
rect 101 319 229 335
rect 19 145 85 285
rect 19 111 35 145
rect 69 111 85 145
rect 19 77 85 111
rect 119 145 161 161
rect 119 111 121 145
rect 155 111 161 145
rect 119 17 161 111
rect 195 122 229 319
rect 263 335 817 347
rect 851 335 853 369
rect 263 329 853 335
rect 263 295 265 329
rect 299 319 853 329
rect 299 313 722 319
rect 299 295 315 313
rect 263 261 315 295
rect 263 227 265 261
rect 299 227 315 261
rect 263 211 315 227
rect 398 261 560 277
rect 398 227 479 261
rect 513 227 560 261
rect 398 211 560 227
rect 602 194 722 313
rect 887 285 943 487
rect 312 143 540 177
rect 602 160 606 194
rect 640 160 722 194
rect 602 144 722 160
rect 771 194 837 210
rect 771 160 787 194
rect 821 160 837 194
rect 195 106 278 122
rect 195 72 228 106
rect 262 72 278 106
rect 195 56 278 72
rect 312 106 354 143
rect 312 72 318 106
rect 352 72 354 106
rect 312 56 354 72
rect 388 106 454 109
rect 388 72 404 106
rect 438 72 454 106
rect 388 17 454 72
rect 488 106 540 143
rect 488 72 490 106
rect 524 72 540 106
rect 488 56 540 72
rect 771 17 837 160
rect 871 181 943 285
rect 871 147 891 181
rect 925 147 943 181
rect 871 75 943 147
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ha_0
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 94 929 128 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6713644
string GDS_START 6704430
<< end >>
