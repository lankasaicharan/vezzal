magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
rect 465 319 693 331
<< pwell >>
rect 32 229 683 235
rect 32 49 1504 229
rect 0 0 1536 49
<< scnmos >>
rect 111 125 141 209
rect 197 125 227 209
rect 269 125 299 209
rect 355 125 385 209
rect 457 125 487 209
rect 574 125 604 209
rect 813 119 843 203
rect 899 119 929 203
rect 985 119 1015 203
rect 1071 119 1101 203
rect 1165 119 1195 203
rect 1237 119 1267 203
rect 1309 119 1339 203
rect 1395 119 1425 203
<< scpmoshvt >>
rect 80 367 110 451
rect 197 367 227 451
rect 269 367 299 451
rect 355 367 385 451
rect 441 367 471 451
rect 574 355 604 439
rect 813 391 843 475
rect 899 391 929 475
rect 985 391 1015 475
rect 1071 391 1101 475
rect 1165 391 1195 475
rect 1237 391 1267 475
rect 1309 391 1339 475
rect 1426 391 1456 475
<< ndiff >>
rect 58 189 111 209
rect 58 155 66 189
rect 100 155 111 189
rect 58 125 111 155
rect 141 171 197 209
rect 141 137 152 171
rect 186 137 197 171
rect 141 125 197 137
rect 227 125 269 209
rect 299 201 355 209
rect 299 167 310 201
rect 344 167 355 201
rect 299 125 355 167
rect 385 201 457 209
rect 385 167 412 201
rect 446 167 457 201
rect 385 125 457 167
rect 487 167 574 209
rect 487 133 519 167
rect 553 133 574 167
rect 487 125 574 133
rect 604 197 657 209
rect 604 163 615 197
rect 649 163 657 197
rect 604 125 657 163
rect 760 165 813 203
rect 760 131 768 165
rect 802 131 813 165
rect 760 119 813 131
rect 843 191 899 203
rect 843 157 854 191
rect 888 157 899 191
rect 843 119 899 157
rect 929 161 985 203
rect 929 127 940 161
rect 974 127 985 161
rect 929 119 985 127
rect 1015 191 1071 203
rect 1015 157 1026 191
rect 1060 157 1071 191
rect 1015 119 1071 157
rect 1101 191 1165 203
rect 1101 157 1120 191
rect 1154 157 1165 191
rect 1101 119 1165 157
rect 1195 119 1237 203
rect 1267 119 1309 203
rect 1339 165 1395 203
rect 1339 131 1350 165
rect 1384 131 1395 165
rect 1339 119 1395 131
rect 1425 185 1478 203
rect 1425 151 1436 185
rect 1470 151 1478 185
rect 1425 119 1478 151
<< pdiff >>
rect 501 451 559 455
rect 27 413 80 451
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 439 197 451
rect 110 405 121 439
rect 155 405 197 439
rect 110 367 197 405
rect 227 367 269 451
rect 299 413 355 451
rect 299 379 310 413
rect 344 379 355 413
rect 299 367 355 379
rect 385 413 441 451
rect 385 379 396 413
rect 430 379 441 413
rect 385 367 441 379
rect 471 447 559 451
rect 471 413 513 447
rect 547 439 559 447
rect 547 413 574 439
rect 471 367 574 413
rect 501 355 574 367
rect 604 401 657 439
rect 604 367 615 401
rect 649 367 657 401
rect 604 355 657 367
rect 760 463 813 475
rect 760 429 768 463
rect 802 429 813 463
rect 760 391 813 429
rect 843 433 899 475
rect 843 399 854 433
rect 888 399 899 433
rect 843 391 899 399
rect 929 463 985 475
rect 929 429 940 463
rect 974 429 985 463
rect 929 391 985 429
rect 1015 433 1071 475
rect 1015 399 1026 433
rect 1060 399 1071 433
rect 1015 391 1071 399
rect 1101 433 1165 475
rect 1101 399 1120 433
rect 1154 399 1165 433
rect 1101 391 1165 399
rect 1195 391 1237 475
rect 1267 391 1309 475
rect 1339 463 1426 475
rect 1339 429 1350 463
rect 1384 429 1426 463
rect 1339 391 1426 429
rect 1456 437 1509 475
rect 1456 403 1467 437
rect 1501 403 1509 437
rect 1456 391 1509 403
<< ndiffc >>
rect 66 155 100 189
rect 152 137 186 171
rect 310 167 344 201
rect 412 167 446 201
rect 519 133 553 167
rect 615 163 649 197
rect 768 131 802 165
rect 854 157 888 191
rect 940 127 974 161
rect 1026 157 1060 191
rect 1120 157 1154 191
rect 1350 131 1384 165
rect 1436 151 1470 185
<< pdiffc >>
rect 35 379 69 413
rect 121 405 155 439
rect 310 379 344 413
rect 396 379 430 413
rect 513 413 547 447
rect 615 367 649 401
rect 768 429 802 463
rect 854 399 888 433
rect 940 429 974 463
rect 1026 399 1060 433
rect 1120 399 1154 433
rect 1350 429 1384 463
rect 1467 403 1501 437
<< poly >>
rect 341 615 1195 645
rect 341 597 407 615
rect 217 575 299 591
rect 217 541 233 575
rect 267 541 299 575
rect 341 563 357 597
rect 391 563 407 597
rect 341 547 407 563
rect 672 557 738 573
rect 217 525 299 541
rect 80 451 110 477
rect 197 451 227 477
rect 269 451 299 525
rect 355 451 385 547
rect 672 523 688 557
rect 722 523 738 557
rect 672 507 738 523
rect 441 451 471 477
rect 574 439 604 465
rect 80 307 110 367
rect 80 291 155 307
rect 80 257 105 291
rect 139 257 155 291
rect 80 241 155 257
rect 111 209 141 241
rect 197 209 227 367
rect 269 209 299 367
rect 355 209 385 367
rect 441 261 471 367
rect 574 333 604 355
rect 672 333 702 507
rect 813 475 843 501
rect 899 475 929 615
rect 985 475 1015 501
rect 1071 475 1101 501
rect 1165 475 1195 615
rect 1237 599 1303 615
rect 1237 565 1253 599
rect 1287 565 1303 599
rect 1237 549 1303 565
rect 1237 475 1267 549
rect 1309 475 1339 501
rect 1426 475 1456 501
rect 813 333 843 391
rect 574 303 843 333
rect 441 231 487 261
rect 457 209 487 231
rect 574 209 604 303
rect 813 203 843 303
rect 899 203 929 391
rect 985 203 1015 391
rect 1071 323 1101 391
rect 1057 307 1123 323
rect 1057 273 1073 307
rect 1107 273 1123 307
rect 1057 257 1123 273
rect 1071 203 1101 257
rect 1165 203 1195 391
rect 1237 203 1267 391
rect 1309 203 1339 391
rect 1426 359 1456 391
rect 1381 343 1456 359
rect 1381 309 1397 343
rect 1431 309 1456 343
rect 1381 275 1456 309
rect 1381 241 1397 275
rect 1431 241 1456 275
rect 1381 225 1456 241
rect 1395 203 1425 225
rect 111 99 141 125
rect 197 51 227 125
rect 269 99 299 125
rect 355 99 385 125
rect 457 103 487 125
rect 433 87 499 103
rect 574 99 604 125
rect 813 93 843 119
rect 899 93 929 119
rect 433 53 449 87
rect 483 53 499 87
rect 433 51 499 53
rect 985 51 1015 119
rect 1071 93 1101 119
rect 1165 93 1195 119
rect 1237 93 1267 119
rect 1309 51 1339 119
rect 1395 93 1425 119
rect 197 21 1339 51
<< polycont >>
rect 233 541 267 575
rect 357 563 391 597
rect 688 523 722 557
rect 105 257 139 291
rect 1253 565 1287 599
rect 1073 273 1107 307
rect 1397 309 1431 343
rect 1397 241 1431 275
rect 449 53 483 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 31 413 69 572
rect 31 379 35 413
rect 105 439 171 649
rect 319 597 391 613
rect 217 541 233 575
rect 267 541 283 575
rect 217 502 283 541
rect 319 563 357 597
rect 319 538 391 563
rect 427 565 1253 599
rect 1287 565 1303 599
rect 427 557 738 565
rect 427 523 688 557
rect 722 523 738 557
rect 427 502 461 523
rect 1366 519 1400 649
rect 217 468 461 502
rect 774 487 1400 519
rect 497 485 1400 487
rect 105 405 121 439
rect 155 405 171 439
rect 497 463 808 485
rect 497 453 768 463
rect 497 447 563 453
rect 105 401 171 405
rect 306 413 348 429
rect 31 205 69 379
rect 306 379 310 413
rect 344 379 348 413
rect 306 307 348 379
rect 392 413 434 429
rect 497 413 513 447
rect 547 413 563 447
rect 764 429 768 453
rect 802 429 808 463
rect 936 463 978 485
rect 392 379 396 413
rect 430 379 434 413
rect 392 377 434 379
rect 611 401 653 417
rect 764 413 808 429
rect 850 433 892 449
rect 611 377 615 401
rect 392 367 615 377
rect 649 367 653 401
rect 392 343 653 367
rect 850 399 854 433
rect 888 399 892 433
rect 936 429 940 463
rect 974 429 978 463
rect 1334 463 1400 485
rect 936 413 978 429
rect 1022 433 1064 449
rect 850 377 892 399
rect 1022 399 1026 433
rect 1060 399 1064 433
rect 1022 377 1064 399
rect 1116 433 1193 449
rect 1116 399 1120 433
rect 1154 399 1193 433
rect 1334 429 1350 463
rect 1384 429 1400 463
rect 1334 425 1400 429
rect 1467 437 1505 572
rect 1116 383 1193 399
rect 850 343 1064 377
rect 105 291 1073 307
rect 139 273 1073 291
rect 1107 273 1123 307
rect 105 241 139 257
rect 31 189 104 205
rect 31 155 66 189
rect 100 155 104 189
rect 294 201 360 273
rect 1159 259 1193 383
rect 1501 403 1505 437
rect 1397 343 1431 359
rect 1397 275 1431 309
rect 1159 241 1397 259
rect 31 139 104 155
rect 148 171 186 187
rect 148 137 152 171
rect 294 167 310 201
rect 344 167 360 201
rect 396 203 653 237
rect 396 201 462 203
rect 396 167 412 201
rect 446 167 462 201
rect 611 197 653 203
rect 148 17 186 137
rect 503 133 519 167
rect 553 133 569 167
rect 611 163 615 197
rect 649 163 653 197
rect 850 201 1064 235
rect 1159 225 1431 241
rect 1159 207 1193 225
rect 850 191 888 201
rect 611 147 653 163
rect 764 165 806 181
rect 503 129 569 133
rect 223 93 449 128
rect 223 87 499 93
rect 223 53 449 87
rect 483 53 499 87
rect 535 17 569 129
rect 764 131 768 165
rect 802 131 806 165
rect 850 157 854 191
rect 1026 191 1064 201
rect 850 141 888 157
rect 924 161 990 165
rect 764 17 806 131
rect 924 127 940 161
rect 974 127 990 161
rect 1060 157 1064 191
rect 1026 141 1064 157
rect 1116 191 1193 207
rect 1116 157 1120 191
rect 1154 157 1193 191
rect 1467 189 1505 403
rect 1420 185 1505 189
rect 1116 141 1193 157
rect 1346 165 1384 181
rect 924 17 990 127
rect 1346 131 1350 165
rect 1420 151 1436 185
rect 1470 151 1505 185
rect 1420 147 1505 151
rect 1346 17 1384 131
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fa_m
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1471 390 1505 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1471 464 1505 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1471 538 1505 572 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2420004
string GDS_START 2408662
<< end >>
