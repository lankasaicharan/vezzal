magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 7 157 390 241
rect 7 49 671 157
rect 0 0 672 49
<< scnmos >>
rect 86 131 116 215
rect 195 47 225 215
rect 281 47 311 215
rect 386 47 416 131
rect 472 47 502 131
rect 562 47 592 131
<< scpmoshvt >>
rect 119 367 149 451
rect 224 367 254 619
rect 310 367 340 619
rect 418 385 448 469
rect 490 385 520 469
rect 562 385 592 469
<< ndiff >>
rect 33 190 86 215
rect 33 156 41 190
rect 75 156 86 190
rect 33 131 86 156
rect 116 179 195 215
rect 116 145 127 179
rect 161 145 195 179
rect 116 131 195 145
rect 138 93 195 131
rect 138 59 146 93
rect 180 59 195 93
rect 138 47 195 59
rect 225 186 281 215
rect 225 152 236 186
rect 270 152 281 186
rect 225 101 281 152
rect 225 67 236 101
rect 270 67 281 101
rect 225 47 281 67
rect 311 179 364 215
rect 311 145 322 179
rect 356 145 364 179
rect 311 131 364 145
rect 311 93 386 131
rect 311 59 341 93
rect 375 59 386 93
rect 311 47 386 59
rect 416 106 472 131
rect 416 72 427 106
rect 461 72 472 106
rect 416 47 472 72
rect 502 106 562 131
rect 502 72 513 106
rect 547 72 562 106
rect 502 47 562 72
rect 592 106 645 131
rect 592 72 603 106
rect 637 72 645 106
rect 592 47 645 72
<< pdiff >>
rect 171 570 224 619
rect 171 536 179 570
rect 213 536 224 570
rect 171 451 224 536
rect 66 428 119 451
rect 66 394 74 428
rect 108 394 119 428
rect 66 367 119 394
rect 149 367 224 451
rect 254 413 310 619
rect 254 379 265 413
rect 299 379 310 413
rect 254 367 310 379
rect 340 570 393 619
rect 340 536 351 570
rect 385 536 393 570
rect 340 469 393 536
rect 340 385 418 469
rect 448 385 490 469
rect 520 385 562 469
rect 592 444 645 469
rect 592 410 603 444
rect 637 410 645 444
rect 592 385 645 410
rect 340 367 393 385
<< ndiffc >>
rect 41 156 75 190
rect 127 145 161 179
rect 146 59 180 93
rect 236 152 270 186
rect 236 67 270 101
rect 322 145 356 179
rect 341 59 375 93
rect 427 72 461 106
rect 513 72 547 106
rect 603 72 637 106
<< pdiffc >>
rect 179 536 213 570
rect 74 394 108 428
rect 265 379 299 413
rect 351 536 385 570
rect 603 410 637 444
<< poly >>
rect 224 619 254 645
rect 310 619 340 645
rect 119 451 149 477
rect 497 593 592 609
rect 497 559 513 593
rect 547 559 592 593
rect 497 543 592 559
rect 418 469 448 495
rect 490 469 520 495
rect 562 469 592 543
rect 119 345 149 367
rect 48 319 149 345
rect 48 285 64 319
rect 98 315 149 319
rect 98 285 116 315
rect 48 269 116 285
rect 86 215 116 269
rect 224 304 254 367
rect 310 304 340 367
rect 418 335 448 385
rect 224 288 340 304
rect 224 267 290 288
rect 195 254 290 267
rect 324 254 340 288
rect 382 319 448 335
rect 382 285 398 319
rect 432 285 448 319
rect 382 269 448 285
rect 490 291 520 385
rect 562 363 592 385
rect 562 333 634 363
rect 490 275 556 291
rect 195 237 340 254
rect 195 215 225 237
rect 281 215 311 237
rect 86 105 116 131
rect 386 131 416 269
rect 490 241 506 275
rect 540 241 556 275
rect 490 225 556 241
rect 490 183 520 225
rect 604 183 634 333
rect 472 153 520 183
rect 562 153 634 183
rect 472 131 502 153
rect 562 131 592 153
rect 195 21 225 47
rect 281 21 311 47
rect 386 21 416 47
rect 472 21 502 47
rect 562 21 592 47
<< polycont >>
rect 513 559 547 593
rect 64 285 98 319
rect 290 254 324 288
rect 398 285 432 319
rect 506 241 540 275
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 163 570 229 649
rect 163 536 179 570
rect 213 536 229 570
rect 163 528 229 536
rect 335 570 401 649
rect 335 536 351 570
rect 385 536 401 570
rect 335 528 401 536
rect 497 559 513 593
rect 547 559 563 593
rect 497 492 563 559
rect 58 458 563 492
rect 58 428 186 458
rect 58 394 74 428
rect 108 394 186 428
rect 597 444 653 460
rect 58 384 186 394
rect 17 319 116 350
rect 17 285 64 319
rect 98 285 116 319
rect 17 281 116 285
rect 150 247 186 384
rect 25 213 186 247
rect 220 413 315 424
rect 220 379 265 413
rect 299 379 315 413
rect 220 363 315 379
rect 25 190 77 213
rect 25 156 41 190
rect 75 156 77 190
rect 220 202 254 363
rect 382 319 461 424
rect 288 288 344 304
rect 288 254 290 288
rect 324 254 344 288
rect 382 285 398 319
rect 432 285 461 319
rect 288 247 344 254
rect 495 275 563 424
rect 288 238 461 247
rect 310 213 461 238
rect 495 241 506 275
rect 540 241 563 275
rect 495 225 563 241
rect 597 410 603 444
rect 637 410 653 444
rect 220 186 272 202
rect 25 140 77 156
rect 111 145 127 179
rect 161 145 186 179
rect 111 93 186 145
rect 111 59 146 93
rect 180 59 186 93
rect 111 17 186 59
rect 220 152 236 186
rect 270 152 272 186
rect 420 191 461 213
rect 597 191 653 410
rect 220 101 272 152
rect 220 67 236 101
rect 270 67 272 101
rect 220 51 272 67
rect 306 145 322 179
rect 356 145 386 179
rect 306 93 386 145
rect 306 59 341 93
rect 375 59 386 93
rect 306 17 386 59
rect 420 157 653 191
rect 420 106 463 157
rect 420 72 427 106
rect 461 72 463 106
rect 420 56 463 72
rect 497 106 563 123
rect 497 72 513 106
rect 547 72 563 106
rect 497 17 563 72
rect 597 106 653 157
rect 597 72 603 106
rect 637 72 653 106
rect 597 56 653 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or3b_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 593916
string GDS_START 587566
<< end >>
