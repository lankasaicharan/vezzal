magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 283 241 651 245
rect 7 49 651 241
rect 0 0 672 49
<< scnmos >>
rect 86 47 116 215
rect 172 47 202 215
rect 362 51 392 219
rect 448 51 478 219
rect 542 51 572 219
<< scpmoshvt >>
rect 86 367 116 619
rect 172 367 202 619
rect 362 367 392 619
rect 448 367 478 619
rect 542 367 572 619
<< ndiff >>
rect 33 203 86 215
rect 33 169 41 203
rect 75 169 86 203
rect 33 93 86 169
rect 33 59 41 93
rect 75 59 86 93
rect 33 47 86 59
rect 116 203 172 215
rect 116 169 127 203
rect 161 169 172 203
rect 116 101 172 169
rect 116 67 127 101
rect 161 67 172 101
rect 116 47 172 67
rect 202 181 255 215
rect 202 147 213 181
rect 247 147 255 181
rect 202 93 255 147
rect 202 59 213 93
rect 247 59 255 93
rect 202 47 255 59
rect 309 207 362 219
rect 309 173 317 207
rect 351 173 362 207
rect 309 101 362 173
rect 309 67 317 101
rect 351 67 362 101
rect 309 51 362 67
rect 392 207 448 219
rect 392 173 403 207
rect 437 173 448 207
rect 392 101 448 173
rect 392 67 403 101
rect 437 67 448 101
rect 392 51 448 67
rect 478 173 542 219
rect 478 139 493 173
rect 527 139 542 173
rect 478 97 542 139
rect 478 63 493 97
rect 527 63 542 97
rect 478 51 542 63
rect 572 207 625 219
rect 572 173 583 207
rect 617 173 625 207
rect 572 101 625 173
rect 572 67 583 101
rect 617 67 625 101
rect 572 51 625 67
<< pdiff >>
rect 33 607 86 619
rect 33 573 41 607
rect 75 573 86 607
rect 33 502 86 573
rect 33 468 41 502
rect 75 468 86 502
rect 33 413 86 468
rect 33 379 41 413
rect 75 379 86 413
rect 33 367 86 379
rect 116 599 172 619
rect 116 565 127 599
rect 161 565 172 599
rect 116 501 172 565
rect 116 467 127 501
rect 161 467 172 501
rect 116 413 172 467
rect 116 379 127 413
rect 161 379 172 413
rect 116 367 172 379
rect 202 607 362 619
rect 202 573 213 607
rect 247 573 317 607
rect 351 573 362 607
rect 202 495 362 573
rect 202 461 213 495
rect 247 461 317 495
rect 351 461 362 495
rect 202 367 362 461
rect 392 599 448 619
rect 392 565 403 599
rect 437 565 448 599
rect 392 507 448 565
rect 392 473 403 507
rect 437 473 448 507
rect 392 418 448 473
rect 392 384 403 418
rect 437 384 448 418
rect 392 367 448 384
rect 478 367 542 619
rect 572 607 625 619
rect 572 573 583 607
rect 617 573 625 607
rect 572 507 625 573
rect 572 473 583 507
rect 617 473 625 507
rect 572 418 625 473
rect 572 384 583 418
rect 617 384 625 418
rect 572 367 625 384
<< ndiffc >>
rect 41 169 75 203
rect 41 59 75 93
rect 127 169 161 203
rect 127 67 161 101
rect 213 147 247 181
rect 213 59 247 93
rect 317 173 351 207
rect 317 67 351 101
rect 403 173 437 207
rect 403 67 437 101
rect 493 139 527 173
rect 493 63 527 97
rect 583 173 617 207
rect 583 67 617 101
<< pdiffc >>
rect 41 573 75 607
rect 41 468 75 502
rect 41 379 75 413
rect 127 565 161 599
rect 127 467 161 501
rect 127 379 161 413
rect 213 573 247 607
rect 317 573 351 607
rect 213 461 247 495
rect 317 461 351 495
rect 403 565 437 599
rect 403 473 437 507
rect 403 384 437 418
rect 583 573 617 607
rect 583 473 617 507
rect 583 384 617 418
<< poly >>
rect 86 619 116 645
rect 172 619 202 645
rect 362 619 392 645
rect 448 619 478 645
rect 542 619 572 645
rect 86 267 116 367
rect 172 303 202 367
rect 362 335 392 367
rect 448 335 478 367
rect 313 319 392 335
rect 172 287 263 303
rect 172 267 213 287
rect 86 253 213 267
rect 247 253 263 287
rect 313 285 329 319
rect 363 285 392 319
rect 313 269 392 285
rect 434 319 500 335
rect 434 285 450 319
rect 484 285 500 319
rect 434 269 500 285
rect 542 325 572 367
rect 542 309 647 325
rect 542 275 597 309
rect 631 275 647 309
rect 86 237 263 253
rect 86 215 116 237
rect 172 215 202 237
rect 362 219 392 269
rect 448 219 478 269
rect 542 259 647 275
rect 542 219 572 259
rect 86 21 116 47
rect 172 21 202 47
rect 362 25 392 51
rect 448 25 478 51
rect 542 25 572 51
<< polycont >>
rect 213 253 247 287
rect 329 285 363 319
rect 450 285 484 319
rect 597 275 631 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 25 607 79 649
rect 25 573 41 607
rect 75 573 79 607
rect 25 502 79 573
rect 25 468 41 502
rect 75 468 79 502
rect 25 413 79 468
rect 25 379 41 413
rect 75 379 79 413
rect 25 363 79 379
rect 113 599 163 615
rect 113 565 127 599
rect 161 565 163 599
rect 113 501 163 565
rect 113 467 127 501
rect 161 467 163 501
rect 113 413 163 467
rect 197 607 367 649
rect 197 573 213 607
rect 247 573 317 607
rect 351 573 367 607
rect 197 495 367 573
rect 197 461 213 495
rect 247 461 317 495
rect 351 461 367 495
rect 197 452 367 461
rect 401 599 453 615
rect 401 565 403 599
rect 437 565 453 599
rect 401 507 453 565
rect 401 473 403 507
rect 437 473 453 507
rect 401 418 453 473
rect 113 379 127 413
rect 161 379 163 413
rect 25 203 79 219
rect 25 169 41 203
rect 75 169 79 203
rect 25 93 79 169
rect 25 59 41 93
rect 75 59 79 93
rect 25 17 79 59
rect 113 203 163 379
rect 229 384 403 418
rect 437 384 453 418
rect 567 607 633 649
rect 567 573 583 607
rect 617 573 633 607
rect 567 507 633 573
rect 567 473 583 507
rect 617 473 633 507
rect 567 418 633 473
rect 567 384 583 418
rect 617 384 633 418
rect 229 304 263 384
rect 197 287 263 304
rect 197 253 213 287
rect 247 253 263 287
rect 297 319 379 350
rect 297 285 329 319
rect 363 285 379 319
rect 297 283 379 285
rect 413 319 547 350
rect 413 285 450 319
rect 484 285 547 319
rect 413 275 547 285
rect 581 309 655 350
rect 581 275 597 309
rect 631 275 655 309
rect 197 249 263 253
rect 197 215 360 249
rect 113 169 127 203
rect 161 169 163 203
rect 301 207 360 215
rect 113 101 163 169
rect 113 67 127 101
rect 161 67 163 101
rect 113 51 163 67
rect 197 147 213 181
rect 247 147 263 181
rect 197 93 263 147
rect 197 59 213 93
rect 247 59 263 93
rect 197 17 263 59
rect 301 173 317 207
rect 351 173 360 207
rect 301 101 360 173
rect 301 67 317 101
rect 351 67 360 101
rect 301 51 360 67
rect 394 207 633 241
rect 394 173 403 207
rect 437 173 443 207
rect 577 173 583 207
rect 617 173 633 207
rect 394 101 443 173
rect 394 67 403 101
rect 437 67 443 101
rect 394 51 443 67
rect 477 139 493 173
rect 527 139 543 173
rect 477 97 543 139
rect 477 63 493 97
rect 527 63 543 97
rect 477 17 543 63
rect 577 101 633 173
rect 577 67 583 101
rect 617 67 633 101
rect 577 51 633 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21a_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 825932
string GDS_START 818758
<< end >>
