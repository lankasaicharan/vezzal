magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 210 157 754 161
rect 1 49 754 157
rect 0 0 768 49
<< scnmos >>
rect 80 47 110 131
rect 289 51 319 135
rect 375 51 405 135
rect 465 51 495 135
rect 551 51 581 135
rect 645 51 675 135
<< scpmoshvt >>
rect 117 483 147 611
rect 203 483 233 611
rect 393 483 423 611
rect 483 483 513 611
rect 573 483 603 611
rect 645 483 675 611
<< ndiff >>
rect 27 105 80 131
rect 27 71 35 105
rect 69 71 80 105
rect 27 47 80 71
rect 110 106 163 131
rect 110 72 121 106
rect 155 72 163 106
rect 110 47 163 72
rect 236 110 289 135
rect 236 76 244 110
rect 278 76 289 110
rect 236 51 289 76
rect 319 110 375 135
rect 319 76 330 110
rect 364 76 375 110
rect 319 51 375 76
rect 405 110 465 135
rect 405 76 419 110
rect 453 76 465 110
rect 405 51 465 76
rect 495 110 551 135
rect 495 76 506 110
rect 540 76 551 110
rect 495 51 551 76
rect 581 100 645 135
rect 581 66 596 100
rect 630 66 645 100
rect 581 51 645 66
rect 675 110 728 135
rect 675 76 686 110
rect 720 76 728 110
rect 675 51 728 76
<< pdiff >>
rect 64 597 117 611
rect 64 563 72 597
rect 106 563 117 597
rect 64 529 117 563
rect 64 495 72 529
rect 106 495 117 529
rect 64 483 117 495
rect 147 599 203 611
rect 147 565 158 599
rect 192 565 203 599
rect 147 529 203 565
rect 147 495 158 529
rect 192 495 203 529
rect 147 483 203 495
rect 233 599 393 611
rect 233 565 244 599
rect 278 565 348 599
rect 382 565 393 599
rect 233 529 393 565
rect 233 495 244 529
rect 278 495 348 529
rect 382 495 393 529
rect 233 483 393 495
rect 423 483 483 611
rect 513 483 573 611
rect 603 483 645 611
rect 675 599 728 611
rect 675 565 686 599
rect 720 565 728 599
rect 675 529 728 565
rect 675 495 686 529
rect 720 495 728 529
rect 675 483 728 495
<< ndiffc >>
rect 35 71 69 105
rect 121 72 155 106
rect 244 76 278 110
rect 330 76 364 110
rect 419 76 453 110
rect 506 76 540 110
rect 596 66 630 100
rect 686 76 720 110
<< pdiffc >>
rect 72 563 106 597
rect 72 495 106 529
rect 158 565 192 599
rect 158 495 192 529
rect 244 565 278 599
rect 348 565 382 599
rect 244 495 278 529
rect 348 495 382 529
rect 686 565 720 599
rect 686 495 720 529
<< poly >>
rect 117 611 147 637
rect 203 611 233 637
rect 393 611 423 637
rect 483 611 513 637
rect 573 611 603 637
rect 645 611 675 637
rect 117 287 147 483
rect 203 350 233 483
rect 393 428 423 483
rect 483 441 513 483
rect 357 412 423 428
rect 357 378 373 412
rect 407 378 423 412
rect 203 334 269 350
rect 203 300 219 334
rect 253 300 269 334
rect 80 271 155 287
rect 80 237 105 271
rect 139 237 155 271
rect 80 203 155 237
rect 203 266 269 300
rect 357 344 423 378
rect 357 310 373 344
rect 407 310 423 344
rect 357 294 423 310
rect 203 232 219 266
rect 253 246 269 266
rect 367 259 423 294
rect 465 425 531 441
rect 465 391 481 425
rect 515 391 531 425
rect 465 357 531 391
rect 465 323 481 357
rect 515 323 531 357
rect 465 307 531 323
rect 573 383 603 483
rect 645 461 675 483
rect 645 431 711 461
rect 573 367 639 383
rect 573 333 589 367
rect 623 333 639 367
rect 253 232 319 246
rect 203 216 319 232
rect 367 229 405 259
rect 80 169 105 203
rect 139 169 155 203
rect 80 153 155 169
rect 80 131 110 153
rect 289 135 319 216
rect 375 135 405 229
rect 465 135 495 307
rect 573 299 639 333
rect 573 265 589 299
rect 623 265 639 299
rect 573 249 639 265
rect 681 325 711 431
rect 681 309 747 325
rect 681 275 697 309
rect 731 275 747 309
rect 573 187 603 249
rect 681 241 747 275
rect 681 207 697 241
rect 731 207 747 241
rect 681 201 747 207
rect 551 157 603 187
rect 645 171 747 201
rect 551 135 581 157
rect 645 135 675 171
rect 80 21 110 47
rect 289 25 319 51
rect 375 25 405 51
rect 465 25 495 51
rect 551 25 581 51
rect 645 25 675 51
<< polycont >>
rect 373 378 407 412
rect 219 300 253 334
rect 105 237 139 271
rect 373 310 407 344
rect 219 232 253 266
rect 481 391 515 425
rect 481 323 515 357
rect 589 333 623 367
rect 105 169 139 203
rect 589 265 623 299
rect 697 275 731 309
rect 697 207 731 241
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 597 108 613
rect 17 563 72 597
rect 106 563 108 597
rect 17 529 108 563
rect 17 495 72 529
rect 106 495 108 529
rect 17 479 108 495
rect 142 599 208 649
rect 142 565 158 599
rect 192 565 208 599
rect 142 529 208 565
rect 142 495 158 529
rect 192 495 208 529
rect 142 479 208 495
rect 242 599 398 615
rect 242 565 244 599
rect 278 565 348 599
rect 382 565 398 599
rect 675 599 738 649
rect 242 529 398 565
rect 242 495 244 529
rect 278 495 348 529
rect 382 495 398 529
rect 242 479 398 495
rect 17 105 71 479
rect 242 443 285 479
rect 105 409 285 443
rect 319 412 447 442
rect 493 441 555 572
rect 105 271 155 409
rect 319 378 373 412
rect 407 378 447 412
rect 139 237 155 271
rect 105 203 155 237
rect 203 334 269 370
rect 203 300 219 334
rect 253 300 269 334
rect 203 266 269 300
rect 203 232 219 266
rect 253 232 269 266
rect 203 216 269 232
rect 319 344 447 378
rect 319 310 373 344
rect 407 310 447 344
rect 319 228 447 310
rect 481 425 555 441
rect 515 391 555 425
rect 481 357 555 391
rect 515 323 555 357
rect 481 228 555 323
rect 589 367 641 572
rect 675 565 686 599
rect 720 565 738 599
rect 675 529 738 565
rect 675 495 686 529
rect 720 495 738 529
rect 675 479 738 495
rect 623 333 641 367
rect 589 299 641 333
rect 623 265 641 299
rect 589 228 641 265
rect 681 309 747 436
rect 681 275 697 309
rect 731 275 747 309
rect 681 241 747 275
rect 681 207 697 241
rect 731 207 747 241
rect 139 182 155 203
rect 139 169 288 182
rect 105 148 288 169
rect 17 71 35 105
rect 69 71 71 105
rect 17 53 71 71
rect 105 106 171 114
rect 105 72 121 106
rect 155 72 171 106
rect 105 17 171 72
rect 228 110 288 148
rect 228 76 244 110
rect 278 76 288 110
rect 228 60 288 76
rect 322 173 540 194
rect 322 160 741 173
rect 322 110 373 160
rect 497 139 741 160
rect 322 76 330 110
rect 364 76 373 110
rect 322 60 373 76
rect 407 110 463 126
rect 407 76 419 110
rect 453 76 463 110
rect 407 17 463 76
rect 497 110 546 139
rect 497 76 506 110
rect 540 76 546 110
rect 680 110 741 139
rect 497 60 546 76
rect 580 100 646 105
rect 580 66 596 100
rect 630 66 646 100
rect 580 17 646 66
rect 680 76 686 110
rect 720 76 741 110
rect 680 60 741 76
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o41a_0
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 362706
string GDS_START 353208
<< end >>
