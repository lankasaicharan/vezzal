magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 597 157 1029 167
rect 1 49 1029 157
rect 0 0 1056 49
<< scnmos >>
rect 84 47 114 131
rect 162 47 192 131
rect 248 47 278 131
rect 320 47 350 131
rect 406 47 436 131
rect 478 47 508 131
rect 680 57 710 141
rect 752 57 782 141
rect 838 57 868 141
rect 916 57 946 141
<< scpmoshvt >>
rect 84 409 134 609
rect 182 409 232 609
rect 428 390 478 590
rect 689 409 739 609
rect 795 409 845 609
rect 916 409 966 609
<< ndiff >>
rect 27 106 84 131
rect 27 72 39 106
rect 73 72 84 106
rect 27 47 84 72
rect 114 47 162 131
rect 192 111 248 131
rect 192 77 203 111
rect 237 77 248 111
rect 192 47 248 77
rect 278 47 320 131
rect 350 103 406 131
rect 350 69 361 103
rect 395 69 406 103
rect 350 47 406 69
rect 436 47 478 131
rect 508 108 565 131
rect 508 74 519 108
rect 553 74 565 108
rect 508 47 565 74
rect 623 116 680 141
rect 623 82 635 116
rect 669 82 680 116
rect 623 57 680 82
rect 710 57 752 141
rect 782 108 838 141
rect 782 74 793 108
rect 827 74 838 108
rect 782 57 838 74
rect 868 57 916 141
rect 946 116 1003 141
rect 946 82 957 116
rect 991 82 1003 116
rect 946 57 1003 82
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 409 182 609
rect 232 597 289 609
rect 232 563 243 597
rect 277 563 289 597
rect 632 597 689 609
rect 232 526 289 563
rect 232 492 243 526
rect 277 492 289 526
rect 232 455 289 492
rect 232 421 243 455
rect 277 421 289 455
rect 232 409 289 421
rect 371 577 428 590
rect 371 543 383 577
rect 417 543 428 577
rect 371 390 428 543
rect 478 436 535 590
rect 478 402 489 436
rect 523 402 535 436
rect 632 563 644 597
rect 678 563 689 597
rect 632 526 689 563
rect 632 492 644 526
rect 678 492 689 526
rect 632 455 689 492
rect 632 421 644 455
rect 678 421 689 455
rect 632 409 689 421
rect 739 597 795 609
rect 739 563 750 597
rect 784 563 795 597
rect 739 526 795 563
rect 739 492 750 526
rect 784 492 795 526
rect 739 455 795 492
rect 739 421 750 455
rect 784 421 795 455
rect 739 409 795 421
rect 845 597 916 609
rect 845 563 856 597
rect 890 563 916 597
rect 845 525 916 563
rect 845 491 856 525
rect 890 491 916 525
rect 845 409 916 491
rect 966 597 1023 609
rect 966 563 977 597
rect 1011 563 1023 597
rect 966 526 1023 563
rect 966 492 977 526
rect 1011 492 1023 526
rect 966 455 1023 492
rect 966 421 977 455
rect 1011 421 1023 455
rect 966 409 1023 421
rect 478 390 535 402
<< ndiffc >>
rect 39 72 73 106
rect 203 77 237 111
rect 361 69 395 103
rect 519 74 553 108
rect 635 82 669 116
rect 793 74 827 108
rect 957 82 991 116
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 243 563 277 597
rect 243 492 277 526
rect 243 421 277 455
rect 383 543 417 577
rect 489 402 523 436
rect 644 563 678 597
rect 644 492 678 526
rect 644 421 678 455
rect 750 563 784 597
rect 750 492 784 526
rect 750 421 784 455
rect 856 563 890 597
rect 856 491 890 525
rect 977 563 1011 597
rect 977 492 1011 526
rect 977 421 1011 455
<< poly >>
rect 84 609 134 635
rect 182 609 232 635
rect 428 590 478 616
rect 689 609 739 635
rect 795 609 845 635
rect 916 609 966 635
rect 84 305 134 409
rect 40 289 134 305
rect 40 255 56 289
rect 90 275 134 289
rect 182 369 232 409
rect 182 353 278 369
rect 428 358 478 390
rect 689 369 739 409
rect 795 369 845 409
rect 916 369 966 409
rect 182 319 228 353
rect 262 319 278 353
rect 182 285 278 319
rect 90 255 114 275
rect 40 221 114 255
rect 182 251 228 285
rect 262 251 278 285
rect 182 235 278 251
rect 40 187 56 221
rect 90 187 114 221
rect 40 157 192 187
rect 84 131 114 157
rect 162 131 192 157
rect 248 176 278 235
rect 345 342 478 358
rect 345 308 361 342
rect 395 308 478 342
rect 345 299 478 308
rect 673 353 739 369
rect 673 319 689 353
rect 723 319 739 353
rect 345 283 583 299
rect 345 274 533 283
rect 345 240 361 274
rect 395 249 533 274
rect 567 249 583 283
rect 395 240 583 249
rect 345 224 583 240
rect 673 285 739 319
rect 673 251 689 285
rect 723 251 739 285
rect 673 235 739 251
rect 787 353 868 369
rect 787 319 803 353
rect 837 319 868 353
rect 787 285 868 319
rect 787 251 803 285
rect 837 251 868 285
rect 787 235 868 251
rect 248 146 350 176
rect 248 131 278 146
rect 320 131 350 146
rect 406 131 436 224
rect 478 215 583 224
rect 478 181 533 215
rect 567 181 583 215
rect 478 165 583 181
rect 680 186 710 235
rect 478 131 508 165
rect 680 156 782 186
rect 680 141 710 156
rect 752 141 782 156
rect 838 141 868 235
rect 916 353 982 369
rect 916 319 932 353
rect 966 319 982 353
rect 916 285 982 319
rect 916 251 932 285
rect 966 251 982 285
rect 916 235 982 251
rect 916 141 946 235
rect 84 21 114 47
rect 162 21 192 47
rect 248 21 278 47
rect 320 21 350 47
rect 406 21 436 47
rect 478 21 508 47
rect 680 31 710 57
rect 752 31 782 57
rect 838 31 868 57
rect 916 31 946 57
<< polycont >>
rect 56 255 90 289
rect 228 319 262 353
rect 228 251 262 285
rect 56 187 90 221
rect 361 308 395 342
rect 689 319 723 353
rect 361 240 395 274
rect 533 249 567 283
rect 689 251 723 285
rect 803 319 837 353
rect 803 251 837 285
rect 533 181 567 215
rect 932 319 966 353
rect 932 251 966 285
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 526 89 563
rect 23 492 39 526
rect 73 492 89 526
rect 23 455 89 492
rect 23 421 39 455
rect 73 439 89 455
rect 227 597 293 613
rect 227 563 243 597
rect 277 563 293 597
rect 227 526 293 563
rect 367 577 433 649
rect 367 543 383 577
rect 417 543 433 577
rect 367 542 433 543
rect 628 597 694 613
rect 628 563 644 597
rect 678 563 694 597
rect 227 492 243 526
rect 277 506 293 526
rect 628 526 694 563
rect 628 506 644 526
rect 277 492 644 506
rect 678 492 694 526
rect 227 472 694 492
rect 227 455 293 472
rect 73 421 176 439
rect 23 405 176 421
rect 227 421 243 455
rect 277 421 293 455
rect 628 455 694 472
rect 227 405 293 421
rect 25 289 106 356
rect 25 255 56 289
rect 90 255 106 289
rect 25 221 106 255
rect 25 187 56 221
rect 90 187 106 221
rect 25 171 106 187
rect 142 199 176 405
rect 447 402 489 436
rect 523 402 551 436
rect 628 421 644 455
rect 678 421 694 455
rect 628 405 694 421
rect 734 597 800 613
rect 734 563 750 597
rect 784 563 800 597
rect 734 526 800 563
rect 734 492 750 526
rect 784 492 800 526
rect 734 455 800 492
rect 840 597 906 649
rect 840 563 856 597
rect 890 563 906 597
rect 840 525 906 563
rect 840 491 856 525
rect 890 491 906 525
rect 840 475 906 491
rect 961 597 1027 613
rect 961 563 977 597
rect 1011 563 1027 597
rect 961 526 1027 563
rect 961 492 977 526
rect 1011 492 1027 526
rect 734 421 750 455
rect 784 439 800 455
rect 961 455 1027 492
rect 961 439 977 455
rect 784 421 977 439
rect 1011 421 1027 455
rect 734 405 1027 421
rect 447 384 551 402
rect 212 353 278 369
rect 212 319 228 353
rect 262 319 278 353
rect 212 285 278 319
rect 212 251 228 285
rect 262 251 278 285
rect 212 235 278 251
rect 345 342 411 358
rect 345 308 361 342
rect 395 308 411 342
rect 345 274 411 308
rect 345 240 361 274
rect 395 240 411 274
rect 345 199 411 240
rect 142 165 411 199
rect 23 106 89 135
rect 23 72 39 106
rect 73 72 89 106
rect 23 17 89 72
rect 142 111 253 165
rect 447 129 481 384
rect 673 353 743 369
rect 673 319 689 353
rect 723 319 743 353
rect 517 283 583 299
rect 517 249 533 283
rect 567 249 583 283
rect 517 215 583 249
rect 673 285 743 319
rect 673 251 689 285
rect 723 251 743 285
rect 673 235 743 251
rect 787 353 853 369
rect 787 319 803 353
rect 837 319 853 353
rect 787 285 853 319
rect 787 251 803 285
rect 837 251 853 285
rect 787 235 853 251
rect 889 353 1031 369
rect 889 319 932 353
rect 966 319 1031 353
rect 889 285 1031 319
rect 889 251 932 285
rect 966 251 1031 285
rect 889 235 1031 251
rect 517 181 533 215
rect 567 199 583 215
rect 567 181 1007 199
rect 517 165 1007 181
rect 142 77 203 111
rect 237 77 253 111
rect 142 53 253 77
rect 345 103 411 129
rect 345 69 361 103
rect 395 69 411 103
rect 345 17 411 69
rect 447 108 569 129
rect 447 74 519 108
rect 553 74 569 108
rect 447 53 569 74
rect 619 116 685 165
rect 619 82 635 116
rect 669 82 685 116
rect 619 53 685 82
rect 777 108 843 129
rect 777 74 793 108
rect 827 74 843 108
rect 777 17 843 74
rect 941 116 1007 165
rect 941 82 957 116
rect 991 82 1007 116
rect 941 53 1007 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2111o_lp
flabel comment s 424 277 424 277 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1063778
string GDS_START 1054244
<< end >>
