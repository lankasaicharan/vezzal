magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 331 1958 704
<< pwell >>
rect 1 49 1913 241
rect 0 0 1920 49
<< scnmos >>
rect 84 47 114 215
rect 170 47 200 215
rect 256 47 286 215
rect 342 47 372 215
rect 428 47 458 215
rect 514 47 544 215
rect 600 47 630 215
rect 686 47 716 215
rect 772 47 802 215
rect 858 47 888 215
rect 944 47 974 215
rect 1030 47 1060 215
rect 1116 47 1146 215
rect 1202 47 1232 215
rect 1288 47 1318 215
rect 1374 47 1404 215
rect 1628 47 1658 215
rect 1714 47 1744 215
rect 1800 47 1830 215
<< scpmoshvt >>
rect 84 367 114 619
rect 170 367 200 619
rect 256 367 286 619
rect 342 367 372 619
rect 428 367 458 619
rect 514 367 544 619
rect 600 367 630 619
rect 686 367 716 619
rect 772 367 802 619
rect 858 367 888 619
rect 944 367 974 619
rect 1030 367 1060 619
rect 1116 367 1146 619
rect 1202 367 1232 619
rect 1288 367 1318 619
rect 1374 367 1404 619
rect 1628 367 1658 619
rect 1714 367 1744 619
rect 1800 367 1830 619
<< ndiff >>
rect 27 186 84 215
rect 27 152 39 186
rect 73 152 84 186
rect 27 101 84 152
rect 27 67 39 101
rect 73 67 84 101
rect 27 47 84 67
rect 114 178 170 215
rect 114 144 125 178
rect 159 144 170 178
rect 114 47 170 144
rect 200 123 256 215
rect 200 89 211 123
rect 245 89 256 123
rect 200 47 256 89
rect 286 178 342 215
rect 286 144 297 178
rect 331 144 342 178
rect 286 47 342 144
rect 372 123 428 215
rect 372 89 383 123
rect 417 89 428 123
rect 372 47 428 89
rect 458 178 514 215
rect 458 144 469 178
rect 503 144 514 178
rect 458 47 514 144
rect 544 123 600 215
rect 544 89 555 123
rect 589 89 600 123
rect 544 47 600 89
rect 630 178 686 215
rect 630 144 641 178
rect 675 144 686 178
rect 630 47 686 144
rect 716 203 772 215
rect 716 169 727 203
rect 761 169 772 203
rect 716 101 772 169
rect 716 67 727 101
rect 761 67 772 101
rect 716 47 772 67
rect 802 177 858 215
rect 802 143 813 177
rect 847 143 858 177
rect 802 93 858 143
rect 802 59 813 93
rect 847 59 858 93
rect 802 47 858 59
rect 888 203 944 215
rect 888 169 899 203
rect 933 169 944 203
rect 888 101 944 169
rect 888 67 899 101
rect 933 67 944 101
rect 888 47 944 67
rect 974 177 1030 215
rect 974 143 985 177
rect 1019 143 1030 177
rect 974 93 1030 143
rect 974 59 985 93
rect 1019 59 1030 93
rect 974 47 1030 59
rect 1060 203 1116 215
rect 1060 169 1071 203
rect 1105 169 1116 203
rect 1060 93 1116 169
rect 1060 59 1071 93
rect 1105 59 1116 93
rect 1060 47 1116 59
rect 1146 177 1202 215
rect 1146 143 1157 177
rect 1191 143 1202 177
rect 1146 93 1202 143
rect 1146 59 1157 93
rect 1191 59 1202 93
rect 1146 47 1202 59
rect 1232 203 1288 215
rect 1232 169 1243 203
rect 1277 169 1288 203
rect 1232 101 1288 169
rect 1232 67 1243 101
rect 1277 67 1288 101
rect 1232 47 1288 67
rect 1318 177 1374 215
rect 1318 143 1329 177
rect 1363 143 1374 177
rect 1318 93 1374 143
rect 1318 59 1329 93
rect 1363 59 1374 93
rect 1318 47 1374 59
rect 1404 203 1461 215
rect 1404 169 1415 203
rect 1449 169 1461 203
rect 1404 101 1461 169
rect 1404 67 1415 101
rect 1449 67 1461 101
rect 1404 47 1461 67
rect 1571 186 1628 215
rect 1571 152 1583 186
rect 1617 152 1628 186
rect 1571 101 1628 152
rect 1571 67 1583 101
rect 1617 67 1628 101
rect 1571 47 1628 67
rect 1658 105 1714 215
rect 1658 71 1669 105
rect 1703 71 1714 105
rect 1658 47 1714 71
rect 1744 186 1800 215
rect 1744 152 1755 186
rect 1789 152 1800 186
rect 1744 101 1800 152
rect 1744 67 1755 101
rect 1789 67 1800 101
rect 1744 47 1800 67
rect 1830 203 1887 215
rect 1830 169 1841 203
rect 1875 169 1887 203
rect 1830 93 1887 169
rect 1830 59 1841 93
rect 1875 59 1887 93
rect 1830 47 1887 59
<< pdiff >>
rect 27 599 84 619
rect 27 565 39 599
rect 73 565 84 599
rect 27 506 84 565
rect 27 472 39 506
rect 73 472 84 506
rect 27 413 84 472
rect 27 379 39 413
rect 73 379 84 413
rect 27 367 84 379
rect 114 531 170 619
rect 114 497 125 531
rect 159 497 170 531
rect 114 413 170 497
rect 114 379 125 413
rect 159 379 170 413
rect 114 367 170 379
rect 200 599 256 619
rect 200 565 211 599
rect 245 565 256 599
rect 200 481 256 565
rect 200 447 211 481
rect 245 447 256 481
rect 200 367 256 447
rect 286 531 342 619
rect 286 497 297 531
rect 331 497 342 531
rect 286 413 342 497
rect 286 379 297 413
rect 331 379 342 413
rect 286 367 342 379
rect 372 599 428 619
rect 372 565 383 599
rect 417 565 428 599
rect 372 481 428 565
rect 372 447 383 481
rect 417 447 428 481
rect 372 367 428 447
rect 458 531 514 619
rect 458 497 469 531
rect 503 497 514 531
rect 458 413 514 497
rect 458 379 469 413
rect 503 379 514 413
rect 458 367 514 379
rect 544 599 600 619
rect 544 565 555 599
rect 589 565 600 599
rect 544 481 600 565
rect 544 447 555 481
rect 589 447 600 481
rect 544 367 600 447
rect 630 531 686 619
rect 630 497 641 531
rect 675 497 686 531
rect 630 413 686 497
rect 630 379 641 413
rect 675 379 686 413
rect 630 367 686 379
rect 716 599 772 619
rect 716 565 727 599
rect 761 565 772 599
rect 716 506 772 565
rect 716 472 727 506
rect 761 472 772 506
rect 716 413 772 472
rect 716 379 727 413
rect 761 379 772 413
rect 716 367 772 379
rect 802 607 858 619
rect 802 573 813 607
rect 847 573 858 607
rect 802 481 858 573
rect 802 447 813 481
rect 847 447 858 481
rect 802 367 858 447
rect 888 599 944 619
rect 888 565 899 599
rect 933 565 944 599
rect 888 506 944 565
rect 888 472 899 506
rect 933 472 944 506
rect 888 413 944 472
rect 888 379 899 413
rect 933 379 944 413
rect 888 367 944 379
rect 974 607 1030 619
rect 974 573 985 607
rect 1019 573 1030 607
rect 974 481 1030 573
rect 974 447 985 481
rect 1019 447 1030 481
rect 974 367 1030 447
rect 1060 599 1116 619
rect 1060 565 1071 599
rect 1105 565 1116 599
rect 1060 506 1116 565
rect 1060 472 1071 506
rect 1105 472 1116 506
rect 1060 413 1116 472
rect 1060 379 1071 413
rect 1105 379 1116 413
rect 1060 367 1116 379
rect 1146 607 1202 619
rect 1146 573 1157 607
rect 1191 573 1202 607
rect 1146 481 1202 573
rect 1146 447 1157 481
rect 1191 447 1202 481
rect 1146 367 1202 447
rect 1232 599 1288 619
rect 1232 565 1243 599
rect 1277 565 1288 599
rect 1232 506 1288 565
rect 1232 472 1243 506
rect 1277 472 1288 506
rect 1232 413 1288 472
rect 1232 379 1243 413
rect 1277 379 1288 413
rect 1232 367 1288 379
rect 1318 599 1374 619
rect 1318 565 1329 599
rect 1363 565 1374 599
rect 1318 367 1374 565
rect 1404 599 1461 619
rect 1404 565 1415 599
rect 1449 565 1461 599
rect 1404 523 1461 565
rect 1404 489 1415 523
rect 1449 489 1461 523
rect 1404 367 1461 489
rect 1571 413 1628 619
rect 1571 379 1583 413
rect 1617 379 1628 413
rect 1571 367 1628 379
rect 1658 594 1714 619
rect 1658 560 1669 594
rect 1703 560 1714 594
rect 1658 367 1714 560
rect 1744 599 1800 619
rect 1744 565 1755 599
rect 1789 565 1800 599
rect 1744 506 1800 565
rect 1744 472 1755 506
rect 1789 472 1800 506
rect 1744 413 1800 472
rect 1744 379 1755 413
rect 1789 379 1800 413
rect 1744 367 1800 379
rect 1830 607 1887 619
rect 1830 573 1841 607
rect 1875 573 1887 607
rect 1830 510 1887 573
rect 1830 476 1841 510
rect 1875 476 1887 510
rect 1830 413 1887 476
rect 1830 379 1841 413
rect 1875 379 1887 413
rect 1830 367 1887 379
<< ndiffc >>
rect 39 152 73 186
rect 39 67 73 101
rect 125 144 159 178
rect 211 89 245 123
rect 297 144 331 178
rect 383 89 417 123
rect 469 144 503 178
rect 555 89 589 123
rect 641 144 675 178
rect 727 169 761 203
rect 727 67 761 101
rect 813 143 847 177
rect 813 59 847 93
rect 899 169 933 203
rect 899 67 933 101
rect 985 143 1019 177
rect 985 59 1019 93
rect 1071 169 1105 203
rect 1071 59 1105 93
rect 1157 143 1191 177
rect 1157 59 1191 93
rect 1243 169 1277 203
rect 1243 67 1277 101
rect 1329 143 1363 177
rect 1329 59 1363 93
rect 1415 169 1449 203
rect 1415 67 1449 101
rect 1583 152 1617 186
rect 1583 67 1617 101
rect 1669 71 1703 105
rect 1755 152 1789 186
rect 1755 67 1789 101
rect 1841 169 1875 203
rect 1841 59 1875 93
<< pdiffc >>
rect 39 565 73 599
rect 39 472 73 506
rect 39 379 73 413
rect 125 497 159 531
rect 125 379 159 413
rect 211 565 245 599
rect 211 447 245 481
rect 297 497 331 531
rect 297 379 331 413
rect 383 565 417 599
rect 383 447 417 481
rect 469 497 503 531
rect 469 379 503 413
rect 555 565 589 599
rect 555 447 589 481
rect 641 497 675 531
rect 641 379 675 413
rect 727 565 761 599
rect 727 472 761 506
rect 727 379 761 413
rect 813 573 847 607
rect 813 447 847 481
rect 899 565 933 599
rect 899 472 933 506
rect 899 379 933 413
rect 985 573 1019 607
rect 985 447 1019 481
rect 1071 565 1105 599
rect 1071 472 1105 506
rect 1071 379 1105 413
rect 1157 573 1191 607
rect 1157 447 1191 481
rect 1243 565 1277 599
rect 1243 472 1277 506
rect 1243 379 1277 413
rect 1329 565 1363 599
rect 1415 565 1449 599
rect 1415 489 1449 523
rect 1583 379 1617 413
rect 1669 560 1703 594
rect 1755 565 1789 599
rect 1755 472 1789 506
rect 1755 379 1789 413
rect 1841 573 1875 607
rect 1841 476 1875 510
rect 1841 379 1875 413
<< poly >>
rect 84 619 114 645
rect 170 619 200 645
rect 256 619 286 645
rect 342 619 372 645
rect 428 619 458 645
rect 514 619 544 645
rect 600 619 630 645
rect 686 619 716 645
rect 772 619 802 645
rect 858 619 888 645
rect 944 619 974 645
rect 1030 619 1060 645
rect 1116 619 1146 645
rect 1202 619 1232 645
rect 1288 619 1318 645
rect 1374 619 1404 645
rect 1628 619 1658 645
rect 1714 619 1744 645
rect 1800 619 1830 645
rect 84 329 114 367
rect 170 329 200 367
rect 256 329 286 367
rect 342 329 372 367
rect 428 329 458 367
rect 514 329 544 367
rect 600 329 630 367
rect 686 329 716 367
rect 84 313 716 329
rect 772 345 802 367
rect 858 345 888 367
rect 944 345 974 367
rect 1030 345 1060 367
rect 1116 345 1146 367
rect 1202 345 1232 367
rect 1288 345 1318 367
rect 1374 345 1404 367
rect 1628 345 1658 367
rect 772 315 1658 345
rect 84 279 235 313
rect 269 279 303 313
rect 337 279 371 313
rect 405 279 439 313
rect 473 279 507 313
rect 541 279 575 313
rect 609 279 643 313
rect 677 279 716 313
rect 84 263 716 279
rect 1573 287 1658 315
rect 84 215 114 263
rect 170 215 200 263
rect 256 215 286 263
rect 342 215 372 263
rect 428 215 458 263
rect 514 215 544 263
rect 600 215 630 263
rect 686 215 716 263
rect 772 237 1513 267
rect 1573 253 1589 287
rect 1623 253 1658 287
rect 1573 237 1658 253
rect 772 215 802 237
rect 858 215 888 237
rect 944 215 974 237
rect 1030 215 1060 237
rect 1116 215 1146 237
rect 1202 215 1232 237
rect 1288 215 1318 237
rect 1374 215 1404 237
rect 1483 185 1513 237
rect 1628 215 1658 237
rect 1714 303 1744 367
rect 1800 303 1830 367
rect 1714 287 1830 303
rect 1714 253 1757 287
rect 1791 253 1830 287
rect 1714 237 1830 253
rect 1714 215 1744 237
rect 1800 215 1830 237
rect 1483 169 1549 185
rect 1483 135 1499 169
rect 1533 135 1549 169
rect 1483 101 1549 135
rect 1483 67 1499 101
rect 1533 67 1549 101
rect 1483 51 1549 67
rect 84 21 114 47
rect 170 21 200 47
rect 256 21 286 47
rect 342 21 372 47
rect 428 21 458 47
rect 514 21 544 47
rect 600 21 630 47
rect 686 21 716 47
rect 772 21 802 47
rect 858 21 888 47
rect 944 21 974 47
rect 1030 21 1060 47
rect 1116 21 1146 47
rect 1202 21 1232 47
rect 1288 21 1318 47
rect 1374 21 1404 47
rect 1628 21 1658 47
rect 1714 21 1744 47
rect 1800 21 1830 47
<< polycont >>
rect 235 279 269 313
rect 303 279 337 313
rect 371 279 405 313
rect 439 279 473 313
rect 507 279 541 313
rect 575 279 609 313
rect 643 279 677 313
rect 1589 253 1623 287
rect 1757 253 1791 287
rect 1499 135 1533 169
rect 1499 67 1533 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 23 599 761 615
rect 23 565 39 599
rect 73 581 211 599
rect 73 565 89 581
rect 23 506 89 565
rect 195 565 211 581
rect 245 581 383 599
rect 23 472 39 506
rect 73 472 89 506
rect 23 413 89 472
rect 23 379 39 413
rect 73 379 89 413
rect 23 363 89 379
rect 125 531 159 547
rect 125 413 159 497
rect 195 481 245 565
rect 417 581 555 599
rect 195 447 211 481
rect 195 431 245 447
rect 281 531 347 547
rect 281 497 297 531
rect 331 497 347 531
rect 281 413 347 497
rect 383 481 417 565
rect 589 581 727 599
rect 383 431 417 447
rect 453 531 519 547
rect 453 497 469 531
rect 503 497 519 531
rect 281 397 297 413
rect 159 379 297 397
rect 331 397 347 413
rect 453 413 519 497
rect 555 481 589 565
rect 555 431 589 447
rect 625 531 691 547
rect 625 497 641 531
rect 675 497 691 531
rect 453 397 469 413
rect 331 379 469 397
rect 503 397 519 413
rect 625 413 691 497
rect 625 397 641 413
rect 503 379 641 397
rect 675 379 691 413
rect 125 363 691 379
rect 727 506 761 565
rect 727 413 761 472
rect 797 607 847 649
rect 797 573 813 607
rect 797 481 847 573
rect 797 447 813 481
rect 797 431 847 447
rect 883 599 949 615
rect 883 565 899 599
rect 933 565 949 599
rect 883 506 949 565
rect 883 472 899 506
rect 933 472 949 506
rect 883 413 949 472
rect 985 607 1019 649
rect 985 481 1019 573
rect 985 431 1019 447
rect 1055 599 1121 615
rect 1055 565 1071 599
rect 1105 565 1121 599
rect 1055 506 1121 565
rect 1055 472 1071 506
rect 1105 472 1121 506
rect 883 397 899 413
rect 761 379 899 397
rect 933 397 949 413
rect 1055 413 1121 472
rect 1157 607 1191 649
rect 1157 481 1191 573
rect 1157 431 1191 447
rect 1227 599 1277 615
rect 1227 565 1243 599
rect 1227 507 1277 565
rect 1313 599 1363 649
rect 1313 565 1329 599
rect 1313 541 1363 565
rect 1399 599 1465 615
rect 1399 565 1415 599
rect 1449 565 1465 599
rect 1399 523 1465 565
rect 1653 594 1703 649
rect 1653 560 1669 594
rect 1653 531 1703 560
rect 1739 599 1805 615
rect 1739 565 1755 599
rect 1789 565 1805 599
rect 1399 507 1415 523
rect 1227 506 1415 507
rect 1227 472 1243 506
rect 1277 489 1415 506
rect 1449 489 1465 523
rect 1739 506 1805 565
rect 1739 497 1755 506
rect 1277 473 1465 489
rect 1055 397 1071 413
rect 933 379 1071 397
rect 1105 397 1121 413
rect 1227 413 1277 472
rect 1499 472 1755 497
rect 1789 472 1805 506
rect 1499 463 1805 472
rect 1499 439 1533 463
rect 1227 397 1243 413
rect 1105 379 1243 397
rect 727 363 1277 379
rect 1311 405 1533 439
rect 1567 413 1633 429
rect 125 282 159 363
rect 1311 329 1345 405
rect 1567 379 1583 413
rect 1617 379 1633 413
rect 1567 371 1633 379
rect 219 313 1345 329
rect 25 236 167 282
rect 219 279 235 313
rect 269 279 303 313
rect 337 279 371 313
rect 405 279 439 313
rect 473 279 507 313
rect 541 279 575 313
rect 609 279 643 313
rect 677 295 1345 313
rect 1483 337 1633 371
rect 1673 413 1805 463
rect 1673 379 1755 413
rect 1789 379 1805 413
rect 1673 363 1805 379
rect 1841 607 1891 649
rect 1875 573 1891 607
rect 1841 510 1891 573
rect 1875 476 1891 510
rect 1841 413 1891 476
rect 1875 379 1891 413
rect 1841 363 1891 379
rect 677 279 693 295
rect 219 263 693 279
rect 109 229 167 236
rect 23 186 73 202
rect 23 152 39 186
rect 23 101 73 152
rect 109 195 691 229
rect 109 178 175 195
rect 109 144 125 178
rect 159 144 175 178
rect 281 178 347 195
rect 109 119 175 144
rect 211 123 245 161
rect 23 67 39 101
rect 281 144 297 178
rect 331 144 347 178
rect 453 178 519 195
rect 281 119 347 144
rect 383 123 417 161
rect 211 85 245 89
rect 453 144 469 178
rect 503 144 519 178
rect 625 178 691 195
rect 453 119 519 144
rect 555 123 589 161
rect 383 85 417 89
rect 625 144 641 178
rect 675 144 691 178
rect 625 119 691 144
rect 727 227 1449 261
rect 727 203 761 227
rect 883 203 949 227
rect 555 85 589 89
rect 727 101 761 169
rect 73 67 727 85
rect 23 51 761 67
rect 797 177 847 193
rect 797 143 813 177
rect 797 93 847 143
rect 797 59 813 93
rect 797 17 847 59
rect 883 169 899 203
rect 933 169 949 203
rect 1055 203 1121 227
rect 883 101 949 169
rect 883 67 899 101
rect 933 67 949 101
rect 883 51 949 67
rect 985 177 1019 193
rect 985 93 1019 143
rect 1055 169 1071 203
rect 1105 169 1121 203
rect 1227 203 1293 227
rect 1055 93 1121 169
rect 1055 59 1071 93
rect 1105 59 1121 93
rect 1157 177 1191 193
rect 1157 93 1191 143
rect 985 17 1019 59
rect 1157 17 1191 59
rect 1227 169 1243 203
rect 1277 169 1293 203
rect 1399 203 1449 227
rect 1227 101 1293 169
rect 1227 67 1243 101
rect 1277 67 1293 101
rect 1227 51 1293 67
rect 1329 177 1363 193
rect 1329 93 1363 143
rect 1329 17 1363 59
rect 1399 169 1415 203
rect 1399 101 1449 169
rect 1399 67 1415 101
rect 1399 51 1449 67
rect 1483 202 1527 337
rect 1561 287 1639 303
rect 1561 253 1589 287
rect 1623 253 1639 287
rect 1561 236 1639 253
rect 1673 202 1707 363
rect 1741 287 1807 303
rect 1741 253 1757 287
rect 1791 253 1807 287
rect 1741 236 1807 253
rect 1841 203 1891 219
rect 1483 186 1633 202
rect 1483 169 1583 186
rect 1483 135 1499 169
rect 1533 152 1583 169
rect 1617 152 1633 186
rect 1673 186 1805 202
rect 1673 168 1755 186
rect 1533 135 1633 152
rect 1483 101 1633 135
rect 1739 152 1755 168
rect 1789 152 1805 186
rect 1483 67 1499 101
rect 1533 67 1583 101
rect 1617 67 1633 101
rect 1483 51 1633 67
rect 1669 105 1703 134
rect 1669 17 1703 71
rect 1739 101 1805 152
rect 1739 67 1755 101
rect 1789 67 1805 101
rect 1739 51 1805 67
rect 1875 169 1891 203
rect 1841 93 1891 169
rect 1875 59 1891 93
rect 1841 17 1891 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ebufn_8
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3324676
string GDS_START 3310924
<< end >>
