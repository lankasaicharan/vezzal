magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 29 49 718 162
rect 0 0 768 49
<< scnmos >>
rect 108 52 138 136
rect 194 52 224 136
rect 417 52 447 136
rect 503 52 533 136
rect 609 52 639 136
<< scpmoshvt >>
rect 81 482 111 610
rect 186 526 216 610
rect 437 458 467 586
rect 523 458 553 586
rect 609 458 639 586
<< ndiff >>
rect 55 111 108 136
rect 55 77 63 111
rect 97 77 108 111
rect 55 52 108 77
rect 138 111 194 136
rect 138 77 149 111
rect 183 77 194 111
rect 138 52 194 77
rect 224 111 277 136
rect 224 77 235 111
rect 269 77 277 111
rect 224 52 277 77
rect 364 111 417 136
rect 364 77 372 111
rect 406 77 417 111
rect 364 52 417 77
rect 447 111 503 136
rect 447 77 458 111
rect 492 77 503 111
rect 447 52 503 77
rect 533 52 609 136
rect 639 111 692 136
rect 639 77 650 111
rect 684 77 692 111
rect 639 52 692 77
<< pdiff >>
rect 28 596 81 610
rect 28 562 36 596
rect 70 562 81 596
rect 28 528 81 562
rect 28 494 36 528
rect 70 494 81 528
rect 28 482 81 494
rect 111 598 186 610
rect 111 564 132 598
rect 166 564 186 598
rect 111 530 186 564
rect 111 496 122 530
rect 156 526 186 530
rect 216 585 269 610
rect 216 551 227 585
rect 261 551 269 585
rect 216 526 269 551
rect 384 572 437 586
rect 384 538 392 572
rect 426 538 437 572
rect 156 496 164 526
rect 111 482 164 496
rect 384 504 437 538
rect 384 470 392 504
rect 426 470 437 504
rect 384 458 437 470
rect 467 572 523 586
rect 467 538 478 572
rect 512 538 523 572
rect 467 504 523 538
rect 467 470 478 504
rect 512 470 523 504
rect 467 458 523 470
rect 553 574 609 586
rect 553 540 564 574
rect 598 540 609 574
rect 553 506 609 540
rect 553 472 564 506
rect 598 472 609 506
rect 553 458 609 472
rect 639 572 692 586
rect 639 538 650 572
rect 684 538 692 572
rect 639 504 692 538
rect 639 470 650 504
rect 684 470 692 504
rect 639 458 692 470
<< ndiffc >>
rect 63 77 97 111
rect 149 77 183 111
rect 235 77 269 111
rect 372 77 406 111
rect 458 77 492 111
rect 650 77 684 111
<< pdiffc >>
rect 36 562 70 596
rect 36 494 70 528
rect 132 564 166 598
rect 122 496 156 530
rect 227 551 261 585
rect 392 538 426 572
rect 392 470 426 504
rect 478 538 512 572
rect 478 470 512 504
rect 564 540 598 574
rect 564 472 598 506
rect 650 538 684 572
rect 650 470 684 504
<< poly >>
rect 81 610 111 636
rect 186 610 216 636
rect 437 586 467 612
rect 523 586 553 612
rect 609 586 639 612
rect 81 346 111 482
rect 72 330 138 346
rect 72 296 88 330
rect 122 296 138 330
rect 72 262 138 296
rect 72 228 88 262
rect 122 228 138 262
rect 72 212 138 228
rect 108 136 138 212
rect 186 292 216 526
rect 264 416 330 432
rect 264 382 280 416
rect 314 382 330 416
rect 264 366 330 382
rect 437 380 467 458
rect 300 292 330 366
rect 417 350 467 380
rect 186 276 252 292
rect 186 242 202 276
rect 236 242 252 276
rect 186 208 252 242
rect 186 174 202 208
rect 236 174 252 208
rect 186 158 252 174
rect 300 276 366 292
rect 300 242 316 276
rect 350 242 366 276
rect 300 208 366 242
rect 300 174 316 208
rect 350 188 366 208
rect 417 188 447 350
rect 523 302 553 458
rect 609 302 639 458
rect 350 174 447 188
rect 300 158 447 174
rect 495 286 561 302
rect 495 252 511 286
rect 545 252 561 286
rect 495 218 561 252
rect 495 184 511 218
rect 545 184 561 218
rect 495 168 561 184
rect 609 286 675 302
rect 609 252 625 286
rect 659 252 675 286
rect 609 218 675 252
rect 609 184 625 218
rect 659 184 675 218
rect 609 168 675 184
rect 194 136 224 158
rect 417 136 447 158
rect 503 136 533 168
rect 609 136 639 168
rect 108 26 138 52
rect 194 26 224 52
rect 417 26 447 52
rect 503 26 533 52
rect 609 26 639 52
<< polycont >>
rect 88 296 122 330
rect 88 228 122 262
rect 280 382 314 416
rect 202 242 236 276
rect 202 174 236 208
rect 316 242 350 276
rect 316 174 350 208
rect 511 252 545 286
rect 511 184 545 218
rect 625 252 659 286
rect 625 184 659 218
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 18 596 84 612
rect 18 562 36 596
rect 70 562 84 596
rect 18 528 84 562
rect 18 494 36 528
rect 70 494 84 528
rect 18 390 84 494
rect 118 598 177 649
rect 118 564 132 598
rect 166 564 177 598
rect 118 530 177 564
rect 118 496 122 530
rect 156 496 177 530
rect 118 480 177 496
rect 211 585 277 601
rect 211 551 227 585
rect 261 551 277 585
rect 211 432 277 551
rect 376 572 434 588
rect 376 538 392 572
rect 426 538 434 572
rect 376 504 434 538
rect 376 470 392 504
rect 426 470 434 504
rect 211 416 330 432
rect 18 127 52 390
rect 211 382 280 416
rect 314 382 330 416
rect 211 380 330 382
rect 376 346 434 470
rect 468 572 520 588
rect 468 538 478 572
rect 512 538 520 572
rect 468 504 520 538
rect 468 470 478 504
rect 512 470 520 504
rect 468 420 520 470
rect 554 574 607 649
rect 554 540 564 574
rect 598 540 607 574
rect 554 506 607 540
rect 554 472 564 506
rect 598 472 607 506
rect 554 456 607 472
rect 641 572 700 588
rect 641 538 650 572
rect 684 538 700 572
rect 641 504 700 538
rect 641 470 650 504
rect 684 470 700 504
rect 641 420 700 470
rect 468 386 700 420
rect 86 330 475 346
rect 86 296 88 330
rect 122 312 475 330
rect 122 296 139 312
rect 86 262 139 296
rect 86 228 88 262
rect 122 228 139 262
rect 86 212 139 228
rect 186 276 266 278
rect 186 242 202 276
rect 236 242 266 276
rect 186 208 266 242
rect 186 174 202 208
rect 236 174 266 208
rect 186 166 266 174
rect 300 242 316 276
rect 350 242 366 276
rect 300 208 366 242
rect 300 174 316 208
rect 350 174 366 208
rect 300 127 334 174
rect 441 127 475 312
rect 509 286 559 351
rect 509 252 511 286
rect 545 252 559 286
rect 509 218 559 252
rect 509 184 511 218
rect 545 184 559 218
rect 509 161 559 184
rect 593 286 675 352
rect 593 252 625 286
rect 659 252 675 286
rect 593 218 675 252
rect 593 184 625 218
rect 659 184 675 218
rect 593 161 675 184
rect 18 111 107 127
rect 18 77 63 111
rect 97 77 107 111
rect 18 61 107 77
rect 141 111 191 127
rect 141 77 149 111
rect 183 77 191 111
rect 141 17 191 77
rect 225 111 334 127
rect 225 77 235 111
rect 269 77 334 111
rect 225 61 334 77
rect 368 111 407 127
rect 368 77 372 111
rect 406 77 407 111
rect 368 17 407 77
rect 441 111 508 127
rect 441 77 458 111
rect 492 77 508 111
rect 441 61 508 77
rect 634 111 700 127
rect 634 77 650 111
rect 684 77 700 111
rect 634 17 700 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21bo_0
flabel comment s 313 317 313 317 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3778520
string GDS_START 3770724
<< end >>
