magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 17 49 667 259
rect 0 0 672 49
<< scnmos >>
rect 96 65 126 233
rect 182 65 212 233
rect 268 65 298 233
rect 362 65 392 233
rect 472 65 502 233
rect 558 65 588 233
<< scpmoshvt >>
rect 96 367 126 619
rect 182 367 212 619
rect 276 367 306 619
rect 362 367 392 619
rect 458 367 488 619
rect 544 367 574 619
<< ndiff >>
rect 43 192 96 233
rect 43 158 51 192
rect 85 158 96 192
rect 43 111 96 158
rect 43 77 51 111
rect 85 77 96 111
rect 43 65 96 77
rect 126 225 182 233
rect 126 191 137 225
rect 171 191 182 225
rect 126 153 182 191
rect 126 119 137 153
rect 171 119 182 153
rect 126 65 182 119
rect 212 225 268 233
rect 212 191 223 225
rect 257 191 268 225
rect 212 111 268 191
rect 212 77 223 111
rect 257 77 268 111
rect 212 65 268 77
rect 298 183 362 233
rect 298 149 313 183
rect 347 149 362 183
rect 298 107 362 149
rect 298 73 313 107
rect 347 73 362 107
rect 298 65 362 73
rect 392 107 472 233
rect 392 73 413 107
rect 447 73 472 107
rect 392 65 472 73
rect 502 183 558 233
rect 502 149 513 183
rect 547 149 558 183
rect 502 107 558 149
rect 502 73 513 107
rect 547 73 558 107
rect 502 65 558 73
rect 588 221 641 233
rect 588 187 599 221
rect 633 187 641 221
rect 588 111 641 187
rect 588 77 599 111
rect 633 77 641 111
rect 588 65 641 77
<< pdiff >>
rect 43 607 96 619
rect 43 573 51 607
rect 85 573 96 607
rect 43 513 96 573
rect 43 479 51 513
rect 85 479 96 513
rect 43 418 96 479
rect 43 384 51 418
rect 85 384 96 418
rect 43 367 96 384
rect 126 599 182 619
rect 126 565 137 599
rect 171 565 182 599
rect 126 505 182 565
rect 126 471 137 505
rect 171 471 182 505
rect 126 409 182 471
rect 126 375 137 409
rect 171 375 182 409
rect 126 367 182 375
rect 212 568 276 619
rect 212 534 227 568
rect 261 534 276 568
rect 212 367 276 534
rect 306 599 362 619
rect 306 565 317 599
rect 351 565 362 599
rect 306 492 362 565
rect 306 458 317 492
rect 351 458 362 492
rect 306 367 362 458
rect 392 574 458 619
rect 392 540 407 574
rect 441 540 458 574
rect 392 367 458 540
rect 488 599 544 619
rect 488 565 499 599
rect 533 565 544 599
rect 488 492 544 565
rect 488 458 499 492
rect 533 458 544 492
rect 488 367 544 458
rect 574 607 627 619
rect 574 573 585 607
rect 619 573 627 607
rect 574 506 627 573
rect 574 472 585 506
rect 619 472 627 506
rect 574 413 627 472
rect 574 379 585 413
rect 619 379 627 413
rect 574 367 627 379
<< ndiffc >>
rect 51 158 85 192
rect 51 77 85 111
rect 137 191 171 225
rect 137 119 171 153
rect 223 191 257 225
rect 223 77 257 111
rect 313 149 347 183
rect 313 73 347 107
rect 413 73 447 107
rect 513 149 547 183
rect 513 73 547 107
rect 599 187 633 221
rect 599 77 633 111
<< pdiffc >>
rect 51 573 85 607
rect 51 479 85 513
rect 51 384 85 418
rect 137 565 171 599
rect 137 471 171 505
rect 137 375 171 409
rect 227 534 261 568
rect 317 565 351 599
rect 317 458 351 492
rect 407 540 441 574
rect 499 565 533 599
rect 499 458 533 492
rect 585 573 619 607
rect 585 472 619 506
rect 585 379 619 413
<< poly >>
rect 96 619 126 645
rect 182 619 212 645
rect 276 619 306 645
rect 362 619 392 645
rect 458 619 488 645
rect 544 619 574 645
rect 96 321 126 367
rect 35 305 126 321
rect 35 271 51 305
rect 85 285 126 305
rect 182 285 212 367
rect 276 335 306 367
rect 362 335 392 367
rect 458 335 488 367
rect 85 271 212 285
rect 35 255 212 271
rect 254 319 320 335
rect 254 285 270 319
rect 304 285 320 319
rect 254 269 320 285
rect 362 319 488 335
rect 362 285 378 319
rect 412 299 488 319
rect 544 335 574 367
rect 544 319 610 335
rect 412 285 502 299
rect 362 269 502 285
rect 544 285 560 319
rect 594 285 610 319
rect 544 269 610 285
rect 96 233 126 255
rect 182 233 212 255
rect 268 233 298 269
rect 362 233 392 269
rect 472 233 502 269
rect 558 233 588 269
rect 96 39 126 65
rect 182 39 212 65
rect 268 39 298 65
rect 362 39 392 65
rect 472 39 502 65
rect 558 39 588 65
<< polycont >>
rect 51 271 85 305
rect 270 285 304 319
rect 378 285 412 319
rect 560 285 594 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 35 607 101 649
rect 35 573 51 607
rect 85 573 101 607
rect 35 513 101 573
rect 35 479 51 513
rect 85 479 101 513
rect 35 418 101 479
rect 35 384 51 418
rect 85 384 101 418
rect 135 599 177 615
rect 135 565 137 599
rect 171 565 177 599
rect 135 505 177 565
rect 211 568 277 649
rect 211 534 227 568
rect 261 534 277 568
rect 211 526 277 534
rect 311 599 357 615
rect 311 565 317 599
rect 351 565 357 599
rect 135 471 137 505
rect 171 492 177 505
rect 311 498 357 565
rect 391 574 457 649
rect 391 540 407 574
rect 441 540 457 574
rect 391 532 457 540
rect 491 599 549 615
rect 491 565 499 599
rect 533 565 549 599
rect 491 498 549 565
rect 311 492 549 498
rect 171 471 317 492
rect 135 458 317 471
rect 351 458 499 492
rect 533 458 549 492
rect 583 607 635 649
rect 583 573 585 607
rect 619 573 635 607
rect 583 506 635 573
rect 583 472 585 506
rect 619 472 635 506
rect 135 409 187 458
rect 135 375 137 409
rect 171 375 187 409
rect 17 305 101 350
rect 17 271 51 305
rect 85 271 101 305
rect 17 242 101 271
rect 135 225 187 375
rect 221 384 549 424
rect 221 319 320 384
rect 221 285 270 319
rect 304 285 320 319
rect 362 319 464 350
rect 362 285 378 319
rect 412 285 464 319
rect 498 329 549 384
rect 583 413 635 472
rect 583 379 585 413
rect 619 379 635 413
rect 583 363 635 379
rect 498 319 610 329
rect 498 285 560 319
rect 594 285 610 319
rect 135 214 137 225
rect 35 192 87 208
rect 35 158 51 192
rect 85 158 87 192
rect 35 111 87 158
rect 121 191 137 214
rect 171 191 187 225
rect 121 153 187 191
rect 121 119 137 153
rect 171 119 187 153
rect 221 225 649 251
rect 221 191 223 225
rect 257 221 649 225
rect 257 217 599 221
rect 257 191 263 217
rect 35 77 51 111
rect 85 85 87 111
rect 221 111 263 191
rect 597 187 599 217
rect 633 187 649 221
rect 221 85 223 111
rect 85 77 223 85
rect 257 77 263 111
rect 35 51 263 77
rect 297 149 313 183
rect 347 149 513 183
rect 547 149 563 183
rect 297 107 363 149
rect 297 73 313 107
rect 347 73 363 107
rect 297 57 363 73
rect 397 107 463 115
rect 397 73 413 107
rect 447 73 463 107
rect 397 17 463 73
rect 497 107 563 149
rect 497 73 513 107
rect 547 73 563 107
rect 497 57 563 73
rect 597 111 649 187
rect 597 77 599 111
rect 633 77 649 111
rect 597 61 649 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand3_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 401686
string GDS_START 394936
<< end >>
