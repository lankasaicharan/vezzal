magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1490 1975
<< nwell >>
rect -38 331 230 704
<< pwell >>
rect 3 49 191 180
rect 0 0 192 49
<< scnmos >>
rect 82 70 112 154
<< scpmoshvt >>
rect 82 462 112 546
<< ndiff >>
rect 29 116 82 154
rect 29 82 37 116
rect 71 82 82 116
rect 29 70 82 82
rect 112 139 165 154
rect 112 105 123 139
rect 157 105 165 139
rect 112 70 165 105
<< pdiff >>
rect 29 522 82 546
rect 29 488 37 522
rect 71 488 82 522
rect 29 462 82 488
rect 112 520 165 546
rect 112 486 123 520
rect 157 486 165 520
rect 112 462 165 486
<< ndiffc >>
rect 37 82 71 116
rect 123 105 157 139
<< pdiffc >>
rect 37 488 71 522
rect 123 486 157 520
<< poly >>
rect 82 546 112 572
rect 82 325 112 462
rect 21 309 112 325
rect 21 275 37 309
rect 71 275 112 309
rect 21 241 112 275
rect 21 207 37 241
rect 71 207 112 241
rect 21 191 112 207
rect 82 154 112 191
rect 82 44 112 70
<< polycont >>
rect 37 275 71 309
rect 37 207 71 241
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 33 522 75 649
rect 33 488 37 522
rect 71 488 75 522
rect 33 460 75 488
rect 119 520 161 592
rect 119 486 123 520
rect 157 486 161 520
rect 31 309 71 424
rect 31 275 37 309
rect 31 241 71 275
rect 31 207 37 241
rect 31 191 71 207
rect 31 168 65 191
rect 119 139 161 486
rect 33 116 71 132
rect 33 82 37 116
rect 119 105 123 139
rect 157 105 161 139
rect 119 89 161 105
rect 33 17 71 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 31 -17 65 17
rect 127 -17 161 17
<< metal1 >>
rect 0 683 192 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 0 617 192 649
rect 0 17 192 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
rect 0 -49 192 -17
<< labels >>
flabel pwell s 0 0 192 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 192 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 inv_0
flabel metal1 s 0 617 192 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 192 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 192 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4479126
string GDS_START 4475486
<< end >>
