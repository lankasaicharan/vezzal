magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
rect 181 329 647 331
<< pwell >>
rect 1 49 860 241
rect 0 0 960 49
<< scnmos >>
rect 80 131 110 215
rect 282 47 312 215
rect 389 47 419 215
rect 493 47 523 215
rect 579 47 609 215
rect 665 47 695 215
rect 751 47 781 215
<< scpmoshvt >>
rect 80 508 110 592
rect 270 365 300 617
rect 356 365 386 617
rect 442 365 472 617
rect 528 365 558 617
rect 763 367 793 619
rect 849 367 879 619
<< ndiff >>
rect 27 190 80 215
rect 27 156 35 190
rect 69 156 80 190
rect 27 131 80 156
rect 110 184 282 215
rect 110 150 121 184
rect 155 172 282 184
rect 155 150 237 172
rect 110 138 237 150
rect 271 138 282 172
rect 110 131 282 138
rect 229 93 282 131
rect 229 59 237 93
rect 271 59 282 93
rect 229 47 282 59
rect 312 207 389 215
rect 312 173 335 207
rect 369 173 389 207
rect 312 101 389 173
rect 312 67 335 101
rect 369 67 389 101
rect 312 47 389 67
rect 419 163 493 215
rect 419 129 440 163
rect 474 129 493 163
rect 419 89 493 129
rect 419 55 440 89
rect 474 55 493 89
rect 419 47 493 55
rect 523 203 579 215
rect 523 169 534 203
rect 568 169 579 203
rect 523 101 579 169
rect 523 67 534 101
rect 568 67 579 101
rect 523 47 579 67
rect 609 165 665 215
rect 609 131 620 165
rect 654 131 665 165
rect 609 89 665 131
rect 609 55 620 89
rect 654 55 665 89
rect 609 47 665 55
rect 695 203 751 215
rect 695 169 706 203
rect 740 169 751 203
rect 695 101 751 169
rect 695 67 706 101
rect 740 67 751 101
rect 695 47 751 67
rect 781 203 834 215
rect 781 169 792 203
rect 826 169 834 203
rect 781 93 834 169
rect 781 59 792 93
rect 826 59 834 93
rect 781 47 834 59
<< pdiff >>
rect 217 599 270 617
rect 27 567 80 592
rect 27 533 35 567
rect 69 533 80 567
rect 27 508 80 533
rect 110 570 163 592
rect 110 536 121 570
rect 155 536 163 570
rect 110 508 163 536
rect 217 565 225 599
rect 259 565 270 599
rect 217 502 270 565
rect 217 468 225 502
rect 259 468 270 502
rect 217 411 270 468
rect 217 377 225 411
rect 259 377 270 411
rect 217 365 270 377
rect 300 547 356 617
rect 300 513 311 547
rect 345 513 356 547
rect 300 477 356 513
rect 300 443 311 477
rect 345 443 356 477
rect 300 407 356 443
rect 300 373 311 407
rect 345 373 356 407
rect 300 365 356 373
rect 386 599 442 617
rect 386 565 397 599
rect 431 565 442 599
rect 386 502 442 565
rect 386 468 397 502
rect 431 468 442 502
rect 386 411 442 468
rect 386 377 397 411
rect 431 377 442 411
rect 386 365 442 377
rect 472 547 528 617
rect 472 513 483 547
rect 517 513 528 547
rect 472 477 528 513
rect 472 443 483 477
rect 517 443 528 477
rect 472 407 528 443
rect 472 373 483 407
rect 517 373 528 407
rect 472 365 528 373
rect 558 599 611 617
rect 558 565 569 599
rect 603 565 611 599
rect 558 502 611 565
rect 558 468 569 502
rect 603 468 611 502
rect 558 365 611 468
rect 710 607 763 619
rect 710 573 718 607
rect 752 573 763 607
rect 710 490 763 573
rect 710 456 718 490
rect 752 456 763 490
rect 710 367 763 456
rect 793 599 849 619
rect 793 565 804 599
rect 838 565 849 599
rect 793 515 849 565
rect 793 481 804 515
rect 838 481 849 515
rect 793 434 849 481
rect 793 400 804 434
rect 838 400 849 434
rect 793 367 849 400
rect 879 607 932 619
rect 879 573 890 607
rect 924 573 932 607
rect 879 511 932 573
rect 879 477 890 511
rect 924 477 932 511
rect 879 418 932 477
rect 879 384 890 418
rect 924 384 932 418
rect 879 367 932 384
<< ndiffc >>
rect 35 156 69 190
rect 121 150 155 184
rect 237 138 271 172
rect 237 59 271 93
rect 335 173 369 207
rect 335 67 369 101
rect 440 129 474 163
rect 440 55 474 89
rect 534 169 568 203
rect 534 67 568 101
rect 620 131 654 165
rect 620 55 654 89
rect 706 169 740 203
rect 706 67 740 101
rect 792 169 826 203
rect 792 59 826 93
<< pdiffc >>
rect 35 533 69 567
rect 121 536 155 570
rect 225 565 259 599
rect 225 468 259 502
rect 225 377 259 411
rect 311 513 345 547
rect 311 443 345 477
rect 311 373 345 407
rect 397 565 431 599
rect 397 468 431 502
rect 397 377 431 411
rect 483 513 517 547
rect 483 443 517 477
rect 483 373 517 407
rect 569 565 603 599
rect 569 468 603 502
rect 718 573 752 607
rect 718 456 752 490
rect 804 565 838 599
rect 804 481 838 515
rect 804 400 838 434
rect 890 573 924 607
rect 890 477 924 511
rect 890 384 924 418
<< poly >>
rect 80 592 110 618
rect 270 617 300 643
rect 356 617 386 643
rect 442 617 472 643
rect 528 617 558 643
rect 763 619 793 645
rect 849 619 879 645
rect 80 424 110 508
rect 44 408 110 424
rect 44 374 60 408
rect 94 374 110 408
rect 44 340 110 374
rect 44 306 60 340
rect 94 306 110 340
rect 44 290 110 306
rect 270 303 300 365
rect 356 303 386 365
rect 442 333 472 365
rect 528 333 558 365
rect 763 335 793 367
rect 849 335 879 367
rect 442 317 622 333
rect 442 303 504 317
rect 80 215 110 290
rect 158 287 386 303
rect 158 253 174 287
rect 208 253 251 287
rect 285 267 386 287
rect 488 283 504 303
rect 538 283 572 317
rect 606 283 622 317
rect 488 267 622 283
rect 665 319 879 335
rect 665 285 693 319
rect 727 285 761 319
rect 795 285 829 319
rect 863 285 879 319
rect 665 269 879 285
rect 285 253 419 267
rect 158 237 419 253
rect 282 215 312 237
rect 389 215 419 237
rect 493 215 523 267
rect 579 215 609 267
rect 665 215 695 269
rect 751 215 781 269
rect 80 105 110 131
rect 282 21 312 47
rect 389 21 419 47
rect 493 21 523 47
rect 579 21 609 47
rect 665 21 695 47
rect 751 21 781 47
<< polycont >>
rect 60 374 94 408
rect 60 306 94 340
rect 174 253 208 287
rect 251 253 285 287
rect 504 283 538 317
rect 572 283 606 317
rect 693 285 727 319
rect 761 285 795 319
rect 829 285 863 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 19 567 71 583
rect 19 533 35 567
rect 69 533 71 567
rect 19 494 71 533
rect 105 570 171 649
rect 105 536 121 570
rect 155 536 171 570
rect 105 528 171 536
rect 219 599 619 615
rect 219 565 225 599
rect 259 581 397 599
rect 259 565 261 581
rect 219 502 261 565
rect 395 565 397 581
rect 431 581 569 599
rect 431 565 433 581
rect 19 460 185 494
rect 17 408 94 426
rect 17 374 60 408
rect 17 340 94 374
rect 17 306 60 340
rect 17 290 94 306
rect 151 303 185 460
rect 219 468 225 502
rect 259 468 261 502
rect 219 411 261 468
rect 219 377 225 411
rect 259 377 261 411
rect 219 361 261 377
rect 295 513 311 547
rect 345 513 361 547
rect 295 477 361 513
rect 295 443 311 477
rect 345 443 361 477
rect 295 407 361 443
rect 295 373 311 407
rect 345 373 361 407
rect 295 369 361 373
rect 151 287 285 303
rect 151 256 174 287
rect 19 253 174 256
rect 208 253 251 287
rect 19 237 285 253
rect 19 222 185 237
rect 319 233 361 369
rect 395 502 433 565
rect 567 565 569 581
rect 603 565 619 599
rect 395 468 397 502
rect 431 468 433 502
rect 395 411 433 468
rect 395 377 397 411
rect 431 377 433 411
rect 395 361 433 377
rect 467 513 483 547
rect 517 513 533 547
rect 467 477 533 513
rect 467 443 483 477
rect 517 443 533 477
rect 567 502 619 565
rect 567 468 569 502
rect 603 468 619 502
rect 567 452 619 468
rect 702 607 768 649
rect 702 573 718 607
rect 752 573 768 607
rect 702 490 768 573
rect 702 456 718 490
rect 752 456 768 490
rect 702 452 768 456
rect 802 599 838 615
rect 802 565 804 599
rect 802 515 838 565
rect 802 481 804 515
rect 467 418 533 443
rect 802 434 838 481
rect 802 418 804 434
rect 467 407 804 418
rect 467 373 483 407
rect 517 400 804 407
rect 517 384 838 400
rect 874 607 940 649
rect 874 573 890 607
rect 924 573 940 607
rect 874 511 940 573
rect 874 477 890 511
rect 924 477 940 511
rect 874 418 940 477
rect 874 384 890 418
rect 924 384 940 418
rect 517 373 533 384
rect 467 369 533 373
rect 572 333 643 350
rect 488 317 643 333
rect 488 283 504 317
rect 538 283 572 317
rect 606 283 643 317
rect 488 267 643 283
rect 677 319 943 350
rect 677 285 693 319
rect 727 285 761 319
rect 795 285 829 319
rect 863 285 943 319
rect 677 267 943 285
rect 19 190 71 222
rect 19 156 35 190
rect 69 156 71 190
rect 319 207 750 233
rect 19 140 71 156
rect 105 184 285 188
rect 105 150 121 184
rect 155 172 285 184
rect 155 150 237 172
rect 105 138 237 150
rect 271 138 285 172
rect 105 93 285 138
rect 105 59 237 93
rect 271 59 285 93
rect 105 17 285 59
rect 319 173 335 207
rect 369 203 750 207
rect 369 197 534 203
rect 369 173 385 197
rect 319 101 385 173
rect 524 169 534 197
rect 568 199 706 203
rect 568 169 570 199
rect 319 67 335 101
rect 369 67 385 101
rect 319 51 385 67
rect 424 129 440 163
rect 474 129 490 163
rect 424 89 490 129
rect 424 55 440 89
rect 474 55 490 89
rect 424 17 490 55
rect 524 101 570 169
rect 704 169 706 199
rect 740 169 750 203
rect 524 67 534 101
rect 568 67 570 101
rect 524 51 570 67
rect 604 131 620 165
rect 654 131 670 165
rect 604 89 670 131
rect 604 55 620 89
rect 654 55 670 89
rect 604 17 670 55
rect 704 101 750 169
rect 704 67 706 101
rect 740 67 750 101
rect 704 51 750 67
rect 784 203 842 219
rect 784 169 792 203
rect 826 169 842 203
rect 784 93 842 169
rect 784 59 792 93
rect 826 59 842 93
rect 784 17 842 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor3b_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1163340
string GDS_START 1153986
<< end >>
