magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3602 1975
<< nwell >>
rect -38 331 2342 704
rect 366 323 1011 331
<< pwell >>
rect 363 273 804 281
rect 10 244 804 273
rect 10 204 1057 244
rect 1407 204 2303 241
rect 10 49 2303 204
rect 0 0 2304 49
<< scnmos >>
rect 93 79 123 247
rect 251 119 281 247
rect 337 119 367 247
rect 446 127 476 255
rect 537 127 567 255
rect 691 127 721 255
rect 944 50 974 218
rect 1134 50 1164 178
rect 1220 50 1250 178
rect 1361 50 1391 178
rect 1511 87 1541 215
rect 1619 47 1649 215
rect 1728 87 1758 215
rect 1866 87 1896 215
rect 2016 87 2046 215
rect 2190 47 2220 215
<< scpmoshvt >>
rect 90 367 120 619
rect 217 367 247 567
rect 329 367 359 535
rect 459 359 489 527
rect 545 359 575 527
rect 670 359 700 527
rect 872 359 902 611
rect 1004 380 1034 580
rect 1118 412 1148 580
rect 1310 412 1340 580
rect 1439 367 1469 567
rect 1541 367 1571 619
rect 1788 411 1818 579
rect 1874 411 1904 579
rect 2086 403 2116 603
rect 2193 367 2223 619
<< ndiff >>
rect 389 247 446 255
rect 36 217 93 247
rect 36 183 48 217
rect 82 183 93 217
rect 36 125 93 183
rect 36 91 48 125
rect 82 91 93 125
rect 36 79 93 91
rect 123 136 251 247
rect 123 102 134 136
rect 168 119 251 136
rect 281 202 337 247
rect 281 168 292 202
rect 326 168 337 202
rect 281 119 337 168
rect 367 243 446 247
rect 367 209 401 243
rect 435 209 446 243
rect 367 173 446 209
rect 367 139 401 173
rect 435 139 446 173
rect 367 127 446 139
rect 476 243 537 255
rect 476 209 491 243
rect 525 209 537 243
rect 476 173 537 209
rect 476 139 491 173
rect 525 139 537 173
rect 476 127 537 139
rect 567 217 691 255
rect 567 183 602 217
rect 636 183 691 217
rect 567 127 691 183
rect 721 243 778 255
rect 721 209 732 243
rect 766 209 778 243
rect 721 173 778 209
rect 721 139 732 173
rect 766 139 778 173
rect 721 127 778 139
rect 871 184 944 218
rect 871 150 883 184
rect 917 150 944 184
rect 367 119 417 127
rect 168 102 180 119
rect 123 79 180 102
rect 871 103 944 150
rect 871 69 883 103
rect 917 69 944 103
rect 871 50 944 69
rect 974 184 1031 218
rect 974 150 985 184
rect 1019 178 1031 184
rect 1433 203 1511 215
rect 1433 178 1445 203
rect 1019 150 1134 178
rect 974 96 1134 150
rect 974 62 985 96
rect 1019 62 1134 96
rect 974 50 1134 62
rect 1164 106 1220 178
rect 1164 72 1175 106
rect 1209 72 1220 106
rect 1164 50 1220 72
rect 1250 108 1361 178
rect 1250 74 1277 108
rect 1311 74 1361 108
rect 1250 50 1361 74
rect 1391 169 1445 178
rect 1479 169 1511 203
rect 1391 103 1511 169
rect 1391 69 1445 103
rect 1479 87 1511 103
rect 1541 184 1619 215
rect 1541 150 1573 184
rect 1607 150 1619 184
rect 1541 93 1619 150
rect 1541 87 1573 93
rect 1479 69 1489 87
rect 1391 50 1489 69
rect 1563 59 1573 87
rect 1607 59 1619 93
rect 1563 47 1619 59
rect 1649 193 1728 215
rect 1649 159 1660 193
rect 1694 159 1728 193
rect 1649 103 1728 159
rect 1649 69 1660 103
rect 1694 87 1728 103
rect 1758 163 1866 215
rect 1758 129 1769 163
rect 1803 129 1866 163
rect 1758 87 1866 129
rect 1896 188 2016 215
rect 1896 154 1971 188
rect 2005 154 2016 188
rect 1896 87 2016 154
rect 2046 93 2190 215
rect 2046 87 2122 93
rect 1694 69 1706 87
rect 1649 47 1706 69
rect 2110 59 2122 87
rect 2156 59 2190 93
rect 2110 47 2190 59
rect 2220 203 2277 215
rect 2220 169 2231 203
rect 2265 169 2277 203
rect 2220 103 2277 169
rect 2220 69 2231 103
rect 2265 69 2277 103
rect 2220 47 2277 69
<< pdiff >>
rect 33 597 90 619
rect 33 563 45 597
rect 79 563 90 597
rect 33 519 90 563
rect 33 485 45 519
rect 79 485 90 519
rect 33 442 90 485
rect 33 408 45 442
rect 79 408 90 442
rect 33 367 90 408
rect 120 607 193 619
rect 120 573 147 607
rect 181 573 193 607
rect 120 567 193 573
rect 120 524 217 567
rect 120 490 147 524
rect 181 490 217 524
rect 120 442 217 490
rect 120 408 147 442
rect 181 408 217 442
rect 120 367 217 408
rect 247 555 304 567
rect 247 521 258 555
rect 292 535 304 555
rect 292 521 329 535
rect 247 421 329 521
rect 247 387 258 421
rect 292 387 329 421
rect 247 367 329 387
rect 359 527 409 535
rect 590 543 648 555
rect 590 527 602 543
rect 359 431 459 527
rect 359 397 414 431
rect 448 397 459 431
rect 359 367 459 397
rect 402 359 459 367
rect 489 403 545 527
rect 489 369 500 403
rect 534 369 545 403
rect 489 359 545 369
rect 575 509 602 527
rect 636 527 648 543
rect 636 509 670 527
rect 575 359 670 509
rect 700 515 756 527
rect 700 481 711 515
rect 745 481 756 515
rect 700 405 756 481
rect 700 371 711 405
rect 745 371 756 405
rect 700 359 756 371
rect 816 597 872 611
rect 816 563 827 597
rect 861 563 872 597
rect 816 501 872 563
rect 816 467 827 501
rect 861 467 872 501
rect 816 405 872 467
rect 816 371 827 405
rect 861 371 872 405
rect 816 359 872 371
rect 902 599 975 611
rect 902 565 929 599
rect 963 580 975 599
rect 963 565 1004 580
rect 902 502 1004 565
rect 902 468 929 502
rect 963 468 1004 502
rect 902 405 1004 468
rect 902 371 929 405
rect 963 380 1004 405
rect 1034 568 1118 580
rect 1034 534 1045 568
rect 1079 534 1118 568
rect 1034 497 1118 534
rect 1034 463 1045 497
rect 1079 463 1118 497
rect 1034 426 1118 463
rect 1034 392 1045 426
rect 1079 412 1118 426
rect 1148 568 1310 580
rect 1148 534 1191 568
rect 1225 534 1310 568
rect 1148 458 1310 534
rect 1148 424 1191 458
rect 1225 424 1310 458
rect 1148 412 1310 424
rect 1340 568 1417 580
rect 1340 534 1372 568
rect 1406 567 1417 568
rect 1491 567 1541 619
rect 1406 534 1439 567
rect 1340 490 1439 534
rect 1340 456 1372 490
rect 1406 456 1439 490
rect 1340 413 1439 456
rect 1340 412 1372 413
rect 1079 392 1091 412
rect 1034 380 1091 392
rect 963 371 975 380
rect 902 359 975 371
rect 1362 379 1372 412
rect 1406 379 1439 413
rect 1362 367 1439 379
rect 1469 555 1541 567
rect 1469 521 1480 555
rect 1514 521 1541 555
rect 1469 422 1541 521
rect 1469 388 1480 422
rect 1514 388 1541 422
rect 1469 367 1541 388
rect 1571 597 1628 619
rect 1571 563 1582 597
rect 1616 563 1628 597
rect 1571 505 1628 563
rect 1571 471 1582 505
rect 1616 471 1628 505
rect 1571 413 1628 471
rect 1571 379 1582 413
rect 1616 379 1628 413
rect 1708 613 1766 625
rect 1708 579 1720 613
rect 1754 579 1766 613
rect 2138 603 2193 619
rect 2029 591 2086 603
rect 1708 411 1788 579
rect 1818 457 1874 579
rect 1818 423 1829 457
rect 1863 423 1874 457
rect 1818 411 1874 423
rect 1904 527 1961 579
rect 1904 493 1915 527
rect 1949 493 1961 527
rect 1904 457 1961 493
rect 1904 423 1915 457
rect 1949 423 1961 457
rect 1904 411 1961 423
rect 2029 557 2041 591
rect 2075 557 2086 591
rect 2029 520 2086 557
rect 2029 486 2041 520
rect 2075 486 2086 520
rect 2029 449 2086 486
rect 2029 415 2041 449
rect 2075 415 2086 449
rect 1571 367 1628 379
rect 2029 403 2086 415
rect 2116 591 2193 603
rect 2116 557 2148 591
rect 2182 557 2193 591
rect 2116 507 2193 557
rect 2116 473 2148 507
rect 2182 473 2193 507
rect 2116 403 2193 473
rect 2138 367 2193 403
rect 2223 597 2277 619
rect 2223 563 2234 597
rect 2268 563 2277 597
rect 2223 505 2277 563
rect 2223 471 2234 505
rect 2268 471 2277 505
rect 2223 413 2277 471
rect 2223 379 2234 413
rect 2268 379 2277 413
rect 2223 367 2277 379
<< ndiffc >>
rect 48 183 82 217
rect 48 91 82 125
rect 134 102 168 136
rect 292 168 326 202
rect 401 209 435 243
rect 401 139 435 173
rect 491 209 525 243
rect 491 139 525 173
rect 602 183 636 217
rect 732 209 766 243
rect 732 139 766 173
rect 883 150 917 184
rect 883 69 917 103
rect 985 150 1019 184
rect 985 62 1019 96
rect 1175 72 1209 106
rect 1277 74 1311 108
rect 1445 169 1479 203
rect 1445 69 1479 103
rect 1573 150 1607 184
rect 1573 59 1607 93
rect 1660 159 1694 193
rect 1660 69 1694 103
rect 1769 129 1803 163
rect 1971 154 2005 188
rect 2122 59 2156 93
rect 2231 169 2265 203
rect 2231 69 2265 103
<< pdiffc >>
rect 45 563 79 597
rect 45 485 79 519
rect 45 408 79 442
rect 147 573 181 607
rect 147 490 181 524
rect 147 408 181 442
rect 258 521 292 555
rect 258 387 292 421
rect 414 397 448 431
rect 500 369 534 403
rect 602 509 636 543
rect 711 481 745 515
rect 711 371 745 405
rect 827 563 861 597
rect 827 467 861 501
rect 827 371 861 405
rect 929 565 963 599
rect 929 468 963 502
rect 929 371 963 405
rect 1045 534 1079 568
rect 1045 463 1079 497
rect 1045 392 1079 426
rect 1191 534 1225 568
rect 1191 424 1225 458
rect 1372 534 1406 568
rect 1372 456 1406 490
rect 1372 379 1406 413
rect 1480 521 1514 555
rect 1480 388 1514 422
rect 1582 563 1616 597
rect 1582 471 1616 505
rect 1582 379 1616 413
rect 1720 579 1754 613
rect 1829 423 1863 457
rect 1915 493 1949 527
rect 1915 423 1949 457
rect 2041 557 2075 591
rect 2041 486 2075 520
rect 2041 415 2075 449
rect 2148 557 2182 591
rect 2148 473 2182 507
rect 2234 563 2268 597
rect 2234 471 2268 505
rect 2234 379 2268 413
<< poly >>
rect 90 619 120 645
rect 459 601 801 631
rect 872 611 902 637
rect 1541 619 1571 645
rect 217 567 247 593
rect 329 535 359 561
rect 459 527 489 601
rect 545 527 575 553
rect 90 335 120 367
rect 217 335 247 367
rect 77 319 143 335
rect 77 285 93 319
rect 127 285 143 319
rect 77 269 143 285
rect 185 319 281 335
rect 185 285 201 319
rect 235 285 281 319
rect 185 269 281 285
rect 329 299 359 367
rect 670 527 700 601
rect 459 337 489 359
rect 446 307 489 337
rect 545 307 575 359
rect 670 337 700 359
rect 670 307 721 337
rect 329 269 367 299
rect 93 247 123 269
rect 251 247 281 269
rect 337 247 367 269
rect 446 255 476 307
rect 537 277 575 307
rect 537 255 567 277
rect 691 255 721 307
rect 771 306 801 601
rect 1004 580 1034 606
rect 1118 580 1148 606
rect 1310 580 1340 606
rect 1439 567 1469 593
rect 872 306 902 359
rect 1004 306 1034 380
rect 771 290 1034 306
rect 771 276 960 290
rect 944 256 960 276
rect 994 270 1034 290
rect 1118 348 1148 412
rect 1310 380 1340 412
rect 1253 364 1340 380
rect 1788 579 1818 605
rect 1874 579 1904 605
rect 2086 603 2116 629
rect 2193 619 2223 645
rect 1788 379 1818 411
rect 1118 332 1184 348
rect 1118 298 1134 332
rect 1168 298 1184 332
rect 1118 282 1184 298
rect 1253 330 1280 364
rect 1314 330 1340 364
rect 1253 314 1340 330
rect 994 256 1076 270
rect 944 240 1076 256
rect 944 218 974 240
rect 1046 234 1076 240
rect 251 93 281 119
rect 93 53 123 79
rect 337 53 367 119
rect 446 101 476 127
rect 537 105 567 127
rect 537 89 643 105
rect 691 101 721 127
rect 537 55 593 89
rect 627 55 643 89
rect 537 53 643 55
rect 337 23 643 53
rect 1046 204 1164 234
rect 1253 230 1283 314
rect 1439 303 1469 367
rect 1541 303 1571 367
rect 1698 363 1818 379
rect 1698 329 1714 363
rect 1748 349 1818 363
rect 1874 371 1904 411
rect 2086 381 2116 403
rect 1874 355 1950 371
rect 1748 329 1764 349
rect 1439 287 1649 303
rect 1439 273 1557 287
rect 1134 178 1164 204
rect 1220 200 1283 230
rect 1331 250 1397 266
rect 1331 216 1347 250
rect 1381 216 1397 250
rect 1331 200 1397 216
rect 1511 253 1557 273
rect 1591 253 1649 287
rect 1511 237 1649 253
rect 1698 295 1764 329
rect 1698 261 1714 295
rect 1748 261 1764 295
rect 1874 321 1900 355
rect 1934 321 1950 355
rect 1874 287 1950 321
rect 1874 267 1900 287
rect 1698 245 1764 261
rect 1866 253 1900 267
rect 1934 253 1950 287
rect 1992 351 2116 381
rect 1992 335 2058 351
rect 1992 301 2008 335
rect 2042 301 2058 335
rect 2193 303 2223 367
rect 1992 285 2058 301
rect 2140 287 2223 303
rect 1511 215 1541 237
rect 1619 215 1649 237
rect 1728 215 1758 245
rect 1866 237 1950 253
rect 1866 215 1896 237
rect 2016 215 2046 285
rect 2140 253 2156 287
rect 2190 253 2223 287
rect 2140 237 2223 253
rect 2190 215 2220 237
rect 1220 178 1250 200
rect 1361 178 1391 200
rect 1511 61 1541 87
rect 944 24 974 50
rect 1134 24 1164 50
rect 1220 24 1250 50
rect 1361 24 1391 50
rect 1728 61 1758 87
rect 1866 61 1896 87
rect 2016 61 2046 87
rect 1619 21 1649 47
rect 2190 21 2220 47
<< polycont >>
rect 93 285 127 319
rect 201 285 235 319
rect 960 256 994 290
rect 1134 298 1168 332
rect 1280 330 1314 364
rect 593 55 627 89
rect 1714 329 1748 363
rect 1347 216 1381 250
rect 1557 253 1591 287
rect 1714 261 1748 295
rect 1900 321 1934 355
rect 1900 253 1934 287
rect 2008 301 2042 335
rect 2156 253 2190 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 18 597 95 613
rect 18 563 45 597
rect 79 563 95 597
rect 18 519 95 563
rect 18 485 45 519
rect 79 485 95 519
rect 18 442 95 485
rect 18 408 45 442
rect 79 408 95 442
rect 18 392 95 408
rect 131 607 197 649
rect 131 573 147 607
rect 181 573 197 607
rect 131 524 197 573
rect 131 490 147 524
rect 181 490 197 524
rect 131 442 197 490
rect 131 408 147 442
rect 181 408 197 442
rect 131 392 197 408
rect 242 579 761 613
rect 242 555 308 579
rect 242 521 258 555
rect 292 521 308 555
rect 242 421 308 521
rect 18 233 52 392
rect 242 387 258 421
rect 292 387 308 421
rect 242 371 308 387
rect 88 319 161 356
rect 88 285 93 319
rect 127 285 161 319
rect 88 269 161 285
rect 197 319 238 335
rect 197 285 201 319
rect 235 285 238 319
rect 197 269 238 285
rect 204 233 238 269
rect 18 217 238 233
rect 18 183 48 217
rect 82 199 238 217
rect 82 183 98 199
rect 18 125 98 183
rect 18 91 48 125
rect 82 91 98 125
rect 18 75 98 91
rect 134 136 168 163
rect 134 17 168 102
rect 204 87 238 199
rect 274 247 308 371
rect 344 509 602 543
rect 636 509 652 543
rect 695 515 761 579
rect 344 317 378 509
rect 695 481 711 515
rect 745 481 761 515
rect 414 439 652 473
rect 414 431 448 439
rect 586 424 652 439
rect 414 355 448 397
rect 484 369 500 403
rect 534 369 550 403
rect 484 353 550 369
rect 586 390 607 424
rect 641 390 652 424
rect 344 283 455 317
rect 274 202 342 247
rect 274 168 292 202
rect 326 168 342 202
rect 274 123 342 168
rect 378 243 455 283
rect 378 209 401 243
rect 435 209 455 243
rect 378 202 455 209
rect 378 173 415 202
rect 378 139 401 173
rect 449 168 455 202
rect 435 139 455 168
rect 378 123 455 139
rect 491 243 541 353
rect 525 209 541 243
rect 491 173 541 209
rect 525 139 541 173
rect 586 217 652 390
rect 586 183 602 217
rect 636 183 652 217
rect 586 141 652 183
rect 695 405 761 481
rect 695 371 711 405
rect 745 371 761 405
rect 695 259 761 371
rect 811 597 877 613
rect 811 563 827 597
rect 861 563 877 597
rect 811 501 877 563
rect 811 467 827 501
rect 861 467 877 501
rect 811 405 877 467
rect 811 371 827 405
rect 861 371 877 405
rect 811 355 877 371
rect 913 599 979 649
rect 913 565 929 599
rect 963 565 979 599
rect 913 502 979 565
rect 913 468 929 502
rect 963 468 979 502
rect 913 405 979 468
rect 913 371 929 405
rect 963 371 979 405
rect 1029 568 1095 584
rect 1029 534 1045 568
rect 1079 534 1095 568
rect 1029 497 1095 534
rect 1029 463 1045 497
rect 1079 463 1095 497
rect 1029 426 1095 463
rect 1029 392 1045 426
rect 1079 392 1095 426
rect 1175 568 1241 584
rect 1175 534 1191 568
rect 1225 534 1241 568
rect 1175 458 1241 534
rect 1175 424 1191 458
rect 1225 424 1241 458
rect 1372 568 1422 584
rect 1406 534 1422 568
rect 1372 490 1422 534
rect 1406 456 1422 490
rect 1175 408 1241 424
rect 1029 376 1095 392
rect 913 355 979 371
rect 695 243 782 259
rect 695 209 732 243
rect 766 209 782 243
rect 695 173 782 209
rect 491 87 541 139
rect 695 139 732 173
rect 766 139 782 173
rect 695 123 782 139
rect 819 200 853 355
rect 889 290 1010 306
rect 889 256 960 290
rect 994 256 1010 290
rect 889 236 1010 256
rect 819 184 933 200
rect 819 150 883 184
rect 917 150 933 184
rect 204 53 541 87
rect 577 89 643 105
rect 577 55 593 89
rect 627 87 643 89
rect 819 103 933 150
rect 819 87 883 103
rect 627 69 883 87
rect 917 69 933 103
rect 627 55 933 69
rect 577 53 933 55
rect 969 184 1019 200
rect 969 150 985 184
rect 969 96 1019 150
rect 969 62 985 96
rect 1061 126 1095 376
rect 1131 332 1171 348
rect 1131 298 1134 332
rect 1168 298 1171 332
rect 1131 208 1171 298
rect 1207 278 1241 408
rect 1277 424 1330 430
rect 1277 390 1279 424
rect 1313 390 1330 424
rect 1277 364 1330 390
rect 1277 330 1280 364
rect 1314 330 1330 364
rect 1277 314 1330 330
rect 1372 413 1422 456
rect 1406 379 1422 413
rect 1372 336 1422 379
rect 1464 555 1530 649
rect 1464 521 1480 555
rect 1514 521 1530 555
rect 1464 422 1530 521
rect 1464 388 1480 422
rect 1514 388 1530 422
rect 1464 372 1530 388
rect 1566 597 1632 613
rect 1566 563 1582 597
rect 1616 563 1632 597
rect 1704 579 1720 613
rect 1754 591 2091 613
rect 1754 579 2041 591
rect 1566 543 1632 563
rect 2075 557 2091 591
rect 1566 527 2005 543
rect 1566 509 1915 527
rect 1566 505 1677 509
rect 1566 471 1582 505
rect 1616 471 1677 505
rect 1899 493 1915 509
rect 1949 493 2005 527
rect 1566 413 1677 471
rect 1829 457 1863 473
rect 1566 379 1582 413
rect 1616 379 1677 413
rect 1753 424 1793 430
rect 1753 390 1759 424
rect 1753 379 1793 390
rect 1566 363 1677 379
rect 1372 302 1495 336
rect 1207 244 1295 278
rect 1131 202 1223 208
rect 1131 168 1183 202
rect 1217 168 1223 202
rect 1131 162 1223 168
rect 1261 130 1295 244
rect 1331 250 1409 266
rect 1331 216 1347 250
rect 1381 216 1409 250
rect 1331 202 1409 216
rect 1331 168 1375 202
rect 1331 166 1409 168
rect 1445 203 1495 302
rect 1541 287 1607 303
rect 1541 253 1557 287
rect 1591 253 1607 287
rect 1541 236 1607 253
rect 1479 169 1495 203
rect 1643 209 1677 363
rect 1713 363 1793 379
rect 1713 329 1714 363
rect 1748 345 1793 363
rect 1748 329 1749 345
rect 1713 295 1749 329
rect 1713 261 1714 295
rect 1748 261 1749 295
rect 1829 278 1863 423
rect 1899 457 2005 493
rect 1899 423 1915 457
rect 1949 423 2005 457
rect 1899 407 2005 423
rect 1713 245 1749 261
rect 1785 244 1863 278
rect 1899 355 1935 371
rect 1899 321 1900 355
rect 1934 321 1935 355
rect 1899 287 1935 321
rect 1899 253 1900 287
rect 1934 253 1935 287
rect 1971 351 2005 407
rect 2041 520 2091 557
rect 2075 486 2091 520
rect 2041 449 2091 486
rect 2132 591 2182 649
rect 2132 557 2148 591
rect 2132 507 2182 557
rect 2132 473 2148 507
rect 2132 457 2182 473
rect 2231 597 2284 613
rect 2231 563 2234 597
rect 2268 563 2284 597
rect 2231 505 2284 563
rect 2231 471 2234 505
rect 2268 471 2284 505
rect 2075 421 2091 449
rect 2075 415 2116 421
rect 2041 387 2116 415
rect 1971 335 2046 351
rect 1971 301 2008 335
rect 2042 301 2046 335
rect 1971 285 2046 301
rect 1785 209 1819 244
rect 1061 106 1225 126
rect 1061 92 1175 106
rect 969 17 1019 62
rect 1159 72 1175 92
rect 1209 72 1225 106
rect 1159 53 1225 72
rect 1261 108 1327 130
rect 1261 74 1277 108
rect 1311 74 1327 108
rect 1261 53 1327 74
rect 1445 103 1495 169
rect 1479 69 1495 103
rect 1445 53 1495 69
rect 1557 184 1607 200
rect 1557 150 1573 184
rect 1557 93 1607 150
rect 1557 59 1573 93
rect 1557 17 1607 59
rect 1643 193 1710 209
rect 1643 159 1660 193
rect 1694 159 1710 193
rect 1643 103 1710 159
rect 1643 69 1660 103
rect 1694 69 1710 103
rect 1643 53 1710 69
rect 1753 163 1819 209
rect 1899 208 1935 253
rect 2082 249 2116 387
rect 2231 413 2284 471
rect 2231 379 2234 413
rect 2268 379 2284 413
rect 1753 129 1769 163
rect 1803 129 1819 163
rect 1855 202 1935 208
rect 1889 168 1935 202
rect 1855 162 1935 168
rect 1971 215 2116 249
rect 2152 287 2195 303
rect 2152 253 2156 287
rect 2190 253 2195 287
rect 1971 188 2005 215
rect 1753 87 1819 129
rect 2152 179 2195 253
rect 1971 123 2005 154
rect 2041 145 2195 179
rect 2231 203 2284 379
rect 2265 169 2284 203
rect 2041 87 2075 145
rect 1753 53 2075 87
rect 2122 93 2172 109
rect 2156 59 2172 93
rect 2122 17 2172 59
rect 2231 103 2284 169
rect 2265 69 2284 103
rect 2231 53 2284 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 607 390 641 424
rect 415 173 449 202
rect 415 168 435 173
rect 435 168 449 173
rect 1279 390 1313 424
rect 1759 390 1793 424
rect 1183 168 1217 202
rect 1375 168 1409 202
rect 1855 168 1889 202
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 595 424 653 430
rect 595 390 607 424
rect 641 421 653 424
rect 1267 424 1325 430
rect 1267 421 1279 424
rect 641 393 1279 421
rect 641 390 653 393
rect 595 384 653 390
rect 1267 390 1279 393
rect 1313 421 1325 424
rect 1747 424 1805 430
rect 1747 421 1759 424
rect 1313 393 1759 421
rect 1313 390 1325 393
rect 1267 384 1325 390
rect 1747 390 1759 393
rect 1793 390 1805 424
rect 1747 384 1805 390
rect 403 202 461 208
rect 403 168 415 202
rect 449 199 461 202
rect 1171 202 1229 208
rect 1171 199 1183 202
rect 449 171 1183 199
rect 449 168 461 171
rect 403 162 461 168
rect 1171 168 1183 171
rect 1217 199 1229 202
rect 1363 202 1421 208
rect 1363 199 1375 202
rect 1217 171 1375 199
rect 1217 168 1229 171
rect 1171 162 1229 168
rect 1363 168 1375 171
rect 1409 199 1421 202
rect 1843 202 1901 208
rect 1843 199 1855 202
rect 1409 171 1855 199
rect 1409 168 1421 171
rect 1363 162 1421 168
rect 1843 168 1855 171
rect 1889 168 1901 202
rect 1843 162 1901 168
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
flabel pwell s 0 0 2304 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2304 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fahcon_1
flabel metal1 s 0 617 2304 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2304 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 2239 94 2273 128 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2239 168 2273 202 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2239 242 2273 276 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2239 316 2273 350 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2239 390 2273 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2239 464 2273 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2239 538 2273 572 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1279 94 1313 128 0 FreeSans 340 0 0 0 COUT_N
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 CI
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2304 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6936476
string GDS_START 6918530
<< end >>
