magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 2 49 864 248
rect 0 0 960 49
<< scnmos >>
rect 81 138 111 222
rect 179 74 209 222
rect 369 138 399 222
rect 467 74 497 222
rect 657 138 687 222
rect 755 74 785 222
<< scpmoshvt >>
rect 83 368 113 452
rect 186 368 216 592
rect 380 368 410 452
rect 483 368 513 592
rect 677 368 707 452
rect 781 368 811 592
<< ndiff >>
rect 28 190 81 222
rect 28 156 36 190
rect 70 156 81 190
rect 28 138 81 156
rect 111 161 179 222
rect 111 138 134 161
rect 126 127 134 138
rect 168 127 179 161
rect 126 74 179 127
rect 209 199 262 222
rect 209 165 220 199
rect 254 165 262 199
rect 209 131 262 165
rect 316 190 369 222
rect 316 156 324 190
rect 358 156 369 190
rect 316 138 369 156
rect 399 161 467 222
rect 399 138 422 161
rect 209 97 220 131
rect 254 97 262 131
rect 414 127 422 138
rect 456 127 467 161
rect 209 74 262 97
rect 414 74 467 127
rect 497 199 550 222
rect 497 165 508 199
rect 542 165 550 199
rect 497 131 550 165
rect 604 190 657 222
rect 604 156 612 190
rect 646 156 657 190
rect 604 138 657 156
rect 687 161 755 222
rect 687 138 710 161
rect 497 97 508 131
rect 542 97 550 131
rect 702 127 710 138
rect 744 127 755 161
rect 497 74 550 97
rect 702 74 755 127
rect 785 199 838 222
rect 785 165 796 199
rect 830 165 838 199
rect 785 131 838 165
rect 785 97 796 131
rect 830 97 838 131
rect 785 74 838 97
<< pdiff >>
rect 131 580 186 592
rect 131 546 139 580
rect 173 546 186 580
rect 131 512 186 546
rect 131 478 139 512
rect 173 478 186 512
rect 131 452 186 478
rect 28 429 83 452
rect 28 395 36 429
rect 70 395 83 429
rect 28 368 83 395
rect 113 368 186 452
rect 216 580 271 592
rect 216 546 229 580
rect 263 546 271 580
rect 216 511 271 546
rect 216 477 229 511
rect 263 477 271 511
rect 428 580 483 592
rect 428 546 436 580
rect 470 546 483 580
rect 428 512 483 546
rect 428 478 436 512
rect 470 478 483 512
rect 216 417 271 477
rect 428 452 483 478
rect 216 383 229 417
rect 263 383 271 417
rect 216 368 271 383
rect 325 429 380 452
rect 325 395 333 429
rect 367 395 380 429
rect 325 368 380 395
rect 410 368 483 452
rect 513 580 568 592
rect 513 546 526 580
rect 560 546 568 580
rect 513 511 568 546
rect 513 477 526 511
rect 560 477 568 511
rect 725 580 781 592
rect 725 546 733 580
rect 767 546 781 580
rect 725 512 781 546
rect 725 478 733 512
rect 767 478 781 512
rect 513 417 568 477
rect 725 452 781 478
rect 513 383 526 417
rect 560 383 568 417
rect 513 368 568 383
rect 622 429 677 452
rect 622 395 630 429
rect 664 395 677 429
rect 622 368 677 395
rect 707 368 781 452
rect 811 580 866 592
rect 811 546 824 580
rect 858 546 866 580
rect 811 511 866 546
rect 811 477 824 511
rect 858 477 866 511
rect 811 417 866 477
rect 811 383 824 417
rect 858 383 866 417
rect 811 368 866 383
<< ndiffc >>
rect 36 156 70 190
rect 134 127 168 161
rect 220 165 254 199
rect 324 156 358 190
rect 220 97 254 131
rect 422 127 456 161
rect 508 165 542 199
rect 612 156 646 190
rect 508 97 542 131
rect 710 127 744 161
rect 796 165 830 199
rect 796 97 830 131
<< pdiffc >>
rect 139 546 173 580
rect 139 478 173 512
rect 36 395 70 429
rect 229 546 263 580
rect 229 477 263 511
rect 436 546 470 580
rect 436 478 470 512
rect 229 383 263 417
rect 333 395 367 429
rect 526 546 560 580
rect 526 477 560 511
rect 733 546 767 580
rect 733 478 767 512
rect 526 383 560 417
rect 630 395 664 429
rect 824 546 858 580
rect 824 477 858 511
rect 824 383 858 417
<< poly >>
rect 186 592 216 618
rect 483 592 513 618
rect 781 592 811 618
rect 83 452 113 478
rect 380 452 410 478
rect 677 452 707 478
rect 83 353 113 368
rect 186 353 216 368
rect 380 353 410 368
rect 483 353 513 368
rect 677 353 707 368
rect 781 353 811 368
rect 80 321 116 353
rect 183 321 219 353
rect 377 321 413 353
rect 480 321 516 353
rect 674 321 710 353
rect 778 321 814 353
rect 45 305 116 321
rect 45 271 61 305
rect 95 271 116 305
rect 45 255 116 271
rect 158 305 224 321
rect 158 271 174 305
rect 208 271 224 305
rect 81 222 111 255
rect 158 252 224 271
rect 333 305 413 321
rect 333 271 349 305
rect 383 271 413 305
rect 333 255 413 271
rect 455 305 521 321
rect 455 271 471 305
rect 505 271 521 305
rect 179 222 209 252
rect 369 222 399 255
rect 455 252 521 271
rect 621 305 710 321
rect 621 271 637 305
rect 671 271 710 305
rect 621 255 710 271
rect 752 305 818 321
rect 752 271 768 305
rect 802 271 818 305
rect 467 222 497 252
rect 657 222 687 255
rect 752 252 818 271
rect 755 222 785 252
rect 81 112 111 138
rect 369 112 399 138
rect 657 112 687 138
rect 179 48 209 74
rect 467 48 497 74
rect 755 48 785 74
<< polycont >>
rect 61 271 95 305
rect 174 271 208 305
rect 349 271 383 305
rect 471 271 505 305
rect 637 271 671 305
rect 768 271 802 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 118 580 177 649
rect 118 546 139 580
rect 173 546 177 580
rect 118 512 177 546
rect 118 478 139 512
rect 173 478 177 512
rect 118 462 177 478
rect 213 580 276 615
rect 213 546 229 580
rect 263 546 276 580
rect 213 511 276 546
rect 213 477 229 511
rect 263 477 276 511
rect 20 429 86 445
rect 20 395 36 429
rect 70 428 86 429
rect 70 395 179 428
rect 20 387 179 395
rect 21 305 111 353
rect 21 271 61 305
rect 95 271 111 305
rect 145 321 179 387
rect 213 424 276 477
rect 420 580 479 649
rect 420 546 436 580
rect 470 546 479 580
rect 420 512 479 546
rect 420 478 436 512
rect 470 478 479 512
rect 420 462 479 478
rect 513 580 573 615
rect 513 546 526 580
rect 560 546 573 580
rect 513 511 573 546
rect 513 477 526 511
rect 560 477 573 511
rect 213 390 223 424
rect 257 417 276 424
rect 213 383 229 390
rect 263 383 276 417
rect 213 367 276 383
rect 310 429 374 445
rect 513 432 573 477
rect 717 580 776 649
rect 717 546 733 580
rect 767 546 776 580
rect 717 512 776 546
rect 717 478 733 512
rect 767 478 776 512
rect 717 462 776 478
rect 810 580 870 615
rect 810 546 824 580
rect 858 546 870 580
rect 810 511 870 546
rect 810 477 824 511
rect 858 477 870 511
rect 310 395 333 429
rect 367 428 374 429
rect 367 395 467 428
rect 310 379 467 395
rect 242 321 276 367
rect 433 321 467 379
rect 501 424 573 432
rect 501 390 511 424
rect 545 417 573 424
rect 501 383 526 390
rect 560 383 573 417
rect 501 367 573 383
rect 614 429 680 445
rect 810 432 870 477
rect 614 395 630 429
rect 664 428 680 429
rect 664 395 761 428
rect 614 379 761 395
rect 539 321 573 367
rect 721 321 761 379
rect 795 424 870 432
rect 795 390 799 424
rect 833 417 870 424
rect 795 383 824 390
rect 858 383 870 417
rect 795 367 870 383
rect 145 305 208 321
rect 145 271 174 305
rect 145 255 208 271
rect 242 305 399 321
rect 242 271 349 305
rect 383 271 399 305
rect 242 263 399 271
rect 433 305 505 321
rect 433 271 471 305
rect 145 229 179 255
rect 20 195 179 229
rect 242 215 276 263
rect 433 255 505 271
rect 539 305 687 321
rect 539 271 637 305
rect 671 271 687 305
rect 539 263 687 271
rect 721 305 802 321
rect 721 271 768 305
rect 433 229 467 255
rect 218 199 276 215
rect 20 190 79 195
rect 20 156 36 190
rect 70 156 79 190
rect 218 165 220 199
rect 254 165 276 199
rect 20 140 79 156
rect 118 127 134 161
rect 168 127 184 161
rect 118 17 184 127
rect 218 131 276 165
rect 310 195 467 229
rect 539 215 573 263
rect 721 255 802 271
rect 721 229 755 255
rect 506 199 573 215
rect 310 190 367 195
rect 310 156 324 190
rect 358 156 367 190
rect 506 165 508 199
rect 542 165 573 199
rect 310 140 367 156
rect 218 97 220 131
rect 254 97 276 131
rect 218 51 276 97
rect 406 127 422 161
rect 456 127 472 161
rect 406 17 472 127
rect 506 131 573 165
rect 612 195 755 229
rect 836 215 870 367
rect 794 199 870 215
rect 612 190 655 195
rect 646 156 655 190
rect 794 165 796 199
rect 830 165 870 199
rect 612 140 655 156
rect 506 97 508 131
rect 542 97 573 131
rect 506 51 573 97
rect 694 127 710 161
rect 744 127 760 161
rect 694 17 760 127
rect 794 131 870 165
rect 794 97 796 131
rect 830 97 870 131
rect 794 51 870 97
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 223 417 257 424
rect 223 390 229 417
rect 229 390 257 417
rect 511 417 545 424
rect 511 390 526 417
rect 526 390 545 417
rect 799 417 833 424
rect 799 390 824 417
rect 824 390 833 417
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 193 464 845 498
rect 193 424 269 430
rect 193 390 223 424
rect 257 390 269 424
rect 193 384 269 390
rect 481 424 557 430
rect 481 390 511 424
rect 545 390 557 424
rect 481 384 557 390
rect 769 424 845 464
rect 769 390 799 424
rect 833 390 845 424
rect 769 384 845 390
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlymetal6s6s_1
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 193 464 842 498 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel locali s 32 316 66 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 2447422
string GDS_START 2439326
<< end >>
