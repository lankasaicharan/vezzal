magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 1 49 863 248
rect 0 0 864 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 263 368 299 592
rect 353 368 389 592
rect 443 368 479 592
rect 533 368 569 592
rect 633 368 669 592
rect 733 368 769 592
<< nmoslvt >>
rect 89 74 119 222
rect 347 74 377 222
rect 443 74 473 222
rect 533 74 563 222
<< ndiff >>
rect 27 188 89 222
rect 27 154 44 188
rect 78 154 89 188
rect 27 120 89 154
rect 27 86 44 120
rect 78 86 89 120
rect 27 74 89 86
rect 119 186 347 222
rect 119 152 130 186
rect 164 152 213 186
rect 247 152 302 186
rect 336 152 347 186
rect 119 118 347 152
rect 119 84 130 118
rect 164 84 213 118
rect 247 84 302 118
rect 336 84 347 118
rect 119 74 347 84
rect 377 127 443 222
rect 377 93 388 127
rect 422 93 443 127
rect 377 74 443 93
rect 473 210 533 222
rect 473 176 488 210
rect 522 176 533 210
rect 473 120 533 176
rect 473 86 488 120
rect 522 86 533 120
rect 473 74 533 86
rect 563 186 837 222
rect 563 152 574 186
rect 608 152 689 186
rect 723 152 791 186
rect 825 152 837 186
rect 563 118 837 152
rect 563 84 574 118
rect 608 84 689 118
rect 723 84 791 118
rect 825 84 837 118
rect 563 74 837 84
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 462 173 546
rect 119 428 129 462
rect 163 428 173 462
rect 119 368 173 428
rect 209 580 263 592
rect 209 546 219 580
rect 253 546 263 580
rect 209 497 263 546
rect 209 463 219 497
rect 253 463 263 497
rect 209 414 263 463
rect 209 380 219 414
rect 253 380 263 414
rect 209 368 263 380
rect 299 580 353 592
rect 299 546 309 580
rect 343 546 353 580
rect 299 462 353 546
rect 299 428 309 462
rect 343 428 353 462
rect 299 368 353 428
rect 389 580 443 592
rect 389 546 399 580
rect 433 546 443 580
rect 389 497 443 546
rect 389 463 399 497
rect 433 463 443 497
rect 389 414 443 463
rect 389 380 399 414
rect 433 380 443 414
rect 389 368 443 380
rect 479 547 533 592
rect 479 513 489 547
rect 523 513 533 547
rect 479 479 533 513
rect 479 445 489 479
rect 523 445 533 479
rect 479 411 533 445
rect 479 377 489 411
rect 523 377 533 411
rect 479 368 533 377
rect 569 582 633 592
rect 569 548 589 582
rect 623 548 633 582
rect 569 514 633 548
rect 569 480 589 514
rect 623 480 633 514
rect 569 446 633 480
rect 569 412 589 446
rect 623 412 633 446
rect 569 368 633 412
rect 669 547 733 592
rect 669 513 689 547
rect 723 513 733 547
rect 669 479 733 513
rect 669 445 689 479
rect 723 445 733 479
rect 669 411 733 445
rect 669 377 689 411
rect 723 377 733 411
rect 669 368 733 377
rect 769 580 837 592
rect 769 546 779 580
rect 813 546 837 580
rect 769 497 837 546
rect 769 463 779 497
rect 813 463 837 497
rect 769 414 837 463
rect 769 380 779 414
rect 813 380 837 414
rect 769 368 837 380
<< ndiffc >>
rect 44 154 78 188
rect 44 86 78 120
rect 130 152 164 186
rect 213 152 247 186
rect 302 152 336 186
rect 130 84 164 118
rect 213 84 247 118
rect 302 84 336 118
rect 388 93 422 127
rect 488 176 522 210
rect 488 86 522 120
rect 574 152 608 186
rect 689 152 723 186
rect 791 152 825 186
rect 574 84 608 118
rect 689 84 723 118
rect 791 84 825 118
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 428 163 462
rect 219 546 253 580
rect 219 463 253 497
rect 219 380 253 414
rect 309 546 343 580
rect 309 428 343 462
rect 399 546 433 580
rect 399 463 433 497
rect 399 380 433 414
rect 489 513 523 547
rect 489 445 523 479
rect 489 377 523 411
rect 589 548 623 582
rect 589 480 623 514
rect 589 412 623 446
rect 689 513 723 547
rect 689 445 723 479
rect 689 377 723 411
rect 779 546 813 580
rect 779 463 813 497
rect 779 380 813 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 263 592 299 618
rect 353 592 389 618
rect 443 592 479 618
rect 533 592 569 618
rect 633 592 669 618
rect 733 592 769 618
rect 83 310 119 368
rect 173 310 209 368
rect 263 310 299 368
rect 353 310 389 368
rect 83 294 389 310
rect 83 260 105 294
rect 139 260 173 294
rect 207 260 241 294
rect 275 260 309 294
rect 343 280 389 294
rect 443 310 479 368
rect 533 310 569 368
rect 633 310 669 368
rect 733 310 769 368
rect 443 294 835 310
rect 343 260 377 280
rect 83 244 377 260
rect 89 222 119 244
rect 347 222 377 244
rect 443 260 649 294
rect 683 260 717 294
rect 751 260 785 294
rect 819 260 835 294
rect 443 244 835 260
rect 443 222 473 244
rect 533 222 563 244
rect 89 48 119 74
rect 347 48 377 74
rect 443 48 473 74
rect 533 48 563 74
<< polycont >>
rect 105 260 139 294
rect 173 260 207 294
rect 241 260 275 294
rect 309 260 343 294
rect 649 260 683 294
rect 717 260 751 294
rect 785 260 819 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 497 89 546
rect 23 463 39 497
rect 73 463 89 497
rect 23 414 89 463
rect 23 380 39 414
rect 73 380 89 414
rect 129 580 163 649
rect 129 462 163 546
rect 129 412 163 428
rect 203 580 269 596
rect 203 546 219 580
rect 253 546 269 580
rect 203 497 269 546
rect 203 463 219 497
rect 253 463 269 497
rect 203 414 269 463
rect 23 378 89 380
rect 203 380 219 414
rect 253 380 269 414
rect 309 580 343 649
rect 309 462 343 546
rect 309 412 343 428
rect 383 582 829 615
rect 383 581 589 582
rect 383 580 439 581
rect 383 546 399 580
rect 433 546 439 580
rect 573 548 589 581
rect 623 581 829 582
rect 623 548 639 581
rect 383 497 439 546
rect 383 463 399 497
rect 433 463 439 497
rect 383 414 439 463
rect 203 378 269 380
rect 383 380 399 414
rect 433 380 439 414
rect 383 378 439 380
rect 23 344 439 378
rect 473 513 489 547
rect 523 513 539 547
rect 473 479 539 513
rect 473 445 489 479
rect 523 445 539 479
rect 473 411 539 445
rect 573 514 639 548
rect 773 580 829 581
rect 573 480 589 514
rect 623 480 639 514
rect 573 446 639 480
rect 573 412 589 446
rect 623 412 639 446
rect 673 513 689 547
rect 723 513 739 547
rect 673 479 739 513
rect 673 445 689 479
rect 723 445 739 479
rect 473 377 489 411
rect 523 378 539 411
rect 673 411 739 445
rect 673 378 689 411
rect 523 377 689 378
rect 723 377 739 411
rect 473 344 739 377
rect 773 546 779 580
rect 813 546 829 580
rect 773 497 829 546
rect 773 463 779 497
rect 813 463 829 497
rect 773 414 829 463
rect 773 380 779 414
rect 813 380 829 414
rect 773 364 829 380
rect 25 294 359 310
rect 25 260 105 294
rect 139 260 173 294
rect 207 260 241 294
rect 275 260 309 294
rect 343 260 359 294
rect 25 236 359 260
rect 473 282 539 344
rect 601 294 839 310
rect 473 236 551 282
rect 601 260 649 294
rect 683 260 717 294
rect 751 260 785 294
rect 819 260 839 294
rect 601 236 839 260
rect 473 226 538 236
rect 472 210 538 226
rect 472 202 488 210
rect 23 188 94 202
rect 23 154 44 188
rect 78 154 94 188
rect 23 120 94 154
rect 23 86 44 120
rect 78 86 94 120
rect 23 17 94 86
rect 128 186 488 202
rect 128 152 130 186
rect 164 152 213 186
rect 247 152 302 186
rect 336 176 488 186
rect 522 176 538 210
rect 336 168 538 176
rect 336 152 338 168
rect 128 118 338 152
rect 128 84 130 118
rect 164 84 213 118
rect 247 84 302 118
rect 336 84 338 118
rect 128 68 338 84
rect 372 127 438 134
rect 372 93 388 127
rect 422 93 438 127
rect 372 17 438 93
rect 472 120 538 168
rect 472 86 488 120
rect 522 86 538 120
rect 472 70 538 86
rect 572 186 841 202
rect 572 152 574 186
rect 608 152 689 186
rect 723 152 791 186
rect 825 152 841 186
rect 572 118 841 152
rect 572 84 574 118
rect 608 84 689 118
rect 723 84 791 118
rect 825 84 841 118
rect 572 17 841 84
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor2_4
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 3203868
string GDS_START 3195968
<< end >>
