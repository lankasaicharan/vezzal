magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 1 170 261 287
rect 1 49 634 170
rect 0 0 672 49
<< scnmos >>
rect 80 177 110 261
rect 152 177 182 261
rect 353 60 383 144
rect 439 60 469 144
rect 525 60 555 144
<< scpmoshvt >>
rect 113 487 143 615
rect 199 487 229 615
rect 353 487 383 615
rect 425 487 455 615
rect 515 487 545 615
<< ndiff >>
rect 27 236 80 261
rect 27 202 35 236
rect 69 202 80 236
rect 27 177 80 202
rect 110 177 152 261
rect 182 236 235 261
rect 182 202 193 236
rect 227 202 235 236
rect 182 177 235 202
rect 300 119 353 144
rect 300 85 308 119
rect 342 85 353 119
rect 300 60 353 85
rect 383 119 439 144
rect 383 85 394 119
rect 428 85 439 119
rect 383 60 439 85
rect 469 119 525 144
rect 469 85 480 119
rect 514 85 525 119
rect 469 60 525 85
rect 555 119 608 144
rect 555 85 566 119
rect 600 85 608 119
rect 555 60 608 85
<< pdiff >>
rect 60 603 113 615
rect 60 569 68 603
rect 102 569 113 603
rect 60 533 113 569
rect 60 499 68 533
rect 102 499 113 533
rect 60 487 113 499
rect 143 597 199 615
rect 143 563 154 597
rect 188 563 199 597
rect 143 529 199 563
rect 143 495 154 529
rect 188 495 199 529
rect 143 487 199 495
rect 229 571 353 615
rect 229 537 240 571
rect 274 537 308 571
rect 342 537 353 571
rect 229 487 353 537
rect 383 487 425 615
rect 455 601 515 615
rect 455 567 470 601
rect 504 567 515 601
rect 455 533 515 567
rect 455 499 470 533
rect 504 499 515 533
rect 455 487 515 499
rect 545 599 598 615
rect 545 565 556 599
rect 590 565 598 599
rect 545 487 598 565
<< ndiffc >>
rect 35 202 69 236
rect 193 202 227 236
rect 308 85 342 119
rect 394 85 428 119
rect 480 85 514 119
rect 566 85 600 119
<< pdiffc >>
rect 68 569 102 603
rect 68 499 102 533
rect 154 563 188 597
rect 154 495 188 529
rect 240 537 274 571
rect 308 537 342 571
rect 470 567 504 601
rect 470 499 504 533
rect 556 565 590 599
<< poly >>
rect 113 615 143 641
rect 199 615 229 641
rect 353 615 383 641
rect 425 615 455 641
rect 515 615 545 641
rect 113 449 143 487
rect 44 433 143 449
rect 44 399 60 433
rect 94 419 143 433
rect 199 419 229 487
rect 94 399 110 419
rect 44 365 110 399
rect 44 331 60 365
rect 94 331 110 365
rect 44 315 110 331
rect 199 403 311 419
rect 199 369 261 403
rect 295 369 311 403
rect 199 335 311 369
rect 199 315 261 335
rect 80 261 110 315
rect 152 301 261 315
rect 295 301 311 335
rect 152 285 311 301
rect 152 261 182 285
rect 353 196 383 487
rect 425 378 455 487
rect 515 456 545 487
rect 515 431 600 456
rect 515 426 550 431
rect 534 397 550 426
rect 584 397 600 431
rect 425 362 491 378
rect 425 328 441 362
rect 475 328 491 362
rect 425 294 491 328
rect 425 260 441 294
rect 475 260 491 294
rect 425 244 491 260
rect 534 363 600 397
rect 534 329 550 363
rect 584 329 600 363
rect 80 151 110 177
rect 152 151 182 177
rect 250 166 383 196
rect 250 103 280 166
rect 353 144 383 166
rect 439 144 469 244
rect 534 196 600 329
rect 525 166 600 196
rect 525 144 555 166
rect 202 87 280 103
rect 202 53 218 87
rect 252 53 280 87
rect 202 37 280 53
rect 353 34 383 60
rect 439 34 469 60
rect 525 34 555 60
<< polycont >>
rect 60 399 94 433
rect 60 331 94 365
rect 261 369 295 403
rect 261 301 295 335
rect 550 397 584 431
rect 441 328 475 362
rect 441 260 475 294
rect 550 329 584 363
rect 218 53 252 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 52 603 114 649
rect 52 569 68 603
rect 102 569 114 603
rect 52 533 114 569
rect 52 499 68 533
rect 102 499 114 533
rect 52 483 114 499
rect 148 597 198 613
rect 148 563 154 597
rect 188 563 198 597
rect 148 529 198 563
rect 148 495 154 529
rect 188 495 198 529
rect 232 571 358 649
rect 232 537 240 571
rect 274 537 308 571
rect 342 537 358 571
rect 232 521 358 537
rect 454 601 520 605
rect 454 567 470 601
rect 504 567 520 601
rect 454 533 520 567
rect 554 599 612 649
rect 554 565 556 599
rect 590 565 612 599
rect 554 549 612 565
rect 148 487 198 495
rect 454 499 470 533
rect 504 515 520 533
rect 504 499 654 515
rect 148 453 420 487
rect 454 481 654 499
rect 17 433 114 449
rect 17 399 60 433
rect 94 419 114 433
rect 94 399 143 419
rect 17 365 143 399
rect 17 331 60 365
rect 94 331 143 365
rect 17 286 143 331
rect 19 236 75 252
rect 19 202 35 236
rect 69 202 75 236
rect 19 17 75 202
rect 109 103 143 286
rect 177 252 225 453
rect 386 447 420 453
rect 386 431 586 447
rect 261 403 314 419
rect 386 413 550 431
rect 295 379 314 403
rect 534 397 550 413
rect 584 397 586 431
rect 295 369 491 379
rect 261 362 491 369
rect 261 335 441 362
rect 295 328 441 335
rect 475 328 491 362
rect 295 301 491 328
rect 534 363 586 397
rect 534 329 550 363
rect 584 329 586 363
rect 534 313 586 329
rect 261 294 491 301
rect 261 285 441 294
rect 319 260 441 285
rect 475 260 491 294
rect 620 276 654 481
rect 177 236 243 252
rect 319 244 491 260
rect 177 202 193 236
rect 227 202 243 236
rect 177 186 243 202
rect 302 169 516 207
rect 302 119 351 169
rect 109 87 268 103
rect 109 53 218 87
rect 252 53 268 87
rect 302 85 308 119
rect 342 85 351 119
rect 302 69 351 85
rect 385 119 436 135
rect 385 85 394 119
rect 428 85 436 119
rect 109 51 268 53
rect 385 17 436 85
rect 470 119 516 169
rect 470 85 480 119
rect 514 85 516 119
rect 470 69 516 85
rect 550 119 654 276
rect 550 85 566 119
rect 600 85 654 119
rect 550 69 654 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xnor2_0
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4359994
string GDS_START 4353578
<< end >>
