magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 2 49 763 241
rect 0 0 768 49
<< scnmos >>
rect 81 131 111 215
rect 186 47 216 215
rect 272 47 302 215
rect 462 47 492 215
rect 548 47 578 215
rect 650 47 680 215
<< scpmoshvt >>
rect 114 367 144 451
rect 243 367 273 619
rect 329 367 359 619
rect 446 367 476 619
rect 534 367 564 619
rect 649 367 679 619
<< ndiff >>
rect 28 190 81 215
rect 28 156 36 190
rect 70 156 81 190
rect 28 131 81 156
rect 111 192 186 215
rect 111 158 122 192
rect 156 158 186 192
rect 111 131 186 158
rect 133 93 186 131
rect 133 59 141 93
rect 175 59 186 93
rect 133 47 186 59
rect 216 203 272 215
rect 216 169 227 203
rect 261 169 272 203
rect 216 101 272 169
rect 216 67 227 101
rect 261 67 272 101
rect 216 47 272 67
rect 302 167 355 215
rect 302 133 313 167
rect 347 133 355 167
rect 302 93 355 133
rect 302 59 313 93
rect 347 59 355 93
rect 302 47 355 59
rect 409 203 462 215
rect 409 169 417 203
rect 451 169 462 203
rect 409 101 462 169
rect 409 67 417 101
rect 451 67 462 101
rect 409 47 462 67
rect 492 167 548 215
rect 492 133 503 167
rect 537 133 548 167
rect 492 91 548 133
rect 492 57 503 91
rect 537 57 548 91
rect 492 47 548 57
rect 578 93 650 215
rect 578 59 603 93
rect 637 59 650 93
rect 578 47 650 59
rect 680 203 737 215
rect 680 169 691 203
rect 725 169 737 203
rect 680 101 737 169
rect 680 67 691 101
rect 725 67 737 101
rect 680 47 737 67
<< pdiff >>
rect 190 568 243 619
rect 190 534 198 568
rect 232 534 243 568
rect 190 451 243 534
rect 61 434 114 451
rect 61 400 69 434
rect 103 400 114 434
rect 61 367 114 400
rect 144 367 243 451
rect 273 420 329 619
rect 273 386 284 420
rect 318 386 329 420
rect 273 367 329 386
rect 359 568 446 619
rect 359 534 384 568
rect 418 534 446 568
rect 359 367 446 534
rect 476 599 534 619
rect 476 565 487 599
rect 521 565 534 599
rect 476 506 534 565
rect 476 472 487 506
rect 521 472 534 506
rect 476 421 534 472
rect 476 387 487 421
rect 521 387 534 421
rect 476 367 534 387
rect 564 367 649 619
rect 679 607 732 619
rect 679 573 690 607
rect 724 573 732 607
rect 679 521 732 573
rect 679 487 690 521
rect 724 487 732 521
rect 679 434 732 487
rect 679 400 690 434
rect 724 400 732 434
rect 679 367 732 400
<< ndiffc >>
rect 36 156 70 190
rect 122 158 156 192
rect 141 59 175 93
rect 227 169 261 203
rect 227 67 261 101
rect 313 133 347 167
rect 313 59 347 93
rect 417 169 451 203
rect 417 67 451 101
rect 503 133 537 167
rect 503 57 537 91
rect 603 59 637 93
rect 691 169 725 203
rect 691 67 725 101
<< pdiffc >>
rect 198 534 232 568
rect 69 400 103 434
rect 284 386 318 420
rect 384 534 418 568
rect 487 565 521 599
rect 487 472 521 506
rect 487 387 521 421
rect 690 573 724 607
rect 690 487 724 521
rect 690 400 724 434
<< poly >>
rect 243 619 273 645
rect 329 619 359 645
rect 446 619 476 645
rect 534 619 564 645
rect 649 619 679 645
rect 114 451 144 477
rect 114 308 144 367
rect 243 345 273 367
rect 329 345 359 367
rect 78 292 144 308
rect 78 258 94 292
rect 128 258 144 292
rect 78 242 144 258
rect 186 287 359 345
rect 446 335 476 367
rect 186 253 309 287
rect 343 253 359 287
rect 401 319 476 335
rect 401 285 417 319
rect 451 299 476 319
rect 534 308 564 367
rect 649 308 679 367
rect 451 285 492 299
rect 401 269 492 285
rect 81 215 111 242
rect 186 237 359 253
rect 186 215 216 237
rect 272 215 302 237
rect 462 215 492 269
rect 534 292 607 308
rect 534 258 557 292
rect 591 258 607 292
rect 534 242 607 258
rect 649 292 727 308
rect 649 258 677 292
rect 711 258 727 292
rect 649 242 727 258
rect 548 215 578 242
rect 650 215 680 242
rect 81 105 111 131
rect 186 21 216 47
rect 272 21 302 47
rect 462 21 492 47
rect 548 21 578 47
rect 650 21 680 47
<< polycont >>
rect 94 258 128 292
rect 309 253 343 287
rect 417 285 451 319
rect 557 258 591 292
rect 677 258 711 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 182 568 248 649
rect 182 534 198 568
rect 232 534 248 568
rect 182 526 248 534
rect 368 568 434 649
rect 368 534 384 568
rect 418 534 434 568
rect 368 526 434 534
rect 481 599 523 615
rect 481 565 487 599
rect 521 565 523 599
rect 481 506 523 565
rect 677 607 740 649
rect 677 573 690 607
rect 724 573 740 607
rect 677 521 740 573
rect 17 458 447 492
rect 17 434 119 458
rect 17 400 69 434
rect 103 400 119 434
rect 17 384 119 400
rect 213 420 334 424
rect 213 386 284 420
rect 318 386 334 420
rect 17 206 54 384
rect 213 370 334 386
rect 88 292 179 350
rect 88 258 94 292
rect 128 258 179 292
rect 88 242 179 258
rect 17 190 72 206
rect 17 156 36 190
rect 70 156 72 190
rect 17 140 72 156
rect 106 192 179 208
rect 106 158 122 192
rect 156 158 179 192
rect 106 93 179 158
rect 106 59 141 93
rect 175 59 179 93
rect 106 17 179 59
rect 213 203 263 370
rect 401 335 447 458
rect 481 472 487 506
rect 521 472 523 506
rect 481 421 523 472
rect 481 387 487 421
rect 521 387 523 421
rect 481 371 523 387
rect 401 319 453 335
rect 213 169 227 203
rect 261 169 263 203
rect 297 287 359 303
rect 297 253 309 287
rect 343 253 359 287
rect 401 285 417 319
rect 451 285 453 319
rect 401 269 453 285
rect 297 235 359 253
rect 487 235 523 371
rect 557 292 643 521
rect 677 487 690 521
rect 724 487 740 521
rect 677 434 740 487
rect 677 400 690 434
rect 724 400 740 434
rect 677 384 740 400
rect 591 258 643 292
rect 557 242 643 258
rect 677 292 751 350
rect 711 258 751 292
rect 677 242 751 258
rect 297 203 523 235
rect 297 201 417 203
rect 213 101 263 169
rect 401 169 417 201
rect 451 201 523 203
rect 675 203 741 208
rect 451 169 453 201
rect 213 67 227 101
rect 261 67 263 101
rect 213 51 263 67
rect 297 133 313 167
rect 347 133 363 167
rect 297 93 363 133
rect 297 59 313 93
rect 347 59 363 93
rect 297 17 363 59
rect 401 101 453 169
rect 675 169 691 203
rect 725 169 741 203
rect 675 167 741 169
rect 401 67 417 101
rect 451 67 453 101
rect 401 51 453 67
rect 487 133 503 167
rect 537 133 741 167
rect 487 131 741 133
rect 487 91 553 131
rect 687 101 741 131
rect 487 57 503 91
rect 537 57 553 91
rect 487 51 553 57
rect 587 93 653 97
rect 587 59 603 93
rect 637 59 653 93
rect 587 17 653 59
rect 687 67 691 101
rect 725 67 741 101
rect 687 51 741 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21ba_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6549682
string GDS_START 6542026
<< end >>
