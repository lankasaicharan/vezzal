magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 496 263 598 267
rect 278 241 598 263
rect 893 241 1343 261
rect 1 49 1343 241
rect 0 0 1344 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 252 47 282 215
rect 384 47 414 215
rect 470 47 500 215
rect 594 47 624 215
rect 696 47 726 215
rect 782 47 812 215
rect 976 67 1006 235
rect 1062 67 1092 235
rect 1148 67 1178 235
rect 1234 67 1264 235
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 452 367 482 619
rect 538 367 568 619
rect 624 367 654 619
rect 710 367 740 619
rect 796 367 826 619
rect 882 367 912 619
rect 976 367 1006 619
rect 1062 367 1092 619
rect 1148 367 1178 619
rect 1234 367 1264 619
<< ndiff >>
rect 304 229 362 237
rect 304 215 316 229
rect 27 192 80 215
rect 27 158 35 192
rect 69 158 80 192
rect 27 93 80 158
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 190 166 215
rect 110 156 121 190
rect 155 156 166 190
rect 110 101 166 156
rect 110 67 121 101
rect 155 67 166 101
rect 110 47 166 67
rect 196 89 252 215
rect 196 55 207 89
rect 241 55 252 89
rect 196 47 252 55
rect 282 195 316 215
rect 350 215 362 229
rect 522 229 572 241
rect 522 215 530 229
rect 350 195 384 215
rect 282 47 384 195
rect 414 89 470 215
rect 414 55 425 89
rect 459 55 470 89
rect 414 47 470 55
rect 500 195 530 215
rect 564 215 572 229
rect 564 195 594 215
rect 500 47 594 195
rect 624 89 696 215
rect 624 55 635 89
rect 669 55 696 89
rect 624 47 696 55
rect 726 175 782 215
rect 726 141 737 175
rect 771 141 782 175
rect 726 107 782 141
rect 726 73 737 107
rect 771 73 782 107
rect 726 47 782 73
rect 812 93 865 215
rect 812 59 823 93
rect 857 59 865 93
rect 919 109 976 235
rect 919 75 931 109
rect 965 75 976 109
rect 919 67 976 75
rect 1006 179 1062 235
rect 1006 145 1017 179
rect 1051 145 1062 179
rect 1006 67 1062 145
rect 1092 109 1148 235
rect 1092 75 1103 109
rect 1137 75 1148 109
rect 1092 67 1148 75
rect 1178 227 1234 235
rect 1178 193 1189 227
rect 1223 193 1234 227
rect 1178 159 1234 193
rect 1178 125 1189 159
rect 1223 125 1234 159
rect 1178 67 1234 125
rect 1264 223 1317 235
rect 1264 189 1275 223
rect 1309 189 1317 223
rect 1264 113 1317 189
rect 1264 79 1275 113
rect 1309 79 1317 113
rect 1264 67 1317 79
rect 812 47 865 59
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 514 80 565
rect 27 480 35 514
rect 69 480 80 514
rect 27 436 80 480
rect 27 402 35 436
rect 69 402 80 436
rect 27 367 80 402
rect 110 531 166 619
rect 110 497 121 531
rect 155 497 166 531
rect 110 413 166 497
rect 110 379 121 413
rect 155 379 166 413
rect 110 367 166 379
rect 196 599 249 619
rect 196 565 207 599
rect 241 565 249 599
rect 196 514 249 565
rect 196 480 207 514
rect 241 480 249 514
rect 196 436 249 480
rect 196 402 207 436
rect 241 402 249 436
rect 196 367 249 402
rect 399 600 452 619
rect 399 566 407 600
rect 441 566 452 600
rect 399 367 452 566
rect 482 436 538 619
rect 482 402 493 436
rect 527 402 538 436
rect 482 367 538 402
rect 568 600 624 619
rect 568 566 579 600
rect 613 566 624 600
rect 568 367 624 566
rect 654 436 710 619
rect 654 402 665 436
rect 699 402 710 436
rect 654 367 710 402
rect 740 600 796 619
rect 740 566 751 600
rect 785 566 796 600
rect 740 367 796 566
rect 826 599 882 619
rect 826 565 837 599
rect 871 565 882 599
rect 826 525 882 565
rect 826 491 837 525
rect 871 491 882 525
rect 826 436 882 491
rect 826 402 837 436
rect 871 402 882 436
rect 826 367 882 402
rect 912 607 976 619
rect 912 573 927 607
rect 961 573 976 607
rect 912 494 976 573
rect 912 460 927 494
rect 961 460 976 494
rect 912 367 976 460
rect 1006 599 1062 619
rect 1006 565 1017 599
rect 1051 565 1062 599
rect 1006 525 1062 565
rect 1006 491 1017 525
rect 1051 491 1062 525
rect 1006 436 1062 491
rect 1006 402 1017 436
rect 1051 402 1062 436
rect 1006 367 1062 402
rect 1092 607 1148 619
rect 1092 573 1103 607
rect 1137 573 1148 607
rect 1092 494 1148 573
rect 1092 460 1103 494
rect 1137 460 1148 494
rect 1092 367 1148 460
rect 1178 599 1234 619
rect 1178 565 1189 599
rect 1223 565 1234 599
rect 1178 525 1234 565
rect 1178 491 1189 525
rect 1223 491 1234 525
rect 1178 436 1234 491
rect 1178 402 1189 436
rect 1223 402 1234 436
rect 1178 367 1234 402
rect 1264 607 1317 619
rect 1264 573 1275 607
rect 1309 573 1317 607
rect 1264 506 1317 573
rect 1264 472 1275 506
rect 1309 472 1317 506
rect 1264 420 1317 472
rect 1264 386 1275 420
rect 1309 386 1317 420
rect 1264 367 1317 386
<< ndiffc >>
rect 35 158 69 192
rect 35 59 69 93
rect 121 156 155 190
rect 121 67 155 101
rect 207 55 241 89
rect 316 195 350 229
rect 425 55 459 89
rect 530 195 564 229
rect 635 55 669 89
rect 737 141 771 175
rect 737 73 771 107
rect 823 59 857 93
rect 931 75 965 109
rect 1017 145 1051 179
rect 1103 75 1137 109
rect 1189 193 1223 227
rect 1189 125 1223 159
rect 1275 189 1309 223
rect 1275 79 1309 113
<< pdiffc >>
rect 35 565 69 599
rect 35 480 69 514
rect 35 402 69 436
rect 121 497 155 531
rect 121 379 155 413
rect 207 565 241 599
rect 207 480 241 514
rect 207 402 241 436
rect 407 566 441 600
rect 493 402 527 436
rect 579 566 613 600
rect 665 402 699 436
rect 751 566 785 600
rect 837 565 871 599
rect 837 491 871 525
rect 837 402 871 436
rect 927 573 961 607
rect 927 460 961 494
rect 1017 565 1051 599
rect 1017 491 1051 525
rect 1017 402 1051 436
rect 1103 573 1137 607
rect 1103 460 1137 494
rect 1189 565 1223 599
rect 1189 491 1223 525
rect 1189 402 1223 436
rect 1275 573 1309 607
rect 1275 472 1309 506
rect 1275 386 1309 420
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 452 619 482 645
rect 538 619 568 645
rect 624 619 654 645
rect 710 619 740 645
rect 796 619 826 645
rect 882 619 912 645
rect 976 619 1006 645
rect 1062 619 1092 645
rect 1148 619 1178 645
rect 1234 619 1264 645
rect 80 308 110 367
rect 166 308 196 367
rect 452 345 482 367
rect 538 345 568 367
rect 624 345 654 367
rect 710 345 740 367
rect 452 329 740 345
rect 796 335 826 367
rect 882 335 912 367
rect 35 292 196 308
rect 378 315 740 329
rect 782 319 912 335
rect 378 313 648 315
rect 378 293 394 313
rect 35 258 51 292
rect 85 278 196 292
rect 85 258 110 278
rect 35 242 110 258
rect 80 215 110 242
rect 166 215 196 278
rect 252 279 394 293
rect 428 279 462 313
rect 496 279 530 313
rect 564 279 598 313
rect 632 279 648 313
rect 252 263 648 279
rect 782 285 798 319
rect 832 305 912 319
rect 976 335 1006 367
rect 1062 335 1092 367
rect 976 319 1092 335
rect 832 285 848 305
rect 782 267 848 285
rect 252 215 282 263
rect 384 215 414 263
rect 470 215 500 263
rect 594 215 624 263
rect 696 237 848 267
rect 976 285 1042 319
rect 1076 285 1092 319
rect 976 269 1092 285
rect 696 215 726 237
rect 782 215 812 237
rect 976 235 1006 269
rect 1062 235 1092 269
rect 1148 335 1178 367
rect 1234 335 1264 367
rect 1148 319 1264 335
rect 1148 285 1214 319
rect 1248 285 1264 319
rect 1148 269 1264 285
rect 1148 235 1178 269
rect 1234 235 1264 269
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 384 21 414 47
rect 470 21 500 47
rect 594 21 624 47
rect 696 21 726 47
rect 782 21 812 47
rect 976 41 1006 67
rect 1062 41 1092 67
rect 1148 41 1178 67
rect 1234 41 1264 67
<< polycont >>
rect 51 258 85 292
rect 394 279 428 313
rect 462 279 496 313
rect 530 279 564 313
rect 598 279 632 313
rect 798 285 832 319
rect 1042 285 1076 319
rect 1214 285 1248 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 19 599 257 615
rect 19 565 35 599
rect 69 581 207 599
rect 69 565 85 581
rect 19 514 85 565
rect 205 565 207 581
rect 241 565 257 599
rect 19 480 35 514
rect 69 480 85 514
rect 19 436 85 480
rect 19 402 35 436
rect 69 402 85 436
rect 19 386 85 402
rect 119 531 171 547
rect 119 497 121 531
rect 155 497 171 531
rect 119 413 171 497
rect 119 379 121 413
rect 155 379 171 413
rect 205 522 257 565
rect 391 600 457 649
rect 391 566 407 600
rect 441 566 457 600
rect 391 556 457 566
rect 563 600 629 649
rect 563 566 579 600
rect 613 566 629 600
rect 563 556 629 566
rect 735 600 801 649
rect 735 566 751 600
rect 785 566 801 600
rect 735 556 801 566
rect 835 599 877 615
rect 835 565 837 599
rect 871 565 877 599
rect 835 525 877 565
rect 835 522 837 525
rect 205 514 837 522
rect 205 480 207 514
rect 241 491 837 514
rect 871 491 877 525
rect 241 488 877 491
rect 241 480 247 488
rect 205 436 247 480
rect 205 402 207 436
rect 241 402 247 436
rect 205 386 247 402
rect 281 436 715 452
rect 281 402 493 436
rect 527 402 665 436
rect 699 402 715 436
rect 281 386 715 402
rect 821 436 877 488
rect 911 607 977 649
rect 911 573 927 607
rect 961 573 977 607
rect 911 494 977 573
rect 911 460 927 494
rect 961 460 977 494
rect 911 454 977 460
rect 1011 599 1053 615
rect 1011 565 1017 599
rect 1051 565 1053 599
rect 1011 525 1053 565
rect 1011 491 1017 525
rect 1051 491 1053 525
rect 821 402 837 436
rect 871 420 877 436
rect 1011 436 1053 491
rect 1087 607 1153 649
rect 1087 573 1103 607
rect 1137 573 1153 607
rect 1087 494 1153 573
rect 1087 460 1103 494
rect 1137 460 1153 494
rect 1087 454 1153 460
rect 1187 599 1225 615
rect 1187 565 1189 599
rect 1223 565 1225 599
rect 1187 525 1225 565
rect 1187 491 1189 525
rect 1223 491 1225 525
rect 1011 420 1017 436
rect 871 402 1017 420
rect 1051 420 1053 436
rect 1187 436 1225 491
rect 1187 420 1189 436
rect 1051 402 1189 420
rect 1223 402 1225 436
rect 821 386 1225 402
rect 1259 607 1325 649
rect 1259 573 1275 607
rect 1309 573 1325 607
rect 1259 506 1325 573
rect 1259 472 1275 506
rect 1309 472 1325 506
rect 1259 420 1325 472
rect 1259 386 1275 420
rect 1309 386 1325 420
rect 31 292 85 352
rect 31 258 51 292
rect 31 242 85 258
rect 19 192 85 208
rect 19 158 35 192
rect 69 158 85 192
rect 19 93 85 158
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 119 190 171 379
rect 281 352 338 386
rect 205 237 338 352
rect 378 313 650 329
rect 378 279 394 313
rect 428 279 462 313
rect 496 279 530 313
rect 564 279 598 313
rect 632 279 650 313
rect 703 319 929 350
rect 703 285 798 319
rect 832 285 929 319
rect 703 283 929 285
rect 991 319 1121 352
rect 991 285 1042 319
rect 1076 285 1121 319
rect 991 283 1121 285
rect 1183 319 1313 352
rect 1183 285 1214 319
rect 1248 285 1313 319
rect 1183 283 1313 285
rect 378 271 650 279
rect 616 249 650 271
rect 205 229 580 237
rect 205 195 316 229
rect 350 195 530 229
rect 564 195 580 229
rect 616 227 1239 249
rect 616 215 1189 227
rect 119 156 121 190
rect 155 161 171 190
rect 616 161 650 215
rect 1173 193 1189 215
rect 1223 193 1239 227
rect 155 156 650 161
rect 119 127 650 156
rect 721 179 1067 181
rect 721 175 1017 179
rect 721 141 737 175
rect 771 145 1017 175
rect 1051 145 1067 179
rect 1173 159 1239 193
rect 771 141 787 145
rect 119 101 157 127
rect 119 67 121 101
rect 155 67 157 101
rect 721 107 787 141
rect 1103 111 1139 129
rect 1173 125 1189 159
rect 1223 125 1239 159
rect 1173 123 1239 125
rect 1273 223 1325 239
rect 1273 189 1275 223
rect 1309 189 1325 223
rect 915 109 1139 111
rect 119 51 157 67
rect 191 89 257 93
rect 191 55 207 89
rect 241 55 257 89
rect 191 17 257 55
rect 409 89 475 93
rect 409 55 425 89
rect 459 55 475 89
rect 409 17 475 55
rect 619 89 685 93
rect 619 55 635 89
rect 669 55 685 89
rect 721 73 737 107
rect 771 73 787 107
rect 721 69 787 73
rect 821 93 861 109
rect 619 17 685 55
rect 821 59 823 93
rect 857 59 861 93
rect 821 17 861 59
rect 915 75 931 109
rect 965 75 1103 109
rect 1137 89 1139 109
rect 1273 113 1325 189
rect 1273 89 1275 113
rect 1137 79 1275 89
rect 1309 79 1325 113
rect 1137 75 1325 79
rect 915 55 1325 75
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a31o_4
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2607920
string GDS_START 2597082
<< end >>
