magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 331 1958 704
rect 238 323 563 331
<< pwell >>
rect 521 254 795 277
rect 242 180 795 254
rect 1551 241 1879 256
rect 3 179 795 180
rect 1102 179 1879 241
rect 3 49 1879 179
rect 0 0 1920 49
<< scnmos >>
rect 82 70 112 154
rect 321 144 351 228
rect 407 144 437 228
rect 600 167 630 251
rect 686 167 716 251
rect 905 69 935 153
rect 991 69 1021 153
rect 1181 47 1211 215
rect 1253 47 1283 215
rect 1406 131 1436 215
rect 1630 62 1660 230
rect 1766 62 1796 230
<< scpmoshvt >>
rect 91 473 121 601
rect 327 359 357 487
rect 444 359 474 487
rect 678 377 708 461
rect 783 377 813 505
rect 855 377 885 505
rect 960 377 990 461
rect 1173 367 1203 619
rect 1259 367 1289 619
rect 1364 367 1394 495
rect 1630 367 1660 619
rect 1716 367 1746 619
<< ndiff >>
rect 268 202 321 228
rect 268 168 276 202
rect 310 168 321 202
rect 29 125 82 154
rect 29 91 37 125
rect 71 91 82 125
rect 29 70 82 91
rect 112 118 165 154
rect 268 144 321 168
rect 351 192 407 228
rect 351 158 362 192
rect 396 158 407 192
rect 351 144 407 158
rect 437 192 490 228
rect 437 158 448 192
rect 482 158 490 192
rect 547 226 600 251
rect 547 192 555 226
rect 589 192 600 226
rect 547 167 600 192
rect 630 239 686 251
rect 630 205 641 239
rect 675 205 686 239
rect 630 167 686 205
rect 716 227 769 251
rect 716 193 727 227
rect 761 193 769 227
rect 716 167 769 193
rect 437 144 490 158
rect 112 84 123 118
rect 157 84 165 118
rect 112 70 165 84
rect 1128 196 1181 215
rect 1128 162 1136 196
rect 1170 162 1181 196
rect 852 128 905 153
rect 852 94 860 128
rect 894 94 905 128
rect 852 69 905 94
rect 935 128 991 153
rect 935 94 946 128
rect 980 94 991 128
rect 935 69 991 94
rect 1021 128 1074 153
rect 1021 94 1032 128
rect 1066 94 1074 128
rect 1021 69 1074 94
rect 1128 95 1181 162
rect 1128 61 1136 95
rect 1170 61 1181 95
rect 1128 47 1181 61
rect 1211 47 1253 215
rect 1283 131 1406 215
rect 1436 191 1508 215
rect 1436 157 1466 191
rect 1500 157 1508 191
rect 1436 131 1508 157
rect 1577 169 1630 230
rect 1577 135 1585 169
rect 1619 135 1630 169
rect 1283 125 1336 131
rect 1283 91 1294 125
rect 1328 91 1336 125
rect 1283 47 1336 91
rect 1577 62 1630 135
rect 1660 202 1766 230
rect 1660 168 1721 202
rect 1755 168 1766 202
rect 1660 108 1766 168
rect 1660 74 1721 108
rect 1755 74 1766 108
rect 1660 62 1766 74
rect 1796 212 1853 230
rect 1796 178 1807 212
rect 1841 178 1853 212
rect 1796 108 1853 178
rect 1796 74 1807 108
rect 1841 74 1853 108
rect 1796 62 1853 74
<< pdiff >>
rect 38 589 91 601
rect 38 555 46 589
rect 80 555 91 589
rect 38 519 91 555
rect 38 485 46 519
rect 80 485 91 519
rect 38 473 91 485
rect 121 589 174 601
rect 121 555 132 589
rect 166 555 174 589
rect 121 521 174 555
rect 121 487 132 521
rect 166 487 174 521
rect 121 473 174 487
rect 274 475 327 487
rect 274 441 282 475
rect 316 441 327 475
rect 274 405 327 441
rect 274 371 282 405
rect 316 371 327 405
rect 274 359 327 371
rect 357 475 444 487
rect 357 441 383 475
rect 417 441 444 475
rect 357 405 444 441
rect 357 371 383 405
rect 417 371 444 405
rect 357 359 444 371
rect 474 473 527 487
rect 474 439 485 473
rect 519 439 527 473
rect 474 405 527 439
rect 474 371 485 405
rect 519 371 527 405
rect 474 359 527 371
rect 730 489 783 505
rect 730 461 738 489
rect 625 436 678 461
rect 625 402 633 436
rect 667 402 678 436
rect 625 377 678 402
rect 708 455 738 461
rect 772 455 783 489
rect 708 377 783 455
rect 813 377 855 505
rect 885 479 938 505
rect 885 445 896 479
rect 930 461 938 479
rect 930 445 960 461
rect 885 377 960 445
rect 990 436 1043 461
rect 990 402 1001 436
rect 1035 402 1043 436
rect 990 377 1043 402
rect 1120 607 1173 619
rect 1120 573 1128 607
rect 1162 573 1173 607
rect 1120 492 1173 573
rect 1120 458 1128 492
rect 1162 458 1173 492
rect 1120 367 1173 458
rect 1203 599 1259 619
rect 1203 565 1214 599
rect 1248 565 1259 599
rect 1203 516 1259 565
rect 1203 482 1214 516
rect 1248 482 1259 516
rect 1203 436 1259 482
rect 1203 402 1214 436
rect 1248 402 1259 436
rect 1203 367 1259 402
rect 1289 607 1342 619
rect 1289 573 1300 607
rect 1334 573 1342 607
rect 1289 515 1342 573
rect 1577 599 1630 619
rect 1577 565 1585 599
rect 1619 565 1630 599
rect 1289 481 1300 515
rect 1334 495 1342 515
rect 1577 504 1630 565
rect 1334 481 1364 495
rect 1289 420 1364 481
rect 1289 386 1312 420
rect 1346 386 1364 420
rect 1289 367 1364 386
rect 1394 481 1447 495
rect 1394 447 1405 481
rect 1439 447 1447 481
rect 1577 470 1585 504
rect 1619 470 1630 504
rect 1394 413 1447 447
rect 1394 379 1405 413
rect 1439 379 1447 413
rect 1394 367 1447 379
rect 1577 420 1630 470
rect 1577 386 1585 420
rect 1619 386 1630 420
rect 1577 367 1630 386
rect 1660 607 1716 619
rect 1660 573 1671 607
rect 1705 573 1716 607
rect 1660 507 1716 573
rect 1660 473 1671 507
rect 1705 473 1716 507
rect 1660 413 1716 473
rect 1660 379 1671 413
rect 1705 379 1716 413
rect 1660 367 1716 379
rect 1746 599 1799 619
rect 1746 565 1757 599
rect 1791 565 1799 599
rect 1746 504 1799 565
rect 1746 470 1757 504
rect 1791 470 1799 504
rect 1746 413 1799 470
rect 1746 379 1757 413
rect 1791 379 1799 413
rect 1746 367 1799 379
<< ndiffc >>
rect 276 168 310 202
rect 37 91 71 125
rect 362 158 396 192
rect 448 158 482 192
rect 555 192 589 226
rect 641 205 675 239
rect 727 193 761 227
rect 123 84 157 118
rect 1136 162 1170 196
rect 860 94 894 128
rect 946 94 980 128
rect 1032 94 1066 128
rect 1136 61 1170 95
rect 1466 157 1500 191
rect 1585 135 1619 169
rect 1294 91 1328 125
rect 1721 168 1755 202
rect 1721 74 1755 108
rect 1807 178 1841 212
rect 1807 74 1841 108
<< pdiffc >>
rect 46 555 80 589
rect 46 485 80 519
rect 132 555 166 589
rect 132 487 166 521
rect 282 441 316 475
rect 282 371 316 405
rect 383 441 417 475
rect 383 371 417 405
rect 485 439 519 473
rect 485 371 519 405
rect 633 402 667 436
rect 738 455 772 489
rect 896 445 930 479
rect 1001 402 1035 436
rect 1128 573 1162 607
rect 1128 458 1162 492
rect 1214 565 1248 599
rect 1214 482 1248 516
rect 1214 402 1248 436
rect 1300 573 1334 607
rect 1585 565 1619 599
rect 1300 481 1334 515
rect 1312 386 1346 420
rect 1405 447 1439 481
rect 1585 470 1619 504
rect 1405 379 1439 413
rect 1585 386 1619 420
rect 1671 573 1705 607
rect 1671 473 1705 507
rect 1671 379 1705 413
rect 1757 565 1791 599
rect 1757 470 1791 504
rect 1757 379 1791 413
<< poly >>
rect 91 601 121 627
rect 281 605 572 621
rect 281 571 297 605
rect 331 591 572 605
rect 331 571 347 591
rect 281 555 347 571
rect 542 513 572 591
rect 669 605 1099 621
rect 1173 619 1203 645
rect 1259 619 1289 645
rect 1630 619 1660 645
rect 1716 619 1746 645
rect 669 571 685 605
rect 719 591 1099 605
rect 719 571 735 591
rect 669 555 735 571
rect 327 487 357 513
rect 444 487 474 513
rect 91 377 121 473
rect 46 361 121 377
rect 46 327 62 361
rect 96 327 121 361
rect 46 293 121 327
rect 163 419 229 435
rect 163 385 179 419
rect 213 385 229 419
rect 163 351 229 385
rect 542 483 708 513
rect 783 505 813 531
rect 855 505 885 531
rect 542 362 572 483
rect 678 461 708 483
rect 960 461 990 487
rect 163 317 179 351
rect 213 331 229 351
rect 327 331 357 359
rect 213 317 357 331
rect 163 301 357 317
rect 444 316 474 359
rect 542 332 630 362
rect 678 351 708 377
rect 46 259 62 293
rect 96 259 121 293
rect 46 243 121 259
rect 82 154 112 243
rect 321 228 351 301
rect 399 300 474 316
rect 399 266 415 300
rect 449 266 474 300
rect 399 250 474 266
rect 600 251 630 332
rect 783 303 813 377
rect 686 273 813 303
rect 686 251 716 273
rect 407 228 437 250
rect 855 205 885 377
rect 960 337 990 377
rect 1069 345 1099 591
rect 1364 495 1394 521
rect 1479 433 1545 449
rect 1479 399 1495 433
rect 1529 399 1545 433
rect 1173 345 1203 367
rect 955 321 1021 337
rect 955 287 971 321
rect 1005 287 1021 321
rect 1069 315 1211 345
rect 955 271 1021 287
rect 794 175 935 205
rect 321 118 351 144
rect 407 118 437 144
rect 600 141 630 167
rect 207 90 273 106
rect 82 44 112 70
rect 207 56 223 90
rect 257 70 273 90
rect 686 70 716 167
rect 794 103 824 175
rect 905 153 935 175
rect 991 153 1021 271
rect 1181 215 1211 315
rect 1259 308 1289 367
rect 1253 292 1319 308
rect 1253 258 1269 292
rect 1303 258 1319 292
rect 1253 242 1319 258
rect 1364 303 1394 367
rect 1479 365 1545 399
rect 1479 331 1495 365
rect 1529 345 1545 365
rect 1630 345 1660 367
rect 1529 331 1660 345
rect 1479 315 1660 331
rect 1364 287 1430 303
rect 1364 253 1380 287
rect 1414 267 1430 287
rect 1414 253 1436 267
rect 1253 215 1283 242
rect 1364 237 1436 253
rect 1406 215 1436 237
rect 1630 230 1660 315
rect 1716 318 1746 367
rect 1716 302 1796 318
rect 1716 268 1732 302
rect 1766 268 1796 302
rect 1716 252 1796 268
rect 1766 230 1796 252
rect 257 56 716 70
rect 207 40 716 56
rect 758 87 824 103
rect 758 53 774 87
rect 808 53 824 87
rect 758 37 824 53
rect 905 43 935 69
rect 991 43 1021 69
rect 1406 105 1436 131
rect 1181 21 1211 47
rect 1253 21 1283 47
rect 1630 36 1660 62
rect 1766 36 1796 62
<< polycont >>
rect 297 571 331 605
rect 685 571 719 605
rect 62 327 96 361
rect 179 385 213 419
rect 179 317 213 351
rect 62 259 96 293
rect 415 266 449 300
rect 1495 399 1529 433
rect 971 287 1005 321
rect 223 56 257 90
rect 1269 258 1303 292
rect 1495 331 1529 365
rect 1380 253 1414 287
rect 1732 268 1766 302
rect 774 53 808 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 30 589 96 649
rect 30 555 46 589
rect 80 555 96 589
rect 30 519 96 555
rect 30 485 46 519
rect 80 485 96 519
rect 30 469 96 485
rect 132 605 347 615
rect 132 589 297 605
rect 166 571 297 589
rect 331 571 347 605
rect 166 555 347 571
rect 132 521 170 555
rect 381 521 449 649
rect 669 605 735 615
rect 669 571 685 605
rect 719 571 735 605
rect 669 542 735 571
rect 166 487 170 521
rect 132 435 170 487
rect 249 475 332 491
rect 249 441 282 475
rect 316 441 332 475
rect 17 361 96 435
rect 17 327 62 361
rect 17 293 96 327
rect 17 259 62 293
rect 17 168 96 259
rect 132 419 213 435
rect 132 385 179 419
rect 132 351 213 385
rect 132 317 179 351
rect 132 301 213 317
rect 249 405 332 441
rect 249 371 282 405
rect 316 371 332 405
rect 249 355 332 371
rect 367 487 449 521
rect 559 541 735 542
rect 559 489 788 541
rect 367 475 433 487
rect 367 441 383 475
rect 417 441 433 475
rect 367 405 433 441
rect 367 371 383 405
rect 417 371 433 405
rect 367 355 433 371
rect 485 473 525 489
rect 519 439 525 473
rect 485 405 525 439
rect 519 371 525 405
rect 485 355 525 371
rect 559 486 738 489
rect 132 134 166 301
rect 249 208 283 355
rect 317 300 451 316
rect 317 266 415 300
rect 449 266 451 300
rect 317 242 451 266
rect 485 208 519 355
rect 559 337 593 486
rect 722 455 738 486
rect 772 455 788 489
rect 627 436 671 452
rect 722 439 788 455
rect 880 479 946 649
rect 880 445 896 479
rect 930 445 946 479
rect 1112 607 1178 649
rect 1112 573 1128 607
rect 1162 573 1178 607
rect 1112 492 1178 573
rect 1112 458 1128 492
rect 1162 458 1178 492
rect 1112 454 1178 458
rect 1212 599 1257 615
rect 1212 565 1214 599
rect 1248 565 1257 599
rect 1212 516 1257 565
rect 1212 482 1214 516
rect 1248 482 1257 516
rect 880 439 946 445
rect 627 402 633 436
rect 667 405 671 436
rect 985 436 1051 452
rect 985 405 1001 436
rect 667 402 1001 405
rect 1035 402 1051 436
rect 1212 436 1257 482
rect 1212 420 1214 436
rect 627 371 1051 402
rect 1085 402 1214 420
rect 1248 402 1257 436
rect 1085 386 1257 402
rect 1291 607 1362 649
rect 1291 573 1300 607
rect 1334 573 1362 607
rect 1291 515 1362 573
rect 1291 481 1300 515
rect 1334 481 1362 515
rect 1567 599 1623 615
rect 1567 565 1585 599
rect 1619 565 1623 599
rect 1567 504 1623 565
rect 1291 420 1362 481
rect 1291 386 1312 420
rect 1346 386 1362 420
rect 1396 481 1533 497
rect 1396 447 1405 481
rect 1439 447 1533 481
rect 1396 433 1533 447
rect 1396 413 1495 433
rect 1085 337 1147 386
rect 1396 379 1405 413
rect 1439 399 1495 413
rect 1529 399 1533 433
rect 1439 379 1533 399
rect 1396 365 1533 379
rect 1396 363 1495 365
rect 559 303 677 337
rect 249 206 326 208
rect 21 125 87 134
rect 21 91 37 125
rect 71 91 87 125
rect 21 17 87 91
rect 121 118 166 134
rect 121 84 123 118
rect 157 84 166 118
rect 121 68 166 84
rect 207 202 326 206
rect 207 168 276 202
rect 310 168 326 202
rect 207 152 326 168
rect 360 192 404 208
rect 360 158 362 192
rect 396 158 404 192
rect 207 90 273 152
rect 207 56 223 90
rect 257 56 273 90
rect 360 17 404 158
rect 438 192 519 208
rect 438 158 448 192
rect 482 158 519 192
rect 438 142 519 158
rect 485 87 519 142
rect 553 226 598 242
rect 553 192 555 226
rect 589 192 598 226
rect 553 155 598 192
rect 632 239 677 303
rect 955 321 1147 337
rect 955 287 971 321
rect 1005 287 1147 321
rect 955 271 1147 287
rect 632 205 641 239
rect 675 205 677 239
rect 632 189 677 205
rect 711 227 1074 235
rect 711 193 727 227
rect 761 193 1074 227
rect 711 189 1074 193
rect 553 128 903 155
rect 553 121 860 128
rect 858 94 860 121
rect 894 94 903 128
rect 485 53 774 87
rect 808 53 824 87
rect 858 78 903 94
rect 937 128 984 144
rect 937 94 946 128
rect 980 94 984 128
rect 937 17 984 94
rect 1028 128 1074 189
rect 1028 94 1032 128
rect 1066 94 1074 128
rect 1028 78 1074 94
rect 1108 200 1147 271
rect 1181 292 1330 352
rect 1479 331 1495 363
rect 1529 331 1533 365
rect 1181 258 1269 292
rect 1303 258 1330 292
rect 1181 234 1330 258
rect 1364 287 1416 303
rect 1364 253 1380 287
rect 1414 253 1416 287
rect 1364 200 1416 253
rect 1479 207 1533 331
rect 1108 196 1416 200
rect 1108 162 1136 196
rect 1170 166 1416 196
rect 1170 162 1186 166
rect 1108 95 1186 162
rect 1108 61 1136 95
rect 1170 61 1186 95
rect 1108 51 1186 61
rect 1278 125 1344 132
rect 1278 91 1294 125
rect 1328 91 1344 125
rect 1278 17 1344 91
rect 1380 85 1416 166
rect 1450 191 1533 207
rect 1450 157 1466 191
rect 1500 157 1533 191
rect 1450 141 1533 157
rect 1567 470 1585 504
rect 1619 470 1623 504
rect 1567 420 1623 470
rect 1567 386 1585 420
rect 1619 386 1623 420
rect 1567 370 1623 386
rect 1657 607 1709 649
rect 1657 573 1671 607
rect 1705 573 1709 607
rect 1657 507 1709 573
rect 1657 473 1671 507
rect 1705 473 1709 507
rect 1657 413 1709 473
rect 1657 379 1671 413
rect 1705 379 1709 413
rect 1567 169 1619 370
rect 1657 363 1709 379
rect 1753 599 1903 615
rect 1753 565 1757 599
rect 1791 565 1903 599
rect 1753 504 1903 565
rect 1753 470 1757 504
rect 1791 470 1903 504
rect 1753 413 1903 470
rect 1753 379 1757 413
rect 1791 379 1903 413
rect 1753 363 1903 379
rect 1567 135 1585 169
rect 1567 119 1619 135
rect 1653 302 1777 318
rect 1653 268 1732 302
rect 1766 268 1777 302
rect 1653 252 1777 268
rect 1653 85 1687 252
rect 1811 228 1903 363
rect 1380 51 1687 85
rect 1721 202 1768 218
rect 1755 168 1768 202
rect 1721 108 1768 168
rect 1755 74 1768 108
rect 1721 17 1768 74
rect 1802 212 1903 228
rect 1802 178 1807 212
rect 1841 178 1903 212
rect 1802 108 1903 178
rect 1802 74 1807 108
rect 1841 74 1903 108
rect 1802 58 1903 74
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrbn_1
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1855 94 1889 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 168 1889 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 390 1889 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 464 1889 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 538 1889 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6234122
string GDS_START 6217974
<< end >>
