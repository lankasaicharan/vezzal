magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1778 1975
<< nwell >>
rect -38 331 518 704
<< pwell >>
rect 197 157 471 241
rect 20 49 471 157
rect 0 0 480 49
<< scnmos >>
rect 99 47 129 131
rect 171 47 201 131
rect 276 47 306 215
rect 362 47 392 215
<< scpmoshvt >>
rect 85 397 115 481
rect 171 397 201 481
rect 276 367 306 619
rect 362 367 392 619
<< ndiff >>
rect 223 131 276 215
rect 46 106 99 131
rect 46 72 54 106
rect 88 72 99 106
rect 46 47 99 72
rect 129 47 171 131
rect 201 97 276 131
rect 201 63 222 97
rect 256 63 276 97
rect 201 47 276 63
rect 306 202 362 215
rect 306 168 317 202
rect 351 168 362 202
rect 306 101 362 168
rect 306 67 317 101
rect 351 67 362 101
rect 306 47 362 67
rect 392 202 445 215
rect 392 168 403 202
rect 437 168 445 202
rect 392 93 445 168
rect 392 59 403 93
rect 437 59 445 93
rect 392 47 445 59
<< pdiff >>
rect 223 607 276 619
rect 223 573 231 607
rect 265 573 276 607
rect 223 526 276 573
rect 223 492 231 526
rect 265 492 276 526
rect 223 481 276 492
rect 32 456 85 481
rect 32 422 40 456
rect 74 422 85 456
rect 32 397 85 422
rect 115 456 171 481
rect 115 422 126 456
rect 160 422 171 456
rect 115 397 171 422
rect 201 439 276 481
rect 201 405 212 439
rect 246 405 276 439
rect 201 397 276 405
rect 223 367 276 397
rect 306 599 362 619
rect 306 565 317 599
rect 351 565 362 599
rect 306 515 362 565
rect 306 481 317 515
rect 351 481 362 515
rect 306 438 362 481
rect 306 404 317 438
rect 351 404 362 438
rect 306 367 362 404
rect 392 607 445 619
rect 392 573 403 607
rect 437 573 445 607
rect 392 507 445 573
rect 392 473 403 507
rect 437 473 445 507
rect 392 413 445 473
rect 392 379 403 413
rect 437 379 445 413
rect 392 367 445 379
<< ndiffc >>
rect 54 72 88 106
rect 222 63 256 97
rect 317 168 351 202
rect 317 67 351 101
rect 403 168 437 202
rect 403 59 437 93
<< pdiffc >>
rect 231 573 265 607
rect 231 492 265 526
rect 40 422 74 456
rect 126 422 160 456
rect 212 405 246 439
rect 317 565 351 599
rect 317 481 351 515
rect 317 404 351 438
rect 403 573 437 607
rect 403 473 437 507
rect 403 379 437 413
<< poly >>
rect 276 619 306 645
rect 362 619 392 645
rect 85 481 115 507
rect 171 481 201 507
rect 85 375 115 397
rect 57 345 115 375
rect 57 325 87 345
rect 21 309 87 325
rect 21 275 37 309
rect 71 275 87 309
rect 171 297 201 397
rect 276 320 306 367
rect 21 241 87 275
rect 21 207 37 241
rect 71 207 87 241
rect 135 281 201 297
rect 135 247 151 281
rect 185 247 201 281
rect 243 304 309 320
rect 243 270 259 304
rect 293 284 309 304
rect 362 284 392 367
rect 293 270 392 284
rect 243 254 392 270
rect 135 231 201 247
rect 21 191 87 207
rect 57 183 87 191
rect 57 153 129 183
rect 99 131 129 153
rect 171 131 201 231
rect 276 215 306 254
rect 362 215 392 254
rect 99 21 129 47
rect 171 21 201 47
rect 276 21 306 47
rect 362 21 392 47
<< polycont >>
rect 37 275 71 309
rect 37 207 71 241
rect 151 247 185 281
rect 259 270 293 304
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 24 456 90 649
rect 203 607 272 649
rect 203 573 231 607
rect 265 573 272 607
rect 203 526 272 573
rect 203 492 231 526
rect 265 492 272 526
rect 24 422 40 456
rect 74 422 90 456
rect 24 406 90 422
rect 124 456 169 472
rect 124 422 126 456
rect 160 422 169 456
rect 21 309 87 372
rect 124 354 169 422
rect 203 439 272 492
rect 203 405 212 439
rect 246 405 272 439
rect 203 389 272 405
rect 306 599 363 615
rect 306 565 317 599
rect 351 565 363 599
rect 306 515 363 565
rect 306 481 317 515
rect 351 481 363 515
rect 306 438 363 481
rect 306 404 317 438
rect 351 404 363 438
rect 306 388 363 404
rect 124 320 293 354
rect 21 275 37 309
rect 71 275 87 309
rect 247 304 293 320
rect 21 241 87 275
rect 21 207 37 241
rect 71 207 87 241
rect 121 281 201 286
rect 121 247 151 281
rect 185 247 201 281
rect 121 225 201 247
rect 247 270 259 304
rect 247 254 293 270
rect 247 173 281 254
rect 327 218 363 388
rect 397 607 453 649
rect 397 573 403 607
rect 437 573 453 607
rect 397 507 453 573
rect 397 473 403 507
rect 437 473 453 507
rect 397 413 453 473
rect 397 379 403 413
rect 437 379 453 413
rect 397 363 453 379
rect 38 139 281 173
rect 315 202 363 218
rect 315 168 317 202
rect 351 168 363 202
rect 38 106 104 139
rect 38 72 54 106
rect 88 72 104 106
rect 38 56 104 72
rect 206 97 272 105
rect 206 63 222 97
rect 256 63 272 97
rect 206 17 272 63
rect 315 101 363 168
rect 315 67 317 101
rect 351 67 363 101
rect 315 51 363 67
rect 397 202 453 218
rect 397 168 403 202
rect 437 168 453 202
rect 397 93 453 168
rect 397 59 403 93
rect 437 59 453 93
rect 397 17 453 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and2_2
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3537652
string GDS_START 3532436
<< end >>
