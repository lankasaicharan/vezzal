magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 1 49 863 157
rect 0 0 864 49
<< scnmos >>
rect 84 47 114 131
rect 156 47 186 131
rect 246 47 276 131
rect 324 47 354 131
rect 402 47 432 131
rect 480 47 510 131
rect 678 47 708 131
rect 750 47 780 131
<< scpmoshvt >>
rect 94 409 144 609
rect 200 409 250 609
rect 306 409 356 609
rect 416 409 466 609
rect 522 409 572 609
rect 684 409 734 609
<< ndiff >>
rect 27 111 84 131
rect 27 77 39 111
rect 73 77 84 111
rect 27 47 84 77
rect 114 47 156 131
rect 186 106 246 131
rect 186 72 197 106
rect 231 72 246 106
rect 186 47 246 72
rect 276 47 324 131
rect 354 47 402 131
rect 432 47 480 131
rect 510 106 567 131
rect 510 72 521 106
rect 555 72 567 106
rect 510 47 567 72
rect 621 101 678 131
rect 621 67 633 101
rect 667 67 678 101
rect 621 47 678 67
rect 708 47 750 131
rect 780 111 837 131
rect 780 77 791 111
rect 825 77 837 111
rect 780 47 837 77
<< pdiff >>
rect 37 597 94 609
rect 37 563 49 597
rect 83 563 94 597
rect 37 514 94 563
rect 37 480 49 514
rect 83 480 94 514
rect 37 409 94 480
rect 144 597 200 609
rect 144 563 155 597
rect 189 563 200 597
rect 144 514 200 563
rect 144 480 155 514
rect 189 480 200 514
rect 144 409 200 480
rect 250 597 306 609
rect 250 563 261 597
rect 295 563 306 597
rect 250 526 306 563
rect 250 492 261 526
rect 295 492 306 526
rect 250 455 306 492
rect 250 421 261 455
rect 295 421 306 455
rect 250 409 306 421
rect 356 597 416 609
rect 356 563 367 597
rect 401 563 416 597
rect 356 514 416 563
rect 356 480 367 514
rect 401 480 416 514
rect 356 409 416 480
rect 466 597 522 609
rect 466 563 477 597
rect 511 563 522 597
rect 466 526 522 563
rect 466 492 477 526
rect 511 492 522 526
rect 466 455 522 492
rect 466 421 477 455
rect 511 421 522 455
rect 466 409 522 421
rect 572 597 684 609
rect 572 563 591 597
rect 625 563 684 597
rect 572 526 684 563
rect 572 492 591 526
rect 625 492 684 526
rect 572 455 684 492
rect 572 421 591 455
rect 625 421 684 455
rect 572 409 684 421
rect 734 597 791 609
rect 734 563 745 597
rect 779 563 791 597
rect 734 526 791 563
rect 734 492 745 526
rect 779 492 791 526
rect 734 455 791 492
rect 734 421 745 455
rect 779 421 791 455
rect 734 409 791 421
<< ndiffc >>
rect 39 77 73 111
rect 197 72 231 106
rect 521 72 555 106
rect 633 67 667 101
rect 791 77 825 111
<< pdiffc >>
rect 49 563 83 597
rect 49 480 83 514
rect 155 563 189 597
rect 155 480 189 514
rect 261 563 295 597
rect 261 492 295 526
rect 261 421 295 455
rect 367 563 401 597
rect 367 480 401 514
rect 477 563 511 597
rect 477 492 511 526
rect 477 421 511 455
rect 591 563 625 597
rect 591 492 625 526
rect 591 421 625 455
rect 745 563 779 597
rect 745 492 779 526
rect 745 421 779 455
<< poly >>
rect 94 609 144 635
rect 200 609 250 635
rect 306 609 356 635
rect 416 609 466 635
rect 522 609 572 635
rect 684 609 734 635
rect 94 367 144 409
rect 84 351 150 367
rect 200 358 250 409
rect 306 358 356 409
rect 416 358 466 409
rect 84 317 100 351
rect 134 317 150 351
rect 84 283 150 317
rect 84 249 100 283
rect 134 249 150 283
rect 84 233 150 249
rect 192 342 258 358
rect 192 308 208 342
rect 242 308 258 342
rect 192 274 258 308
rect 192 240 208 274
rect 242 240 258 274
rect 84 176 114 233
rect 192 224 258 240
rect 300 342 366 358
rect 300 308 316 342
rect 350 308 366 342
rect 300 274 366 308
rect 300 240 316 274
rect 350 240 366 274
rect 300 224 366 240
rect 408 342 474 358
rect 408 308 424 342
rect 458 308 474 342
rect 522 339 572 409
rect 408 274 474 308
rect 408 240 424 274
rect 458 240 474 274
rect 408 224 474 240
rect 542 323 636 339
rect 542 289 586 323
rect 620 289 636 323
rect 228 176 258 224
rect 84 146 186 176
rect 228 146 276 176
rect 84 131 114 146
rect 156 131 186 146
rect 246 131 276 146
rect 324 131 354 224
rect 408 176 438 224
rect 542 176 636 289
rect 684 237 734 409
rect 402 146 438 176
rect 480 146 636 176
rect 678 221 780 237
rect 678 187 720 221
rect 754 187 780 221
rect 678 171 780 187
rect 402 131 432 146
rect 480 131 510 146
rect 678 131 708 171
rect 750 131 780 171
rect 84 21 114 47
rect 156 21 186 47
rect 246 21 276 47
rect 324 21 354 47
rect 402 21 432 47
rect 480 21 510 47
rect 678 21 708 47
rect 750 21 780 47
<< polycont >>
rect 100 317 134 351
rect 100 249 134 283
rect 208 308 242 342
rect 208 240 242 274
rect 316 308 350 342
rect 316 240 350 274
rect 424 308 458 342
rect 424 240 458 274
rect 586 289 620 323
rect 720 187 754 221
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 18 597 99 613
rect 18 563 49 597
rect 83 563 99 597
rect 18 514 99 563
rect 18 480 49 514
rect 83 480 99 514
rect 18 464 99 480
rect 139 597 205 649
rect 139 563 155 597
rect 189 563 205 597
rect 139 514 205 563
rect 139 480 155 514
rect 189 480 205 514
rect 139 464 205 480
rect 245 597 311 613
rect 245 563 261 597
rect 295 563 311 597
rect 245 526 311 563
rect 245 492 261 526
rect 295 492 311 526
rect 18 135 52 464
rect 245 455 311 492
rect 351 597 417 649
rect 351 563 367 597
rect 401 563 417 597
rect 351 514 417 563
rect 351 480 367 514
rect 401 480 417 514
rect 351 464 417 480
rect 461 597 539 613
rect 461 563 477 597
rect 511 563 539 597
rect 461 526 539 563
rect 461 492 477 526
rect 511 492 539 526
rect 245 428 261 455
rect 88 421 261 428
rect 295 428 311 455
rect 461 455 539 492
rect 461 428 477 455
rect 295 421 477 428
rect 511 421 539 455
rect 88 394 539 421
rect 575 597 641 649
rect 575 563 591 597
rect 625 563 641 597
rect 575 526 641 563
rect 575 492 591 526
rect 625 492 641 526
rect 575 455 641 492
rect 575 421 591 455
rect 625 421 641 455
rect 575 405 641 421
rect 729 597 795 613
rect 729 563 745 597
rect 779 563 795 597
rect 729 526 795 563
rect 729 492 745 526
rect 779 492 795 526
rect 729 455 795 492
rect 729 421 745 455
rect 779 421 795 455
rect 88 351 150 394
rect 88 317 100 351
rect 134 317 150 351
rect 88 283 150 317
rect 88 249 100 283
rect 134 249 150 283
rect 88 233 150 249
rect 192 342 263 358
rect 192 308 208 342
rect 242 308 263 342
rect 192 274 263 308
rect 192 240 208 274
rect 242 240 263 274
rect 192 224 263 240
rect 300 342 366 358
rect 300 308 316 342
rect 350 308 366 342
rect 300 274 366 308
rect 300 240 316 274
rect 350 240 366 274
rect 18 111 89 135
rect 18 77 39 111
rect 73 77 89 111
rect 18 53 89 77
rect 181 106 247 135
rect 181 72 197 106
rect 231 72 247 106
rect 300 88 366 240
rect 408 342 469 358
rect 408 308 424 342
rect 458 308 469 342
rect 408 274 469 308
rect 408 240 424 274
rect 458 240 469 274
rect 408 88 469 240
rect 505 126 539 394
rect 729 339 795 421
rect 575 323 795 339
rect 575 289 586 323
rect 620 307 795 323
rect 620 289 841 307
rect 575 273 841 289
rect 601 221 770 237
rect 601 187 720 221
rect 754 187 770 221
rect 601 171 770 187
rect 601 162 647 171
rect 807 135 841 273
rect 505 106 571 126
rect 181 17 247 72
rect 505 72 521 106
rect 555 72 571 106
rect 505 53 571 72
rect 617 101 683 126
rect 617 67 633 101
rect 667 67 683 101
rect 617 17 683 67
rect 775 111 841 135
rect 775 77 791 111
rect 825 77 841 111
rect 775 53 841 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4b_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5354008
string GDS_START 5345824
<< end >>
