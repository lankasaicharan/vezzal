magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2402 1852
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1082 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 287 47 317 177
rect 381 47 411 177
rect 475 47 505 177
rect 569 47 599 177
rect 656 47 686 177
rect 750 47 780 177
rect 844 47 874 177
rect 948 47 978 177
<< scpmoshvt >>
rect 81 297 117 497
rect 279 297 315 497
rect 373 297 409 497
rect 467 297 503 497
rect 561 297 597 497
rect 658 297 694 497
rect 752 297 788 497
rect 846 297 882 497
rect 940 297 976 497
<< ndiff >>
rect 27 161 89 177
rect 27 127 35 161
rect 69 127 89 161
rect 27 93 89 127
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 93 171 177
rect 119 59 129 93
rect 163 59 171 93
rect 119 47 171 59
rect 225 161 287 177
rect 225 127 233 161
rect 267 127 287 161
rect 225 93 287 127
rect 225 59 233 93
rect 267 59 287 93
rect 225 47 287 59
rect 317 161 381 177
rect 317 127 327 161
rect 361 127 381 161
rect 317 47 381 127
rect 411 93 475 177
rect 411 59 421 93
rect 455 59 475 93
rect 411 47 475 59
rect 505 161 569 177
rect 505 127 515 161
rect 549 127 569 161
rect 505 47 569 127
rect 599 161 656 177
rect 599 127 612 161
rect 646 127 656 161
rect 599 93 656 127
rect 599 59 612 93
rect 646 59 656 93
rect 599 47 656 59
rect 686 93 750 177
rect 686 59 706 93
rect 740 59 750 93
rect 686 47 750 59
rect 780 161 844 177
rect 780 127 800 161
rect 834 127 844 161
rect 780 93 844 127
rect 780 59 800 93
rect 834 59 844 93
rect 780 47 844 59
rect 874 93 948 177
rect 874 59 894 93
rect 928 59 948 93
rect 874 47 948 59
rect 978 161 1056 177
rect 978 127 1010 161
rect 1044 127 1056 161
rect 978 93 1056 127
rect 978 59 1010 93
rect 1044 59 1056 93
rect 978 47 1056 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 171 497
rect 117 451 129 485
rect 163 451 171 485
rect 117 417 171 451
rect 117 383 129 417
rect 163 383 171 417
rect 117 297 171 383
rect 225 485 279 497
rect 225 451 233 485
rect 267 451 279 485
rect 225 417 279 451
rect 225 383 233 417
rect 267 383 279 417
rect 225 349 279 383
rect 225 315 233 349
rect 267 315 279 349
rect 225 297 279 315
rect 315 485 373 497
rect 315 451 327 485
rect 361 451 373 485
rect 315 417 373 451
rect 315 383 327 417
rect 361 383 373 417
rect 315 349 373 383
rect 315 315 327 349
rect 361 315 373 349
rect 315 297 373 315
rect 409 485 467 497
rect 409 451 421 485
rect 455 451 467 485
rect 409 417 467 451
rect 409 383 421 417
rect 455 383 467 417
rect 409 297 467 383
rect 503 485 561 497
rect 503 451 515 485
rect 549 451 561 485
rect 503 417 561 451
rect 503 383 515 417
rect 549 383 561 417
rect 503 349 561 383
rect 503 315 515 349
rect 549 315 561 349
rect 503 297 561 315
rect 597 485 658 497
rect 597 451 612 485
rect 646 451 658 485
rect 597 417 658 451
rect 597 383 612 417
rect 646 383 658 417
rect 597 297 658 383
rect 694 485 752 497
rect 694 451 706 485
rect 740 451 752 485
rect 694 417 752 451
rect 694 383 706 417
rect 740 383 752 417
rect 694 349 752 383
rect 694 315 706 349
rect 740 315 752 349
rect 694 297 752 315
rect 788 485 846 497
rect 788 451 800 485
rect 834 451 846 485
rect 788 417 846 451
rect 788 383 800 417
rect 834 383 846 417
rect 788 297 846 383
rect 882 485 940 497
rect 882 451 894 485
rect 928 451 940 485
rect 882 417 940 451
rect 882 383 894 417
rect 928 383 940 417
rect 882 349 940 383
rect 882 315 894 349
rect 928 315 940 349
rect 882 297 940 315
rect 976 485 1056 497
rect 976 451 1010 485
rect 1044 451 1056 485
rect 976 417 1056 451
rect 976 383 1010 417
rect 1044 383 1056 417
rect 976 349 1056 383
rect 976 315 1010 349
rect 1044 315 1056 349
rect 976 297 1056 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 59 163 93
rect 233 127 267 161
rect 233 59 267 93
rect 327 127 361 161
rect 421 59 455 93
rect 515 127 549 161
rect 612 127 646 161
rect 612 59 646 93
rect 706 59 740 93
rect 800 127 834 161
rect 800 59 834 93
rect 894 59 928 93
rect 1010 127 1044 161
rect 1010 59 1044 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 233 451 267 485
rect 233 383 267 417
rect 233 315 267 349
rect 327 451 361 485
rect 327 383 361 417
rect 327 315 361 349
rect 421 451 455 485
rect 421 383 455 417
rect 515 451 549 485
rect 515 383 549 417
rect 515 315 549 349
rect 612 451 646 485
rect 612 383 646 417
rect 706 451 740 485
rect 706 383 740 417
rect 706 315 740 349
rect 800 451 834 485
rect 800 383 834 417
rect 894 451 928 485
rect 894 383 928 417
rect 894 315 928 349
rect 1010 451 1044 485
rect 1010 383 1044 417
rect 1010 315 1044 349
<< poly >>
rect 81 497 117 523
rect 279 497 315 523
rect 373 497 409 523
rect 467 497 503 523
rect 561 497 597 523
rect 658 497 694 523
rect 752 497 788 523
rect 846 497 882 523
rect 940 497 976 523
rect 81 282 117 297
rect 279 282 315 297
rect 373 282 409 297
rect 467 282 503 297
rect 561 282 597 297
rect 658 282 694 297
rect 752 282 788 297
rect 846 282 882 297
rect 940 282 976 297
rect 79 261 119 282
rect 22 249 119 261
rect 277 259 317 282
rect 371 259 411 282
rect 465 259 505 282
rect 559 259 599 282
rect 22 215 38 249
rect 72 215 119 249
rect 22 203 119 215
rect 211 249 599 259
rect 211 215 227 249
rect 261 215 327 249
rect 361 215 421 249
rect 455 215 599 249
rect 211 205 599 215
rect 89 177 119 203
rect 287 177 317 205
rect 381 177 411 205
rect 475 177 505 205
rect 569 177 599 205
rect 656 259 696 282
rect 750 259 790 282
rect 844 259 884 282
rect 938 259 978 282
rect 656 249 1044 259
rect 656 215 707 249
rect 741 215 800 249
rect 834 215 893 249
rect 927 215 994 249
rect 1028 215 1044 249
rect 656 205 1044 215
rect 656 177 686 205
rect 750 177 780 205
rect 844 177 874 205
rect 948 177 978 205
rect 89 21 119 47
rect 287 21 317 47
rect 381 21 411 47
rect 475 21 505 47
rect 569 21 599 47
rect 656 21 686 47
rect 750 21 780 47
rect 844 21 874 47
rect 948 21 978 47
<< polycont >>
rect 38 215 72 249
rect 227 215 261 249
rect 327 215 361 249
rect 421 215 455 249
rect 707 215 741 249
rect 800 215 834 249
rect 893 215 927 249
rect 994 215 1028 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 18 485 85 493
rect 18 451 35 485
rect 69 451 85 485
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 18 349 85 383
rect 129 485 267 527
rect 163 451 233 485
rect 129 417 267 451
rect 163 383 233 417
rect 129 367 267 383
rect 18 315 35 349
rect 69 333 85 349
rect 204 349 267 367
rect 69 315 166 333
rect 18 289 166 315
rect 204 315 233 349
rect 204 289 267 315
rect 301 485 377 493
rect 301 451 327 485
rect 361 451 377 485
rect 301 417 377 451
rect 301 383 327 417
rect 361 383 377 417
rect 301 349 377 383
rect 421 485 455 527
rect 421 417 455 451
rect 421 367 455 383
rect 489 485 568 493
rect 489 451 515 485
rect 549 451 568 485
rect 489 417 568 451
rect 489 383 515 417
rect 549 383 568 417
rect 301 315 327 349
rect 361 333 377 349
rect 489 349 568 383
rect 612 485 646 527
rect 612 417 646 451
rect 612 367 646 383
rect 680 485 756 493
rect 680 451 706 485
rect 740 451 756 485
rect 680 417 756 451
rect 680 383 706 417
rect 740 383 756 417
rect 489 333 515 349
rect 361 315 515 333
rect 549 333 568 349
rect 680 349 756 383
rect 800 485 834 527
rect 800 417 834 451
rect 800 367 834 383
rect 868 485 944 493
rect 868 451 894 485
rect 928 451 944 485
rect 868 417 944 451
rect 868 383 894 417
rect 928 383 944 417
rect 680 333 706 349
rect 549 315 706 333
rect 740 333 756 349
rect 868 349 944 383
rect 868 333 894 349
rect 740 315 894 333
rect 928 315 944 349
rect 301 289 944 315
rect 994 485 1060 527
rect 994 451 1010 485
rect 1044 451 1060 485
rect 994 417 1060 451
rect 994 383 1010 417
rect 1044 383 1060 417
rect 994 349 1060 383
rect 994 315 1010 349
rect 1044 315 1060 349
rect 994 299 1060 315
rect 132 255 166 289
rect 22 249 88 255
rect 22 215 38 249
rect 72 215 88 249
rect 132 249 471 255
rect 132 215 227 249
rect 261 215 327 249
rect 361 215 421 249
rect 455 215 471 249
rect 132 181 166 215
rect 515 181 568 289
rect 681 249 1078 255
rect 681 215 707 249
rect 741 215 800 249
rect 834 215 893 249
rect 927 215 994 249
rect 1028 215 1078 249
rect 18 161 166 181
rect 18 127 35 161
rect 69 143 166 161
rect 217 161 267 181
rect 69 127 85 143
rect 18 93 85 127
rect 217 127 233 161
rect 301 161 568 181
rect 301 127 327 161
rect 361 127 515 161
rect 549 127 568 161
rect 612 161 1060 181
rect 646 143 800 161
rect 646 127 662 143
rect 18 59 35 93
rect 69 59 85 93
rect 18 51 85 59
rect 129 93 168 109
rect 163 59 168 93
rect 129 17 168 59
rect 217 93 267 127
rect 612 93 662 127
rect 774 127 800 143
rect 834 143 1010 161
rect 834 127 850 143
rect 217 59 233 93
rect 267 59 421 93
rect 455 59 612 93
rect 646 59 662 93
rect 217 51 662 59
rect 706 93 740 109
rect 706 17 740 59
rect 774 93 850 127
rect 994 127 1010 143
rect 1044 127 1060 161
rect 774 59 800 93
rect 834 59 850 93
rect 774 51 850 59
rect 894 93 942 109
rect 928 59 942 93
rect 894 17 942 59
rect 994 93 1060 127
rect 994 59 1010 93
rect 1044 59 1060 93
rect 994 51 1060 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 681 215 1078 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 949 238 949 238 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel locali s 858 221 892 255 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel locali s 695 238 695 238 0 FreeSans 250 0 0 0 B
port 2 nsew
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel locali s 868 333 944 493 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 548 377 548 377 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel locali s 548 445 548 445 0 FreeSans 250 0 0 0 Y
port 7 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2b_4
rlabel locali s 680 333 756 493 1 Y
port 7 nsew signal output
rlabel locali s 515 181 568 289 1 Y
port 7 nsew signal output
rlabel locali s 489 333 568 493 1 Y
port 7 nsew signal output
rlabel locali s 301 333 377 493 1 Y
port 7 nsew signal output
rlabel locali s 301 289 944 333 1 Y
port 7 nsew signal output
rlabel locali s 301 127 568 181 1 Y
port 7 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2223138
string GDS_START 2213762
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
