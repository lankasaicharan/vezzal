magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 54 49 652 167
rect 0 0 672 49
<< scnmos >>
rect 137 57 167 141
rect 215 57 245 141
rect 317 57 347 141
rect 431 57 461 141
rect 539 57 569 141
<< scpmoshvt >>
rect 111 409 161 609
rect 217 409 267 609
rect 327 409 377 609
rect 433 409 483 609
rect 533 409 583 609
<< ndiff >>
rect 80 116 137 141
rect 80 82 92 116
rect 126 82 137 116
rect 80 57 137 82
rect 167 57 215 141
rect 245 57 317 141
rect 347 116 431 141
rect 347 82 376 116
rect 410 82 431 116
rect 347 57 431 82
rect 461 103 539 141
rect 461 69 478 103
rect 512 69 539 103
rect 461 57 539 69
rect 569 116 626 141
rect 569 82 580 116
rect 614 82 626 116
rect 569 57 626 82
<< pdiff >>
rect 54 597 111 609
rect 54 563 66 597
rect 100 563 111 597
rect 54 473 111 563
rect 54 439 66 473
rect 100 439 111 473
rect 54 409 111 439
rect 161 597 217 609
rect 161 563 172 597
rect 206 563 217 597
rect 161 526 217 563
rect 161 492 172 526
rect 206 492 217 526
rect 161 455 217 492
rect 161 421 172 455
rect 206 421 217 455
rect 161 409 217 421
rect 267 597 327 609
rect 267 563 278 597
rect 312 563 327 597
rect 267 515 327 563
rect 267 481 278 515
rect 312 481 327 515
rect 267 409 327 481
rect 377 597 433 609
rect 377 563 388 597
rect 422 563 433 597
rect 377 526 433 563
rect 377 492 388 526
rect 422 492 433 526
rect 377 455 433 492
rect 377 421 388 455
rect 422 421 433 455
rect 377 409 433 421
rect 483 409 533 609
rect 583 597 640 609
rect 583 563 594 597
rect 628 563 640 597
rect 583 526 640 563
rect 583 492 594 526
rect 628 492 640 526
rect 583 455 640 492
rect 583 421 594 455
rect 628 421 640 455
rect 583 409 640 421
<< ndiffc >>
rect 92 82 126 116
rect 376 82 410 116
rect 478 69 512 103
rect 580 82 614 116
<< pdiffc >>
rect 66 563 100 597
rect 66 439 100 473
rect 172 563 206 597
rect 172 492 206 526
rect 172 421 206 455
rect 278 563 312 597
rect 278 481 312 515
rect 388 563 422 597
rect 388 492 422 526
rect 388 421 422 455
rect 594 563 628 597
rect 594 492 628 526
rect 594 421 628 455
<< poly >>
rect 111 609 161 635
rect 217 609 267 635
rect 327 609 377 635
rect 433 609 483 635
rect 533 609 583 635
rect 111 315 161 409
rect 217 317 267 409
rect 327 359 377 409
rect 433 359 483 409
rect 317 343 383 359
rect 101 299 167 315
rect 101 265 117 299
rect 151 265 167 299
rect 101 231 167 265
rect 101 197 117 231
rect 151 197 167 231
rect 101 181 167 197
rect 209 301 275 317
rect 209 267 225 301
rect 259 267 275 301
rect 209 233 275 267
rect 209 199 225 233
rect 259 199 275 233
rect 209 183 275 199
rect 317 309 333 343
rect 367 309 383 343
rect 317 275 383 309
rect 317 241 333 275
rect 367 241 383 275
rect 317 225 383 241
rect 425 343 491 359
rect 425 309 441 343
rect 475 309 491 343
rect 425 275 491 309
rect 425 241 441 275
rect 475 241 491 275
rect 425 225 491 241
rect 533 302 583 409
rect 533 286 651 302
rect 533 252 601 286
rect 635 252 651 286
rect 533 236 651 252
rect 137 141 167 181
rect 215 141 245 183
rect 317 141 347 225
rect 431 141 461 225
rect 539 141 569 236
rect 137 31 167 57
rect 215 31 245 57
rect 317 31 347 57
rect 431 31 461 57
rect 539 31 569 57
<< polycont >>
rect 117 265 151 299
rect 117 197 151 231
rect 225 267 259 301
rect 225 199 259 233
rect 333 309 367 343
rect 333 241 367 275
rect 441 309 475 343
rect 441 241 475 275
rect 601 252 635 286
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 50 597 116 649
rect 50 563 66 597
rect 100 563 116 597
rect 50 473 116 563
rect 50 439 66 473
rect 100 439 116 473
rect 50 423 116 439
rect 156 597 222 613
rect 156 563 172 597
rect 206 563 222 597
rect 156 526 222 563
rect 156 492 172 526
rect 206 492 222 526
rect 156 455 222 492
rect 262 597 328 649
rect 262 563 278 597
rect 312 563 328 597
rect 262 515 328 563
rect 262 481 278 515
rect 312 481 328 515
rect 262 465 328 481
rect 372 597 438 613
rect 372 563 388 597
rect 422 563 438 597
rect 372 526 438 563
rect 372 492 388 526
rect 422 492 438 526
rect 156 421 172 455
rect 206 429 222 455
rect 372 455 438 492
rect 372 429 388 455
rect 206 421 388 429
rect 422 421 438 455
rect 156 395 438 421
rect 578 597 644 649
rect 578 563 594 597
rect 628 563 644 597
rect 578 526 644 563
rect 578 492 594 526
rect 628 492 644 526
rect 578 455 644 492
rect 578 421 594 455
rect 628 421 644 455
rect 578 405 644 421
rect 156 387 222 395
rect 25 353 222 387
rect 25 145 67 353
rect 313 343 381 359
rect 103 299 167 315
rect 103 265 117 299
rect 151 265 167 299
rect 103 231 167 265
rect 103 197 117 231
rect 151 197 167 231
rect 103 181 167 197
rect 209 301 275 317
rect 209 267 225 301
rect 259 267 275 301
rect 209 233 275 267
rect 209 199 225 233
rect 259 199 275 233
rect 313 309 333 343
rect 367 309 381 343
rect 313 275 381 309
rect 313 241 333 275
rect 367 241 381 275
rect 313 225 381 241
rect 425 343 549 359
rect 425 309 441 343
rect 475 309 549 343
rect 425 275 549 309
rect 425 241 441 275
rect 475 241 549 275
rect 425 225 549 241
rect 585 286 651 356
rect 585 252 601 286
rect 635 252 651 286
rect 585 236 651 252
rect 25 116 142 145
rect 25 82 92 116
rect 126 82 142 116
rect 209 88 275 199
rect 360 155 630 189
rect 360 116 426 155
rect 25 53 142 82
rect 360 82 376 116
rect 410 82 426 116
rect 360 53 426 82
rect 462 103 528 119
rect 462 69 478 103
rect 512 69 528 103
rect 462 17 528 69
rect 564 116 630 155
rect 564 82 580 116
rect 614 82 630 116
rect 564 53 630 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2111ai_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4709982
string GDS_START 4702778
<< end >>
