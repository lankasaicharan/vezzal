magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3602 1975
<< nwell >>
rect -38 332 2342 704
rect 250 329 1007 332
<< pwell >>
rect 363 274 784 287
rect 1 248 784 274
rect 1 228 1053 248
rect 1536 228 2303 248
rect 1 49 2303 228
rect 0 0 2304 49
<< scpmos >>
rect 91 368 127 592
rect 208 368 244 568
rect 336 365 372 533
rect 450 365 486 533
rect 540 365 576 533
rect 662 365 698 533
rect 869 365 905 589
rect 990 389 1026 589
rect 1097 421 1133 589
rect 1228 421 1264 589
rect 1472 392 1508 592
rect 1573 368 1609 592
rect 1792 368 1828 536
rect 1882 368 1918 536
rect 2084 392 2120 592
rect 2185 368 2221 592
<< nmoslvt >>
rect 84 100 114 248
rect 258 120 288 248
rect 344 120 374 248
rect 462 133 492 261
rect 550 133 580 261
rect 671 133 701 261
rect 947 74 977 222
rect 1042 74 1072 202
rect 1228 74 1258 202
rect 1370 74 1400 202
rect 1510 74 1540 202
rect 1612 74 1642 222
rect 1714 94 1744 222
rect 1876 94 1906 222
rect 2008 94 2038 222
rect 2190 74 2220 222
<< ndiff >>
rect 389 248 462 261
rect 27 220 84 248
rect 27 186 39 220
rect 73 186 84 220
rect 27 146 84 186
rect 27 112 39 146
rect 73 112 84 146
rect 27 100 84 112
rect 114 146 258 248
rect 114 112 128 146
rect 162 120 258 146
rect 288 237 344 248
rect 288 203 299 237
rect 333 203 344 237
rect 288 169 344 203
rect 288 135 299 169
rect 333 135 344 169
rect 288 120 344 135
rect 374 244 462 248
rect 374 210 401 244
rect 435 210 462 244
rect 374 169 462 210
rect 374 135 401 169
rect 435 135 462 169
rect 374 133 462 135
rect 492 247 550 261
rect 492 213 505 247
rect 539 213 550 247
rect 492 179 550 213
rect 492 145 505 179
rect 539 145 550 179
rect 492 133 550 145
rect 580 247 671 261
rect 580 213 605 247
rect 639 213 671 247
rect 580 179 671 213
rect 580 145 605 179
rect 639 145 671 179
rect 580 133 671 145
rect 701 249 758 261
rect 701 215 712 249
rect 746 215 758 249
rect 701 179 758 215
rect 701 145 712 179
rect 746 145 758 179
rect 701 133 758 145
rect 821 196 947 222
rect 821 162 897 196
rect 931 162 947 196
rect 374 120 447 133
rect 162 112 177 120
rect 114 100 177 112
rect 821 120 947 162
rect 821 86 829 120
rect 863 86 902 120
rect 936 86 947 120
rect 821 74 947 86
rect 977 202 1027 222
rect 1562 202 1612 222
rect 977 148 1042 202
rect 977 114 997 148
rect 1031 114 1042 148
rect 977 74 1042 114
rect 1072 128 1228 202
rect 1072 94 1083 128
rect 1117 94 1180 128
rect 1214 94 1228 128
rect 1072 74 1228 94
rect 1258 190 1370 202
rect 1258 156 1280 190
rect 1314 156 1370 190
rect 1258 120 1370 156
rect 1258 86 1280 120
rect 1314 86 1370 120
rect 1258 74 1370 86
rect 1400 188 1510 202
rect 1400 154 1465 188
rect 1499 154 1510 188
rect 1400 120 1510 154
rect 1400 86 1465 120
rect 1499 86 1510 120
rect 1400 74 1510 86
rect 1540 186 1612 202
rect 1540 152 1565 186
rect 1599 152 1612 186
rect 1540 116 1612 152
rect 1540 82 1565 116
rect 1599 82 1612 116
rect 1540 74 1612 82
rect 1642 210 1714 222
rect 1642 176 1653 210
rect 1687 176 1714 210
rect 1642 120 1714 176
rect 1642 86 1653 120
rect 1687 94 1714 120
rect 1744 210 1876 222
rect 1744 176 1771 210
rect 1805 176 1876 210
rect 1744 140 1876 176
rect 1744 106 1771 140
rect 1805 106 1876 140
rect 1744 94 1876 106
rect 1906 185 2008 222
rect 1906 151 1963 185
rect 1997 151 2008 185
rect 1906 94 2008 151
rect 2038 94 2190 222
rect 1687 86 1699 94
rect 1642 74 1699 86
rect 2103 82 2190 94
rect 2103 48 2122 82
rect 2156 74 2190 82
rect 2220 210 2277 222
rect 2220 176 2231 210
rect 2265 176 2277 210
rect 2220 120 2277 176
rect 2220 86 2231 120
rect 2265 86 2277 120
rect 2220 74 2277 86
rect 2156 48 2175 74
rect 2103 36 2175 48
<< pdiff >>
rect 35 580 91 592
rect 35 546 47 580
rect 81 546 91 580
rect 35 510 91 546
rect 35 476 47 510
rect 81 476 91 510
rect 35 440 91 476
rect 35 406 47 440
rect 81 406 91 440
rect 35 368 91 406
rect 127 580 193 592
rect 127 546 147 580
rect 181 568 193 580
rect 181 546 208 568
rect 127 510 208 546
rect 127 476 147 510
rect 181 476 208 510
rect 127 440 208 476
rect 127 406 147 440
rect 181 406 208 440
rect 127 368 208 406
rect 244 556 300 568
rect 244 522 254 556
rect 288 533 300 556
rect 591 547 647 559
rect 591 533 602 547
rect 288 522 336 533
rect 244 488 336 522
rect 244 454 254 488
rect 288 454 336 488
rect 244 420 336 454
rect 244 386 254 420
rect 288 386 336 420
rect 244 368 336 386
rect 286 365 336 368
rect 372 456 450 533
rect 372 422 406 456
rect 440 422 450 456
rect 372 365 450 422
rect 486 411 540 533
rect 486 377 496 411
rect 530 377 540 411
rect 486 365 540 377
rect 576 513 602 533
rect 636 533 647 547
rect 636 513 662 533
rect 576 365 662 513
rect 698 521 753 533
rect 698 487 708 521
rect 742 487 753 521
rect 698 411 753 487
rect 698 377 708 411
rect 742 377 753 411
rect 698 365 753 377
rect 1422 589 1472 592
rect 813 577 869 589
rect 813 543 825 577
rect 859 543 869 577
rect 813 494 869 543
rect 813 460 825 494
rect 859 460 869 494
rect 813 411 869 460
rect 813 377 825 411
rect 859 377 869 411
rect 813 365 869 377
rect 905 577 990 589
rect 905 543 925 577
rect 959 543 990 577
rect 905 494 990 543
rect 905 460 925 494
rect 959 460 990 494
rect 905 411 990 460
rect 905 377 925 411
rect 959 389 990 411
rect 1026 577 1097 589
rect 1026 543 1036 577
rect 1070 543 1097 577
rect 1026 509 1097 543
rect 1026 475 1036 509
rect 1070 475 1097 509
rect 1026 441 1097 475
rect 1026 407 1036 441
rect 1070 421 1097 441
rect 1133 577 1228 589
rect 1133 543 1174 577
rect 1208 543 1228 577
rect 1133 467 1228 543
rect 1133 433 1174 467
rect 1208 433 1228 467
rect 1133 421 1228 433
rect 1264 577 1472 589
rect 1264 543 1274 577
rect 1308 543 1351 577
rect 1385 543 1428 577
rect 1462 543 1472 577
rect 1264 467 1472 543
rect 1264 433 1274 467
rect 1308 433 1351 467
rect 1385 433 1428 467
rect 1462 433 1472 467
rect 1264 421 1472 433
rect 1070 407 1082 421
rect 1026 389 1082 407
rect 959 377 971 389
rect 905 365 971 377
rect 1422 392 1472 421
rect 1508 580 1573 592
rect 1508 546 1529 580
rect 1563 546 1573 580
rect 1508 509 1573 546
rect 1508 475 1529 509
rect 1563 475 1573 509
rect 1508 438 1573 475
rect 1508 404 1529 438
rect 1563 404 1573 438
rect 1508 392 1573 404
rect 1523 368 1573 392
rect 1609 580 1665 592
rect 1609 546 1619 580
rect 1653 546 1665 580
rect 1609 497 1665 546
rect 1609 463 1619 497
rect 1653 463 1665 497
rect 1609 414 1665 463
rect 1609 380 1619 414
rect 1653 380 1665 414
rect 1609 368 1665 380
rect 1719 582 1777 594
rect 1719 548 1731 582
rect 1765 548 1777 582
rect 2028 580 2084 592
rect 1719 536 1777 548
rect 2028 546 2040 580
rect 2074 546 2084 580
rect 1719 368 1792 536
rect 1828 414 1882 536
rect 1828 380 1838 414
rect 1872 380 1882 414
rect 1828 368 1882 380
rect 1918 524 1974 536
rect 1918 490 1928 524
rect 1962 490 1974 524
rect 1918 414 1974 490
rect 1918 380 1928 414
rect 1962 380 1974 414
rect 2028 509 2084 546
rect 2028 475 2040 509
rect 2074 475 2084 509
rect 2028 438 2084 475
rect 2028 404 2040 438
rect 2074 404 2084 438
rect 2028 392 2084 404
rect 2120 580 2185 592
rect 2120 546 2130 580
rect 2164 546 2185 580
rect 2120 470 2185 546
rect 2120 436 2130 470
rect 2164 436 2185 470
rect 2120 392 2185 436
rect 1918 368 1974 380
rect 2135 368 2185 392
rect 2221 580 2277 592
rect 2221 546 2231 580
rect 2265 546 2277 580
rect 2221 497 2277 546
rect 2221 463 2231 497
rect 2265 463 2277 497
rect 2221 414 2277 463
rect 2221 380 2231 414
rect 2265 380 2277 414
rect 2221 368 2277 380
<< ndiffc >>
rect 39 186 73 220
rect 39 112 73 146
rect 128 112 162 146
rect 299 203 333 237
rect 299 135 333 169
rect 401 210 435 244
rect 401 135 435 169
rect 505 213 539 247
rect 505 145 539 179
rect 605 213 639 247
rect 605 145 639 179
rect 712 215 746 249
rect 712 145 746 179
rect 897 162 931 196
rect 829 86 863 120
rect 902 86 936 120
rect 997 114 1031 148
rect 1083 94 1117 128
rect 1180 94 1214 128
rect 1280 156 1314 190
rect 1280 86 1314 120
rect 1465 154 1499 188
rect 1465 86 1499 120
rect 1565 152 1599 186
rect 1565 82 1599 116
rect 1653 176 1687 210
rect 1653 86 1687 120
rect 1771 176 1805 210
rect 1771 106 1805 140
rect 1963 151 1997 185
rect 2122 48 2156 82
rect 2231 176 2265 210
rect 2231 86 2265 120
<< pdiffc >>
rect 47 546 81 580
rect 47 476 81 510
rect 47 406 81 440
rect 147 546 181 580
rect 147 476 181 510
rect 147 406 181 440
rect 254 522 288 556
rect 254 454 288 488
rect 254 386 288 420
rect 406 422 440 456
rect 496 377 530 411
rect 602 513 636 547
rect 708 487 742 521
rect 708 377 742 411
rect 825 543 859 577
rect 825 460 859 494
rect 825 377 859 411
rect 925 543 959 577
rect 925 460 959 494
rect 925 377 959 411
rect 1036 543 1070 577
rect 1036 475 1070 509
rect 1036 407 1070 441
rect 1174 543 1208 577
rect 1174 433 1208 467
rect 1274 543 1308 577
rect 1351 543 1385 577
rect 1428 543 1462 577
rect 1274 433 1308 467
rect 1351 433 1385 467
rect 1428 433 1462 467
rect 1529 546 1563 580
rect 1529 475 1563 509
rect 1529 404 1563 438
rect 1619 546 1653 580
rect 1619 463 1653 497
rect 1619 380 1653 414
rect 1731 548 1765 582
rect 2040 546 2074 580
rect 1838 380 1872 414
rect 1928 490 1962 524
rect 1928 380 1962 414
rect 2040 475 2074 509
rect 2040 404 2074 438
rect 2130 546 2164 580
rect 2130 436 2164 470
rect 2231 546 2265 580
rect 2231 463 2265 497
rect 2231 380 2265 414
<< poly >>
rect 91 592 127 618
rect 450 607 798 637
rect 208 568 244 594
rect 336 533 372 559
rect 450 533 486 607
rect 540 533 576 559
rect 91 336 127 368
rect 208 336 244 368
rect 662 533 698 607
rect 75 320 141 336
rect 75 286 91 320
rect 125 286 141 320
rect 75 270 141 286
rect 183 320 288 336
rect 183 286 199 320
rect 233 286 288 320
rect 183 270 288 286
rect 84 248 114 270
rect 258 248 288 270
rect 336 293 372 365
rect 450 323 486 365
rect 450 293 492 323
rect 336 263 374 293
rect 344 248 374 263
rect 462 261 492 293
rect 540 306 576 365
rect 662 350 698 365
rect 662 320 701 350
rect 540 276 580 306
rect 550 261 580 276
rect 671 261 701 320
rect 768 310 798 607
rect 869 589 905 615
rect 990 589 1026 615
rect 1097 589 1133 615
rect 1228 589 1264 615
rect 1472 592 1508 618
rect 1573 592 1609 618
rect 869 310 905 365
rect 990 310 1026 389
rect 1097 361 1133 421
rect 1228 376 1264 421
rect 1097 345 1180 361
rect 1097 331 1130 345
rect 768 294 1026 310
rect 1114 311 1130 331
rect 1164 311 1180 345
rect 1114 295 1180 311
rect 1228 360 1322 376
rect 1228 326 1272 360
rect 1306 326 1322 360
rect 1228 310 1322 326
rect 1364 344 1430 360
rect 1364 310 1380 344
rect 1414 310 1430 344
rect 768 280 963 294
rect 947 260 963 280
rect 997 274 1026 294
rect 997 260 1072 274
rect 947 244 1072 260
rect 947 222 977 244
rect 84 74 114 100
rect 258 94 288 120
rect 344 59 374 120
rect 462 107 492 133
rect 550 111 580 133
rect 550 95 623 111
rect 671 107 701 133
rect 550 61 573 95
rect 607 61 623 95
rect 1042 202 1072 244
rect 1228 202 1258 310
rect 1364 276 1430 310
rect 1472 358 1508 392
rect 2084 592 2120 618
rect 2185 592 2221 618
rect 1792 536 1828 562
rect 1882 536 1918 562
rect 1472 310 1502 358
rect 1573 322 1609 368
rect 1792 326 1828 368
rect 1573 310 1603 322
rect 1472 294 1603 310
rect 1472 280 1551 294
rect 1364 242 1380 276
rect 1414 242 1430 276
rect 1364 226 1430 242
rect 1510 260 1551 280
rect 1585 274 1603 294
rect 1695 310 1828 326
rect 1882 318 1918 368
rect 2084 318 2120 392
rect 2185 326 2221 368
rect 1695 276 1711 310
rect 1745 296 1828 310
rect 1876 302 1949 318
rect 1745 276 1761 296
rect 1585 260 1642 274
rect 1695 260 1761 276
rect 1876 268 1899 302
rect 1933 268 1949 302
rect 1510 244 1642 260
rect 1370 202 1400 226
rect 1510 202 1540 244
rect 1612 222 1642 244
rect 1714 222 1744 260
rect 1876 252 1949 268
rect 1991 302 2120 318
rect 1991 268 2007 302
rect 2041 288 2120 302
rect 2162 310 2228 326
rect 2041 268 2057 288
rect 1991 252 2057 268
rect 2162 276 2178 310
rect 2212 276 2228 310
rect 2162 260 2228 276
rect 1876 222 1906 252
rect 2008 222 2038 252
rect 2190 222 2220 260
rect 550 59 623 61
rect 344 29 623 59
rect 947 48 977 74
rect 1042 48 1072 74
rect 1228 48 1258 74
rect 1370 48 1400 74
rect 1510 48 1540 74
rect 1612 48 1642 74
rect 1714 68 1744 94
rect 1876 68 1906 94
rect 2008 68 2038 94
rect 2190 48 2220 74
<< polycont >>
rect 91 286 125 320
rect 199 286 233 320
rect 1130 311 1164 345
rect 1272 326 1306 360
rect 1380 310 1414 344
rect 963 260 997 294
rect 573 61 607 95
rect 1380 242 1414 276
rect 1551 260 1585 294
rect 1711 276 1745 310
rect 1899 268 1933 302
rect 2007 268 2041 302
rect 2178 276 2212 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 17 580 97 596
rect 17 546 47 580
rect 81 546 97 580
rect 17 510 97 546
rect 17 476 47 510
rect 81 476 97 510
rect 17 440 97 476
rect 17 406 47 440
rect 81 406 97 440
rect 17 390 97 406
rect 131 580 197 649
rect 131 546 147 580
rect 181 546 197 580
rect 131 510 197 546
rect 131 476 147 510
rect 181 476 197 510
rect 131 440 197 476
rect 131 406 147 440
rect 181 406 197 440
rect 131 390 197 406
rect 238 581 762 615
rect 238 556 304 581
rect 238 522 254 556
rect 288 522 304 556
rect 238 488 304 522
rect 238 454 254 488
rect 288 454 304 488
rect 238 420 304 454
rect 17 236 51 390
rect 238 386 254 420
rect 288 386 304 420
rect 238 370 304 386
rect 85 320 161 356
rect 85 286 91 320
rect 125 286 161 320
rect 85 270 161 286
rect 195 320 236 336
rect 195 286 199 320
rect 233 286 236 320
rect 195 236 236 286
rect 270 298 304 370
rect 338 513 602 547
rect 636 513 652 547
rect 692 521 762 581
rect 338 366 372 513
rect 692 487 708 521
rect 742 487 762 521
rect 406 456 655 479
rect 440 445 655 456
rect 406 400 440 422
rect 480 377 496 411
rect 530 377 555 411
rect 338 332 419 366
rect 480 361 555 377
rect 270 264 349 298
rect 17 230 236 236
rect 283 237 349 264
rect 17 220 249 230
rect 17 186 39 220
rect 73 196 249 220
rect 17 146 73 186
rect 17 112 39 146
rect 17 96 73 112
rect 109 146 181 162
rect 109 112 128 146
rect 162 112 181 146
rect 109 96 181 112
rect 109 17 143 96
rect 215 85 249 196
rect 283 203 299 237
rect 333 203 349 237
rect 283 169 349 203
rect 283 135 299 169
rect 333 135 349 169
rect 283 119 349 135
rect 385 265 419 332
rect 385 244 455 265
rect 385 210 401 244
rect 435 210 455 244
rect 385 202 455 210
rect 385 169 415 202
rect 385 135 401 169
rect 449 168 455 202
rect 435 135 455 168
rect 385 119 455 135
rect 489 247 555 361
rect 489 213 505 247
rect 539 213 555 247
rect 489 179 555 213
rect 489 145 505 179
rect 539 145 555 179
rect 589 350 655 445
rect 589 316 607 350
rect 641 316 655 350
rect 589 247 655 316
rect 589 213 605 247
rect 639 213 655 247
rect 589 179 655 213
rect 589 145 605 179
rect 639 145 655 179
rect 692 411 762 487
rect 692 377 708 411
rect 742 377 762 411
rect 692 249 762 377
rect 692 215 712 249
rect 746 215 762 249
rect 692 179 762 215
rect 692 145 712 179
rect 746 145 762 179
rect 489 85 523 145
rect 692 129 762 145
rect 808 577 875 593
rect 808 543 825 577
rect 859 543 875 577
rect 808 494 875 543
rect 808 460 825 494
rect 859 460 875 494
rect 808 411 875 460
rect 808 377 825 411
rect 859 377 875 411
rect 808 361 875 377
rect 909 577 975 649
rect 909 543 925 577
rect 959 543 975 577
rect 909 494 975 543
rect 909 460 925 494
rect 959 460 975 494
rect 909 411 975 460
rect 909 377 925 411
rect 959 377 975 411
rect 1020 577 1086 593
rect 1020 543 1036 577
rect 1070 543 1086 577
rect 1020 509 1086 543
rect 1020 475 1036 509
rect 1070 475 1086 509
rect 1020 441 1086 475
rect 1020 407 1036 441
rect 1070 407 1086 441
rect 1158 577 1224 593
rect 1158 543 1174 577
rect 1208 543 1224 577
rect 1158 467 1224 543
rect 1158 433 1174 467
rect 1208 451 1224 467
rect 1269 577 1495 594
rect 1269 543 1274 577
rect 1308 543 1351 577
rect 1385 543 1428 577
rect 1462 543 1495 577
rect 1269 467 1495 543
rect 1208 433 1235 451
rect 1158 417 1235 433
rect 1269 433 1274 467
rect 1308 433 1351 467
rect 1385 433 1428 467
rect 1462 433 1495 467
rect 1269 417 1495 433
rect 1020 395 1086 407
rect 909 361 975 377
rect 808 202 842 361
rect 889 294 1012 310
rect 889 260 963 294
rect 997 260 1012 294
rect 889 236 1012 260
rect 1046 261 1080 395
rect 1114 345 1167 361
rect 1114 311 1130 345
rect 1164 311 1167 345
rect 1114 295 1167 311
rect 1046 227 1099 261
rect 808 196 947 202
rect 808 162 897 196
rect 931 162 947 196
rect 808 120 947 162
rect 215 51 523 85
rect 557 95 623 111
rect 557 61 573 95
rect 607 85 623 95
rect 808 86 829 120
rect 863 86 902 120
rect 936 86 947 120
rect 808 85 947 86
rect 607 61 947 85
rect 557 51 947 61
rect 981 148 1031 193
rect 981 114 997 148
rect 981 17 1031 114
rect 1065 128 1099 227
rect 1133 208 1167 295
rect 1201 276 1235 417
rect 1269 360 1322 376
rect 1269 326 1272 360
rect 1306 350 1322 360
rect 1269 316 1279 326
rect 1313 316 1322 350
rect 1269 310 1322 316
rect 1364 344 1427 360
rect 1364 310 1380 344
rect 1414 310 1427 344
rect 1364 276 1427 310
rect 1201 242 1330 276
rect 1133 202 1223 208
rect 1133 168 1183 202
rect 1217 168 1223 202
rect 1133 162 1223 168
rect 1264 190 1330 242
rect 1264 156 1280 190
rect 1314 156 1330 190
rect 1364 242 1380 276
rect 1414 242 1427 276
rect 1364 226 1427 242
rect 1364 202 1415 226
rect 1364 168 1375 202
rect 1409 168 1415 202
rect 1461 192 1495 417
rect 1529 580 1563 649
rect 1529 509 1563 546
rect 1529 438 1563 475
rect 1529 388 1563 404
rect 1603 580 1669 596
rect 1603 546 1619 580
rect 1653 546 1669 580
rect 1603 498 1669 546
rect 1715 582 2091 608
rect 1715 548 1731 582
rect 1765 580 2091 582
rect 1765 574 2040 580
rect 1765 548 1781 574
rect 1715 532 1781 548
rect 2074 546 2091 580
rect 1912 524 2006 540
rect 1912 498 1928 524
rect 1603 497 1928 498
rect 1603 463 1619 497
rect 1653 490 1928 497
rect 1962 490 2006 524
rect 1653 464 2006 490
rect 1653 463 1669 464
rect 1603 414 1669 463
rect 1603 380 1619 414
rect 1653 380 1669 414
rect 1603 364 1669 380
rect 1535 294 1601 310
rect 1535 260 1551 294
rect 1585 260 1601 294
rect 1535 236 1601 260
rect 1635 226 1669 364
rect 1827 414 1872 430
rect 1827 380 1838 414
rect 1827 364 1872 380
rect 1912 414 2006 464
rect 1912 380 1928 414
rect 1962 380 2006 414
rect 1912 364 2006 380
rect 1703 350 1793 356
rect 1703 316 1759 350
rect 1703 310 1793 316
rect 1703 276 1711 310
rect 1745 276 1753 310
rect 1827 276 1861 364
rect 1972 318 2006 364
rect 2040 509 2091 546
rect 2074 475 2091 509
rect 2040 438 2091 475
rect 2074 404 2091 438
rect 2130 580 2180 649
rect 2164 546 2180 580
rect 2130 470 2180 546
rect 2164 436 2180 470
rect 2130 420 2180 436
rect 2215 580 2287 596
rect 2215 546 2231 580
rect 2265 546 2287 580
rect 2215 497 2287 546
rect 2215 463 2231 497
rect 2265 463 2287 497
rect 2040 386 2091 404
rect 2215 414 2287 463
rect 2040 352 2125 386
rect 2215 380 2231 414
rect 2265 380 2287 414
rect 2215 364 2287 380
rect 1703 260 1753 276
rect 1787 242 1861 276
rect 1895 302 1938 318
rect 1895 268 1899 302
rect 1933 268 1938 302
rect 1895 252 1938 268
rect 1972 302 2057 318
rect 1972 268 2007 302
rect 2041 268 2057 302
rect 1972 252 2057 268
rect 1787 226 1821 242
rect 1635 210 1703 226
rect 1364 162 1415 168
rect 1449 188 1515 192
rect 1065 94 1083 128
rect 1117 94 1180 128
rect 1214 94 1230 128
rect 1065 78 1230 94
rect 1264 120 1330 156
rect 1264 86 1280 120
rect 1314 86 1330 120
rect 1264 70 1330 86
rect 1449 154 1465 188
rect 1499 154 1515 188
rect 1449 120 1515 154
rect 1449 86 1465 120
rect 1499 86 1515 120
rect 1449 70 1515 86
rect 1549 186 1599 202
rect 1549 152 1565 186
rect 1549 116 1599 152
rect 1549 82 1565 116
rect 1549 17 1599 82
rect 1635 176 1653 210
rect 1687 176 1703 210
rect 1635 120 1703 176
rect 1635 86 1653 120
rect 1687 86 1703 120
rect 1635 70 1703 86
rect 1755 210 1821 226
rect 1755 176 1771 210
rect 1805 176 1821 210
rect 1895 208 1929 252
rect 2091 218 2125 352
rect 1755 140 1821 176
rect 1855 202 1929 208
rect 1889 168 1929 202
rect 1855 162 1929 168
rect 1963 185 2125 218
rect 1755 106 1771 140
rect 1805 106 1821 140
rect 1997 184 2125 185
rect 2162 310 2219 326
rect 2162 276 2178 310
rect 2212 276 2219 310
rect 2162 260 2219 276
rect 1963 119 1997 151
rect 2162 150 2196 260
rect 2253 226 2287 364
rect 1755 85 1821 106
rect 2031 116 2196 150
rect 2231 210 2287 226
rect 2265 176 2287 210
rect 2231 120 2287 176
rect 2031 85 2065 116
rect 1755 51 2065 85
rect 2265 86 2287 120
rect 2099 48 2122 82
rect 2156 48 2179 82
rect 2231 70 2287 86
rect 2099 17 2179 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 415 169 449 202
rect 415 168 435 169
rect 435 168 449 169
rect 607 316 641 350
rect 1279 326 1306 350
rect 1306 326 1313 350
rect 1279 316 1313 326
rect 1183 168 1217 202
rect 1375 168 1409 202
rect 1759 316 1793 350
rect 1855 168 1889 202
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 595 350 653 356
rect 595 316 607 350
rect 641 347 653 350
rect 1267 350 1325 356
rect 1267 347 1279 350
rect 641 319 1279 347
rect 641 316 653 319
rect 595 310 653 316
rect 1267 316 1279 319
rect 1313 347 1325 350
rect 1747 350 1805 356
rect 1747 347 1759 350
rect 1313 319 1759 347
rect 1313 316 1325 319
rect 1267 310 1325 316
rect 1747 316 1759 319
rect 1793 316 1805 350
rect 1747 310 1805 316
rect 403 202 461 208
rect 403 168 415 202
rect 449 199 461 202
rect 1171 202 1229 208
rect 1171 199 1183 202
rect 449 171 1183 199
rect 449 168 461 171
rect 403 162 461 168
rect 1171 168 1183 171
rect 1217 199 1229 202
rect 1363 202 1421 208
rect 1363 199 1375 202
rect 1217 171 1375 199
rect 1217 168 1229 171
rect 1171 162 1229 168
rect 1363 168 1375 171
rect 1409 199 1421 202
rect 1843 202 1901 208
rect 1843 199 1855 202
rect 1409 171 1855 199
rect 1409 168 1421 171
rect 1363 162 1421 168
rect 1843 168 1855 171
rect 1889 168 1901 202
rect 1843 162 1901 168
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
flabel pwell s 0 0 2304 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2304 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fahcon_1
flabel metal1 s 0 617 2304 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2304 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 CI
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 2239 390 2273 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2239 464 2273 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2239 538 2273 572 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1279 94 1313 128 0 FreeSans 340 0 0 0 COUT_N
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2304 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 3916918
string GDS_START 3899164
<< end >>
