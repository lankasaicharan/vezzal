magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 4 49 661 241
rect 0 0 672 49
<< scnmos >>
rect 83 47 113 215
rect 169 47 199 215
rect 255 47 285 215
rect 380 47 410 215
rect 466 47 496 215
rect 552 47 582 215
<< scpmoshvt >>
rect 83 367 113 619
rect 169 367 199 619
rect 255 367 285 619
rect 372 367 402 619
rect 466 367 496 619
rect 552 367 582 619
<< ndiff >>
rect 30 203 83 215
rect 30 169 38 203
rect 72 169 83 203
rect 30 101 83 169
rect 30 67 38 101
rect 72 67 83 101
rect 30 47 83 67
rect 113 127 169 215
rect 113 93 124 127
rect 158 93 169 127
rect 113 47 169 93
rect 199 203 255 215
rect 199 169 210 203
rect 244 169 255 203
rect 199 101 255 169
rect 199 67 210 101
rect 244 67 255 101
rect 199 47 255 67
rect 285 161 380 215
rect 285 127 323 161
rect 357 127 380 161
rect 285 93 380 127
rect 285 59 323 93
rect 357 59 380 93
rect 285 47 380 59
rect 410 203 466 215
rect 410 169 421 203
rect 455 169 466 203
rect 410 101 466 169
rect 410 67 421 101
rect 455 67 466 101
rect 410 47 466 67
rect 496 169 552 215
rect 496 135 507 169
rect 541 135 552 169
rect 496 47 552 135
rect 582 192 635 215
rect 582 158 593 192
rect 627 158 635 192
rect 582 101 635 158
rect 582 67 593 101
rect 627 67 635 101
rect 582 47 635 67
<< pdiff >>
rect 30 607 83 619
rect 30 573 38 607
rect 72 573 83 607
rect 30 522 83 573
rect 30 488 38 522
rect 72 488 83 522
rect 30 441 83 488
rect 30 407 38 441
rect 72 407 83 441
rect 30 367 83 407
rect 113 599 169 619
rect 113 565 124 599
rect 158 565 169 599
rect 113 529 169 565
rect 113 495 124 529
rect 158 495 169 529
rect 113 457 169 495
rect 113 423 124 457
rect 158 423 169 457
rect 113 367 169 423
rect 199 531 255 619
rect 199 497 210 531
rect 244 497 255 531
rect 199 457 255 497
rect 199 423 210 457
rect 244 423 255 457
rect 199 367 255 423
rect 285 597 372 619
rect 285 563 311 597
rect 345 563 372 597
rect 285 515 372 563
rect 285 481 311 515
rect 345 481 372 515
rect 285 367 372 481
rect 402 607 466 619
rect 402 573 416 607
rect 450 573 466 607
rect 402 515 466 573
rect 402 481 416 515
rect 450 481 466 515
rect 402 367 466 481
rect 496 599 552 619
rect 496 565 507 599
rect 541 565 552 599
rect 496 505 552 565
rect 496 471 507 505
rect 541 471 552 505
rect 496 413 552 471
rect 496 379 507 413
rect 541 379 552 413
rect 496 367 552 379
rect 582 607 635 619
rect 582 573 593 607
rect 627 573 635 607
rect 582 516 635 573
rect 582 482 593 516
rect 627 482 635 516
rect 582 434 635 482
rect 582 400 593 434
rect 627 400 635 434
rect 582 367 635 400
<< ndiffc >>
rect 38 169 72 203
rect 38 67 72 101
rect 124 93 158 127
rect 210 169 244 203
rect 210 67 244 101
rect 323 127 357 161
rect 323 59 357 93
rect 421 169 455 203
rect 421 67 455 101
rect 507 135 541 169
rect 593 158 627 192
rect 593 67 627 101
<< pdiffc >>
rect 38 573 72 607
rect 38 488 72 522
rect 38 407 72 441
rect 124 565 158 599
rect 124 495 158 529
rect 124 423 158 457
rect 210 497 244 531
rect 210 423 244 457
rect 311 563 345 597
rect 311 481 345 515
rect 416 573 450 607
rect 416 481 450 515
rect 507 565 541 599
rect 507 471 541 505
rect 507 379 541 413
rect 593 573 627 607
rect 593 482 627 516
rect 593 400 627 434
<< poly >>
rect 83 619 113 645
rect 169 619 199 645
rect 255 619 285 645
rect 372 619 402 645
rect 466 619 496 645
rect 552 619 582 645
rect 83 325 113 367
rect 25 309 113 325
rect 25 275 41 309
rect 75 275 113 309
rect 169 303 199 367
rect 255 303 285 367
rect 372 335 402 367
rect 25 259 113 275
rect 83 215 113 259
rect 155 287 285 303
rect 155 253 171 287
rect 205 253 285 287
rect 358 319 424 335
rect 358 285 374 319
rect 408 285 424 319
rect 358 269 424 285
rect 466 303 496 367
rect 552 303 582 367
rect 466 287 647 303
rect 155 237 285 253
rect 169 215 199 237
rect 255 215 285 237
rect 380 215 410 269
rect 466 253 597 287
rect 631 253 647 287
rect 466 242 647 253
rect 466 215 496 242
rect 552 237 647 242
rect 552 215 582 237
rect 83 21 113 47
rect 169 21 199 47
rect 255 21 285 47
rect 380 21 410 47
rect 466 21 496 47
rect 552 21 582 47
<< polycont >>
rect 41 275 75 309
rect 171 253 205 287
rect 374 285 408 319
rect 597 253 631 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 22 607 88 649
rect 22 573 38 607
rect 72 573 88 607
rect 22 522 88 573
rect 22 488 38 522
rect 72 488 88 522
rect 22 441 88 488
rect 22 407 38 441
rect 72 407 88 441
rect 122 599 361 615
rect 122 565 124 599
rect 158 597 361 599
rect 158 581 311 597
rect 158 565 166 581
rect 122 529 166 565
rect 295 563 311 581
rect 345 563 361 597
rect 122 495 124 529
rect 158 495 166 529
rect 122 457 166 495
rect 122 423 124 457
rect 158 423 166 457
rect 122 407 166 423
rect 200 531 260 547
rect 200 497 210 531
rect 244 497 260 531
rect 200 457 260 497
rect 295 515 361 563
rect 295 481 311 515
rect 345 481 361 515
rect 295 475 361 481
rect 400 607 466 649
rect 400 573 416 607
rect 450 573 466 607
rect 400 515 466 573
rect 400 481 416 515
rect 450 481 466 515
rect 400 475 466 481
rect 500 599 547 615
rect 500 565 507 599
rect 541 565 547 599
rect 500 505 547 565
rect 200 423 210 457
rect 244 441 260 457
rect 500 471 507 505
rect 541 471 547 505
rect 500 441 547 471
rect 244 423 547 441
rect 200 413 547 423
rect 200 407 507 413
rect 319 384 507 407
rect 505 379 507 384
rect 541 379 547 413
rect 581 607 643 649
rect 581 573 593 607
rect 627 573 643 607
rect 581 516 643 573
rect 581 482 593 516
rect 627 482 643 516
rect 581 434 643 482
rect 581 400 593 434
rect 627 400 643 434
rect 581 384 643 400
rect 25 350 283 373
rect 25 339 471 350
rect 25 309 91 339
rect 25 275 41 309
rect 75 275 91 309
rect 249 319 471 339
rect 125 287 205 303
rect 125 253 171 287
rect 249 285 374 319
rect 408 285 471 319
rect 249 269 471 285
rect 125 237 205 253
rect 239 203 471 235
rect 22 169 38 203
rect 72 169 210 203
rect 244 201 421 203
rect 244 169 273 201
rect 22 101 74 169
rect 22 67 38 101
rect 72 67 74 101
rect 22 51 74 67
rect 108 127 174 135
rect 108 93 124 127
rect 158 93 174 127
rect 108 17 174 93
rect 208 101 273 169
rect 407 169 421 201
rect 455 169 471 203
rect 208 67 210 101
rect 244 67 273 101
rect 208 51 273 67
rect 307 161 373 165
rect 307 127 323 161
rect 357 127 373 161
rect 307 93 373 127
rect 307 59 323 93
rect 357 59 373 93
rect 307 17 373 59
rect 407 101 471 169
rect 505 169 547 379
rect 581 287 653 350
rect 581 253 597 287
rect 631 253 653 287
rect 581 242 653 253
rect 505 135 507 169
rect 541 135 547 169
rect 505 119 547 135
rect 581 192 643 208
rect 581 158 593 192
rect 627 158 643 192
rect 407 67 421 101
rect 455 85 471 101
rect 581 101 643 158
rect 581 85 593 101
rect 455 67 593 85
rect 627 67 643 101
rect 407 51 643 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21ai_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4532004
string GDS_START 4525078
<< end >>
