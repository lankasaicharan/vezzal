magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 383 1478 704
rect -38 331 768 383
rect 1041 337 1478 383
rect 1307 331 1478 337
<< pwell >>
rect 810 157 1265 295
rect 1 49 1439 157
rect 0 0 1440 49
<< scnmos >>
rect 893 185 923 269
rect 988 185 1018 269
rect 1074 185 1104 269
rect 1152 185 1182 269
rect 80 47 110 131
rect 152 47 182 131
rect 254 47 284 131
rect 332 47 362 131
rect 418 47 448 131
rect 584 47 614 131
rect 670 47 700 131
rect 748 47 778 131
rect 1254 47 1284 131
rect 1326 47 1356 131
<< scpmoshvt >>
rect 90 419 140 619
rect 204 419 254 619
rect 302 419 352 619
rect 476 419 526 619
rect 590 419 640 619
rect 711 419 761 619
rect 991 419 1041 619
rect 1097 419 1147 619
rect 1203 419 1253 619
rect 1309 419 1359 619
<< ndiff >>
rect 836 229 893 269
rect 836 195 848 229
rect 882 195 893 229
rect 836 185 893 195
rect 923 185 988 269
rect 1018 235 1074 269
rect 1018 201 1029 235
rect 1063 201 1074 235
rect 1018 185 1074 201
rect 1104 185 1152 269
rect 1182 244 1239 269
rect 1182 210 1193 244
rect 1227 210 1239 244
rect 1182 185 1239 210
rect 27 111 80 131
rect 27 77 35 111
rect 69 77 80 111
rect 27 47 80 77
rect 110 47 152 131
rect 182 100 254 131
rect 182 66 193 100
rect 227 66 254 100
rect 182 47 254 66
rect 284 47 332 131
rect 362 105 418 131
rect 362 71 373 105
rect 407 71 418 105
rect 362 47 418 71
rect 448 47 584 131
rect 614 102 670 131
rect 614 68 625 102
rect 659 68 670 102
rect 614 47 670 68
rect 700 47 748 131
rect 778 111 835 131
rect 778 77 789 111
rect 823 77 835 111
rect 778 47 835 77
rect 1197 106 1254 131
rect 1197 72 1209 106
rect 1243 72 1254 106
rect 1197 47 1254 72
rect 1284 47 1326 131
rect 1356 111 1413 131
rect 1356 77 1367 111
rect 1401 77 1413 111
rect 1356 47 1413 77
<< pdiff >>
rect 33 597 90 619
rect 33 563 45 597
rect 79 563 90 597
rect 33 516 90 563
rect 33 482 45 516
rect 79 482 90 516
rect 33 419 90 482
rect 140 607 204 619
rect 140 573 151 607
rect 185 573 204 607
rect 140 516 204 573
rect 140 482 151 516
rect 185 482 204 516
rect 140 419 204 482
rect 254 419 302 619
rect 352 466 476 619
rect 352 432 431 466
rect 465 432 476 466
rect 352 419 476 432
rect 526 419 590 619
rect 640 607 711 619
rect 640 573 652 607
rect 686 573 711 607
rect 640 419 711 573
rect 761 466 818 619
rect 761 432 772 466
rect 806 432 818 466
rect 761 419 818 432
rect 934 597 991 619
rect 934 563 946 597
rect 980 563 991 597
rect 934 513 991 563
rect 934 479 946 513
rect 980 479 991 513
rect 934 419 991 479
rect 1041 607 1097 619
rect 1041 573 1052 607
rect 1086 573 1097 607
rect 1041 513 1097 573
rect 1041 479 1052 513
rect 1086 479 1097 513
rect 1041 419 1097 479
rect 1147 597 1203 619
rect 1147 563 1158 597
rect 1192 563 1203 597
rect 1147 513 1203 563
rect 1147 479 1158 513
rect 1192 479 1203 513
rect 1147 419 1203 479
rect 1253 595 1309 619
rect 1253 561 1264 595
rect 1298 561 1309 595
rect 1253 419 1309 561
rect 1359 597 1413 619
rect 1359 563 1370 597
rect 1404 563 1413 597
rect 1359 465 1413 563
rect 1359 431 1370 465
rect 1404 431 1413 465
rect 1359 419 1413 431
<< ndiffc >>
rect 848 195 882 229
rect 1029 201 1063 235
rect 1193 210 1227 244
rect 35 77 69 111
rect 193 66 227 100
rect 373 71 407 105
rect 625 68 659 102
rect 789 77 823 111
rect 1209 72 1243 106
rect 1367 77 1401 111
<< pdiffc >>
rect 45 563 79 597
rect 45 482 79 516
rect 151 573 185 607
rect 151 482 185 516
rect 431 432 465 466
rect 652 573 686 607
rect 772 432 806 466
rect 946 563 980 597
rect 946 479 980 513
rect 1052 573 1086 607
rect 1052 479 1086 513
rect 1158 563 1192 597
rect 1158 479 1192 513
rect 1264 561 1298 595
rect 1370 563 1404 597
rect 1370 431 1404 465
<< poly >>
rect 90 619 140 645
rect 204 619 254 645
rect 302 619 352 645
rect 476 619 526 645
rect 590 619 640 645
rect 711 619 761 645
rect 991 619 1041 645
rect 1097 619 1147 645
rect 1203 619 1253 645
rect 1309 619 1359 645
rect 90 279 140 419
rect 204 387 254 419
rect 188 371 254 387
rect 188 337 204 371
rect 238 337 254 371
rect 302 368 352 419
rect 302 338 434 368
rect 188 321 254 337
rect 80 263 155 279
rect 80 229 105 263
rect 139 243 155 263
rect 139 229 182 243
rect 80 213 182 229
rect 80 131 110 213
rect 152 131 182 213
rect 224 176 254 321
rect 296 274 362 290
rect 296 240 312 274
rect 346 240 362 274
rect 296 224 362 240
rect 224 146 284 176
rect 254 131 284 146
rect 332 131 362 224
rect 404 219 434 338
rect 476 356 526 419
rect 476 340 542 356
rect 590 343 640 419
rect 711 387 761 419
rect 991 392 1041 419
rect 1097 392 1147 419
rect 692 371 761 387
rect 476 306 492 340
rect 526 306 542 340
rect 476 290 542 306
rect 584 327 650 343
rect 584 293 600 327
rect 634 293 650 327
rect 692 337 708 371
rect 742 337 761 371
rect 692 321 761 337
rect 988 362 1147 392
rect 1203 375 1253 419
rect 988 341 1104 362
rect 988 321 1005 341
rect 584 277 650 293
rect 404 203 484 219
rect 404 189 434 203
rect 418 169 434 189
rect 468 169 484 203
rect 418 153 484 169
rect 418 131 448 153
rect 584 131 614 277
rect 698 229 728 321
rect 893 307 1005 321
rect 1039 307 1104 341
rect 1189 359 1255 375
rect 1189 325 1205 359
rect 1239 325 1255 359
rect 1189 314 1255 325
rect 1309 315 1359 419
rect 893 291 1104 307
rect 893 269 923 291
rect 988 269 1018 291
rect 1074 269 1104 291
rect 1152 284 1255 314
rect 1297 299 1363 315
rect 1152 269 1182 284
rect 660 213 728 229
rect 660 179 676 213
rect 710 193 728 213
rect 710 179 778 193
rect 1297 265 1313 299
rect 1347 265 1363 299
rect 1297 231 1363 265
rect 1297 211 1313 231
rect 1254 197 1313 211
rect 1347 197 1363 231
rect 660 163 778 179
rect 670 131 700 163
rect 748 131 778 163
rect 893 159 923 185
rect 988 159 1018 185
rect 1074 159 1104 185
rect 1152 159 1182 185
rect 1254 181 1363 197
rect 1254 131 1284 181
rect 1326 131 1356 181
rect 80 21 110 47
rect 152 21 182 47
rect 254 21 284 47
rect 332 21 362 47
rect 418 21 448 47
rect 584 21 614 47
rect 670 21 700 47
rect 748 21 778 47
rect 1254 21 1284 47
rect 1326 21 1356 47
<< polycont >>
rect 204 337 238 371
rect 105 229 139 263
rect 312 240 346 274
rect 492 306 526 340
rect 600 293 634 327
rect 708 337 742 371
rect 434 169 468 203
rect 1005 307 1039 341
rect 1205 325 1239 359
rect 676 179 710 213
rect 1313 265 1347 299
rect 1313 197 1347 231
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 19 597 95 613
rect 19 563 45 597
rect 79 563 95 597
rect 19 516 95 563
rect 19 482 45 516
rect 79 482 95 516
rect 19 466 95 482
rect 135 607 201 649
rect 135 573 151 607
rect 185 573 201 607
rect 636 607 702 649
rect 636 573 652 607
rect 686 573 702 607
rect 930 597 996 613
rect 135 516 201 573
rect 930 563 946 597
rect 980 563 996 597
rect 930 537 996 563
rect 135 482 151 516
rect 185 482 201 516
rect 135 466 201 482
rect 328 513 996 537
rect 328 503 946 513
rect 19 177 53 466
rect 121 371 254 430
rect 121 337 204 371
rect 238 337 254 371
rect 121 321 254 337
rect 328 356 362 503
rect 864 479 946 503
rect 980 479 996 513
rect 415 466 720 467
rect 415 432 431 466
rect 465 432 720 466
rect 415 415 720 432
rect 756 466 828 467
rect 756 432 772 466
rect 806 432 828 466
rect 756 431 828 432
rect 686 387 720 415
rect 686 371 758 387
rect 328 340 542 356
rect 328 306 492 340
rect 526 306 542 340
rect 328 290 542 306
rect 584 327 650 343
rect 686 337 708 371
rect 742 337 758 371
rect 686 335 758 337
rect 584 293 600 327
rect 634 299 650 327
rect 794 299 828 431
rect 634 293 828 299
rect 296 279 362 290
rect 89 274 362 279
rect 89 263 312 274
rect 89 229 105 263
rect 139 240 312 263
rect 346 240 362 274
rect 584 265 828 293
rect 864 463 996 479
rect 1036 607 1102 649
rect 1036 573 1052 607
rect 1086 573 1102 607
rect 1036 513 1102 573
rect 1036 479 1052 513
rect 1086 479 1102 513
rect 1036 463 1102 479
rect 1142 597 1208 613
rect 1142 563 1158 597
rect 1192 563 1208 597
rect 1142 513 1208 563
rect 1248 595 1314 649
rect 1248 561 1264 595
rect 1298 561 1314 595
rect 1248 533 1314 561
rect 1369 597 1422 613
rect 1369 563 1370 597
rect 1404 563 1422 597
rect 1142 479 1158 513
rect 1192 497 1208 513
rect 1192 479 1331 497
rect 1142 463 1331 479
rect 139 229 362 240
rect 89 213 362 229
rect 418 203 484 219
rect 418 177 434 203
rect 19 169 434 177
rect 468 169 484 203
rect 19 143 484 169
rect 520 213 726 229
rect 520 179 676 213
rect 710 179 726 213
rect 520 163 726 179
rect 19 111 85 143
rect 19 77 35 111
rect 69 77 85 111
rect 520 107 554 163
rect 762 135 796 265
rect 864 229 898 463
rect 832 195 848 229
rect 882 195 898 229
rect 832 179 898 195
rect 934 393 1255 427
rect 934 135 968 393
rect 1189 359 1255 393
rect 1004 341 1127 357
rect 1004 307 1005 341
rect 1039 307 1127 341
rect 1189 325 1205 359
rect 1239 325 1255 359
rect 1189 309 1255 325
rect 1297 315 1331 463
rect 1369 465 1422 563
rect 1369 431 1370 465
rect 1404 431 1422 465
rect 1369 384 1422 431
rect 1004 291 1127 307
rect 1297 299 1352 315
rect 19 53 85 77
rect 177 100 243 107
rect 177 66 193 100
rect 227 66 243 100
rect 177 17 243 66
rect 357 105 554 107
rect 357 71 373 105
rect 407 71 554 105
rect 357 53 554 71
rect 609 102 675 127
rect 609 68 625 102
rect 659 68 675 102
rect 609 17 675 68
rect 762 111 968 135
rect 762 77 789 111
rect 823 101 968 111
rect 1013 235 1079 255
rect 1013 201 1029 235
rect 1063 201 1079 235
rect 823 77 839 101
rect 762 53 839 77
rect 1013 17 1079 201
rect 1177 244 1243 273
rect 1177 210 1193 244
rect 1227 215 1243 244
rect 1297 265 1313 299
rect 1347 265 1352 299
rect 1297 231 1352 265
rect 1297 215 1313 231
rect 1227 210 1313 215
rect 1177 197 1313 210
rect 1347 197 1352 231
rect 1177 181 1352 197
rect 1388 135 1422 384
rect 1193 106 1259 135
rect 1193 72 1209 106
rect 1243 72 1259 106
rect 1193 17 1259 72
rect 1351 111 1422 135
rect 1351 77 1367 111
rect 1401 77 1422 111
rect 1351 53 1422 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlclkp_lp
flabel comment s 710 282 710 282 0 FreeSans 200 270 0 0 no_jumper_check
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1375 390 1409 424 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1375 464 1409 498 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1375 538 1409 572 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3486268
string GDS_START 3476164
<< end >>
