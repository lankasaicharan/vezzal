magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 11 49 738 235
rect 0 0 768 49
<< scnmos >>
rect 94 125 124 209
rect 180 125 210 209
rect 298 125 328 209
rect 384 125 414 209
rect 521 125 551 209
rect 629 125 659 209
<< scpmoshvt >>
rect 107 535 137 619
rect 193 535 223 619
rect 265 535 295 619
rect 449 429 479 513
rect 535 429 565 513
rect 635 429 665 513
<< ndiff >>
rect 37 171 94 209
rect 37 137 45 171
rect 79 137 94 171
rect 37 125 94 137
rect 124 190 180 209
rect 124 156 135 190
rect 169 156 180 190
rect 124 125 180 156
rect 210 136 298 209
rect 210 125 237 136
rect 225 102 237 125
rect 271 125 298 136
rect 328 190 384 209
rect 328 156 339 190
rect 373 156 384 190
rect 328 125 384 156
rect 414 197 521 209
rect 414 163 425 197
rect 459 163 521 197
rect 414 125 521 163
rect 551 125 629 209
rect 659 171 712 209
rect 659 137 670 171
rect 704 137 712 171
rect 659 125 712 137
rect 271 102 283 125
rect 225 94 283 102
<< pdiff >>
rect 50 581 107 619
rect 50 547 58 581
rect 92 547 107 581
rect 50 535 107 547
rect 137 607 193 619
rect 137 573 148 607
rect 182 573 193 607
rect 137 535 193 573
rect 223 535 265 619
rect 295 609 352 619
rect 295 575 306 609
rect 340 575 352 609
rect 295 567 352 575
rect 295 535 345 567
rect 399 481 449 513
rect 392 471 449 481
rect 392 437 404 471
rect 438 437 449 471
rect 392 429 449 437
rect 479 475 535 513
rect 479 441 490 475
rect 524 441 535 475
rect 479 429 535 441
rect 565 505 635 513
rect 565 471 580 505
rect 614 471 635 505
rect 565 429 635 471
rect 665 475 718 513
rect 665 441 676 475
rect 710 441 718 475
rect 665 429 718 441
<< ndiffc >>
rect 45 137 79 171
rect 135 156 169 190
rect 237 102 271 136
rect 339 156 373 190
rect 425 163 459 197
rect 670 137 704 171
<< pdiffc >>
rect 58 547 92 581
rect 148 573 182 607
rect 306 575 340 609
rect 404 437 438 471
rect 490 441 524 475
rect 580 471 614 505
rect 676 441 710 475
<< poly >>
rect 107 619 137 645
rect 193 619 223 645
rect 265 619 295 645
rect 413 597 479 613
rect 413 563 429 597
rect 463 563 479 597
rect 413 547 479 563
rect 107 479 137 535
rect 85 463 151 479
rect 85 429 101 463
rect 135 429 151 463
rect 85 395 151 429
rect 85 361 101 395
rect 135 361 151 395
rect 85 345 151 361
rect 94 209 124 345
rect 193 297 223 535
rect 265 440 295 535
rect 449 513 479 547
rect 535 513 565 539
rect 635 513 665 539
rect 265 424 343 440
rect 265 390 293 424
rect 327 390 343 424
rect 265 374 343 390
rect 180 281 246 297
rect 180 247 196 281
rect 230 247 246 281
rect 180 231 246 247
rect 180 209 210 231
rect 298 209 328 374
rect 449 261 479 429
rect 535 365 565 429
rect 635 365 665 429
rect 384 231 479 261
rect 521 349 587 365
rect 521 315 537 349
rect 571 315 587 349
rect 521 281 587 315
rect 521 247 537 281
rect 571 247 587 281
rect 521 231 587 247
rect 629 349 695 365
rect 629 315 645 349
rect 679 315 695 349
rect 629 281 695 315
rect 629 247 645 281
rect 679 247 695 281
rect 629 231 695 247
rect 384 209 414 231
rect 521 209 551 231
rect 629 209 659 231
rect 94 99 124 125
rect 180 99 210 125
rect 298 99 328 125
rect 384 103 414 125
rect 384 87 450 103
rect 521 99 551 125
rect 629 99 659 125
rect 384 53 400 87
rect 434 53 450 87
rect 384 37 450 53
<< polycont >>
rect 429 563 463 597
rect 101 429 135 463
rect 101 361 135 395
rect 293 390 327 424
rect 196 247 230 281
rect 537 315 571 349
rect 537 247 571 281
rect 645 315 679 349
rect 645 247 679 281
rect 400 53 434 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 132 607 198 649
rect 29 581 96 597
rect 29 547 58 581
rect 92 547 96 581
rect 132 573 148 607
rect 182 573 198 607
rect 132 569 198 573
rect 290 609 463 613
rect 290 575 306 609
rect 340 597 463 609
rect 340 575 429 597
rect 290 563 429 575
rect 290 547 463 563
rect 29 531 96 547
rect 29 175 65 531
rect 564 505 630 649
rect 101 463 135 479
rect 101 395 135 429
rect 223 424 353 498
rect 223 390 293 424
rect 327 390 353 424
rect 400 471 443 487
rect 400 437 404 471
rect 438 437 443 471
rect 101 354 135 361
rect 400 354 443 437
rect 486 475 528 491
rect 486 441 490 475
rect 524 441 528 475
rect 564 471 580 505
rect 614 471 630 505
rect 672 475 714 491
rect 486 435 528 441
rect 672 441 676 475
rect 710 441 714 475
rect 672 435 714 441
rect 486 401 714 435
rect 101 320 443 354
rect 127 247 196 281
rect 230 247 353 281
rect 127 242 353 247
rect 409 276 443 320
rect 511 349 571 365
rect 511 315 537 349
rect 511 281 571 315
rect 131 190 373 206
rect 29 171 95 175
rect 29 137 45 171
rect 79 137 95 171
rect 29 94 95 137
rect 131 156 135 190
rect 169 172 339 190
rect 169 156 173 172
rect 131 17 173 156
rect 335 156 339 172
rect 409 197 475 276
rect 409 163 425 197
rect 459 163 475 197
rect 409 159 475 163
rect 511 247 537 281
rect 335 140 373 156
rect 221 102 237 136
rect 271 102 287 136
rect 221 87 287 102
rect 511 94 571 247
rect 607 349 737 350
rect 607 315 645 349
rect 679 315 737 349
rect 607 281 737 315
rect 607 247 645 281
rect 679 247 737 281
rect 607 242 737 247
rect 654 171 720 175
rect 654 137 670 171
rect 704 137 720 171
rect 221 53 400 87
rect 434 53 450 87
rect 654 17 720 137
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2bb2o_m
flabel comment s 461 363 461 363 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5860686
string GDS_START 5851702
<< end >>
