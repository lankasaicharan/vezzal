magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
<< pwell >>
rect 2 49 2052 241
rect 0 0 2112 49
<< scnmos >>
rect 81 47 111 215
rect 167 47 197 215
rect 253 47 283 215
rect 339 47 369 215
rect 425 47 455 215
rect 511 47 541 215
rect 597 47 627 215
rect 683 47 713 215
rect 893 47 923 215
rect 979 47 1009 215
rect 1065 47 1095 215
rect 1151 47 1181 215
rect 1237 47 1267 215
rect 1323 47 1353 215
rect 1409 47 1439 215
rect 1495 47 1525 215
rect 1685 47 1715 215
rect 1771 47 1801 215
rect 1857 47 1887 215
rect 1943 47 1973 215
<< scpmoshvt >>
rect 95 367 125 619
rect 181 367 211 619
rect 267 367 297 619
rect 353 367 383 619
rect 439 367 469 619
rect 525 367 555 619
rect 611 367 641 619
rect 697 367 727 619
rect 805 367 835 619
rect 891 367 921 619
rect 977 367 1007 619
rect 1131 367 1161 619
rect 1217 367 1247 619
rect 1375 367 1405 619
rect 1461 367 1491 619
rect 1547 367 1577 619
rect 1633 367 1663 619
rect 1719 367 1749 619
rect 1805 367 1835 619
rect 1891 367 1921 619
<< ndiff >>
rect 28 192 81 215
rect 28 158 36 192
rect 70 158 81 192
rect 28 101 81 158
rect 28 67 36 101
rect 70 67 81 101
rect 28 47 81 67
rect 111 129 167 215
rect 111 95 122 129
rect 156 95 167 129
rect 111 47 167 95
rect 197 192 253 215
rect 197 158 208 192
rect 242 158 253 192
rect 197 101 253 158
rect 197 67 208 101
rect 242 67 253 101
rect 197 47 253 67
rect 283 129 339 215
rect 283 95 294 129
rect 328 95 339 129
rect 283 47 339 95
rect 369 192 425 215
rect 369 158 380 192
rect 414 158 425 192
rect 369 101 425 158
rect 369 67 380 101
rect 414 67 425 101
rect 369 47 425 67
rect 455 202 511 215
rect 455 168 466 202
rect 500 168 511 202
rect 455 47 511 168
rect 541 103 597 215
rect 541 69 552 103
rect 586 69 597 103
rect 541 47 597 69
rect 627 202 683 215
rect 627 168 638 202
rect 672 168 683 202
rect 627 47 683 168
rect 713 103 766 215
rect 713 69 724 103
rect 758 69 766 103
rect 713 47 766 69
rect 840 103 893 215
rect 840 69 848 103
rect 882 69 893 103
rect 840 47 893 69
rect 923 202 979 215
rect 923 168 934 202
rect 968 168 979 202
rect 923 47 979 168
rect 1009 103 1065 215
rect 1009 69 1020 103
rect 1054 69 1065 103
rect 1009 47 1065 69
rect 1095 202 1151 215
rect 1095 168 1106 202
rect 1140 168 1151 202
rect 1095 47 1151 168
rect 1181 103 1237 215
rect 1181 69 1192 103
rect 1226 69 1237 103
rect 1181 47 1237 69
rect 1267 193 1323 215
rect 1267 159 1278 193
rect 1312 159 1323 193
rect 1267 47 1323 159
rect 1353 103 1409 215
rect 1353 69 1364 103
rect 1398 69 1409 103
rect 1353 47 1409 69
rect 1439 193 1495 215
rect 1439 159 1450 193
rect 1484 159 1495 193
rect 1439 47 1495 159
rect 1525 103 1578 215
rect 1525 69 1536 103
rect 1570 69 1578 103
rect 1525 47 1578 69
rect 1632 110 1685 215
rect 1632 76 1640 110
rect 1674 76 1685 110
rect 1632 47 1685 76
rect 1715 192 1771 215
rect 1715 158 1726 192
rect 1760 158 1771 192
rect 1715 101 1771 158
rect 1715 67 1726 101
rect 1760 67 1771 101
rect 1715 47 1771 67
rect 1801 110 1857 215
rect 1801 76 1812 110
rect 1846 76 1857 110
rect 1801 47 1857 76
rect 1887 192 1943 215
rect 1887 158 1898 192
rect 1932 158 1943 192
rect 1887 101 1943 158
rect 1887 67 1898 101
rect 1932 67 1943 101
rect 1887 47 1943 67
rect 1973 203 2026 215
rect 1973 169 1984 203
rect 2018 169 2026 203
rect 1973 93 2026 169
rect 1973 59 1984 93
rect 2018 59 2026 93
rect 1973 47 2026 59
<< pdiff >>
rect 42 599 95 619
rect 42 565 50 599
rect 84 565 95 599
rect 42 506 95 565
rect 42 472 50 506
rect 84 472 95 506
rect 42 415 95 472
rect 42 381 50 415
rect 84 381 95 415
rect 42 367 95 381
rect 125 547 181 619
rect 125 513 136 547
rect 170 513 181 547
rect 125 479 181 513
rect 125 445 136 479
rect 170 445 181 479
rect 125 411 181 445
rect 125 377 136 411
rect 170 377 181 411
rect 125 367 181 377
rect 211 599 267 619
rect 211 565 222 599
rect 256 565 267 599
rect 211 529 267 565
rect 211 495 222 529
rect 256 495 267 529
rect 211 459 267 495
rect 211 425 222 459
rect 256 425 267 459
rect 211 367 267 425
rect 297 547 353 619
rect 297 513 308 547
rect 342 513 353 547
rect 297 479 353 513
rect 297 445 308 479
rect 342 445 353 479
rect 297 411 353 445
rect 297 377 308 411
rect 342 377 353 411
rect 297 367 353 377
rect 383 599 439 619
rect 383 565 394 599
rect 428 565 439 599
rect 383 529 439 565
rect 383 495 394 529
rect 428 495 439 529
rect 383 459 439 495
rect 383 425 394 459
rect 428 425 439 459
rect 383 367 439 425
rect 469 547 525 619
rect 469 513 480 547
rect 514 513 525 547
rect 469 479 525 513
rect 469 445 480 479
rect 514 445 525 479
rect 469 411 525 445
rect 469 377 480 411
rect 514 377 525 411
rect 469 367 525 377
rect 555 599 611 619
rect 555 565 566 599
rect 600 565 611 599
rect 555 529 611 565
rect 555 495 566 529
rect 600 495 611 529
rect 555 459 611 495
rect 555 425 566 459
rect 600 425 611 459
rect 555 367 611 425
rect 641 547 697 619
rect 641 513 652 547
rect 686 513 697 547
rect 641 479 697 513
rect 641 445 652 479
rect 686 445 697 479
rect 641 411 697 445
rect 641 377 652 411
rect 686 377 697 411
rect 641 367 697 377
rect 727 599 805 619
rect 727 565 749 599
rect 783 565 805 599
rect 727 529 805 565
rect 727 495 749 529
rect 783 495 805 529
rect 727 459 805 495
rect 727 425 749 459
rect 783 425 805 459
rect 727 367 805 425
rect 835 607 891 619
rect 835 573 846 607
rect 880 573 891 607
rect 835 517 891 573
rect 835 483 846 517
rect 880 483 891 517
rect 835 367 891 483
rect 921 599 977 619
rect 921 565 932 599
rect 966 565 977 599
rect 921 529 977 565
rect 921 495 932 529
rect 966 495 977 529
rect 921 459 977 495
rect 921 425 932 459
rect 966 425 977 459
rect 921 367 977 425
rect 1007 607 1131 619
rect 1007 573 1018 607
rect 1052 573 1086 607
rect 1120 573 1131 607
rect 1007 526 1131 573
rect 1007 492 1018 526
rect 1052 492 1086 526
rect 1120 492 1131 526
rect 1007 367 1131 492
rect 1161 599 1217 619
rect 1161 565 1172 599
rect 1206 565 1217 599
rect 1161 529 1217 565
rect 1161 495 1172 529
rect 1206 495 1217 529
rect 1161 459 1217 495
rect 1161 425 1172 459
rect 1206 425 1217 459
rect 1161 367 1217 425
rect 1247 607 1375 619
rect 1247 573 1258 607
rect 1292 573 1330 607
rect 1364 573 1375 607
rect 1247 517 1375 573
rect 1247 483 1258 517
rect 1292 483 1330 517
rect 1364 483 1375 517
rect 1247 367 1375 483
rect 1405 599 1461 619
rect 1405 565 1416 599
rect 1450 565 1461 599
rect 1405 510 1461 565
rect 1405 476 1416 510
rect 1450 476 1461 510
rect 1405 409 1461 476
rect 1405 375 1416 409
rect 1450 375 1461 409
rect 1405 367 1461 375
rect 1491 607 1547 619
rect 1491 573 1502 607
rect 1536 573 1547 607
rect 1491 519 1547 573
rect 1491 485 1502 519
rect 1536 485 1547 519
rect 1491 423 1547 485
rect 1491 389 1502 423
rect 1536 389 1547 423
rect 1491 367 1547 389
rect 1577 599 1633 619
rect 1577 565 1588 599
rect 1622 565 1633 599
rect 1577 510 1633 565
rect 1577 476 1588 510
rect 1622 476 1633 510
rect 1577 409 1633 476
rect 1577 375 1588 409
rect 1622 375 1633 409
rect 1577 367 1633 375
rect 1663 607 1719 619
rect 1663 573 1674 607
rect 1708 573 1719 607
rect 1663 519 1719 573
rect 1663 485 1674 519
rect 1708 485 1719 519
rect 1663 423 1719 485
rect 1663 389 1674 423
rect 1708 389 1719 423
rect 1663 367 1719 389
rect 1749 599 1805 619
rect 1749 565 1760 599
rect 1794 565 1805 599
rect 1749 510 1805 565
rect 1749 476 1760 510
rect 1794 476 1805 510
rect 1749 413 1805 476
rect 1749 379 1760 413
rect 1794 379 1805 413
rect 1749 367 1805 379
rect 1835 607 1891 619
rect 1835 573 1846 607
rect 1880 573 1891 607
rect 1835 519 1891 573
rect 1835 485 1846 519
rect 1880 485 1891 519
rect 1835 423 1891 485
rect 1835 389 1846 423
rect 1880 389 1891 423
rect 1835 367 1891 389
rect 1921 599 1974 619
rect 1921 565 1932 599
rect 1966 565 1974 599
rect 1921 510 1974 565
rect 1921 476 1932 510
rect 1966 476 1974 510
rect 1921 413 1974 476
rect 1921 379 1932 413
rect 1966 379 1974 413
rect 1921 367 1974 379
<< ndiffc >>
rect 36 158 70 192
rect 36 67 70 101
rect 122 95 156 129
rect 208 158 242 192
rect 208 67 242 101
rect 294 95 328 129
rect 380 158 414 192
rect 380 67 414 101
rect 466 168 500 202
rect 552 69 586 103
rect 638 168 672 202
rect 724 69 758 103
rect 848 69 882 103
rect 934 168 968 202
rect 1020 69 1054 103
rect 1106 168 1140 202
rect 1192 69 1226 103
rect 1278 159 1312 193
rect 1364 69 1398 103
rect 1450 159 1484 193
rect 1536 69 1570 103
rect 1640 76 1674 110
rect 1726 158 1760 192
rect 1726 67 1760 101
rect 1812 76 1846 110
rect 1898 158 1932 192
rect 1898 67 1932 101
rect 1984 169 2018 203
rect 1984 59 2018 93
<< pdiffc >>
rect 50 565 84 599
rect 50 472 84 506
rect 50 381 84 415
rect 136 513 170 547
rect 136 445 170 479
rect 136 377 170 411
rect 222 565 256 599
rect 222 495 256 529
rect 222 425 256 459
rect 308 513 342 547
rect 308 445 342 479
rect 308 377 342 411
rect 394 565 428 599
rect 394 495 428 529
rect 394 425 428 459
rect 480 513 514 547
rect 480 445 514 479
rect 480 377 514 411
rect 566 565 600 599
rect 566 495 600 529
rect 566 425 600 459
rect 652 513 686 547
rect 652 445 686 479
rect 652 377 686 411
rect 749 565 783 599
rect 749 495 783 529
rect 749 425 783 459
rect 846 573 880 607
rect 846 483 880 517
rect 932 565 966 599
rect 932 495 966 529
rect 932 425 966 459
rect 1018 573 1052 607
rect 1086 573 1120 607
rect 1018 492 1052 526
rect 1086 492 1120 526
rect 1172 565 1206 599
rect 1172 495 1206 529
rect 1172 425 1206 459
rect 1258 573 1292 607
rect 1330 573 1364 607
rect 1258 483 1292 517
rect 1330 483 1364 517
rect 1416 565 1450 599
rect 1416 476 1450 510
rect 1416 375 1450 409
rect 1502 573 1536 607
rect 1502 485 1536 519
rect 1502 389 1536 423
rect 1588 565 1622 599
rect 1588 476 1622 510
rect 1588 375 1622 409
rect 1674 573 1708 607
rect 1674 485 1708 519
rect 1674 389 1708 423
rect 1760 565 1794 599
rect 1760 476 1794 510
rect 1760 379 1794 413
rect 1846 573 1880 607
rect 1846 485 1880 519
rect 1846 389 1880 423
rect 1932 565 1966 599
rect 1932 476 1966 510
rect 1932 379 1966 413
<< poly >>
rect 95 619 125 645
rect 181 619 211 645
rect 267 619 297 645
rect 353 619 383 645
rect 439 619 469 645
rect 525 619 555 645
rect 611 619 641 645
rect 697 619 727 645
rect 805 619 835 645
rect 891 619 921 645
rect 977 619 1007 645
rect 1131 619 1161 645
rect 1217 619 1247 645
rect 1375 619 1405 645
rect 1461 619 1491 645
rect 1547 619 1577 645
rect 1633 619 1663 645
rect 1719 619 1749 645
rect 1805 619 1835 645
rect 1891 619 1921 645
rect 95 303 125 367
rect 181 303 211 367
rect 267 303 297 367
rect 353 303 383 367
rect 439 303 469 367
rect 525 303 555 367
rect 611 303 641 367
rect 697 303 727 367
rect 805 333 835 367
rect 891 333 921 367
rect 977 333 1007 367
rect 1131 333 1161 367
rect 31 287 383 303
rect 31 253 47 287
rect 81 253 115 287
rect 149 253 183 287
rect 217 253 251 287
rect 285 253 319 287
rect 353 273 383 287
rect 425 287 763 303
rect 353 253 369 273
rect 31 237 369 253
rect 81 215 111 237
rect 167 215 197 237
rect 253 215 283 237
rect 339 215 369 237
rect 425 253 441 287
rect 475 253 509 287
rect 543 253 577 287
rect 611 253 645 287
rect 679 253 713 287
rect 747 253 763 287
rect 425 237 763 253
rect 805 287 1161 333
rect 1217 345 1247 367
rect 1217 315 1267 345
rect 805 253 821 287
rect 855 253 889 287
rect 923 253 957 287
rect 991 253 1025 287
rect 1059 253 1093 287
rect 1127 267 1161 287
rect 1237 303 1267 315
rect 1375 303 1405 367
rect 1461 303 1491 367
rect 1547 303 1577 367
rect 1633 333 1663 367
rect 1719 333 1749 367
rect 1805 333 1835 367
rect 1891 333 1921 367
rect 1633 303 1921 333
rect 1237 287 1591 303
rect 1127 253 1181 267
rect 805 237 1181 253
rect 425 215 455 237
rect 511 215 541 237
rect 597 215 627 237
rect 683 215 713 237
rect 893 215 923 237
rect 979 215 1009 237
rect 1065 215 1095 237
rect 1151 215 1181 237
rect 1237 253 1269 287
rect 1303 253 1337 287
rect 1371 253 1405 287
rect 1439 253 1473 287
rect 1507 253 1541 287
rect 1575 253 1591 287
rect 1237 237 1591 253
rect 1685 287 2091 303
rect 1685 253 1701 287
rect 1735 253 1769 287
rect 1803 253 1837 287
rect 1871 253 1905 287
rect 1939 253 1973 287
rect 2007 253 2041 287
rect 2075 253 2091 287
rect 1685 237 2091 253
rect 1237 215 1267 237
rect 1323 215 1353 237
rect 1409 215 1439 237
rect 1495 215 1525 237
rect 1685 215 1715 237
rect 1771 215 1801 237
rect 1857 215 1887 237
rect 1943 215 1973 237
rect 81 21 111 47
rect 167 21 197 47
rect 253 21 283 47
rect 339 21 369 47
rect 425 21 455 47
rect 511 21 541 47
rect 597 21 627 47
rect 683 21 713 47
rect 893 21 923 47
rect 979 21 1009 47
rect 1065 21 1095 47
rect 1151 21 1181 47
rect 1237 21 1267 47
rect 1323 21 1353 47
rect 1409 21 1439 47
rect 1495 21 1525 47
rect 1685 21 1715 47
rect 1771 21 1801 47
rect 1857 21 1887 47
rect 1943 21 1973 47
<< polycont >>
rect 47 253 81 287
rect 115 253 149 287
rect 183 253 217 287
rect 251 253 285 287
rect 319 253 353 287
rect 441 253 475 287
rect 509 253 543 287
rect 577 253 611 287
rect 645 253 679 287
rect 713 253 747 287
rect 821 253 855 287
rect 889 253 923 287
rect 957 253 991 287
rect 1025 253 1059 287
rect 1093 253 1127 287
rect 1269 253 1303 287
rect 1337 253 1371 287
rect 1405 253 1439 287
rect 1473 253 1507 287
rect 1541 253 1575 287
rect 1701 253 1735 287
rect 1769 253 1803 287
rect 1837 253 1871 287
rect 1905 253 1939 287
rect 1973 253 2007 287
rect 2041 253 2075 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 34 599 796 615
rect 34 565 50 599
rect 84 581 222 599
rect 84 565 86 581
rect 34 506 86 565
rect 220 565 222 581
rect 256 581 394 599
rect 256 565 258 581
rect 34 472 50 506
rect 84 472 86 506
rect 34 415 86 472
rect 34 381 50 415
rect 84 381 86 415
rect 34 365 86 381
rect 120 513 136 547
rect 170 513 186 547
rect 120 479 186 513
rect 120 445 136 479
rect 170 445 186 479
rect 120 411 186 445
rect 120 377 136 411
rect 170 377 186 411
rect 220 529 258 565
rect 392 565 394 581
rect 428 581 566 599
rect 428 565 430 581
rect 220 495 222 529
rect 256 495 258 529
rect 220 459 258 495
rect 220 425 222 459
rect 256 425 258 459
rect 220 409 258 425
rect 292 513 308 547
rect 342 513 358 547
rect 292 479 358 513
rect 292 445 308 479
rect 342 445 358 479
rect 292 411 358 445
rect 120 375 186 377
rect 292 377 308 411
rect 342 377 358 411
rect 392 529 430 565
rect 564 565 566 581
rect 600 581 749 599
rect 600 565 602 581
rect 392 495 394 529
rect 428 495 430 529
rect 392 459 430 495
rect 392 425 394 459
rect 428 425 430 459
rect 392 409 430 425
rect 464 513 480 547
rect 514 513 530 547
rect 464 479 530 513
rect 464 445 480 479
rect 514 445 530 479
rect 464 411 530 445
rect 292 375 358 377
rect 464 377 480 411
rect 514 377 530 411
rect 564 529 602 565
rect 736 565 749 581
rect 783 565 796 599
rect 564 495 566 529
rect 600 495 602 529
rect 564 459 602 495
rect 564 425 566 459
rect 600 425 602 459
rect 564 409 602 425
rect 636 513 652 547
rect 686 513 702 547
rect 636 479 702 513
rect 636 445 652 479
rect 686 445 702 479
rect 636 411 702 445
rect 464 375 530 377
rect 636 377 652 411
rect 686 377 702 411
rect 736 529 796 565
rect 736 495 749 529
rect 783 495 796 529
rect 736 459 796 495
rect 830 607 896 649
rect 830 573 846 607
rect 880 573 896 607
rect 830 517 896 573
rect 830 483 846 517
rect 880 483 896 517
rect 830 479 896 483
rect 930 599 968 615
rect 930 565 932 599
rect 966 565 968 599
rect 930 529 968 565
rect 930 495 932 529
rect 966 495 968 529
rect 736 425 749 459
rect 783 445 796 459
rect 930 459 968 495
rect 1002 607 1136 649
rect 1002 573 1018 607
rect 1052 573 1086 607
rect 1120 573 1136 607
rect 1002 526 1136 573
rect 1002 492 1018 526
rect 1052 492 1086 526
rect 1120 492 1136 526
rect 1002 489 1136 492
rect 1170 599 1208 615
rect 1170 565 1172 599
rect 1206 565 1208 599
rect 1170 529 1208 565
rect 1170 495 1172 529
rect 1206 495 1208 529
rect 930 445 932 459
rect 783 425 932 445
rect 966 445 968 459
rect 1170 459 1208 495
rect 1242 607 1380 649
rect 1242 573 1258 607
rect 1292 573 1330 607
rect 1364 573 1380 607
rect 1242 517 1380 573
rect 1242 483 1258 517
rect 1292 483 1330 517
rect 1364 483 1380 517
rect 1242 479 1380 483
rect 1414 599 1452 615
rect 1414 565 1416 599
rect 1450 565 1452 599
rect 1414 510 1452 565
rect 1170 445 1172 459
rect 966 425 1172 445
rect 1206 445 1208 459
rect 1414 476 1416 510
rect 1450 476 1452 510
rect 1414 445 1452 476
rect 1206 425 1452 445
rect 736 409 1452 425
rect 636 375 702 377
rect 1400 375 1416 409
rect 1450 375 1452 409
rect 1486 607 1552 649
rect 1486 573 1502 607
rect 1536 573 1552 607
rect 1486 519 1552 573
rect 1486 485 1502 519
rect 1536 485 1552 519
rect 1486 423 1552 485
rect 1486 389 1502 423
rect 1536 389 1552 423
rect 1586 599 1624 615
rect 1586 565 1588 599
rect 1622 565 1624 599
rect 1586 510 1624 565
rect 1586 476 1588 510
rect 1622 476 1624 510
rect 1586 409 1624 476
rect 120 321 1219 375
rect 1400 355 1452 375
rect 1586 375 1588 409
rect 1622 375 1624 409
rect 1658 607 1724 649
rect 1658 573 1674 607
rect 1708 573 1724 607
rect 1658 519 1724 573
rect 1658 485 1674 519
rect 1708 485 1724 519
rect 1658 423 1724 485
rect 1658 389 1674 423
rect 1708 389 1724 423
rect 1758 599 1796 615
rect 1758 565 1760 599
rect 1794 565 1796 599
rect 1758 510 1796 565
rect 1758 476 1760 510
rect 1794 476 1796 510
rect 1758 413 1796 476
rect 1586 355 1624 375
rect 1758 379 1760 413
rect 1794 379 1796 413
rect 1830 607 1896 649
rect 1830 573 1846 607
rect 1880 573 1896 607
rect 1830 519 1896 573
rect 1830 485 1846 519
rect 1880 485 1896 519
rect 1830 423 1896 485
rect 1830 389 1846 423
rect 1880 389 1896 423
rect 1930 599 1982 615
rect 1930 565 1932 599
rect 1966 565 1982 599
rect 1930 510 1982 565
rect 1930 476 1932 510
rect 1966 476 1982 510
rect 1930 413 1982 476
rect 1758 355 1796 379
rect 1930 379 1932 413
rect 1966 379 1982 413
rect 1930 355 1982 379
rect 1400 321 1982 355
rect 31 253 47 287
rect 81 253 115 287
rect 149 253 183 287
rect 217 253 251 287
rect 285 253 319 287
rect 353 253 369 287
rect 31 242 369 253
rect 415 253 441 287
rect 475 253 509 287
rect 543 253 577 287
rect 611 253 645 287
rect 679 253 713 287
rect 747 253 763 287
rect 415 242 763 253
rect 799 253 821 287
rect 855 253 889 287
rect 923 253 957 287
rect 991 253 1025 287
rect 1059 253 1093 287
rect 1127 253 1143 287
rect 799 242 1143 253
rect 1177 208 1219 321
rect 1253 253 1269 287
rect 1303 253 1337 287
rect 1371 253 1405 287
rect 1439 253 1473 287
rect 1507 253 1541 287
rect 1575 253 1601 287
rect 1253 242 1601 253
rect 1663 253 1701 287
rect 1735 253 1769 287
rect 1803 253 1837 287
rect 1871 253 1905 287
rect 1939 253 1973 287
rect 2007 253 2041 287
rect 2075 253 2091 287
rect 1663 242 2091 253
rect 20 192 416 208
rect 20 158 36 192
rect 70 174 208 192
rect 70 158 72 174
rect 20 101 72 158
rect 206 158 208 174
rect 242 174 380 192
rect 242 158 244 174
rect 20 67 36 101
rect 70 67 72 101
rect 20 51 72 67
rect 106 129 172 140
rect 106 95 122 129
rect 156 95 172 129
rect 106 17 172 95
rect 206 101 244 158
rect 378 158 380 174
rect 414 158 416 192
rect 206 67 208 101
rect 242 67 244 101
rect 206 51 244 67
rect 278 129 344 140
rect 278 95 294 129
rect 328 95 344 129
rect 278 17 344 95
rect 378 119 416 158
rect 450 202 1219 208
rect 450 168 466 202
rect 500 168 638 202
rect 672 168 934 202
rect 968 168 1106 202
rect 1140 168 1219 202
rect 450 153 1219 168
rect 1262 193 1934 208
rect 1262 159 1278 193
rect 1312 159 1450 193
rect 1484 192 1934 193
rect 1484 159 1726 192
rect 1262 158 1726 159
rect 1760 163 1898 192
rect 1760 158 1762 163
rect 1262 153 1762 158
rect 378 103 774 119
rect 378 101 552 103
rect 378 67 380 101
rect 414 69 552 101
rect 586 69 724 103
rect 758 69 774 103
rect 414 67 774 69
rect 378 51 774 67
rect 832 103 1586 119
rect 832 69 848 103
rect 882 69 1020 103
rect 1054 69 1192 103
rect 1226 69 1364 103
rect 1398 69 1536 103
rect 1570 69 1586 103
rect 832 53 1586 69
rect 1624 110 1690 119
rect 1624 76 1640 110
rect 1674 76 1690 110
rect 1624 17 1690 76
rect 1724 101 1762 153
rect 1896 158 1898 163
rect 1932 158 1934 192
rect 1724 67 1726 101
rect 1760 67 1762 101
rect 1724 51 1762 67
rect 1796 110 1862 119
rect 1796 76 1812 110
rect 1846 76 1862 110
rect 1796 17 1862 76
rect 1896 101 1934 158
rect 1896 67 1898 101
rect 1932 67 1934 101
rect 1896 51 1934 67
rect 1968 203 2034 208
rect 1968 169 1984 203
rect 2018 169 2034 203
rect 1968 93 2034 169
rect 1968 59 1984 93
rect 2018 59 2034 93
rect 1968 17 2034 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a32oi_4
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 991 168 1025 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1183 168 1217 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 898886
string GDS_START 880428
<< end >>
