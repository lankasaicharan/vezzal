magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 121 49 567 180
rect 0 0 672 49
<< scnmos >>
rect 200 70 230 154
rect 286 70 316 154
rect 372 70 402 154
rect 458 70 488 154
<< scpmoshvt >>
rect 114 367 144 619
rect 200 367 230 619
rect 286 367 316 619
rect 372 367 402 619
rect 458 367 488 619
rect 544 367 574 619
<< ndiff >>
rect 147 118 200 154
rect 147 84 155 118
rect 189 84 200 118
rect 147 70 200 84
rect 230 129 286 154
rect 230 95 241 129
rect 275 95 286 129
rect 230 70 286 95
rect 316 118 372 154
rect 316 84 327 118
rect 361 84 372 118
rect 316 70 372 84
rect 402 129 458 154
rect 402 95 413 129
rect 447 95 458 129
rect 402 70 458 95
rect 488 118 541 154
rect 488 84 499 118
rect 533 84 541 118
rect 488 70 541 84
<< pdiff >>
rect 60 599 114 619
rect 60 565 69 599
rect 103 565 114 599
rect 60 529 114 565
rect 60 495 69 529
rect 103 495 114 529
rect 60 461 114 495
rect 60 427 69 461
rect 103 427 114 461
rect 60 367 114 427
rect 144 593 200 619
rect 144 559 155 593
rect 189 559 200 593
rect 144 505 200 559
rect 144 471 155 505
rect 189 471 200 505
rect 144 417 200 471
rect 144 383 155 417
rect 189 383 200 417
rect 144 367 200 383
rect 230 599 286 619
rect 230 565 241 599
rect 275 565 286 599
rect 230 529 286 565
rect 230 495 241 529
rect 275 495 286 529
rect 230 461 286 495
rect 230 427 241 461
rect 275 427 286 461
rect 230 367 286 427
rect 316 593 372 619
rect 316 559 327 593
rect 361 559 372 593
rect 316 505 372 559
rect 316 471 327 505
rect 361 471 372 505
rect 316 417 372 471
rect 316 383 327 417
rect 361 383 372 417
rect 316 367 372 383
rect 402 599 458 619
rect 402 565 413 599
rect 447 565 458 599
rect 402 529 458 565
rect 402 495 413 529
rect 447 495 458 529
rect 402 461 458 495
rect 402 427 413 461
rect 447 427 458 461
rect 402 367 458 427
rect 488 593 544 619
rect 488 559 499 593
rect 533 559 544 593
rect 488 505 544 559
rect 488 471 499 505
rect 533 471 544 505
rect 488 417 544 471
rect 488 383 499 417
rect 533 383 544 417
rect 488 367 544 383
rect 574 599 627 619
rect 574 565 585 599
rect 619 565 627 599
rect 574 529 627 565
rect 574 495 585 529
rect 619 495 627 529
rect 574 461 627 495
rect 574 427 585 461
rect 619 427 627 461
rect 574 367 627 427
<< ndiffc >>
rect 155 84 189 118
rect 241 95 275 129
rect 327 84 361 118
rect 413 95 447 129
rect 499 84 533 118
<< pdiffc >>
rect 69 565 103 599
rect 69 495 103 529
rect 69 427 103 461
rect 155 559 189 593
rect 155 471 189 505
rect 155 383 189 417
rect 241 565 275 599
rect 241 495 275 529
rect 241 427 275 461
rect 327 559 361 593
rect 327 471 361 505
rect 327 383 361 417
rect 413 565 447 599
rect 413 495 447 529
rect 413 427 447 461
rect 499 559 533 593
rect 499 471 533 505
rect 499 383 533 417
rect 585 565 619 599
rect 585 495 619 529
rect 585 427 619 461
<< poly >>
rect 114 619 144 645
rect 200 619 230 645
rect 286 619 316 645
rect 372 619 402 645
rect 458 619 488 645
rect 544 619 574 645
rect 114 335 144 367
rect 200 335 230 367
rect 286 335 316 367
rect 372 335 402 367
rect 458 335 488 367
rect 544 335 574 367
rect 114 330 574 335
rect 114 309 592 330
rect 114 275 183 309
rect 217 275 251 309
rect 285 275 319 309
rect 353 275 387 309
rect 421 275 455 309
rect 489 275 523 309
rect 557 275 592 309
rect 114 259 592 275
rect 200 154 230 259
rect 286 154 316 259
rect 372 154 402 259
rect 458 154 488 259
rect 200 44 230 70
rect 286 44 316 70
rect 372 44 402 70
rect 458 44 488 70
<< polycont >>
rect 183 275 217 309
rect 251 275 285 309
rect 319 275 353 309
rect 387 275 421 309
rect 455 275 489 309
rect 523 275 557 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 60 599 112 615
rect 60 545 69 599
rect 103 545 112 599
rect 60 529 112 545
rect 60 495 69 529
rect 103 495 112 529
rect 60 461 112 495
rect 60 427 69 461
rect 103 427 112 461
rect 60 411 112 427
rect 147 593 198 609
rect 147 559 155 593
rect 189 559 198 593
rect 147 505 198 559
rect 147 471 155 505
rect 189 471 198 505
rect 147 417 198 471
rect 147 383 155 417
rect 189 383 198 417
rect 232 599 284 615
rect 232 565 241 599
rect 275 579 284 599
rect 232 545 242 565
rect 276 545 284 579
rect 232 529 284 545
rect 232 495 241 529
rect 275 495 284 529
rect 232 461 284 495
rect 232 427 241 461
rect 275 427 284 461
rect 232 411 284 427
rect 319 593 370 609
rect 319 559 327 593
rect 361 559 370 593
rect 319 505 370 559
rect 319 471 327 505
rect 361 471 370 505
rect 319 417 370 471
rect 147 377 198 383
rect 319 383 327 417
rect 361 383 370 417
rect 404 599 456 615
rect 404 579 413 599
rect 404 545 412 579
rect 447 565 456 599
rect 446 545 456 565
rect 404 529 456 545
rect 404 495 413 529
rect 447 495 456 529
rect 404 461 456 495
rect 404 427 413 461
rect 447 427 456 461
rect 404 411 456 427
rect 490 593 542 609
rect 490 559 499 593
rect 533 559 542 593
rect 490 505 542 559
rect 490 471 499 505
rect 533 471 542 505
rect 490 417 542 471
rect 319 377 370 383
rect 490 383 499 417
rect 533 383 542 417
rect 576 599 627 615
rect 576 565 585 599
rect 619 579 627 599
rect 576 545 586 565
rect 620 545 627 579
rect 576 529 627 545
rect 576 495 585 529
rect 619 495 627 529
rect 576 461 627 495
rect 576 427 585 461
rect 619 427 627 461
rect 576 411 627 427
rect 490 377 542 383
rect 46 343 644 377
rect 46 208 80 343
rect 114 275 183 309
rect 217 275 251 309
rect 285 275 319 309
rect 353 275 387 309
rect 421 275 455 309
rect 489 275 523 309
rect 557 275 573 309
rect 114 242 573 275
rect 607 208 644 343
rect 46 168 644 208
rect 139 118 198 134
rect 139 84 155 118
rect 189 84 198 118
rect 139 17 198 84
rect 232 129 284 168
rect 232 95 241 129
rect 275 95 284 129
rect 232 79 284 95
rect 318 118 370 134
rect 318 84 327 118
rect 361 84 370 118
rect 318 17 370 84
rect 404 129 455 168
rect 404 95 413 129
rect 447 95 455 129
rect 404 79 455 95
rect 489 118 549 134
rect 489 84 499 118
rect 533 84 549 118
rect 489 17 549 84
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 69 565 103 579
rect 69 545 103 565
rect 242 565 275 579
rect 275 565 276 579
rect 242 545 276 565
rect 412 565 413 579
rect 413 565 446 579
rect 412 545 446 565
rect 586 565 619 579
rect 619 565 620 579
rect 586 545 620 565
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 14 579 658 589
rect 14 545 69 579
rect 103 545 242 579
rect 276 545 412 579
rect 446 545 586 579
rect 620 545 658 579
rect 14 538 658 545
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 invkapwr_4
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 14 538 658 589 0 FreeSans 200 0 0 0 KAPWR
port 2 nsew power bidirectional
flabel metal1 s 337 564 337 564 0 FreeSans 200 0 0 0 KAPWR
port 2 nsew
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y
string GDS_END 3883072
string GDS_START 3875900
<< end >>
