magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 656 243 758 269
rect 449 241 1323 243
rect 1 49 1323 241
rect 0 0 1344 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 252 47 282 215
rect 338 47 368 215
rect 544 49 574 217
rect 630 49 660 217
rect 754 49 784 217
rect 840 49 870 217
rect 934 49 964 217
rect 1042 49 1072 217
rect 1128 49 1158 217
rect 1214 49 1244 217
<< scpmoshvt >>
rect 158 367 188 619
rect 244 367 274 619
rect 330 367 360 619
rect 416 367 446 619
rect 502 367 532 619
rect 668 367 698 619
rect 754 367 784 619
rect 862 367 892 619
rect 956 367 986 619
rect 1042 367 1072 619
rect 1128 367 1158 619
rect 1214 367 1244 619
<< ndiff >>
rect 682 231 732 243
rect 682 217 690 231
rect 27 171 80 215
rect 27 137 35 171
rect 69 137 80 171
rect 27 93 80 137
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 203 166 215
rect 110 169 121 203
rect 155 169 166 203
rect 110 101 166 169
rect 110 67 121 101
rect 155 67 166 101
rect 110 47 166 67
rect 196 173 252 215
rect 196 139 207 173
rect 241 139 252 173
rect 196 89 252 139
rect 196 55 207 89
rect 241 55 252 89
rect 196 47 252 55
rect 282 203 338 215
rect 282 169 293 203
rect 327 169 338 203
rect 282 101 338 169
rect 282 67 293 101
rect 327 67 338 101
rect 282 47 338 67
rect 368 172 421 215
rect 368 138 379 172
rect 413 138 421 172
rect 368 93 421 138
rect 368 59 379 93
rect 413 59 421 93
rect 368 47 421 59
rect 475 173 544 217
rect 475 139 483 173
rect 517 139 544 173
rect 475 95 544 139
rect 475 61 483 95
rect 517 61 544 95
rect 475 49 544 61
rect 574 91 630 217
rect 574 57 585 91
rect 619 57 630 91
rect 574 49 630 57
rect 660 197 690 217
rect 724 217 732 231
rect 724 197 754 217
rect 660 49 754 197
rect 784 91 840 217
rect 784 57 795 91
rect 829 57 840 91
rect 784 49 840 57
rect 870 189 934 217
rect 870 155 889 189
rect 923 155 934 189
rect 870 103 934 155
rect 870 69 889 103
rect 923 69 934 103
rect 870 49 934 69
rect 964 105 1042 217
rect 964 71 983 105
rect 1017 71 1042 105
rect 964 49 1042 71
rect 1072 178 1128 217
rect 1072 144 1083 178
rect 1117 144 1128 178
rect 1072 101 1128 144
rect 1072 67 1083 101
rect 1117 67 1128 101
rect 1072 49 1128 67
rect 1158 99 1214 217
rect 1158 65 1169 99
rect 1203 65 1214 99
rect 1158 49 1214 65
rect 1244 178 1297 217
rect 1244 144 1255 178
rect 1289 144 1297 178
rect 1244 101 1297 144
rect 1244 67 1255 101
rect 1289 67 1297 101
rect 1244 49 1297 67
<< pdiff >>
rect 105 607 158 619
rect 105 573 113 607
rect 147 573 158 607
rect 105 530 158 573
rect 105 496 113 530
rect 147 496 158 530
rect 105 453 158 496
rect 105 419 113 453
rect 147 419 158 453
rect 105 367 158 419
rect 188 599 244 619
rect 188 565 199 599
rect 233 565 244 599
rect 188 508 244 565
rect 188 474 199 508
rect 233 474 244 508
rect 188 413 244 474
rect 188 379 199 413
rect 233 379 244 413
rect 188 367 244 379
rect 274 607 330 619
rect 274 573 285 607
rect 319 573 330 607
rect 274 530 330 573
rect 274 496 285 530
rect 319 496 330 530
rect 274 453 330 496
rect 274 419 285 453
rect 319 419 330 453
rect 274 367 330 419
rect 360 599 416 619
rect 360 565 371 599
rect 405 565 416 599
rect 360 508 416 565
rect 360 474 371 508
rect 405 474 416 508
rect 360 413 416 474
rect 360 379 371 413
rect 405 379 416 413
rect 360 367 416 379
rect 446 563 502 619
rect 446 529 457 563
rect 491 529 502 563
rect 446 367 502 529
rect 532 599 668 619
rect 532 565 543 599
rect 577 565 623 599
rect 657 565 668 599
rect 532 504 668 565
rect 532 470 543 504
rect 577 470 623 504
rect 657 470 668 504
rect 532 367 668 470
rect 698 572 754 619
rect 698 538 709 572
rect 743 538 754 572
rect 698 367 754 538
rect 784 599 862 619
rect 784 565 809 599
rect 843 565 862 599
rect 784 504 862 565
rect 784 470 809 504
rect 843 470 862 504
rect 784 367 862 470
rect 892 572 956 619
rect 892 538 903 572
rect 937 538 956 572
rect 892 367 956 538
rect 986 594 1042 619
rect 986 560 997 594
rect 1031 560 1042 594
rect 986 367 1042 560
rect 1072 517 1128 619
rect 1072 483 1083 517
rect 1117 483 1128 517
rect 1072 424 1128 483
rect 1072 390 1083 424
rect 1117 390 1128 424
rect 1072 367 1128 390
rect 1158 599 1214 619
rect 1158 565 1169 599
rect 1203 565 1214 599
rect 1158 519 1214 565
rect 1158 485 1169 519
rect 1203 485 1214 519
rect 1158 436 1214 485
rect 1158 402 1169 436
rect 1203 402 1214 436
rect 1158 367 1214 402
rect 1244 607 1297 619
rect 1244 573 1255 607
rect 1289 573 1297 607
rect 1244 513 1297 573
rect 1244 479 1255 513
rect 1289 479 1297 513
rect 1244 420 1297 479
rect 1244 386 1255 420
rect 1289 386 1297 420
rect 1244 367 1297 386
<< ndiffc >>
rect 35 137 69 171
rect 35 59 69 93
rect 121 169 155 203
rect 121 67 155 101
rect 207 139 241 173
rect 207 55 241 89
rect 293 169 327 203
rect 293 67 327 101
rect 379 138 413 172
rect 379 59 413 93
rect 483 139 517 173
rect 483 61 517 95
rect 585 57 619 91
rect 690 197 724 231
rect 795 57 829 91
rect 889 155 923 189
rect 889 69 923 103
rect 983 71 1017 105
rect 1083 144 1117 178
rect 1083 67 1117 101
rect 1169 65 1203 99
rect 1255 144 1289 178
rect 1255 67 1289 101
<< pdiffc >>
rect 113 573 147 607
rect 113 496 147 530
rect 113 419 147 453
rect 199 565 233 599
rect 199 474 233 508
rect 199 379 233 413
rect 285 573 319 607
rect 285 496 319 530
rect 285 419 319 453
rect 371 565 405 599
rect 371 474 405 508
rect 371 379 405 413
rect 457 529 491 563
rect 543 565 577 599
rect 623 565 657 599
rect 543 470 577 504
rect 623 470 657 504
rect 709 538 743 572
rect 809 565 843 599
rect 809 470 843 504
rect 903 538 937 572
rect 997 560 1031 594
rect 1083 483 1117 517
rect 1083 390 1117 424
rect 1169 565 1203 599
rect 1169 485 1203 519
rect 1169 402 1203 436
rect 1255 573 1289 607
rect 1255 479 1289 513
rect 1255 386 1289 420
<< poly >>
rect 158 619 188 645
rect 244 619 274 645
rect 330 619 360 645
rect 416 619 446 645
rect 502 619 532 645
rect 668 619 698 645
rect 754 619 784 645
rect 862 619 892 645
rect 956 619 986 645
rect 1042 619 1072 645
rect 1128 619 1158 645
rect 1214 619 1244 645
rect 158 329 188 367
rect 244 329 274 367
rect 330 329 360 367
rect 416 329 446 367
rect 502 335 532 367
rect 668 335 698 367
rect 754 335 784 367
rect 862 335 892 367
rect 80 313 446 329
rect 80 279 124 313
rect 158 279 192 313
rect 226 279 260 313
rect 294 279 328 313
rect 362 279 396 313
rect 430 279 446 313
rect 80 263 446 279
rect 488 319 575 335
rect 488 285 525 319
rect 559 285 575 319
rect 488 269 575 285
rect 630 319 784 335
rect 630 285 734 319
rect 768 285 784 319
rect 630 269 784 285
rect 826 319 892 335
rect 826 285 842 319
rect 876 285 892 319
rect 956 305 986 367
rect 1042 335 1072 367
rect 1128 335 1158 367
rect 1042 319 1158 335
rect 826 269 892 285
rect 934 289 1000 305
rect 80 215 110 263
rect 166 215 196 263
rect 252 215 282 263
rect 338 215 368 263
rect 544 217 574 269
rect 630 217 660 269
rect 754 217 784 269
rect 840 217 870 269
rect 934 255 950 289
rect 984 255 1000 289
rect 934 239 1000 255
rect 1042 285 1058 319
rect 1092 285 1158 319
rect 1042 269 1158 285
rect 934 217 964 239
rect 1042 217 1072 269
rect 1128 217 1158 269
rect 1214 305 1244 367
rect 1214 289 1323 305
rect 1214 255 1273 289
rect 1307 255 1323 289
rect 1214 239 1323 255
rect 1214 217 1244 239
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 544 23 574 49
rect 630 23 660 49
rect 754 23 784 49
rect 840 23 870 49
rect 934 23 964 49
rect 1042 23 1072 49
rect 1128 23 1158 49
rect 1214 23 1244 49
<< polycont >>
rect 124 279 158 313
rect 192 279 226 313
rect 260 279 294 313
rect 328 279 362 313
rect 396 279 430 313
rect 525 285 559 319
rect 734 285 768 319
rect 842 285 876 319
rect 950 255 984 289
rect 1058 285 1092 319
rect 1273 255 1307 289
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 97 607 163 649
rect 97 573 113 607
rect 147 573 163 607
rect 97 530 163 573
rect 97 496 113 530
rect 147 496 163 530
rect 97 453 163 496
rect 97 419 113 453
rect 147 419 163 453
rect 197 599 233 615
rect 197 565 199 599
rect 197 508 233 565
rect 197 474 199 508
rect 197 413 233 474
rect 269 607 335 649
rect 269 573 285 607
rect 319 573 335 607
rect 269 530 335 573
rect 269 496 285 530
rect 319 496 335 530
rect 269 453 335 496
rect 269 419 285 453
rect 319 419 335 453
rect 369 599 407 615
rect 369 565 371 599
rect 405 565 407 599
rect 369 508 407 565
rect 441 563 507 649
rect 441 529 457 563
rect 491 529 507 563
rect 441 522 507 529
rect 541 599 659 615
rect 541 565 543 599
rect 577 565 623 599
rect 657 565 659 599
rect 369 474 371 508
rect 405 474 407 508
rect 541 504 659 565
rect 693 572 759 649
rect 693 538 709 572
rect 743 538 759 572
rect 693 522 759 538
rect 793 599 860 615
rect 793 565 809 599
rect 843 565 860 599
rect 541 488 543 504
rect 197 385 199 413
rect 17 379 199 385
rect 369 413 407 474
rect 369 385 371 413
rect 233 379 371 385
rect 405 379 407 413
rect 17 351 407 379
rect 441 470 543 488
rect 577 470 623 504
rect 657 488 659 504
rect 793 504 860 565
rect 894 572 947 649
rect 894 538 903 572
rect 937 538 947 572
rect 981 599 1205 615
rect 981 594 1169 599
rect 981 560 997 594
rect 1031 565 1169 594
rect 1203 565 1205 599
rect 1031 560 1205 565
rect 981 556 1205 560
rect 894 522 947 538
rect 793 488 809 504
rect 657 470 809 488
rect 843 488 860 504
rect 1067 517 1133 522
rect 1067 488 1083 517
rect 843 483 1083 488
rect 1117 483 1133 517
rect 843 470 1133 483
rect 441 454 1133 470
rect 17 243 74 351
rect 441 317 475 454
rect 1067 424 1133 454
rect 108 313 475 317
rect 108 279 124 313
rect 158 279 192 313
rect 226 279 260 313
rect 294 279 328 313
rect 362 279 396 313
rect 430 279 475 313
rect 509 386 892 420
rect 1067 390 1083 424
rect 1117 390 1133 424
rect 1067 386 1133 390
rect 1167 519 1205 556
rect 1167 485 1169 519
rect 1203 485 1205 519
rect 1167 436 1205 485
rect 1167 402 1169 436
rect 1203 402 1205 436
rect 1167 386 1205 402
rect 1239 607 1305 649
rect 1239 573 1255 607
rect 1289 573 1305 607
rect 1239 513 1305 573
rect 1239 479 1255 513
rect 1289 479 1305 513
rect 1239 420 1305 479
rect 1239 386 1255 420
rect 1289 386 1305 420
rect 509 319 655 386
rect 509 285 525 319
rect 559 285 655 319
rect 509 281 655 285
rect 689 319 784 352
rect 689 285 734 319
rect 768 285 784 319
rect 689 281 784 285
rect 826 319 892 386
rect 826 285 842 319
rect 876 285 892 319
rect 1042 319 1229 352
rect 108 277 475 279
rect 441 247 475 277
rect 826 269 892 285
rect 934 289 1000 305
rect 934 255 950 289
rect 984 255 1000 289
rect 1042 285 1058 319
rect 1092 285 1229 319
rect 1263 289 1327 352
rect 934 251 1000 255
rect 1263 255 1273 289
rect 1307 255 1327 289
rect 1263 251 1327 255
rect 17 209 331 243
rect 441 231 740 247
rect 934 239 1327 251
rect 441 213 690 231
rect 119 203 157 209
rect 19 171 85 175
rect 19 137 35 171
rect 69 137 85 171
rect 19 93 85 137
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 119 169 121 203
rect 155 169 157 203
rect 291 203 331 209
rect 119 101 157 169
rect 119 67 121 101
rect 155 67 157 101
rect 119 51 157 67
rect 191 173 257 175
rect 191 139 207 173
rect 241 139 257 173
rect 191 89 257 139
rect 191 55 207 89
rect 241 55 257 89
rect 191 17 257 55
rect 291 169 293 203
rect 327 169 331 203
rect 674 197 690 213
rect 724 197 740 231
rect 966 217 1327 239
rect 674 195 740 197
rect 873 189 932 205
rect 291 101 331 169
rect 291 67 293 101
rect 327 67 331 101
rect 291 51 331 67
rect 370 172 417 188
rect 370 138 379 172
rect 413 138 417 172
rect 370 93 417 138
rect 370 59 379 93
rect 413 59 417 93
rect 370 17 417 59
rect 467 173 533 179
rect 467 139 483 173
rect 517 161 533 173
rect 873 161 889 189
rect 517 155 889 161
rect 923 183 932 189
rect 923 178 1305 183
rect 923 155 1083 178
rect 517 149 1083 155
rect 517 139 933 149
rect 467 127 933 139
rect 467 95 533 127
rect 467 61 483 95
rect 517 61 533 95
rect 879 103 933 127
rect 1067 144 1083 149
rect 1117 149 1255 178
rect 1117 144 1133 149
rect 467 51 533 61
rect 569 91 845 93
rect 569 57 585 91
rect 619 57 795 91
rect 829 57 845 91
rect 569 51 845 57
rect 879 69 889 103
rect 923 69 933 103
rect 879 51 933 69
rect 967 105 1033 115
rect 967 71 983 105
rect 1017 71 1033 105
rect 967 17 1033 71
rect 1067 101 1133 144
rect 1239 144 1255 149
rect 1289 144 1305 178
rect 1067 67 1083 101
rect 1117 67 1133 101
rect 1067 51 1133 67
rect 1167 99 1205 115
rect 1167 65 1169 99
rect 1203 65 1205 99
rect 1167 17 1205 65
rect 1239 101 1305 144
rect 1239 67 1255 101
rect 1289 67 1305 101
rect 1239 51 1305 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o211a_4
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2813400
string GDS_START 2802140
<< end >>
