magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 42 49 826 248
rect 0 0 864 49
<< scpmos >>
rect 106 368 136 592
rect 196 368 226 592
rect 300 392 330 592
rect 396 392 426 592
rect 534 392 564 592
rect 630 392 660 592
rect 714 392 744 592
<< nmoslvt >>
rect 121 74 151 222
rect 207 74 237 222
rect 321 74 351 222
rect 393 74 423 222
rect 501 74 531 222
rect 609 74 639 222
rect 717 74 747 222
<< ndiff >>
rect 68 210 121 222
rect 68 176 76 210
rect 110 176 121 210
rect 68 120 121 176
rect 68 86 76 120
rect 110 86 121 120
rect 68 74 121 86
rect 151 214 207 222
rect 151 180 162 214
rect 196 180 207 214
rect 151 116 207 180
rect 151 82 162 116
rect 196 82 207 116
rect 151 74 207 82
rect 237 134 321 222
rect 237 100 269 134
rect 303 100 321 134
rect 237 74 321 100
rect 351 74 393 222
rect 423 74 501 222
rect 531 202 609 222
rect 531 168 546 202
rect 580 168 609 202
rect 531 120 609 168
rect 531 86 546 120
rect 580 86 609 120
rect 531 74 609 86
rect 639 134 717 222
rect 639 100 654 134
rect 688 100 717 134
rect 639 74 717 100
rect 747 202 800 222
rect 747 168 758 202
rect 792 168 800 202
rect 747 120 800 168
rect 747 86 758 120
rect 792 86 800 120
rect 747 74 800 86
<< pdiff >>
rect 51 564 106 592
rect 51 530 59 564
rect 93 530 106 564
rect 51 368 106 530
rect 136 412 196 592
rect 136 378 149 412
rect 183 378 196 412
rect 136 368 196 378
rect 226 564 300 592
rect 226 530 239 564
rect 273 530 300 564
rect 226 392 300 530
rect 330 584 396 592
rect 330 550 343 584
rect 377 550 396 584
rect 330 498 396 550
rect 330 464 343 498
rect 377 464 396 498
rect 330 392 396 464
rect 426 582 534 592
rect 426 548 463 582
rect 497 548 534 582
rect 426 392 534 548
rect 564 584 630 592
rect 564 550 583 584
rect 617 550 630 584
rect 564 498 630 550
rect 564 464 583 498
rect 617 464 630 498
rect 564 392 630 464
rect 660 392 714 592
rect 744 580 799 592
rect 744 546 757 580
rect 791 546 799 580
rect 744 510 799 546
rect 744 476 757 510
rect 791 476 799 510
rect 744 440 799 476
rect 744 406 757 440
rect 791 406 799 440
rect 744 392 799 406
rect 226 368 281 392
<< ndiffc >>
rect 76 176 110 210
rect 76 86 110 120
rect 162 180 196 214
rect 162 82 196 116
rect 269 100 303 134
rect 546 168 580 202
rect 546 86 580 120
rect 654 100 688 134
rect 758 168 792 202
rect 758 86 792 120
<< pdiffc >>
rect 59 530 93 564
rect 149 378 183 412
rect 239 530 273 564
rect 343 550 377 584
rect 343 464 377 498
rect 463 548 497 582
rect 583 550 617 584
rect 583 464 617 498
rect 757 546 791 580
rect 757 476 791 510
rect 757 406 791 440
<< poly >>
rect 106 592 136 618
rect 196 592 226 618
rect 300 592 330 618
rect 396 592 426 618
rect 534 592 564 618
rect 630 592 660 618
rect 714 592 744 618
rect 300 377 330 392
rect 396 377 426 392
rect 534 377 564 392
rect 630 377 660 392
rect 714 377 744 392
rect 106 353 136 368
rect 196 353 226 368
rect 103 336 139 353
rect 21 320 151 336
rect 21 286 37 320
rect 71 300 151 320
rect 193 300 229 353
rect 297 318 333 377
rect 393 356 429 377
rect 531 356 567 377
rect 393 340 459 356
rect 285 302 351 318
rect 71 286 237 300
rect 21 270 237 286
rect 121 222 151 270
rect 207 222 237 270
rect 285 268 301 302
rect 335 268 351 302
rect 285 252 351 268
rect 321 222 351 252
rect 393 306 409 340
rect 443 306 459 340
rect 393 290 459 306
rect 501 340 567 356
rect 501 306 517 340
rect 551 306 567 340
rect 627 318 663 377
rect 711 354 747 377
rect 711 341 843 354
rect 717 338 843 341
rect 501 290 567 306
rect 609 302 675 318
rect 393 222 423 290
rect 501 222 531 290
rect 609 268 625 302
rect 659 268 675 302
rect 609 252 675 268
rect 717 304 793 338
rect 827 304 843 338
rect 717 288 843 304
rect 609 222 639 252
rect 717 222 747 288
rect 121 48 151 74
rect 207 48 237 74
rect 321 48 351 74
rect 393 48 423 74
rect 501 48 531 74
rect 609 48 639 74
rect 717 48 747 74
<< polycont >>
rect 37 286 71 320
rect 301 268 335 302
rect 409 306 443 340
rect 517 306 551 340
rect 625 268 659 302
rect 793 304 827 338
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 43 564 109 649
rect 43 530 59 564
rect 93 530 109 564
rect 43 514 109 530
rect 223 564 289 649
rect 223 530 239 564
rect 273 530 289 564
rect 223 514 289 530
rect 327 584 393 596
rect 327 550 343 584
rect 377 550 393 584
rect 327 514 393 550
rect 427 582 533 649
rect 427 548 463 582
rect 497 548 533 582
rect 567 584 633 596
rect 567 550 583 584
rect 617 550 633 584
rect 567 514 633 550
rect 327 498 633 514
rect 21 446 267 480
rect 327 464 343 498
rect 377 464 583 498
rect 617 464 633 498
rect 327 458 633 464
rect 741 580 807 596
rect 741 546 757 580
rect 791 546 807 580
rect 741 510 807 546
rect 741 476 757 510
rect 791 476 807 510
rect 21 320 87 446
rect 233 424 267 446
rect 741 440 807 476
rect 741 424 757 440
rect 21 286 37 320
rect 71 286 87 320
rect 121 378 149 412
rect 183 378 199 412
rect 121 310 199 378
rect 21 270 87 286
rect 60 210 110 226
rect 60 176 76 210
rect 60 120 110 176
rect 60 86 76 120
rect 60 17 110 86
rect 146 214 199 310
rect 146 180 162 214
rect 196 180 199 214
rect 233 406 757 424
rect 791 406 807 440
rect 233 390 807 406
rect 233 218 267 390
rect 301 302 359 356
rect 335 268 359 302
rect 393 340 459 356
rect 393 306 409 340
rect 443 306 459 340
rect 393 290 459 306
rect 501 340 567 356
rect 501 306 517 340
rect 551 306 567 340
rect 501 290 567 306
rect 601 302 743 356
rect 301 252 359 268
rect 601 268 625 302
rect 659 268 743 302
rect 777 338 843 356
rect 777 304 793 338
rect 827 304 843 338
rect 777 288 843 304
rect 601 252 743 268
rect 233 202 808 218
rect 233 184 546 202
rect 146 150 199 180
rect 526 168 546 184
rect 580 184 758 202
rect 580 168 600 184
rect 146 116 212 150
rect 146 82 162 116
rect 196 82 212 116
rect 146 70 212 82
rect 246 134 326 150
rect 246 100 269 134
rect 303 100 326 134
rect 246 17 326 100
rect 526 120 600 168
rect 742 168 758 184
rect 792 168 808 202
rect 526 86 546 120
rect 580 86 600 120
rect 526 70 600 86
rect 634 134 708 150
rect 634 100 654 134
rect 688 100 708 134
rect 634 17 708 100
rect 742 120 808 168
rect 742 86 758 120
rect 792 86 808 120
rect 742 70 808 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a311o_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 1813012
string GDS_START 1805796
<< end >>
