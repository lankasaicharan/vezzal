magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 331 1958 704
rect 195 323 1061 331
<< pwell >>
rect 482 254 772 265
rect 4 191 772 254
rect 1075 248 1637 254
rect 1075 191 1917 248
rect 4 49 1917 191
rect 0 0 1920 49
<< scnmos >>
rect 83 144 113 228
rect 276 144 306 228
rect 362 144 392 228
rect 561 155 591 239
rect 647 155 677 239
rect 870 81 900 165
rect 956 81 986 165
rect 1154 60 1184 228
rect 1226 60 1256 228
rect 1334 60 1364 228
rect 1420 60 1450 228
rect 1528 144 1558 228
rect 1722 54 1752 222
rect 1808 54 1838 222
<< scpmoshvt >>
rect 89 473 119 601
rect 284 359 314 487
rect 401 359 431 487
rect 659 359 689 443
rect 764 359 794 487
rect 836 359 866 487
rect 942 359 972 443
rect 1154 367 1184 619
rect 1240 367 1270 619
rect 1334 367 1364 619
rect 1420 367 1450 619
rect 1525 367 1555 495
rect 1722 367 1752 619
rect 1808 367 1838 619
<< ndiff >>
rect 30 200 83 228
rect 30 166 38 200
rect 72 166 83 200
rect 30 144 83 166
rect 113 190 166 228
rect 113 156 124 190
rect 158 156 166 190
rect 113 144 166 156
rect 223 203 276 228
rect 223 169 231 203
rect 265 169 276 203
rect 223 144 276 169
rect 306 192 362 228
rect 306 158 317 192
rect 351 158 362 192
rect 306 144 362 158
rect 392 192 445 228
rect 392 158 403 192
rect 437 158 445 192
rect 392 144 445 158
rect 508 214 561 239
rect 508 180 516 214
rect 550 180 561 214
rect 508 155 561 180
rect 591 231 647 239
rect 591 197 602 231
rect 636 197 647 231
rect 591 155 647 197
rect 677 227 746 239
rect 677 193 704 227
rect 738 193 746 227
rect 677 155 746 193
rect 1101 216 1154 228
rect 1101 182 1109 216
rect 1143 182 1154 216
rect 813 157 870 165
rect 813 123 825 157
rect 859 123 870 157
rect 813 81 870 123
rect 900 137 956 165
rect 900 103 911 137
rect 945 103 956 137
rect 900 81 956 103
rect 986 141 1039 165
rect 986 107 997 141
rect 1031 107 1039 141
rect 986 81 1039 107
rect 1101 106 1154 182
rect 1101 72 1109 106
rect 1143 72 1154 106
rect 1101 60 1154 72
rect 1184 60 1226 228
rect 1256 208 1334 228
rect 1256 174 1275 208
rect 1309 174 1334 208
rect 1256 106 1334 174
rect 1256 72 1275 106
rect 1309 72 1334 106
rect 1256 60 1334 72
rect 1364 215 1420 228
rect 1364 181 1375 215
rect 1409 181 1420 215
rect 1364 118 1420 181
rect 1364 84 1375 118
rect 1409 84 1420 118
rect 1364 60 1420 84
rect 1450 215 1528 228
rect 1450 181 1483 215
rect 1517 181 1528 215
rect 1450 144 1528 181
rect 1558 216 1611 228
rect 1558 182 1569 216
rect 1603 182 1611 216
rect 1558 144 1611 182
rect 1450 106 1503 144
rect 1665 135 1722 222
rect 1450 72 1461 106
rect 1495 72 1503 106
rect 1450 60 1503 72
rect 1665 101 1673 135
rect 1707 101 1722 135
rect 1665 54 1722 101
rect 1752 210 1808 222
rect 1752 176 1763 210
rect 1797 176 1808 210
rect 1752 101 1808 176
rect 1752 67 1763 101
rect 1797 67 1808 101
rect 1752 54 1808 67
rect 1838 210 1891 222
rect 1838 176 1849 210
rect 1883 176 1891 210
rect 1838 100 1891 176
rect 1838 66 1849 100
rect 1883 66 1891 100
rect 1838 54 1891 66
<< pdiff >>
rect 36 574 89 601
rect 36 540 44 574
rect 78 540 89 574
rect 36 473 89 540
rect 119 589 172 601
rect 119 555 130 589
rect 164 555 172 589
rect 119 521 172 555
rect 119 487 130 521
rect 164 487 172 521
rect 119 473 172 487
rect 231 473 284 487
rect 231 439 239 473
rect 273 439 284 473
rect 231 405 284 439
rect 231 371 239 405
rect 273 371 284 405
rect 231 359 284 371
rect 314 434 401 487
rect 314 400 338 434
rect 372 400 401 434
rect 314 359 401 400
rect 431 473 484 487
rect 431 439 442 473
rect 476 439 484 473
rect 431 405 484 439
rect 431 371 442 405
rect 476 371 484 405
rect 431 359 484 371
rect 711 461 764 487
rect 711 443 719 461
rect 606 407 659 443
rect 606 373 614 407
rect 648 373 659 407
rect 606 359 659 373
rect 689 427 719 443
rect 753 427 764 461
rect 689 359 764 427
rect 794 359 836 487
rect 866 466 920 487
rect 866 432 878 466
rect 912 443 920 466
rect 912 432 942 443
rect 866 359 942 432
rect 972 418 1025 443
rect 972 384 983 418
rect 1017 384 1025 418
rect 972 359 1025 384
rect 1101 583 1154 619
rect 1101 549 1109 583
rect 1143 549 1154 583
rect 1101 367 1154 549
rect 1184 599 1240 619
rect 1184 565 1195 599
rect 1229 565 1240 599
rect 1184 515 1240 565
rect 1184 481 1195 515
rect 1229 481 1240 515
rect 1184 367 1240 481
rect 1270 571 1334 619
rect 1270 537 1285 571
rect 1319 537 1334 571
rect 1270 367 1334 537
rect 1364 413 1420 619
rect 1364 379 1375 413
rect 1409 379 1420 413
rect 1364 367 1420 379
rect 1450 571 1503 619
rect 1450 537 1461 571
rect 1495 537 1503 571
rect 1450 495 1503 537
rect 1669 607 1722 619
rect 1669 573 1677 607
rect 1711 573 1722 607
rect 1669 539 1722 573
rect 1669 505 1677 539
rect 1711 505 1722 539
rect 1450 367 1525 495
rect 1555 481 1608 495
rect 1555 447 1566 481
rect 1600 447 1608 481
rect 1555 413 1608 447
rect 1555 379 1566 413
rect 1600 379 1608 413
rect 1555 367 1608 379
rect 1669 471 1722 505
rect 1669 437 1677 471
rect 1711 437 1722 471
rect 1669 367 1722 437
rect 1752 599 1808 619
rect 1752 565 1763 599
rect 1797 565 1808 599
rect 1752 500 1808 565
rect 1752 466 1763 500
rect 1797 466 1808 500
rect 1752 413 1808 466
rect 1752 379 1763 413
rect 1797 379 1808 413
rect 1752 367 1808 379
rect 1838 607 1891 619
rect 1838 573 1849 607
rect 1883 573 1891 607
rect 1838 507 1891 573
rect 1838 473 1849 507
rect 1883 473 1891 507
rect 1838 413 1891 473
rect 1838 379 1849 413
rect 1883 379 1891 413
rect 1838 367 1891 379
<< ndiffc >>
rect 38 166 72 200
rect 124 156 158 190
rect 231 169 265 203
rect 317 158 351 192
rect 403 158 437 192
rect 516 180 550 214
rect 602 197 636 231
rect 704 193 738 227
rect 1109 182 1143 216
rect 825 123 859 157
rect 911 103 945 137
rect 997 107 1031 141
rect 1109 72 1143 106
rect 1275 174 1309 208
rect 1275 72 1309 106
rect 1375 181 1409 215
rect 1375 84 1409 118
rect 1483 181 1517 215
rect 1569 182 1603 216
rect 1461 72 1495 106
rect 1673 101 1707 135
rect 1763 176 1797 210
rect 1763 67 1797 101
rect 1849 176 1883 210
rect 1849 66 1883 100
<< pdiffc >>
rect 44 540 78 574
rect 130 555 164 589
rect 130 487 164 521
rect 239 439 273 473
rect 239 371 273 405
rect 338 400 372 434
rect 442 439 476 473
rect 442 371 476 405
rect 614 373 648 407
rect 719 427 753 461
rect 878 432 912 466
rect 983 384 1017 418
rect 1109 549 1143 583
rect 1195 565 1229 599
rect 1195 481 1229 515
rect 1285 537 1319 571
rect 1375 379 1409 413
rect 1461 537 1495 571
rect 1677 573 1711 607
rect 1677 505 1711 539
rect 1566 447 1600 481
rect 1566 379 1600 413
rect 1677 437 1711 471
rect 1763 565 1797 599
rect 1763 466 1797 500
rect 1763 379 1797 413
rect 1849 573 1883 607
rect 1849 473 1883 507
rect 1849 379 1883 413
<< poly >>
rect 89 601 119 627
rect 238 605 304 621
rect 238 571 254 605
rect 288 591 304 605
rect 760 605 1086 621
rect 1154 619 1184 645
rect 1240 619 1270 645
rect 1334 619 1364 645
rect 1420 619 1450 645
rect 1722 619 1752 645
rect 1808 619 1838 645
rect 288 571 689 591
rect 238 561 689 571
rect 238 555 304 561
rect 284 487 314 513
rect 401 487 431 513
rect 89 384 119 473
rect 44 368 119 384
rect 44 334 60 368
rect 94 334 119 368
rect 44 300 119 334
rect 284 316 314 359
rect 401 316 431 359
rect 44 266 60 300
rect 94 266 119 300
rect 44 250 119 266
rect 161 300 314 316
rect 161 266 177 300
rect 211 266 314 300
rect 161 250 314 266
rect 356 300 431 316
rect 356 266 372 300
rect 406 266 431 300
rect 356 250 431 266
rect 83 228 113 250
rect 276 228 306 250
rect 362 228 392 250
rect 561 239 591 561
rect 659 443 689 561
rect 760 571 776 605
rect 810 591 1086 605
rect 810 571 826 591
rect 760 555 826 571
rect 764 487 794 513
rect 836 487 866 513
rect 942 443 972 469
rect 659 333 689 359
rect 764 291 794 359
rect 647 261 794 291
rect 647 239 677 261
rect 836 217 866 359
rect 942 318 972 359
rect 1056 345 1086 591
rect 1525 495 1555 521
rect 1154 345 1184 367
rect 942 302 1008 318
rect 1056 315 1184 345
rect 1240 316 1270 367
rect 1334 331 1364 367
rect 1420 331 1450 367
rect 1525 331 1555 367
rect 942 268 958 302
rect 992 268 1008 302
rect 942 252 1008 268
rect 761 187 900 217
rect 83 118 113 144
rect 276 118 306 144
rect 362 118 392 144
rect 561 129 591 155
rect 162 90 228 106
rect 162 56 178 90
rect 212 70 228 90
rect 647 70 677 155
rect 761 103 791 187
rect 870 165 900 187
rect 956 165 986 252
rect 1154 228 1184 315
rect 1226 300 1292 316
rect 1226 266 1242 300
rect 1276 266 1292 300
rect 1226 250 1292 266
rect 1334 315 1631 331
rect 1722 328 1752 367
rect 1334 281 1445 315
rect 1479 281 1513 315
rect 1547 281 1581 315
rect 1615 281 1631 315
rect 1334 265 1631 281
rect 1673 312 1752 328
rect 1673 278 1689 312
rect 1723 292 1752 312
rect 1808 292 1838 367
rect 1723 278 1838 292
rect 1226 228 1256 250
rect 1334 228 1364 265
rect 1420 228 1450 265
rect 1528 228 1558 265
rect 1673 262 1838 278
rect 212 56 677 70
rect 162 40 677 56
rect 725 87 791 103
rect 725 53 741 87
rect 775 53 791 87
rect 870 55 900 81
rect 956 55 986 81
rect 1722 222 1752 262
rect 1808 222 1838 262
rect 1528 118 1558 144
rect 725 37 791 53
rect 1154 34 1184 60
rect 1226 34 1256 60
rect 1334 34 1364 60
rect 1420 34 1450 60
rect 1722 28 1752 54
rect 1808 28 1838 54
<< polycont >>
rect 254 571 288 605
rect 60 334 94 368
rect 60 266 94 300
rect 177 266 211 300
rect 372 266 406 300
rect 776 571 810 605
rect 958 268 992 302
rect 178 56 212 90
rect 1242 266 1276 300
rect 1445 281 1479 315
rect 1513 281 1547 315
rect 1581 281 1615 315
rect 1689 278 1723 312
rect 741 53 775 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 28 574 94 649
rect 28 540 44 574
rect 78 540 94 574
rect 28 532 94 540
rect 128 605 304 615
rect 128 589 254 605
rect 128 555 130 589
rect 164 571 254 589
rect 288 571 304 605
rect 164 555 304 571
rect 128 521 180 555
rect 17 368 94 498
rect 17 334 60 368
rect 17 300 94 334
rect 17 266 60 300
rect 17 242 94 266
rect 128 487 130 521
rect 164 487 180 521
rect 128 316 180 487
rect 223 473 281 489
rect 223 439 239 473
rect 273 439 281 473
rect 223 405 281 439
rect 223 371 239 405
rect 273 371 281 405
rect 338 434 388 649
rect 760 571 776 605
rect 810 571 826 605
rect 760 519 826 571
rect 372 400 388 434
rect 338 384 388 400
rect 426 473 492 489
rect 426 439 442 473
rect 476 439 492 473
rect 426 405 492 439
rect 426 384 442 405
rect 223 355 281 371
rect 128 300 211 316
rect 128 266 177 300
rect 128 250 211 266
rect 22 200 88 208
rect 128 206 164 250
rect 247 216 281 355
rect 440 371 442 384
rect 476 371 492 405
rect 440 355 492 371
rect 540 461 826 519
rect 540 457 719 461
rect 315 300 406 350
rect 315 266 372 300
rect 315 242 406 266
rect 22 166 38 200
rect 72 166 88 200
rect 22 17 88 166
rect 122 190 164 206
rect 122 156 124 190
rect 158 156 164 190
rect 122 140 164 156
rect 215 203 281 216
rect 440 208 476 355
rect 540 319 574 457
rect 703 427 719 457
rect 753 457 826 461
rect 862 466 928 649
rect 1105 583 1153 649
rect 1105 549 1109 583
rect 1143 549 1153 583
rect 1105 533 1153 549
rect 1187 599 1235 615
rect 1187 565 1195 599
rect 1229 565 1235 599
rect 1187 515 1235 565
rect 1269 571 1335 649
rect 1269 537 1285 571
rect 1319 537 1335 571
rect 1269 533 1335 537
rect 1445 571 1511 649
rect 1445 537 1461 571
rect 1495 537 1511 571
rect 1445 533 1511 537
rect 1661 607 1725 649
rect 1661 573 1677 607
rect 1711 573 1725 607
rect 1661 539 1725 573
rect 1187 499 1195 515
rect 753 427 769 457
rect 703 423 769 427
rect 862 432 878 466
rect 912 432 928 466
rect 1113 481 1195 499
rect 1229 499 1235 515
rect 1661 505 1677 539
rect 1711 505 1725 539
rect 1229 481 1516 499
rect 1113 465 1516 481
rect 862 423 928 432
rect 608 407 664 423
rect 608 373 614 407
rect 648 389 664 407
rect 967 418 1033 434
rect 967 389 983 418
rect 648 384 983 389
rect 1017 384 1033 418
rect 648 373 1033 384
rect 608 355 1033 373
rect 1113 321 1147 465
rect 540 285 652 319
rect 586 231 652 285
rect 942 302 1147 321
rect 942 268 958 302
rect 992 268 1147 302
rect 942 265 1147 268
rect 215 169 231 203
rect 265 169 281 203
rect 215 90 281 169
rect 162 56 178 90
rect 212 56 281 90
rect 315 192 359 208
rect 315 158 317 192
rect 351 158 359 192
rect 315 17 359 158
rect 393 192 476 208
rect 393 158 403 192
rect 437 158 476 192
rect 393 140 476 158
rect 442 89 476 140
rect 510 214 552 230
rect 510 180 516 214
rect 550 180 552 214
rect 586 197 602 231
rect 636 197 652 231
rect 586 193 652 197
rect 688 227 1047 231
rect 688 193 704 227
rect 738 193 1047 227
rect 510 159 552 180
rect 510 157 875 159
rect 510 123 825 157
rect 859 123 875 157
rect 909 137 953 153
rect 909 103 911 137
rect 945 103 953 137
rect 442 87 791 89
rect 442 53 741 87
rect 775 53 791 87
rect 442 51 791 53
rect 909 17 953 103
rect 987 141 1047 193
rect 987 107 997 141
rect 1031 107 1047 141
rect 987 91 1047 107
rect 1093 216 1147 265
rect 1183 300 1325 431
rect 1183 266 1242 300
rect 1276 266 1325 300
rect 1183 242 1325 266
rect 1359 413 1411 431
rect 1359 379 1375 413
rect 1409 379 1411 413
rect 1359 363 1411 379
rect 1093 182 1109 216
rect 1143 182 1147 216
rect 1359 231 1393 363
rect 1445 315 1516 465
rect 1550 481 1604 497
rect 1550 447 1566 481
rect 1600 447 1604 481
rect 1550 413 1604 447
rect 1661 471 1725 505
rect 1661 437 1677 471
rect 1711 437 1725 471
rect 1661 421 1725 437
rect 1759 599 1807 615
rect 1759 565 1763 599
rect 1797 565 1807 599
rect 1759 500 1807 565
rect 1759 466 1763 500
rect 1797 466 1807 500
rect 1550 379 1566 413
rect 1600 385 1604 413
rect 1759 413 1807 466
rect 1600 379 1723 385
rect 1550 351 1723 379
rect 1429 281 1445 315
rect 1479 281 1513 315
rect 1547 281 1581 315
rect 1615 281 1631 315
rect 1673 312 1723 351
rect 1673 278 1689 312
rect 1359 215 1413 231
rect 1093 106 1147 182
rect 1093 72 1109 106
rect 1143 72 1147 106
rect 1093 56 1147 72
rect 1259 174 1275 208
rect 1309 174 1325 208
rect 1259 106 1325 174
rect 1259 72 1275 106
rect 1309 72 1325 106
rect 1259 17 1325 72
rect 1359 181 1375 215
rect 1409 181 1413 215
rect 1359 118 1413 181
rect 1359 84 1375 118
rect 1409 84 1413 118
rect 1359 68 1413 84
rect 1457 215 1519 231
rect 1673 223 1723 278
rect 1457 181 1483 215
rect 1517 181 1519 215
rect 1457 106 1519 181
rect 1553 216 1723 223
rect 1553 182 1569 216
rect 1603 182 1723 216
rect 1553 177 1723 182
rect 1759 379 1763 413
rect 1797 379 1807 413
rect 1759 210 1807 379
rect 1841 607 1899 649
rect 1841 573 1849 607
rect 1883 573 1899 607
rect 1841 507 1899 573
rect 1841 473 1849 507
rect 1883 473 1899 507
rect 1841 413 1899 473
rect 1841 379 1849 413
rect 1883 379 1899 413
rect 1841 363 1899 379
rect 1759 176 1763 210
rect 1797 176 1807 210
rect 1457 72 1461 106
rect 1495 72 1519 106
rect 1457 17 1519 72
rect 1657 135 1723 143
rect 1657 101 1673 135
rect 1707 101 1723 135
rect 1657 17 1723 101
rect 1759 101 1807 176
rect 1759 67 1763 101
rect 1797 67 1807 101
rect 1759 51 1807 67
rect 1841 210 1899 226
rect 1841 176 1849 210
rect 1883 176 1899 210
rect 1841 100 1899 176
rect 1841 66 1849 100
rect 1883 66 1899 100
rect 1841 17 1899 66
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrbn_2
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1375 168 1409 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1759 316 1793 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1759 390 1793 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1759 464 1793 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1759 538 1793 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1183 390 1217 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6217918
string GDS_START 6202534
<< end >>
