magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 47 49 1339 241
rect 0 0 1344 49
<< scnmos >>
rect 126 47 156 215
rect 216 47 246 215
rect 302 47 332 215
rect 388 47 418 215
rect 474 47 504 215
rect 628 47 658 215
rect 714 47 744 215
rect 800 47 830 215
rect 886 47 916 215
rect 972 47 1002 215
rect 1058 47 1088 215
rect 1144 47 1174 215
rect 1230 47 1260 215
<< scpmoshvt >>
rect 86 367 116 619
rect 276 367 306 619
rect 362 367 392 619
rect 448 367 478 619
rect 534 367 564 619
rect 626 367 656 619
rect 714 367 744 619
rect 800 367 830 619
rect 886 367 916 619
rect 972 367 1002 619
rect 1058 367 1088 619
rect 1144 367 1174 619
rect 1230 367 1260 619
<< ndiff >>
rect 73 192 126 215
rect 73 158 81 192
rect 115 158 126 192
rect 73 101 126 158
rect 73 67 81 101
rect 115 67 126 101
rect 73 47 126 67
rect 156 129 216 215
rect 156 95 171 129
rect 205 95 216 129
rect 156 47 216 95
rect 246 124 302 215
rect 246 90 257 124
rect 291 90 302 124
rect 246 47 302 90
rect 332 157 388 215
rect 332 123 343 157
rect 377 123 388 157
rect 332 89 388 123
rect 332 55 343 89
rect 377 55 388 89
rect 332 47 388 55
rect 418 203 474 215
rect 418 169 429 203
rect 463 169 474 203
rect 418 101 474 169
rect 418 67 429 101
rect 463 67 474 101
rect 418 47 474 67
rect 504 89 628 215
rect 504 55 515 89
rect 549 55 583 89
rect 617 55 628 89
rect 504 47 628 55
rect 658 101 714 215
rect 658 67 669 101
rect 703 67 714 101
rect 658 47 714 67
rect 744 175 800 215
rect 744 141 755 175
rect 789 141 800 175
rect 744 47 800 141
rect 830 101 886 215
rect 830 67 841 101
rect 875 67 886 101
rect 830 47 886 67
rect 916 175 972 215
rect 916 141 927 175
rect 961 141 972 175
rect 916 47 972 141
rect 1002 165 1058 215
rect 1002 131 1013 165
rect 1047 131 1058 165
rect 1002 97 1058 131
rect 1002 63 1013 97
rect 1047 63 1058 97
rect 1002 47 1058 63
rect 1088 97 1144 215
rect 1088 63 1099 97
rect 1133 63 1144 97
rect 1088 47 1144 63
rect 1174 192 1230 215
rect 1174 158 1185 192
rect 1219 158 1230 192
rect 1174 101 1230 158
rect 1174 67 1185 101
rect 1219 67 1230 101
rect 1174 47 1230 67
rect 1260 192 1313 215
rect 1260 158 1271 192
rect 1305 158 1313 192
rect 1260 93 1313 158
rect 1260 59 1271 93
rect 1305 59 1313 93
rect 1260 47 1313 59
<< pdiff >>
rect 33 599 86 619
rect 33 565 41 599
rect 75 565 86 599
rect 33 508 86 565
rect 33 474 41 508
rect 75 474 86 508
rect 33 418 86 474
rect 33 384 41 418
rect 75 384 86 418
rect 33 367 86 384
rect 116 607 169 619
rect 116 573 127 607
rect 161 573 169 607
rect 116 486 169 573
rect 116 452 127 486
rect 161 452 169 486
rect 116 367 169 452
rect 223 599 276 619
rect 223 565 231 599
rect 265 565 276 599
rect 223 502 276 565
rect 223 468 231 502
rect 265 468 276 502
rect 223 367 276 468
rect 306 481 362 619
rect 306 447 317 481
rect 351 447 362 481
rect 306 413 362 447
rect 306 379 317 413
rect 351 379 362 413
rect 306 367 362 379
rect 392 611 448 619
rect 392 577 403 611
rect 437 577 448 611
rect 392 543 448 577
rect 392 509 403 543
rect 437 509 448 543
rect 392 475 448 509
rect 392 441 403 475
rect 437 441 448 475
rect 392 367 448 441
rect 478 517 534 619
rect 478 483 489 517
rect 523 483 534 517
rect 478 413 534 483
rect 478 379 489 413
rect 523 379 534 413
rect 478 367 534 379
rect 564 599 626 619
rect 564 565 581 599
rect 615 565 626 599
rect 564 517 626 565
rect 564 483 581 517
rect 615 483 626 517
rect 564 449 626 483
rect 564 415 581 449
rect 615 415 626 449
rect 564 367 626 415
rect 656 587 714 619
rect 656 553 669 587
rect 703 553 714 587
rect 656 492 714 553
rect 656 458 669 492
rect 703 458 714 492
rect 656 367 714 458
rect 744 583 800 619
rect 744 549 755 583
rect 789 549 800 583
rect 744 367 800 549
rect 830 492 886 619
rect 830 458 841 492
rect 875 458 886 492
rect 830 367 886 458
rect 916 597 972 619
rect 916 563 927 597
rect 961 563 972 597
rect 916 517 972 563
rect 916 483 927 517
rect 961 483 972 517
rect 916 434 972 483
rect 916 400 927 434
rect 961 400 972 434
rect 916 367 972 400
rect 1002 607 1058 619
rect 1002 573 1013 607
rect 1047 573 1058 607
rect 1002 492 1058 573
rect 1002 458 1013 492
rect 1047 458 1058 492
rect 1002 367 1058 458
rect 1088 599 1144 619
rect 1088 565 1099 599
rect 1133 565 1144 599
rect 1088 506 1144 565
rect 1088 472 1099 506
rect 1133 472 1144 506
rect 1088 413 1144 472
rect 1088 379 1099 413
rect 1133 379 1144 413
rect 1088 367 1144 379
rect 1174 607 1230 619
rect 1174 573 1185 607
rect 1219 573 1230 607
rect 1174 529 1230 573
rect 1174 495 1185 529
rect 1219 495 1230 529
rect 1174 455 1230 495
rect 1174 421 1185 455
rect 1219 421 1230 455
rect 1174 367 1230 421
rect 1260 599 1313 619
rect 1260 565 1271 599
rect 1305 565 1313 599
rect 1260 512 1313 565
rect 1260 478 1271 512
rect 1305 478 1313 512
rect 1260 413 1313 478
rect 1260 379 1271 413
rect 1305 379 1313 413
rect 1260 367 1313 379
<< ndiffc >>
rect 81 158 115 192
rect 81 67 115 101
rect 171 95 205 129
rect 257 90 291 124
rect 343 123 377 157
rect 343 55 377 89
rect 429 169 463 203
rect 429 67 463 101
rect 515 55 549 89
rect 583 55 617 89
rect 669 67 703 101
rect 755 141 789 175
rect 841 67 875 101
rect 927 141 961 175
rect 1013 131 1047 165
rect 1013 63 1047 97
rect 1099 63 1133 97
rect 1185 158 1219 192
rect 1185 67 1219 101
rect 1271 158 1305 192
rect 1271 59 1305 93
<< pdiffc >>
rect 41 565 75 599
rect 41 474 75 508
rect 41 384 75 418
rect 127 573 161 607
rect 127 452 161 486
rect 231 565 265 599
rect 231 468 265 502
rect 317 447 351 481
rect 317 379 351 413
rect 403 577 437 611
rect 403 509 437 543
rect 403 441 437 475
rect 489 483 523 517
rect 489 379 523 413
rect 581 565 615 599
rect 581 483 615 517
rect 581 415 615 449
rect 669 553 703 587
rect 669 458 703 492
rect 755 549 789 583
rect 841 458 875 492
rect 927 563 961 597
rect 927 483 961 517
rect 927 400 961 434
rect 1013 573 1047 607
rect 1013 458 1047 492
rect 1099 565 1133 599
rect 1099 472 1133 506
rect 1099 379 1133 413
rect 1185 573 1219 607
rect 1185 495 1219 529
rect 1185 421 1219 455
rect 1271 565 1305 599
rect 1271 478 1305 512
rect 1271 379 1305 413
<< poly >>
rect 86 619 116 645
rect 276 619 306 645
rect 362 619 392 645
rect 448 619 478 645
rect 534 619 564 645
rect 626 619 656 645
rect 714 619 744 645
rect 800 619 830 645
rect 886 619 916 645
rect 972 619 1002 645
rect 1058 619 1088 645
rect 1144 619 1174 645
rect 1230 619 1260 645
rect 86 303 116 367
rect 276 325 306 367
rect 362 325 392 367
rect 448 325 478 367
rect 534 325 564 367
rect 205 309 564 325
rect 86 287 156 303
rect 86 253 102 287
rect 136 253 156 287
rect 205 275 221 309
rect 255 275 289 309
rect 323 275 357 309
rect 391 275 425 309
rect 459 291 564 309
rect 626 303 656 367
rect 714 335 744 367
rect 800 335 830 367
rect 886 335 916 367
rect 972 335 1002 367
rect 714 319 1002 335
rect 459 275 504 291
rect 205 255 504 275
rect 86 237 156 253
rect 126 215 156 237
rect 216 215 246 255
rect 302 215 332 255
rect 388 215 418 255
rect 474 215 504 255
rect 606 287 672 303
rect 606 253 622 287
rect 656 253 672 287
rect 606 237 672 253
rect 714 285 748 319
rect 782 285 816 319
rect 850 285 884 319
rect 918 285 952 319
rect 986 285 1002 319
rect 714 269 1002 285
rect 628 215 658 237
rect 714 215 744 269
rect 800 215 830 269
rect 886 215 916 269
rect 972 215 1002 269
rect 1058 303 1088 367
rect 1144 303 1174 367
rect 1230 303 1260 367
rect 1058 287 1289 303
rect 1058 253 1103 287
rect 1137 253 1171 287
rect 1205 253 1239 287
rect 1273 253 1289 287
rect 1058 237 1289 253
rect 1058 215 1088 237
rect 1144 215 1174 237
rect 1230 215 1260 237
rect 126 21 156 47
rect 216 21 246 47
rect 302 21 332 47
rect 388 21 418 47
rect 474 21 504 47
rect 628 21 658 47
rect 714 21 744 47
rect 800 21 830 47
rect 886 21 916 47
rect 972 21 1002 47
rect 1058 21 1088 47
rect 1144 21 1174 47
rect 1230 21 1260 47
<< polycont >>
rect 102 253 136 287
rect 221 275 255 309
rect 289 275 323 309
rect 357 275 391 309
rect 425 275 459 309
rect 622 253 656 287
rect 748 285 782 319
rect 816 285 850 319
rect 884 285 918 319
rect 952 285 986 319
rect 1103 253 1137 287
rect 1171 253 1205 287
rect 1239 253 1273 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 25 599 77 615
rect 25 565 41 599
rect 75 565 77 599
rect 25 508 77 565
rect 25 474 41 508
rect 75 474 77 508
rect 25 418 77 474
rect 111 607 177 649
rect 111 573 127 607
rect 161 573 177 607
rect 111 486 177 573
rect 111 452 127 486
rect 161 452 177 486
rect 215 611 619 615
rect 215 599 403 611
rect 215 565 231 599
rect 265 577 403 599
rect 437 599 619 611
rect 437 577 581 599
rect 265 567 581 577
rect 265 565 453 567
rect 215 543 453 565
rect 215 533 403 543
rect 215 502 267 533
rect 215 468 231 502
rect 265 468 267 502
rect 387 509 403 533
rect 437 509 453 543
rect 579 565 581 567
rect 615 565 619 599
rect 215 452 267 468
rect 301 481 353 497
rect 301 447 317 481
rect 351 447 353 481
rect 25 384 41 418
rect 75 384 239 418
rect 31 287 161 350
rect 31 253 102 287
rect 136 253 161 287
rect 31 242 161 253
rect 195 309 239 384
rect 301 413 353 447
rect 387 475 453 509
rect 387 441 403 475
rect 437 441 453 475
rect 487 517 545 533
rect 487 483 489 517
rect 523 483 545 517
rect 301 379 317 413
rect 351 407 353 413
rect 487 413 545 483
rect 487 407 489 413
rect 351 379 489 407
rect 523 379 545 413
rect 579 517 619 565
rect 579 483 581 517
rect 615 483 619 517
rect 579 449 619 483
rect 653 587 719 649
rect 653 553 669 587
rect 703 553 719 587
rect 653 499 719 553
rect 753 597 963 613
rect 753 583 927 597
rect 753 549 755 583
rect 789 563 927 583
rect 961 563 963 597
rect 789 549 963 563
rect 753 533 963 549
rect 925 517 963 533
rect 653 492 891 499
rect 653 458 669 492
rect 703 458 841 492
rect 875 458 891 492
rect 653 452 891 458
rect 925 483 927 517
rect 961 483 963 517
rect 579 415 581 449
rect 615 418 619 449
rect 925 434 963 483
rect 997 607 1063 649
rect 997 573 1013 607
rect 1047 573 1063 607
rect 997 492 1063 573
rect 997 458 1013 492
rect 1047 458 1063 492
rect 997 452 1063 458
rect 1097 599 1133 615
rect 1097 565 1099 599
rect 1097 506 1133 565
rect 1097 472 1099 506
rect 925 418 927 434
rect 615 415 927 418
rect 579 400 927 415
rect 961 418 963 434
rect 1097 418 1133 472
rect 1169 607 1235 649
rect 1169 573 1185 607
rect 1219 573 1235 607
rect 1169 529 1235 573
rect 1169 495 1185 529
rect 1219 495 1235 529
rect 1169 455 1235 495
rect 1169 421 1185 455
rect 1219 421 1235 455
rect 1269 599 1321 615
rect 1269 565 1271 599
rect 1305 565 1321 599
rect 1269 512 1321 565
rect 1269 478 1271 512
rect 1305 478 1321 512
rect 961 413 1133 418
rect 961 400 1099 413
rect 579 384 1099 400
rect 301 350 545 379
rect 1067 379 1099 384
rect 1269 413 1321 478
rect 1269 385 1271 413
rect 1133 379 1271 385
rect 1305 379 1321 413
rect 301 343 572 350
rect 195 275 221 309
rect 255 275 289 309
rect 323 275 357 309
rect 391 275 425 309
rect 459 275 475 309
rect 195 208 229 275
rect 509 241 572 343
rect 697 319 1033 350
rect 1067 337 1321 379
rect 65 192 229 208
rect 65 158 81 192
rect 115 174 229 192
rect 263 207 572 241
rect 606 287 663 303
rect 606 253 622 287
rect 656 253 663 287
rect 697 285 748 319
rect 782 285 816 319
rect 850 285 884 319
rect 918 285 952 319
rect 986 285 1033 319
rect 697 283 1033 285
rect 1067 287 1321 303
rect 606 249 663 253
rect 1067 253 1103 287
rect 1137 253 1171 287
rect 1205 253 1239 287
rect 1273 253 1321 287
rect 1067 249 1321 253
rect 606 242 1321 249
rect 606 215 1121 242
rect 115 158 121 174
rect 65 101 121 158
rect 263 140 297 207
rect 427 203 572 207
rect 65 67 81 101
rect 115 67 121 101
rect 65 51 121 67
rect 155 129 221 138
rect 155 95 171 129
rect 205 95 221 129
rect 155 17 221 95
rect 255 124 297 140
rect 255 90 257 124
rect 291 90 297 124
rect 255 74 297 90
rect 331 157 393 173
rect 331 123 343 157
rect 377 123 393 157
rect 331 89 393 123
rect 331 55 343 89
rect 377 55 393 89
rect 331 17 393 55
rect 427 169 429 203
rect 463 179 572 203
rect 1181 192 1227 208
rect 1181 181 1185 192
rect 463 175 977 179
rect 463 169 755 175
rect 427 141 755 169
rect 789 141 927 175
rect 961 141 977 175
rect 427 139 977 141
rect 1011 165 1185 181
rect 427 101 473 139
rect 1011 131 1013 165
rect 1047 158 1185 165
rect 1219 158 1227 192
rect 1047 147 1227 158
rect 1047 131 1063 147
rect 1011 105 1063 131
rect 427 67 429 101
rect 463 67 473 101
rect 427 51 473 67
rect 507 89 619 105
rect 507 55 515 89
rect 549 55 583 89
rect 617 55 619 89
rect 507 17 619 55
rect 653 101 1063 105
rect 653 67 669 101
rect 703 67 841 101
rect 875 97 1063 101
rect 875 67 1013 97
rect 653 63 1013 67
rect 1047 63 1063 97
rect 653 51 1063 63
rect 1097 97 1143 113
rect 1097 63 1099 97
rect 1133 63 1143 97
rect 1097 17 1143 63
rect 1177 101 1227 147
rect 1177 67 1185 101
rect 1219 67 1227 101
rect 1177 51 1227 67
rect 1261 192 1321 208
rect 1261 158 1271 192
rect 1305 158 1321 192
rect 1261 93 1321 158
rect 1261 59 1271 93
rect 1305 59 1321 93
rect 1261 17 1321 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21boi_4
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5477584
string GDS_START 5465528
<< end >>
