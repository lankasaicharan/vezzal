magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 157 189 159
rect 568 157 756 241
rect 1 49 756 157
rect 0 0 768 49
<< scnmos >>
rect 80 49 110 133
rect 270 47 300 131
rect 342 47 372 131
rect 414 47 444 131
rect 486 47 516 131
rect 647 47 677 215
<< scpmoshvt >>
rect 91 367 121 451
rect 185 367 215 451
rect 271 367 301 451
rect 459 367 489 451
rect 545 367 575 451
rect 650 367 680 619
<< ndiff >>
rect 27 108 80 133
rect 27 74 35 108
rect 69 74 80 108
rect 27 49 80 74
rect 110 97 163 133
rect 594 187 647 215
rect 594 153 602 187
rect 636 153 647 187
rect 594 131 647 153
rect 110 63 121 97
rect 155 63 163 97
rect 110 49 163 63
rect 217 95 270 131
rect 217 61 225 95
rect 259 61 270 95
rect 217 47 270 61
rect 300 47 342 131
rect 372 47 414 131
rect 444 47 486 131
rect 516 106 647 131
rect 516 72 527 106
rect 561 93 647 106
rect 561 72 602 93
rect 516 59 602 72
rect 636 59 647 93
rect 516 47 647 59
rect 677 172 730 215
rect 677 138 688 172
rect 722 138 730 172
rect 677 98 730 138
rect 677 64 688 98
rect 722 64 730 98
rect 677 47 730 64
<< pdiff >>
rect 597 607 650 619
rect 597 573 605 607
rect 639 573 650 607
rect 597 507 650 573
rect 597 473 605 507
rect 639 473 650 507
rect 597 451 650 473
rect 38 426 91 451
rect 38 392 46 426
rect 80 392 91 426
rect 38 367 91 392
rect 121 441 185 451
rect 121 407 136 441
rect 170 407 185 441
rect 121 367 185 407
rect 215 409 271 451
rect 215 375 226 409
rect 260 375 271 409
rect 215 367 271 375
rect 301 426 459 451
rect 301 392 333 426
rect 367 392 414 426
rect 448 392 459 426
rect 301 367 459 392
rect 489 409 545 451
rect 489 375 500 409
rect 534 375 545 409
rect 489 367 545 375
rect 575 413 650 451
rect 575 379 596 413
rect 630 379 650 413
rect 575 367 650 379
rect 680 599 733 619
rect 680 565 691 599
rect 725 565 733 599
rect 680 507 733 565
rect 680 473 691 507
rect 725 473 733 507
rect 680 413 733 473
rect 680 379 691 413
rect 725 379 733 413
rect 680 367 733 379
<< ndiffc >>
rect 35 74 69 108
rect 602 153 636 187
rect 121 63 155 97
rect 225 61 259 95
rect 527 72 561 106
rect 602 59 636 93
rect 688 138 722 172
rect 688 64 722 98
<< pdiffc >>
rect 605 573 639 607
rect 605 473 639 507
rect 46 392 80 426
rect 136 407 170 441
rect 226 375 260 409
rect 333 392 367 426
rect 414 392 448 426
rect 500 375 534 409
rect 596 379 630 413
rect 691 565 725 599
rect 691 473 725 507
rect 691 379 725 413
<< poly >>
rect 650 619 680 645
rect 495 575 575 591
rect 495 541 511 575
rect 545 541 575 575
rect 495 525 575 541
rect 91 451 121 477
rect 185 451 215 477
rect 271 451 301 477
rect 459 451 489 477
rect 545 451 575 525
rect 91 319 121 367
rect 44 303 121 319
rect 44 269 60 303
rect 94 289 121 303
rect 185 289 215 367
rect 271 308 301 367
rect 459 338 489 367
rect 414 319 489 338
rect 271 292 372 308
rect 94 269 110 289
rect 44 235 110 269
rect 44 201 60 235
rect 94 201 110 235
rect 44 185 110 201
rect 80 133 110 185
rect 163 273 229 289
rect 163 239 179 273
rect 213 239 229 273
rect 271 258 319 292
rect 353 258 372 292
rect 271 242 372 258
rect 163 205 229 239
rect 163 171 179 205
rect 213 185 229 205
rect 213 171 300 185
rect 163 155 300 171
rect 270 131 300 155
rect 342 131 372 242
rect 414 285 430 319
rect 464 308 489 319
rect 464 285 480 308
rect 414 269 480 285
rect 414 131 444 269
rect 545 260 575 367
rect 650 303 680 367
rect 528 230 575 260
rect 617 287 683 303
rect 617 253 633 287
rect 667 253 683 287
rect 617 237 683 253
rect 528 221 558 230
rect 486 191 558 221
rect 647 215 677 237
rect 486 131 516 191
rect 80 23 110 49
rect 270 21 300 47
rect 342 21 372 47
rect 414 21 444 47
rect 486 21 516 47
rect 647 21 677 47
<< polycont >>
rect 511 541 545 575
rect 60 269 94 303
rect 60 201 94 235
rect 179 239 213 273
rect 319 258 353 292
rect 179 171 213 205
rect 430 285 464 319
rect 633 253 667 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 30 426 86 442
rect 30 392 46 426
rect 80 392 86 426
rect 120 441 186 649
rect 120 407 136 441
rect 170 407 186 441
rect 317 426 464 649
rect 589 607 653 649
rect 498 575 555 591
rect 498 541 511 575
rect 545 541 555 575
rect 498 459 555 541
rect 589 573 605 607
rect 639 573 653 607
rect 589 507 653 573
rect 589 473 605 507
rect 639 473 653 507
rect 222 409 281 425
rect 30 373 86 392
rect 222 375 226 409
rect 260 375 281 409
rect 317 392 333 426
rect 367 392 414 426
rect 448 392 464 426
rect 589 425 653 473
rect 317 387 464 392
rect 498 409 546 425
rect 30 339 186 373
rect 222 359 281 375
rect 31 269 60 303
rect 94 269 110 303
rect 31 235 110 269
rect 31 201 60 235
rect 94 201 110 235
rect 152 289 186 339
rect 152 273 213 289
rect 152 239 179 273
rect 152 205 213 239
rect 152 171 179 205
rect 152 165 213 171
rect 19 131 213 165
rect 247 206 281 359
rect 498 375 500 409
rect 534 375 546 409
rect 315 292 372 353
rect 315 258 319 292
rect 353 258 372 292
rect 315 242 372 258
rect 406 319 464 353
rect 406 285 430 319
rect 406 240 464 285
rect 498 303 546 375
rect 580 413 653 425
rect 580 379 596 413
rect 630 379 653 413
rect 580 363 653 379
rect 687 599 751 615
rect 687 565 691 599
rect 725 565 751 599
rect 687 507 751 565
rect 687 473 691 507
rect 725 473 751 507
rect 687 413 751 473
rect 687 379 691 413
rect 725 379 751 413
rect 687 363 751 379
rect 498 287 667 303
rect 498 253 633 287
rect 498 237 667 253
rect 498 206 534 237
rect 247 172 534 206
rect 701 203 751 363
rect 586 187 638 203
rect 19 108 71 131
rect 19 74 35 108
rect 69 74 71 108
rect 247 97 303 172
rect 586 153 602 187
rect 636 153 638 187
rect 586 122 638 153
rect 19 58 71 74
rect 105 63 121 97
rect 155 63 171 97
rect 105 17 171 63
rect 209 95 303 97
rect 209 61 225 95
rect 259 61 303 95
rect 209 51 303 61
rect 511 106 638 122
rect 511 72 527 106
rect 561 93 638 106
rect 561 72 602 93
rect 511 59 602 72
rect 636 59 638 93
rect 511 17 638 59
rect 672 172 751 203
rect 672 138 688 172
rect 722 138 751 172
rect 672 98 751 138
rect 672 64 688 98
rect 722 64 751 98
rect 672 51 751 64
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4b_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5345766
string GDS_START 5337810
<< end >>
