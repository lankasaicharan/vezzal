magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 6002 1975
<< nwell >>
rect -38 331 4742 704
<< pwell >>
rect 1763 241 1866 271
rect 171 157 617 241
rect 1377 194 1972 241
rect 1114 157 1972 194
rect 2493 201 2980 241
rect 1 49 2228 157
rect 2493 49 4356 201
rect 0 0 4704 49
<< scnmos >>
rect 80 47 110 131
rect 152 47 182 131
rect 250 47 280 215
rect 336 47 366 215
rect 422 47 452 215
rect 508 47 538 215
rect 698 47 728 131
rect 1023 47 1053 131
rect 1095 47 1125 131
rect 1456 47 1486 215
rect 1592 47 1622 215
rect 1744 47 1774 215
rect 1866 47 1896 215
rect 2033 47 2063 131
rect 2119 47 2149 131
rect 2572 47 2602 215
rect 2677 47 2707 215
rect 2776 47 2806 215
rect 2862 47 2892 215
rect 3125 47 3155 175
rect 3211 47 3241 175
rect 3297 47 3327 175
rect 3383 47 3413 175
rect 3469 47 3499 175
rect 3555 47 3585 175
rect 3641 47 3671 175
rect 3727 47 3757 175
rect 3813 47 3843 175
rect 3899 47 3929 175
rect 3985 47 4015 175
rect 4071 47 4101 175
rect 4157 47 4187 175
rect 4243 47 4273 175
<< scpmoshvt >>
rect 80 419 130 619
rect 198 491 228 619
rect 270 491 300 619
rect 460 491 490 619
rect 675 367 705 619
rect 780 367 810 619
rect 866 367 896 619
rect 952 367 982 619
rect 1142 451 1172 619
rect 1214 451 1244 619
rect 1300 451 1330 619
rect 1545 367 1575 619
rect 1631 367 1661 619
rect 1717 367 1747 619
rect 1803 367 1833 619
rect 2003 373 2033 541
rect 2075 373 2105 541
rect 2315 367 2345 619
rect 2401 367 2431 619
rect 2591 367 2621 619
rect 2677 367 2707 619
rect 2867 367 2897 619
rect 2953 367 2983 619
rect 3039 367 3069 619
rect 3125 367 3155 619
rect 3211 367 3241 619
rect 3297 367 3327 619
rect 3383 367 3413 619
rect 3469 367 3499 619
rect 3555 367 3585 619
rect 3641 367 3671 619
rect 3727 367 3757 619
rect 3813 367 3843 619
rect 3899 367 3929 619
rect 3985 367 4015 619
rect 4071 367 4101 619
rect 4157 367 4187 619
rect 4243 367 4273 619
rect 4329 367 4359 619
rect 4415 367 4445 619
rect 4501 367 4531 619
<< ndiff >>
rect 197 188 250 215
rect 197 154 205 188
rect 239 154 250 188
rect 197 131 250 154
rect 27 101 80 131
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 47 152 131
rect 182 89 250 131
rect 182 55 205 89
rect 239 55 250 89
rect 182 47 250 55
rect 280 207 336 215
rect 280 173 291 207
rect 325 173 336 207
rect 280 101 336 173
rect 280 67 291 101
rect 325 67 336 101
rect 280 47 336 67
rect 366 122 422 215
rect 366 88 377 122
rect 411 88 422 122
rect 366 47 422 88
rect 452 184 508 215
rect 452 150 463 184
rect 497 150 508 184
rect 452 101 508 150
rect 452 67 463 101
rect 497 67 508 101
rect 452 47 508 67
rect 538 192 591 215
rect 538 158 549 192
rect 583 158 591 192
rect 538 94 591 158
rect 1140 155 1190 168
rect 1789 233 1840 245
rect 1789 215 1798 233
rect 1140 131 1148 155
rect 538 60 549 94
rect 583 60 591 94
rect 538 47 591 60
rect 645 105 698 131
rect 645 71 653 105
rect 687 71 698 105
rect 645 47 698 71
rect 728 89 1023 131
rect 728 55 751 89
rect 785 55 831 89
rect 865 55 902 89
rect 936 55 972 89
rect 1006 55 1023 89
rect 728 47 1023 55
rect 1053 47 1095 131
rect 1125 121 1148 131
rect 1182 121 1190 155
rect 1125 47 1190 121
rect 1403 120 1456 215
rect 1403 86 1411 120
rect 1445 86 1456 120
rect 1403 47 1456 86
rect 1486 181 1592 215
rect 1486 147 1547 181
rect 1581 147 1592 181
rect 1486 47 1592 147
rect 1622 93 1744 215
rect 1622 59 1699 93
rect 1733 59 1744 93
rect 1622 47 1744 59
rect 1774 199 1798 215
rect 1832 215 1840 233
rect 1832 199 1866 215
rect 1774 47 1866 199
rect 1896 131 1946 215
rect 1896 89 2033 131
rect 1896 55 1907 89
rect 1941 55 1988 89
rect 2022 55 2033 89
rect 1896 47 2033 55
rect 2063 111 2119 131
rect 2063 77 2074 111
rect 2108 77 2119 111
rect 2063 47 2119 77
rect 2149 93 2202 131
rect 2149 59 2160 93
rect 2194 59 2202 93
rect 2519 93 2572 215
rect 2149 47 2202 59
rect 2519 59 2527 93
rect 2561 59 2572 93
rect 2519 47 2572 59
rect 2602 135 2677 215
rect 2602 101 2624 135
rect 2658 101 2677 135
rect 2602 47 2677 101
rect 2707 203 2776 215
rect 2707 169 2731 203
rect 2765 169 2776 203
rect 2707 103 2776 169
rect 2707 69 2731 103
rect 2765 69 2776 103
rect 2707 47 2776 69
rect 2806 180 2862 215
rect 2806 146 2817 180
rect 2851 146 2862 180
rect 2806 47 2862 146
rect 2892 203 2954 215
rect 2892 169 2908 203
rect 2942 169 2954 203
rect 2892 103 2954 169
rect 2892 69 2908 103
rect 2942 69 2954 103
rect 2892 47 2954 69
rect 3068 157 3125 175
rect 3068 123 3080 157
rect 3114 123 3125 157
rect 3068 89 3125 123
rect 3068 55 3080 89
rect 3114 55 3125 89
rect 3068 47 3125 55
rect 3155 157 3211 175
rect 3155 123 3166 157
rect 3200 123 3211 157
rect 3155 89 3211 123
rect 3155 55 3166 89
rect 3200 55 3211 89
rect 3155 47 3211 55
rect 3241 157 3297 175
rect 3241 123 3252 157
rect 3286 123 3297 157
rect 3241 89 3297 123
rect 3241 55 3252 89
rect 3286 55 3297 89
rect 3241 47 3297 55
rect 3327 157 3383 175
rect 3327 123 3338 157
rect 3372 123 3383 157
rect 3327 89 3383 123
rect 3327 55 3338 89
rect 3372 55 3383 89
rect 3327 47 3383 55
rect 3413 157 3469 175
rect 3413 123 3424 157
rect 3458 123 3469 157
rect 3413 89 3469 123
rect 3413 55 3424 89
rect 3458 55 3469 89
rect 3413 47 3469 55
rect 3499 157 3555 175
rect 3499 123 3510 157
rect 3544 123 3555 157
rect 3499 89 3555 123
rect 3499 55 3510 89
rect 3544 55 3555 89
rect 3499 47 3555 55
rect 3585 157 3641 175
rect 3585 123 3596 157
rect 3630 123 3641 157
rect 3585 89 3641 123
rect 3585 55 3596 89
rect 3630 55 3641 89
rect 3585 47 3641 55
rect 3671 157 3727 175
rect 3671 123 3682 157
rect 3716 123 3727 157
rect 3671 89 3727 123
rect 3671 55 3682 89
rect 3716 55 3727 89
rect 3671 47 3727 55
rect 3757 157 3813 175
rect 3757 123 3768 157
rect 3802 123 3813 157
rect 3757 89 3813 123
rect 3757 55 3768 89
rect 3802 55 3813 89
rect 3757 47 3813 55
rect 3843 157 3899 175
rect 3843 123 3854 157
rect 3888 123 3899 157
rect 3843 89 3899 123
rect 3843 55 3854 89
rect 3888 55 3899 89
rect 3843 47 3899 55
rect 3929 157 3985 175
rect 3929 123 3940 157
rect 3974 123 3985 157
rect 3929 89 3985 123
rect 3929 55 3940 89
rect 3974 55 3985 89
rect 3929 47 3985 55
rect 4015 157 4071 175
rect 4015 123 4026 157
rect 4060 123 4071 157
rect 4015 89 4071 123
rect 4015 55 4026 89
rect 4060 55 4071 89
rect 4015 47 4071 55
rect 4101 157 4157 175
rect 4101 123 4112 157
rect 4146 123 4157 157
rect 4101 89 4157 123
rect 4101 55 4112 89
rect 4146 55 4157 89
rect 4101 47 4157 55
rect 4187 157 4243 175
rect 4187 123 4198 157
rect 4232 123 4243 157
rect 4187 89 4243 123
rect 4187 55 4198 89
rect 4232 55 4243 89
rect 4187 47 4243 55
rect 4273 157 4330 175
rect 4273 123 4284 157
rect 4318 123 4330 157
rect 4273 89 4330 123
rect 4273 55 4284 89
rect 4318 55 4330 89
rect 4273 47 4330 55
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 531 80 565
rect 27 497 35 531
rect 69 497 80 531
rect 27 419 80 497
rect 130 597 198 619
rect 130 563 141 597
rect 175 563 198 597
rect 130 503 198 563
rect 130 469 141 503
rect 175 491 198 503
rect 228 491 270 619
rect 300 607 353 619
rect 300 573 311 607
rect 345 573 353 607
rect 300 539 353 573
rect 300 505 311 539
rect 345 505 353 539
rect 300 491 353 505
rect 407 607 460 619
rect 407 573 415 607
rect 449 573 460 607
rect 407 539 460 573
rect 407 505 415 539
rect 449 505 460 539
rect 407 491 460 505
rect 490 601 675 619
rect 490 567 515 601
rect 549 567 630 601
rect 664 567 675 601
rect 490 533 675 567
rect 490 499 515 533
rect 549 499 630 533
rect 664 499 675 533
rect 490 491 675 499
rect 175 469 183 491
rect 130 419 183 469
rect 625 367 675 491
rect 705 597 780 619
rect 705 563 735 597
rect 769 563 780 597
rect 705 502 780 563
rect 705 468 735 502
rect 769 468 780 502
rect 705 409 780 468
rect 705 375 735 409
rect 769 375 780 409
rect 705 367 780 375
rect 810 593 866 619
rect 810 559 821 593
rect 855 559 866 593
rect 810 502 866 559
rect 810 468 821 502
rect 855 468 866 502
rect 810 420 866 468
rect 810 386 821 420
rect 855 386 866 420
rect 810 367 866 386
rect 896 598 952 619
rect 896 564 907 598
rect 941 564 952 598
rect 896 530 952 564
rect 896 496 907 530
rect 941 496 952 530
rect 896 462 952 496
rect 896 428 907 462
rect 941 428 952 462
rect 896 367 952 428
rect 982 576 1035 619
rect 982 542 993 576
rect 1027 542 1035 576
rect 982 367 1035 542
rect 1089 583 1142 619
rect 1089 549 1097 583
rect 1131 549 1142 583
rect 1089 451 1142 549
rect 1172 451 1214 619
rect 1244 597 1300 619
rect 1244 563 1255 597
rect 1289 563 1300 597
rect 1244 497 1300 563
rect 1244 463 1255 497
rect 1289 463 1300 497
rect 1244 451 1300 463
rect 1330 607 1383 619
rect 1330 573 1341 607
rect 1375 573 1383 607
rect 1330 537 1383 573
rect 1330 503 1341 537
rect 1375 503 1383 537
rect 1330 451 1383 503
rect 1492 597 1545 619
rect 1492 563 1500 597
rect 1534 563 1545 597
rect 1492 505 1545 563
rect 1492 471 1500 505
rect 1534 471 1545 505
rect 1492 413 1545 471
rect 1492 379 1500 413
rect 1534 379 1545 413
rect 1492 367 1545 379
rect 1575 527 1631 619
rect 1575 493 1586 527
rect 1620 493 1631 527
rect 1575 413 1631 493
rect 1575 379 1586 413
rect 1620 379 1631 413
rect 1575 367 1631 379
rect 1661 597 1717 619
rect 1661 563 1672 597
rect 1706 563 1717 597
rect 1661 505 1717 563
rect 1661 471 1672 505
rect 1706 471 1717 505
rect 1661 413 1717 471
rect 1661 379 1672 413
rect 1706 379 1717 413
rect 1661 367 1717 379
rect 1747 584 1803 619
rect 1747 550 1758 584
rect 1792 550 1803 584
rect 1747 367 1803 550
rect 1833 582 1886 619
rect 1833 548 1844 582
rect 1878 548 1886 582
rect 1833 514 1886 548
rect 1833 480 1844 514
rect 1878 480 1886 514
rect 1833 367 1886 480
rect 1946 529 2003 541
rect 1946 495 1958 529
rect 1992 495 2003 529
rect 1946 419 2003 495
rect 1946 385 1958 419
rect 1992 385 2003 419
rect 1946 373 2003 385
rect 2033 373 2075 541
rect 2105 529 2158 541
rect 2105 495 2116 529
rect 2150 495 2158 529
rect 2105 419 2158 495
rect 2105 385 2116 419
rect 2150 385 2158 419
rect 2105 373 2158 385
rect 2262 597 2315 619
rect 2262 563 2270 597
rect 2304 563 2315 597
rect 2262 514 2315 563
rect 2262 480 2270 514
rect 2304 480 2315 514
rect 2262 367 2315 480
rect 2345 597 2401 619
rect 2345 563 2356 597
rect 2390 563 2401 597
rect 2345 514 2401 563
rect 2345 480 2356 514
rect 2390 480 2401 514
rect 2345 367 2401 480
rect 2431 597 2484 619
rect 2431 563 2442 597
rect 2476 563 2484 597
rect 2431 367 2484 563
rect 2538 599 2591 619
rect 2538 565 2546 599
rect 2580 565 2591 599
rect 2538 487 2591 565
rect 2538 453 2546 487
rect 2580 453 2591 487
rect 2538 367 2591 453
rect 2621 505 2677 619
rect 2621 471 2632 505
rect 2666 471 2677 505
rect 2621 413 2677 471
rect 2621 379 2632 413
rect 2666 379 2677 413
rect 2621 367 2677 379
rect 2707 599 2760 619
rect 2707 565 2718 599
rect 2752 565 2760 599
rect 2707 487 2760 565
rect 2707 453 2718 487
rect 2752 453 2760 487
rect 2707 367 2760 453
rect 2814 607 2867 619
rect 2814 573 2822 607
rect 2856 573 2867 607
rect 2814 539 2867 573
rect 2814 505 2822 539
rect 2856 505 2867 539
rect 2814 471 2867 505
rect 2814 437 2822 471
rect 2856 437 2867 471
rect 2814 367 2867 437
rect 2897 597 2953 619
rect 2897 563 2908 597
rect 2942 563 2953 597
rect 2897 519 2953 563
rect 2897 485 2908 519
rect 2942 485 2953 519
rect 2897 442 2953 485
rect 2897 408 2908 442
rect 2942 408 2953 442
rect 2897 367 2953 408
rect 2983 607 3039 619
rect 2983 573 2994 607
rect 3028 573 3039 607
rect 2983 512 3039 573
rect 2983 478 2994 512
rect 3028 478 3039 512
rect 2983 367 3039 478
rect 3069 597 3125 619
rect 3069 563 3080 597
rect 3114 563 3125 597
rect 3069 517 3125 563
rect 3069 483 3080 517
rect 3114 483 3125 517
rect 3069 438 3125 483
rect 3069 404 3080 438
rect 3114 404 3125 438
rect 3069 367 3125 404
rect 3155 607 3211 619
rect 3155 573 3166 607
rect 3200 573 3211 607
rect 3155 508 3211 573
rect 3155 474 3166 508
rect 3200 474 3211 508
rect 3155 367 3211 474
rect 3241 597 3297 619
rect 3241 563 3252 597
rect 3286 563 3297 597
rect 3241 517 3297 563
rect 3241 483 3252 517
rect 3286 483 3297 517
rect 3241 438 3297 483
rect 3241 404 3252 438
rect 3286 404 3297 438
rect 3241 367 3297 404
rect 3327 607 3383 619
rect 3327 573 3338 607
rect 3372 573 3383 607
rect 3327 508 3383 573
rect 3327 474 3338 508
rect 3372 474 3383 508
rect 3327 367 3383 474
rect 3413 597 3469 619
rect 3413 563 3424 597
rect 3458 563 3469 597
rect 3413 517 3469 563
rect 3413 483 3424 517
rect 3458 483 3469 517
rect 3413 438 3469 483
rect 3413 404 3424 438
rect 3458 404 3469 438
rect 3413 367 3469 404
rect 3499 607 3555 619
rect 3499 573 3510 607
rect 3544 573 3555 607
rect 3499 508 3555 573
rect 3499 474 3510 508
rect 3544 474 3555 508
rect 3499 367 3555 474
rect 3585 597 3641 619
rect 3585 563 3596 597
rect 3630 563 3641 597
rect 3585 517 3641 563
rect 3585 483 3596 517
rect 3630 483 3641 517
rect 3585 438 3641 483
rect 3585 404 3596 438
rect 3630 404 3641 438
rect 3585 367 3641 404
rect 3671 607 3727 619
rect 3671 573 3682 607
rect 3716 573 3727 607
rect 3671 508 3727 573
rect 3671 474 3682 508
rect 3716 474 3727 508
rect 3671 367 3727 474
rect 3757 597 3813 619
rect 3757 563 3768 597
rect 3802 563 3813 597
rect 3757 517 3813 563
rect 3757 483 3768 517
rect 3802 483 3813 517
rect 3757 438 3813 483
rect 3757 404 3768 438
rect 3802 404 3813 438
rect 3757 367 3813 404
rect 3843 607 3899 619
rect 3843 573 3854 607
rect 3888 573 3899 607
rect 3843 508 3899 573
rect 3843 474 3854 508
rect 3888 474 3899 508
rect 3843 367 3899 474
rect 3929 597 3985 619
rect 3929 563 3940 597
rect 3974 563 3985 597
rect 3929 517 3985 563
rect 3929 483 3940 517
rect 3974 483 3985 517
rect 3929 438 3985 483
rect 3929 404 3940 438
rect 3974 404 3985 438
rect 3929 367 3985 404
rect 4015 607 4071 619
rect 4015 573 4026 607
rect 4060 573 4071 607
rect 4015 508 4071 573
rect 4015 474 4026 508
rect 4060 474 4071 508
rect 4015 367 4071 474
rect 4101 597 4157 619
rect 4101 563 4112 597
rect 4146 563 4157 597
rect 4101 517 4157 563
rect 4101 483 4112 517
rect 4146 483 4157 517
rect 4101 438 4157 483
rect 4101 404 4112 438
rect 4146 404 4157 438
rect 4101 367 4157 404
rect 4187 607 4243 619
rect 4187 573 4198 607
rect 4232 573 4243 607
rect 4187 508 4243 573
rect 4187 474 4198 508
rect 4232 474 4243 508
rect 4187 367 4243 474
rect 4273 597 4329 619
rect 4273 563 4284 597
rect 4318 563 4329 597
rect 4273 517 4329 563
rect 4273 483 4284 517
rect 4318 483 4329 517
rect 4273 438 4329 483
rect 4273 404 4284 438
rect 4318 404 4329 438
rect 4273 367 4329 404
rect 4359 607 4415 619
rect 4359 573 4370 607
rect 4404 573 4415 607
rect 4359 508 4415 573
rect 4359 474 4370 508
rect 4404 474 4415 508
rect 4359 367 4415 474
rect 4445 597 4501 619
rect 4445 563 4456 597
rect 4490 563 4501 597
rect 4445 517 4501 563
rect 4445 483 4456 517
rect 4490 483 4501 517
rect 4445 438 4501 483
rect 4445 404 4456 438
rect 4490 404 4501 438
rect 4445 367 4501 404
rect 4531 607 4588 619
rect 4531 573 4542 607
rect 4576 573 4588 607
rect 4531 508 4588 573
rect 4531 474 4542 508
rect 4576 474 4588 508
rect 4531 367 4588 474
<< ndiffc >>
rect 205 154 239 188
rect 35 67 69 101
rect 205 55 239 89
rect 291 173 325 207
rect 291 67 325 101
rect 377 88 411 122
rect 463 150 497 184
rect 463 67 497 101
rect 549 158 583 192
rect 549 60 583 94
rect 653 71 687 105
rect 751 55 785 89
rect 831 55 865 89
rect 902 55 936 89
rect 972 55 1006 89
rect 1148 121 1182 155
rect 1411 86 1445 120
rect 1547 147 1581 181
rect 1699 59 1733 93
rect 1798 199 1832 233
rect 1907 55 1941 89
rect 1988 55 2022 89
rect 2074 77 2108 111
rect 2160 59 2194 93
rect 2527 59 2561 93
rect 2624 101 2658 135
rect 2731 169 2765 203
rect 2731 69 2765 103
rect 2817 146 2851 180
rect 2908 169 2942 203
rect 2908 69 2942 103
rect 3080 123 3114 157
rect 3080 55 3114 89
rect 3166 123 3200 157
rect 3166 55 3200 89
rect 3252 123 3286 157
rect 3252 55 3286 89
rect 3338 123 3372 157
rect 3338 55 3372 89
rect 3424 123 3458 157
rect 3424 55 3458 89
rect 3510 123 3544 157
rect 3510 55 3544 89
rect 3596 123 3630 157
rect 3596 55 3630 89
rect 3682 123 3716 157
rect 3682 55 3716 89
rect 3768 123 3802 157
rect 3768 55 3802 89
rect 3854 123 3888 157
rect 3854 55 3888 89
rect 3940 123 3974 157
rect 3940 55 3974 89
rect 4026 123 4060 157
rect 4026 55 4060 89
rect 4112 123 4146 157
rect 4112 55 4146 89
rect 4198 123 4232 157
rect 4198 55 4232 89
rect 4284 123 4318 157
rect 4284 55 4318 89
<< pdiffc >>
rect 35 565 69 599
rect 35 497 69 531
rect 141 563 175 597
rect 141 469 175 503
rect 311 573 345 607
rect 311 505 345 539
rect 415 573 449 607
rect 415 505 449 539
rect 515 567 549 601
rect 630 567 664 601
rect 515 499 549 533
rect 630 499 664 533
rect 735 563 769 597
rect 735 468 769 502
rect 735 375 769 409
rect 821 559 855 593
rect 821 468 855 502
rect 821 386 855 420
rect 907 564 941 598
rect 907 496 941 530
rect 907 428 941 462
rect 993 542 1027 576
rect 1097 549 1131 583
rect 1255 563 1289 597
rect 1255 463 1289 497
rect 1341 573 1375 607
rect 1341 503 1375 537
rect 1500 563 1534 597
rect 1500 471 1534 505
rect 1500 379 1534 413
rect 1586 493 1620 527
rect 1586 379 1620 413
rect 1672 563 1706 597
rect 1672 471 1706 505
rect 1672 379 1706 413
rect 1758 550 1792 584
rect 1844 548 1878 582
rect 1844 480 1878 514
rect 1958 495 1992 529
rect 1958 385 1992 419
rect 2116 495 2150 529
rect 2116 385 2150 419
rect 2270 563 2304 597
rect 2270 480 2304 514
rect 2356 563 2390 597
rect 2356 480 2390 514
rect 2442 563 2476 597
rect 2546 565 2580 599
rect 2546 453 2580 487
rect 2632 471 2666 505
rect 2632 379 2666 413
rect 2718 565 2752 599
rect 2718 453 2752 487
rect 2822 573 2856 607
rect 2822 505 2856 539
rect 2822 437 2856 471
rect 2908 563 2942 597
rect 2908 485 2942 519
rect 2908 408 2942 442
rect 2994 573 3028 607
rect 2994 478 3028 512
rect 3080 563 3114 597
rect 3080 483 3114 517
rect 3080 404 3114 438
rect 3166 573 3200 607
rect 3166 474 3200 508
rect 3252 563 3286 597
rect 3252 483 3286 517
rect 3252 404 3286 438
rect 3338 573 3372 607
rect 3338 474 3372 508
rect 3424 563 3458 597
rect 3424 483 3458 517
rect 3424 404 3458 438
rect 3510 573 3544 607
rect 3510 474 3544 508
rect 3596 563 3630 597
rect 3596 483 3630 517
rect 3596 404 3630 438
rect 3682 573 3716 607
rect 3682 474 3716 508
rect 3768 563 3802 597
rect 3768 483 3802 517
rect 3768 404 3802 438
rect 3854 573 3888 607
rect 3854 474 3888 508
rect 3940 563 3974 597
rect 3940 483 3974 517
rect 3940 404 3974 438
rect 4026 573 4060 607
rect 4026 474 4060 508
rect 4112 563 4146 597
rect 4112 483 4146 517
rect 4112 404 4146 438
rect 4198 573 4232 607
rect 4198 474 4232 508
rect 4284 563 4318 597
rect 4284 483 4318 517
rect 4284 404 4318 438
rect 4370 573 4404 607
rect 4370 474 4404 508
rect 4456 563 4490 597
rect 4456 483 4490 517
rect 4456 404 4490 438
rect 4542 573 4576 607
rect 4542 474 4576 508
<< poly >>
rect 80 619 130 645
rect 198 619 228 645
rect 270 619 300 645
rect 460 619 490 645
rect 675 619 705 645
rect 780 619 810 645
rect 866 619 896 645
rect 952 619 982 645
rect 1142 619 1172 645
rect 1214 619 1244 645
rect 1300 619 1330 645
rect 1545 619 1575 645
rect 1631 619 1661 645
rect 1717 619 1747 645
rect 1803 619 1833 645
rect 80 316 130 419
rect 198 316 228 491
rect 270 387 300 491
rect 460 459 490 491
rect 460 429 610 459
rect 270 357 446 387
rect 80 315 228 316
rect 416 317 446 357
rect 580 343 610 429
rect 1142 419 1172 451
rect 1069 403 1172 419
rect 1069 369 1085 403
rect 1119 369 1172 403
rect 675 343 705 367
rect 780 343 810 367
rect 580 319 810 343
rect 80 300 366 315
rect 80 266 135 300
rect 169 266 366 300
rect 80 250 366 266
rect 80 131 110 250
rect 152 131 182 250
rect 250 215 280 250
rect 336 215 366 250
rect 416 301 538 317
rect 416 267 432 301
rect 466 267 538 301
rect 416 241 538 267
rect 580 285 596 319
rect 630 285 810 319
rect 580 250 810 285
rect 866 341 896 367
rect 952 341 982 367
rect 1069 353 1172 369
rect 866 331 982 341
rect 866 306 981 331
rect 1214 311 1244 451
rect 1300 382 1330 451
rect 1300 381 1352 382
rect 866 272 913 306
rect 947 272 981 306
rect 866 256 981 272
rect 1023 281 1244 311
rect 1286 365 1352 381
rect 1286 331 1302 365
rect 1336 331 1352 365
rect 1286 315 1352 331
rect 1394 365 1460 381
rect 1901 615 2243 645
rect 2315 619 2345 645
rect 2401 619 2431 645
rect 2591 619 2621 645
rect 2677 619 2707 645
rect 2867 619 2897 645
rect 2953 619 2983 645
rect 3039 619 3069 645
rect 3125 619 3155 645
rect 3211 619 3241 645
rect 3297 619 3327 645
rect 3383 619 3413 645
rect 3469 619 3499 645
rect 3555 619 3585 645
rect 3641 619 3671 645
rect 3727 619 3757 645
rect 3813 619 3843 645
rect 3899 619 3929 645
rect 3985 619 4015 645
rect 4071 619 4101 645
rect 4157 619 4187 645
rect 4243 619 4273 645
rect 4329 619 4359 645
rect 4415 619 4445 645
rect 4501 619 4531 645
rect 1394 331 1410 365
rect 1444 345 1460 365
rect 1545 345 1575 367
rect 1631 345 1661 367
rect 1444 331 1661 345
rect 1394 315 1661 331
rect 1717 343 1747 367
rect 1803 343 1833 367
rect 1901 343 1931 615
rect 2003 541 2033 567
rect 2075 541 2105 567
rect 422 215 452 241
rect 508 215 538 241
rect 698 214 810 250
rect 1023 214 1053 281
rect 1286 239 1316 315
rect 1717 313 1931 343
rect 1717 282 1896 313
rect 698 184 1053 214
rect 698 131 728 184
rect 1023 131 1053 184
rect 1095 209 1316 239
rect 1358 237 1622 267
rect 1095 131 1125 209
rect 1358 167 1388 237
rect 1456 215 1486 237
rect 1592 215 1622 237
rect 1744 215 1774 282
rect 1289 151 1388 167
rect 1289 117 1305 151
rect 1339 117 1388 151
rect 1289 101 1388 117
rect 1866 215 1896 282
rect 2003 266 2033 373
rect 2075 338 2105 373
rect 2213 345 2243 615
rect 2075 317 2171 338
rect 2075 308 2121 317
rect 2105 283 2121 308
rect 2155 283 2171 317
rect 2213 315 2247 345
rect 2315 334 2345 367
rect 2401 334 2431 367
rect 2591 345 2621 367
rect 2677 345 2707 367
rect 2003 265 2063 266
rect 1997 249 2063 265
rect 1997 215 2013 249
rect 2047 215 2063 249
rect 1997 199 2063 215
rect 2105 249 2171 283
rect 2105 215 2121 249
rect 2155 215 2171 249
rect 2105 199 2171 215
rect 2033 131 2063 199
rect 2119 131 2149 199
rect 2217 187 2247 315
rect 2289 306 2431 334
rect 2289 272 2305 306
rect 2339 272 2373 306
rect 2407 272 2431 306
rect 2289 256 2431 272
rect 2473 315 2707 345
rect 2867 345 2897 367
rect 2953 345 2983 367
rect 3039 345 3069 367
rect 3125 345 3155 367
rect 3211 345 3241 367
rect 3297 345 3327 367
rect 3383 345 3413 367
rect 3469 345 3499 367
rect 3555 345 3585 367
rect 3641 345 3671 367
rect 3727 345 3757 367
rect 3813 345 3843 367
rect 3899 345 3929 367
rect 3985 345 4015 367
rect 4071 345 4101 367
rect 4157 345 4187 367
rect 4243 345 4273 367
rect 4329 345 4359 367
rect 4415 345 4445 367
rect 4501 345 4531 367
rect 2473 187 2503 315
rect 2572 215 2602 315
rect 2677 215 2707 315
rect 2749 305 2815 321
rect 2867 319 4531 345
rect 2867 315 3852 319
rect 2749 271 2765 305
rect 2799 271 2815 305
rect 3836 285 3852 315
rect 3886 285 4024 319
rect 4058 285 4196 319
rect 4230 285 4368 319
rect 4402 285 4436 319
rect 4470 285 4531 319
rect 2749 267 2815 271
rect 2749 237 2892 267
rect 2776 215 2806 237
rect 2862 215 2892 237
rect 2969 257 3734 273
rect 3836 269 4531 285
rect 2969 223 2996 257
rect 3030 223 3168 257
rect 3202 223 3336 257
rect 3370 223 3512 257
rect 3546 223 3684 257
rect 3718 227 3734 257
rect 3718 223 4273 227
rect 2217 157 2503 187
rect 2280 138 2503 157
rect 2280 104 2296 138
rect 2330 104 2427 138
rect 2461 104 2503 138
rect 2280 88 2503 104
rect 2969 207 4273 223
rect 3125 175 3155 207
rect 3211 175 3241 207
rect 3297 175 3327 207
rect 3383 175 3413 207
rect 3469 197 4273 207
rect 3469 175 3499 197
rect 3555 175 3585 197
rect 3641 175 3671 197
rect 3727 175 3757 197
rect 3813 175 3843 197
rect 3899 175 3929 197
rect 3985 175 4015 197
rect 4071 175 4101 197
rect 4157 175 4187 197
rect 4243 175 4273 197
rect 80 21 110 47
rect 152 21 182 47
rect 250 21 280 47
rect 336 21 366 47
rect 422 21 452 47
rect 508 21 538 47
rect 698 21 728 47
rect 1023 21 1053 47
rect 1095 21 1125 47
rect 1456 21 1486 47
rect 1592 21 1622 47
rect 1744 21 1774 47
rect 1866 21 1896 47
rect 2033 21 2063 47
rect 2119 21 2149 47
rect 2572 21 2602 47
rect 2677 21 2707 47
rect 2776 21 2806 47
rect 2862 21 2892 47
rect 3125 21 3155 47
rect 3211 21 3241 47
rect 3297 21 3327 47
rect 3383 21 3413 47
rect 3469 21 3499 47
rect 3555 21 3585 47
rect 3641 21 3671 47
rect 3727 21 3757 47
rect 3813 21 3843 47
rect 3899 21 3929 47
rect 3985 21 4015 47
rect 4071 21 4101 47
rect 4157 21 4187 47
rect 4243 21 4273 47
<< polycont >>
rect 1085 369 1119 403
rect 135 266 169 300
rect 432 267 466 301
rect 596 285 630 319
rect 913 272 947 306
rect 1302 331 1336 365
rect 1410 331 1444 365
rect 1305 117 1339 151
rect 2121 283 2155 317
rect 2013 215 2047 249
rect 2121 215 2155 249
rect 2305 272 2339 306
rect 2373 272 2407 306
rect 2765 271 2799 305
rect 3852 285 3886 319
rect 4024 285 4058 319
rect 4196 285 4230 319
rect 4368 285 4402 319
rect 4436 285 4470 319
rect 2996 223 3030 257
rect 3168 223 3202 257
rect 3336 223 3370 257
rect 3512 223 3546 257
rect 3684 223 3718 257
rect 2296 104 2330 138
rect 2427 104 2461 138
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3775 683
rect 3809 649 3871 683
rect 3905 649 3967 683
rect 4001 649 4063 683
rect 4097 649 4159 683
rect 4193 649 4255 683
rect 4289 649 4351 683
rect 4385 649 4447 683
rect 4481 649 4543 683
rect 4577 649 4639 683
rect 4673 649 4704 683
rect 19 599 85 615
rect 19 565 35 599
rect 69 565 85 599
rect 19 531 85 565
rect 19 497 35 531
rect 69 497 85 531
rect 19 350 85 497
rect 125 597 191 649
rect 125 563 141 597
rect 175 563 191 597
rect 125 503 191 563
rect 125 469 141 503
rect 175 469 191 503
rect 125 464 191 469
rect 295 607 361 613
rect 295 573 311 607
rect 345 573 361 607
rect 295 539 361 573
rect 295 505 311 539
rect 345 505 361 539
rect 19 316 31 350
rect 65 316 85 350
rect 19 101 85 316
rect 119 424 185 430
rect 119 390 137 424
rect 171 390 185 424
rect 119 300 185 390
rect 295 386 361 505
rect 399 607 465 615
rect 399 573 415 607
rect 449 573 465 607
rect 399 539 465 573
rect 399 505 415 539
rect 449 505 465 539
rect 399 454 465 505
rect 499 601 680 615
rect 499 577 515 601
rect 549 577 630 601
rect 664 577 680 601
rect 499 543 500 577
rect 549 567 572 577
rect 534 543 572 567
rect 606 567 630 577
rect 606 543 644 567
rect 678 543 680 577
rect 499 533 680 543
rect 499 499 515 533
rect 549 499 630 533
rect 664 499 680 533
rect 499 488 680 499
rect 735 597 779 613
rect 769 563 779 597
rect 735 502 779 563
rect 769 468 779 502
rect 399 420 701 454
rect 119 266 135 300
rect 169 266 185 300
rect 119 240 185 266
rect 284 352 633 386
rect 284 207 325 352
rect 580 319 633 352
rect 407 301 483 318
rect 407 267 432 301
rect 466 267 483 301
rect 580 285 596 319
rect 630 285 633 319
rect 580 269 633 285
rect 407 240 483 267
rect 19 67 35 101
rect 69 67 85 101
rect 19 51 85 67
rect 189 188 250 204
rect 189 154 205 188
rect 239 154 250 188
rect 189 89 250 154
rect 189 55 205 89
rect 239 55 250 89
rect 189 17 250 55
rect 284 173 291 207
rect 325 184 510 206
rect 325 173 463 184
rect 284 172 463 173
rect 284 101 327 172
rect 461 150 463 172
rect 497 150 510 184
rect 284 67 291 101
rect 325 67 327 101
rect 284 51 327 67
rect 361 122 427 138
rect 361 88 377 122
rect 411 88 427 122
rect 361 17 427 88
rect 461 101 510 150
rect 461 67 463 101
rect 497 67 510 101
rect 461 51 510 67
rect 544 192 599 208
rect 544 158 549 192
rect 583 158 599 192
rect 544 94 599 158
rect 667 163 701 420
rect 735 409 779 468
rect 769 375 779 409
rect 735 231 779 375
rect 813 593 863 609
rect 813 543 821 593
rect 855 543 863 593
rect 813 502 863 543
rect 813 468 821 502
rect 855 468 863 502
rect 813 420 863 468
rect 813 386 821 420
rect 855 386 863 420
rect 897 598 943 614
rect 897 564 907 598
rect 941 564 943 598
rect 897 530 943 564
rect 977 577 1043 603
rect 977 543 991 577
rect 1025 576 1043 577
rect 977 542 993 543
rect 1027 542 1043 576
rect 977 533 1043 542
rect 1081 583 1147 649
rect 1081 549 1097 583
rect 1131 549 1147 583
rect 1081 533 1147 549
rect 1239 597 1305 613
rect 1239 563 1255 597
rect 1289 563 1305 597
rect 897 496 907 530
rect 941 499 943 530
rect 1239 499 1305 563
rect 941 497 1305 499
rect 941 496 1255 497
rect 897 465 1255 496
rect 897 462 943 465
rect 897 428 907 462
rect 941 428 943 462
rect 1239 463 1255 465
rect 1289 463 1305 497
rect 1341 607 1391 649
rect 1375 573 1391 607
rect 1341 537 1391 573
rect 1375 503 1391 537
rect 1341 487 1391 503
rect 1500 597 1722 613
rect 1534 579 1672 597
rect 1534 563 1550 579
rect 1500 505 1550 563
rect 1656 563 1672 579
rect 1706 563 1722 597
rect 1239 451 1305 463
rect 1534 471 1550 505
rect 897 412 943 428
rect 1054 424 1135 431
rect 813 370 863 386
rect 1054 390 1083 424
rect 1117 403 1135 424
rect 1239 417 1446 451
rect 1054 369 1085 390
rect 1119 369 1135 403
rect 897 350 963 363
rect 1054 353 1135 369
rect 1267 365 1352 381
rect 897 316 913 350
rect 947 316 963 350
rect 1267 350 1302 365
rect 1267 344 1279 350
rect 897 306 963 316
rect 897 272 913 306
rect 947 272 963 306
rect 897 265 963 272
rect 1169 316 1279 344
rect 1336 331 1352 365
rect 1313 316 1352 331
rect 1169 310 1352 316
rect 1394 365 1446 417
rect 1394 331 1410 365
rect 1444 331 1446 365
rect 1500 413 1550 471
rect 1534 379 1550 413
rect 1500 363 1550 379
rect 1584 527 1622 543
rect 1584 493 1586 527
rect 1620 493 1622 527
rect 1584 413 1622 493
rect 1584 379 1586 413
rect 1620 379 1622 413
rect 1169 231 1203 310
rect 1394 274 1446 331
rect 735 197 1203 231
rect 1237 240 1446 274
rect 1584 245 1622 379
rect 1656 505 1722 563
rect 1756 584 1808 649
rect 1756 550 1758 584
rect 1792 550 1808 584
rect 1756 534 1808 550
rect 1842 582 1894 613
rect 1842 548 1844 582
rect 1878 548 1894 582
rect 1656 471 1672 505
rect 1706 500 1722 505
rect 1842 514 1894 548
rect 1842 500 1844 514
rect 1706 480 1844 500
rect 1878 480 1894 514
rect 1706 471 1894 480
rect 1656 464 1894 471
rect 1942 529 2008 649
rect 2254 597 2306 649
rect 2254 563 2270 597
rect 2304 563 2306 597
rect 1942 495 1958 529
rect 1992 495 2008 529
rect 1656 413 1722 464
rect 1656 379 1672 413
rect 1706 379 1722 413
rect 1656 363 1722 379
rect 1942 419 2008 495
rect 1942 385 1958 419
rect 1992 385 2008 419
rect 1942 369 2008 385
rect 2100 529 2166 545
rect 2100 495 2116 529
rect 2150 495 2166 529
rect 2100 419 2166 495
rect 2254 514 2306 563
rect 2254 480 2270 514
rect 2304 480 2306 514
rect 2254 464 2306 480
rect 2340 597 2406 607
rect 2340 563 2356 597
rect 2390 563 2406 597
rect 2340 514 2406 563
rect 2440 597 2492 649
rect 2440 563 2442 597
rect 2476 563 2492 597
rect 2440 547 2492 563
rect 2530 599 2768 615
rect 2530 565 2546 599
rect 2580 565 2718 599
rect 2752 565 2768 599
rect 2530 555 2768 565
rect 2340 480 2356 514
rect 2390 498 2406 514
rect 2530 498 2596 555
rect 2390 487 2596 498
rect 2390 480 2546 487
rect 2340 464 2546 480
rect 2530 453 2546 464
rect 2580 453 2596 487
rect 2530 437 2596 453
rect 2630 505 2682 521
rect 2630 471 2632 505
rect 2666 471 2682 505
rect 2100 385 2116 419
rect 2150 403 2166 419
rect 2342 424 2411 430
rect 2150 385 2228 403
rect 2100 369 2228 385
rect 2097 317 2160 333
rect 1237 163 1271 240
rect 1547 233 1622 245
rect 1891 276 1949 301
rect 1891 242 1903 276
rect 1937 242 1949 276
rect 2097 283 2121 317
rect 2155 283 2160 317
rect 2097 276 2160 283
rect 1891 233 1949 242
rect 667 129 1091 163
rect 667 121 701 129
rect 544 60 549 94
rect 583 60 599 94
rect 544 17 599 60
rect 637 105 701 121
rect 637 71 653 105
rect 687 71 701 105
rect 637 55 701 71
rect 735 89 1022 95
rect 735 55 751 89
rect 785 55 831 89
rect 865 55 902 89
rect 936 55 972 89
rect 1006 55 1022 89
rect 735 17 1022 55
rect 1057 87 1091 129
rect 1132 155 1271 163
rect 1132 121 1148 155
rect 1182 121 1271 155
rect 1305 170 1513 204
rect 1305 151 1339 170
rect 1305 87 1339 117
rect 1057 53 1339 87
rect 1395 120 1445 136
rect 1395 86 1411 120
rect 1395 17 1445 86
rect 1479 87 1513 170
rect 1547 199 1798 233
rect 1832 199 1949 233
rect 1997 249 2063 265
rect 1997 215 2013 249
rect 2047 215 2063 249
rect 1997 199 2063 215
rect 2131 249 2160 276
rect 2097 215 2121 242
rect 2155 215 2160 249
rect 2097 199 2160 215
rect 2194 226 2228 369
rect 2342 390 2356 424
rect 2390 390 2411 424
rect 2342 323 2411 390
rect 2630 413 2682 471
rect 2718 487 2768 555
rect 2752 453 2768 487
rect 2718 437 2768 453
rect 2805 607 2872 649
rect 2805 573 2822 607
rect 2856 573 2872 607
rect 2805 539 2872 573
rect 2805 505 2822 539
rect 2856 505 2872 539
rect 2805 471 2872 505
rect 2805 437 2822 471
rect 2856 437 2872 471
rect 2805 427 2872 437
rect 2908 597 2942 613
rect 2908 519 2942 563
rect 2908 442 2942 485
rect 2978 607 3028 649
rect 2978 573 2994 607
rect 2978 512 3028 573
rect 2978 478 2994 512
rect 2978 462 3028 478
rect 3064 597 3130 613
rect 3064 563 3080 597
rect 3114 563 3130 597
rect 3064 517 3130 563
rect 3064 483 3080 517
rect 3114 483 3130 517
rect 2630 379 2632 413
rect 2666 391 2682 413
rect 3064 438 3130 483
rect 3166 607 3200 649
rect 3166 508 3200 573
rect 3166 458 3200 474
rect 3236 597 3302 613
rect 3236 563 3252 597
rect 3286 563 3302 597
rect 3236 517 3302 563
rect 3236 483 3252 517
rect 3286 483 3302 517
rect 3064 426 3080 438
rect 2666 379 2874 391
rect 2942 390 3080 426
rect 3114 390 3130 438
rect 2630 357 2874 379
rect 2840 356 2874 357
rect 2840 350 2972 356
rect 2289 306 2423 323
rect 2289 272 2305 306
rect 2339 272 2373 306
rect 2407 272 2423 306
rect 2289 265 2423 272
rect 2457 305 2806 321
rect 2457 271 2765 305
rect 2799 271 2806 305
rect 2457 255 2806 271
rect 2840 316 2919 350
rect 2953 316 2972 350
rect 2840 310 2972 316
rect 2457 226 2491 255
rect 1547 181 1581 199
rect 1997 165 2031 199
rect 1547 121 1581 147
rect 1615 131 2031 165
rect 2194 191 2491 226
rect 2840 219 2874 310
rect 2992 276 3030 282
rect 2992 223 2996 276
rect 2536 203 2781 219
rect 2194 163 2228 191
rect 1615 87 1649 131
rect 2072 129 2228 163
rect 2536 185 2731 203
rect 2280 138 2477 154
rect 2072 111 2110 129
rect 1479 53 1649 87
rect 1683 59 1699 93
rect 1733 59 1757 93
rect 1683 17 1757 59
rect 1891 89 2038 97
rect 1891 55 1907 89
rect 1941 55 1988 89
rect 2022 55 2038 89
rect 1891 17 2038 55
rect 2072 77 2074 111
rect 2108 77 2110 111
rect 2280 104 2296 138
rect 2330 104 2427 138
rect 2461 104 2477 138
rect 2072 53 2110 77
rect 2144 59 2160 93
rect 2194 59 2210 93
rect 2280 88 2477 104
rect 2536 93 2577 185
rect 2715 169 2731 185
rect 2765 169 2781 203
rect 2511 59 2527 93
rect 2561 59 2577 93
rect 2611 135 2673 151
rect 2611 101 2624 135
rect 2658 101 2673 135
rect 2144 17 2210 59
rect 2611 17 2673 101
rect 2715 103 2781 169
rect 2815 180 2874 219
rect 2815 146 2817 180
rect 2851 146 2874 180
rect 2815 123 2874 146
rect 2908 203 2958 219
rect 2992 207 3030 223
rect 2942 169 2958 203
rect 2715 69 2731 103
rect 2765 87 2781 103
rect 2908 103 2958 169
rect 2765 69 2908 87
rect 2942 69 2958 103
rect 2715 53 2958 69
rect 3064 157 3130 390
rect 3236 438 3302 483
rect 3338 607 3372 649
rect 3338 508 3372 573
rect 3338 458 3372 474
rect 3408 597 3474 613
rect 3408 563 3424 597
rect 3458 563 3474 597
rect 3408 517 3474 563
rect 3408 483 3424 517
rect 3458 483 3474 517
rect 3236 390 3252 438
rect 3286 390 3302 438
rect 3164 276 3202 282
rect 3164 223 3168 276
rect 3164 207 3202 223
rect 3064 123 3080 157
rect 3114 123 3130 157
rect 3064 89 3130 123
rect 3064 55 3080 89
rect 3114 55 3130 89
rect 3064 51 3130 55
rect 3166 157 3200 173
rect 3166 89 3200 123
rect 3166 17 3200 55
rect 3236 157 3302 390
rect 3408 438 3474 483
rect 3510 607 3544 649
rect 3510 508 3544 573
rect 3510 458 3544 474
rect 3580 597 3646 613
rect 3580 563 3596 597
rect 3630 563 3646 597
rect 3580 517 3646 563
rect 3580 483 3596 517
rect 3630 483 3646 517
rect 3408 390 3424 438
rect 3458 390 3474 438
rect 3336 276 3374 282
rect 3336 257 3340 276
rect 3370 223 3374 242
rect 3336 207 3374 223
rect 3236 123 3252 157
rect 3286 123 3302 157
rect 3236 89 3302 123
rect 3236 55 3252 89
rect 3286 55 3302 89
rect 3236 51 3302 55
rect 3338 157 3372 173
rect 3338 89 3372 123
rect 3338 17 3372 55
rect 3408 157 3474 390
rect 3580 438 3646 483
rect 3682 607 3716 649
rect 3682 508 3716 573
rect 3682 458 3716 474
rect 3752 597 3818 613
rect 3752 563 3768 597
rect 3802 563 3818 597
rect 3752 517 3818 563
rect 3752 483 3768 517
rect 3802 483 3818 517
rect 3580 390 3596 438
rect 3630 390 3646 438
rect 3508 276 3546 282
rect 3508 223 3512 276
rect 3508 207 3546 223
rect 3408 123 3424 157
rect 3458 123 3474 157
rect 3408 89 3474 123
rect 3408 55 3424 89
rect 3458 55 3474 89
rect 3408 51 3474 55
rect 3510 157 3544 173
rect 3510 89 3544 123
rect 3510 17 3544 55
rect 3580 157 3646 390
rect 3752 438 3818 483
rect 3854 607 3888 649
rect 3854 508 3888 573
rect 3854 458 3888 474
rect 3924 597 3990 613
rect 3924 563 3940 597
rect 3974 563 3990 597
rect 3924 517 3990 563
rect 3924 483 3940 517
rect 3974 483 3990 517
rect 3752 390 3768 438
rect 3802 390 3818 438
rect 3680 276 3718 282
rect 3680 223 3684 276
rect 3680 207 3718 223
rect 3580 123 3596 157
rect 3630 123 3646 157
rect 3580 89 3646 123
rect 3580 55 3596 89
rect 3630 55 3646 89
rect 3580 51 3646 55
rect 3682 157 3716 173
rect 3682 89 3716 123
rect 3682 17 3716 55
rect 3752 157 3818 390
rect 3924 438 3990 483
rect 4026 607 4060 649
rect 4026 508 4060 573
rect 4026 458 4060 474
rect 4096 597 4162 613
rect 4096 563 4112 597
rect 4146 563 4162 597
rect 4096 517 4162 563
rect 4096 483 4112 517
rect 4146 483 4162 517
rect 3924 390 3940 438
rect 3974 390 3990 438
rect 3852 350 3890 352
rect 3886 285 3890 350
rect 3852 269 3890 285
rect 3752 123 3768 157
rect 3802 123 3818 157
rect 3752 89 3818 123
rect 3752 55 3768 89
rect 3802 55 3818 89
rect 3752 51 3818 55
rect 3854 157 3888 173
rect 3854 89 3888 123
rect 3854 17 3888 55
rect 3924 157 3990 390
rect 4096 438 4162 483
rect 4198 607 4232 649
rect 4198 508 4232 573
rect 4198 458 4232 474
rect 4268 597 4334 613
rect 4268 563 4284 597
rect 4318 563 4334 597
rect 4268 517 4334 563
rect 4268 483 4284 517
rect 4318 483 4334 517
rect 4096 390 4112 438
rect 4146 390 4162 438
rect 4024 350 4062 352
rect 4058 285 4062 350
rect 4024 269 4062 285
rect 3924 123 3940 157
rect 3974 123 3990 157
rect 3924 89 3990 123
rect 3924 55 3940 89
rect 3974 55 3990 89
rect 3924 51 3990 55
rect 4026 157 4060 173
rect 4026 89 4060 123
rect 4026 17 4060 55
rect 4096 157 4162 390
rect 4268 438 4334 483
rect 4370 607 4404 649
rect 4370 508 4404 573
rect 4370 458 4404 474
rect 4440 597 4506 613
rect 4440 563 4456 597
rect 4490 563 4506 597
rect 4440 517 4506 563
rect 4440 483 4456 517
rect 4490 483 4506 517
rect 4268 390 4284 438
rect 4318 390 4334 438
rect 4196 350 4234 352
rect 4230 285 4234 350
rect 4196 269 4234 285
rect 4096 123 4112 157
rect 4146 123 4162 157
rect 4096 89 4162 123
rect 4096 55 4112 89
rect 4146 55 4162 89
rect 4096 52 4162 55
rect 4198 157 4232 173
rect 4198 89 4232 123
rect 4198 17 4232 55
rect 4268 157 4334 390
rect 4440 438 4506 483
rect 4542 607 4592 649
rect 4576 573 4592 607
rect 4542 508 4592 573
rect 4576 474 4592 508
rect 4542 458 4592 474
rect 4440 390 4456 438
rect 4490 390 4506 438
rect 4440 388 4506 390
rect 4368 350 4486 352
rect 4402 319 4440 350
rect 4402 285 4436 319
rect 4474 316 4486 350
rect 4470 285 4486 316
rect 4368 269 4486 285
rect 4268 123 4284 157
rect 4318 123 4334 157
rect 4268 89 4334 123
rect 4268 55 4284 89
rect 4318 55 4334 89
rect 4268 51 4334 55
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4704 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 3583 649 3617 683
rect 3679 649 3713 683
rect 3775 649 3809 683
rect 3871 649 3905 683
rect 3967 649 4001 683
rect 4063 649 4097 683
rect 4159 649 4193 683
rect 4255 649 4289 683
rect 4351 649 4385 683
rect 4447 649 4481 683
rect 4543 649 4577 683
rect 4639 649 4673 683
rect 31 316 65 350
rect 137 390 171 424
rect 500 567 515 577
rect 515 567 534 577
rect 500 543 534 567
rect 572 543 606 577
rect 644 567 664 577
rect 664 567 678 577
rect 644 543 678 567
rect 821 559 855 577
rect 821 543 855 559
rect 991 576 1025 577
rect 991 543 993 576
rect 993 543 1025 576
rect 1083 403 1117 424
rect 1083 390 1085 403
rect 1085 390 1117 403
rect 913 316 947 350
rect 1279 331 1302 350
rect 1302 331 1313 350
rect 1279 316 1313 331
rect 1903 242 1937 276
rect 2097 249 2131 276
rect 2097 242 2121 249
rect 2121 242 2131 249
rect 2356 390 2390 424
rect 2908 408 2942 424
rect 2908 390 2942 408
rect 3080 404 3114 424
rect 3080 390 3114 404
rect 2919 316 2953 350
rect 2996 257 3030 276
rect 2996 242 3030 257
rect 3252 404 3286 424
rect 3252 390 3286 404
rect 3168 257 3202 276
rect 3168 242 3202 257
rect 3424 404 3458 424
rect 3424 390 3458 404
rect 3340 257 3374 276
rect 3340 242 3370 257
rect 3370 242 3374 257
rect 3596 404 3630 424
rect 3596 390 3630 404
rect 3512 257 3546 276
rect 3512 242 3546 257
rect 3768 404 3802 424
rect 3768 390 3802 404
rect 3684 257 3718 276
rect 3684 242 3718 257
rect 3940 404 3974 424
rect 3940 390 3974 404
rect 3852 319 3886 350
rect 3852 316 3886 319
rect 4112 404 4146 424
rect 4112 390 4146 404
rect 4024 319 4058 350
rect 4024 316 4058 319
rect 4284 404 4318 424
rect 4284 390 4318 404
rect 4196 319 4230 350
rect 4196 316 4230 319
rect 4456 404 4490 424
rect 4456 390 4490 404
rect 4368 319 4402 350
rect 4440 319 4474 350
rect 4368 316 4402 319
rect 4440 316 4470 319
rect 4470 316 4474 319
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
rect 4063 -17 4097 17
rect 4159 -17 4193 17
rect 4255 -17 4289 17
rect 4351 -17 4385 17
rect 4447 -17 4481 17
rect 4543 -17 4577 17
rect 4639 -17 4673 17
<< metal1 >>
rect 0 683 4704 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3775 683
rect 3809 649 3871 683
rect 3905 649 3967 683
rect 4001 649 4063 683
rect 4097 649 4159 683
rect 4193 649 4255 683
rect 4289 649 4351 683
rect 4385 649 4447 683
rect 4481 649 4543 683
rect 4577 649 4639 683
rect 4673 649 4704 683
rect 0 617 4704 649
rect 14 577 4690 589
rect 14 543 500 577
rect 534 543 572 577
rect 606 543 644 577
rect 678 543 821 577
rect 855 543 991 577
rect 1025 543 4690 577
rect 14 535 4690 543
rect 125 424 183 430
rect 1071 424 1129 430
rect 2344 424 2402 430
rect 125 390 137 424
rect 171 390 1083 424
rect 1117 390 2356 424
rect 2390 390 2402 424
rect 125 384 183 390
rect 1071 384 1129 390
rect 2344 384 2402 390
rect 2896 424 4502 430
rect 2896 390 2908 424
rect 2942 390 3080 424
rect 3114 390 3252 424
rect 3286 390 3424 424
rect 3458 390 3596 424
rect 3630 390 3768 424
rect 3802 390 3940 424
rect 3974 390 4112 424
rect 4146 390 4284 424
rect 4318 390 4456 424
rect 4490 390 4502 424
rect 2896 384 4502 390
rect 19 350 77 356
rect 19 316 31 350
rect 65 347 77 350
rect 901 350 959 356
rect 901 347 913 350
rect 65 319 913 347
rect 65 316 77 319
rect 19 310 77 316
rect 901 316 913 319
rect 947 316 959 350
rect 901 310 959 316
rect 1267 350 1325 356
rect 1267 316 1279 350
rect 1313 347 1325 350
rect 2900 350 4493 356
rect 2900 347 2919 350
rect 1313 319 2919 347
rect 1313 316 1325 319
rect 1267 310 1325 316
rect 2901 316 2919 319
rect 2953 316 3852 350
rect 3886 316 4024 350
rect 4058 316 4196 350
rect 4230 316 4368 350
rect 4402 316 4440 350
rect 4474 316 4493 350
rect 2901 310 4493 316
rect 1891 276 1949 282
rect 1891 242 1903 276
rect 1937 273 1949 276
rect 2085 276 2143 282
rect 2085 273 2097 276
rect 1937 245 2097 273
rect 1937 242 1949 245
rect 1891 236 1949 242
rect 2085 242 2097 245
rect 2131 273 2143 276
rect 2984 276 3739 282
rect 2984 273 2996 276
rect 2131 245 2996 273
rect 2131 242 2143 245
rect 2085 236 2143 242
rect 2984 242 2996 245
rect 3030 242 3168 276
rect 3202 242 3340 276
rect 3374 242 3512 276
rect 3546 242 3684 276
rect 3718 242 3739 276
rect 2984 236 3739 242
rect 0 17 4704 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4704 17
rect 0 -49 4704 -17
<< labels >>
flabel pwell s 0 0 4704 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 4704 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sky130_fd_sc_lp__busdrivernovlp_20_sleep
flabel metal1 s 2896 384 4502 430 0 FreeSans 200 0 0 0 Z
port 9 nsew signal output
flabel metal1 s 0 617 4704 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 4704 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 14 535 4690 589 0 FreeSans 200 0 0 0 KAPWR
port 4 nsew power bidirectional
flabel metal1 s 127 390 161 424 0 FreeSans 200 0 0 0 SLEEP
port 2 nsew signal input
flabel locali s 430 242 464 276 0 FreeSans 200 0 0 0 TE_B
port 3 nsew signal input
flabel locali s 2431 94 2465 128 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 2335 94 2369 128 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 4704 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y
string GDS_END 6005516
string GDS_START 5972320
<< end >>
