magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 23 49 915 243
rect 0 0 960 49
<< scnmos >>
rect 102 133 132 217
rect 253 49 283 217
rect 339 49 369 217
rect 425 49 455 217
rect 511 49 541 217
rect 613 49 643 217
rect 699 49 729 217
rect 806 49 836 217
<< scpmoshvt >>
rect 102 367 132 451
rect 260 367 290 619
rect 346 367 376 619
rect 432 367 462 619
rect 518 367 548 619
rect 626 367 656 619
rect 698 367 728 619
rect 806 367 836 619
<< ndiff >>
rect 49 192 102 217
rect 49 158 57 192
rect 91 158 102 192
rect 49 133 102 158
rect 132 165 253 217
rect 132 133 208 165
rect 200 131 208 133
rect 242 131 253 165
rect 200 95 253 131
rect 200 61 208 95
rect 242 61 253 95
rect 200 49 253 61
rect 283 205 339 217
rect 283 171 294 205
rect 328 171 339 205
rect 283 101 339 171
rect 283 67 294 101
rect 328 67 339 101
rect 283 49 339 67
rect 369 181 425 217
rect 369 147 380 181
rect 414 147 425 181
rect 369 95 425 147
rect 369 61 380 95
rect 414 61 425 95
rect 369 49 425 61
rect 455 205 511 217
rect 455 171 466 205
rect 500 171 511 205
rect 455 101 511 171
rect 455 67 466 101
rect 500 67 511 101
rect 455 49 511 67
rect 541 167 613 217
rect 541 133 560 167
rect 594 133 613 167
rect 541 91 613 133
rect 541 57 560 91
rect 594 57 613 91
rect 541 49 613 57
rect 643 205 699 217
rect 643 171 654 205
rect 688 171 699 205
rect 643 101 699 171
rect 643 67 654 101
rect 688 67 699 101
rect 643 49 699 67
rect 729 167 806 217
rect 729 133 751 167
rect 785 133 806 167
rect 729 91 806 133
rect 729 57 751 91
rect 785 57 806 91
rect 729 49 806 57
rect 836 205 889 217
rect 836 171 847 205
rect 881 171 889 205
rect 836 101 889 171
rect 836 67 847 101
rect 881 67 889 101
rect 836 49 889 67
<< pdiff >>
rect 207 573 260 619
rect 207 539 215 573
rect 249 539 260 573
rect 207 451 260 539
rect 49 426 102 451
rect 49 392 57 426
rect 91 392 102 426
rect 49 367 102 392
rect 132 367 260 451
rect 290 413 346 619
rect 290 379 301 413
rect 335 379 346 413
rect 290 367 346 379
rect 376 573 432 619
rect 376 539 387 573
rect 421 539 432 573
rect 376 367 432 539
rect 462 413 518 619
rect 462 379 473 413
rect 507 379 518 413
rect 462 367 518 379
rect 548 573 626 619
rect 548 539 570 573
rect 604 539 626 573
rect 548 367 626 539
rect 656 367 698 619
rect 728 367 806 619
rect 836 599 896 619
rect 836 565 847 599
rect 881 565 896 599
rect 836 503 896 565
rect 836 469 852 503
rect 886 469 896 503
rect 836 413 896 469
rect 836 379 852 413
rect 886 379 896 413
rect 836 367 896 379
<< ndiffc >>
rect 57 158 91 192
rect 208 131 242 165
rect 208 61 242 95
rect 294 171 328 205
rect 294 67 328 101
rect 380 147 414 181
rect 380 61 414 95
rect 466 171 500 205
rect 466 67 500 101
rect 560 133 594 167
rect 560 57 594 91
rect 654 171 688 205
rect 654 67 688 101
rect 751 133 785 167
rect 751 57 785 91
rect 847 171 881 205
rect 847 67 881 101
<< pdiffc >>
rect 215 539 249 573
rect 57 392 91 426
rect 301 379 335 413
rect 387 539 421 573
rect 473 379 507 413
rect 570 539 604 573
rect 847 565 881 599
rect 852 469 886 503
rect 852 379 886 413
<< poly >>
rect 260 619 290 645
rect 346 619 376 645
rect 432 619 462 645
rect 518 619 548 645
rect 626 619 656 645
rect 698 619 728 645
rect 806 619 836 645
rect 102 451 132 477
rect 102 305 132 367
rect 260 335 290 367
rect 346 335 376 367
rect 432 335 462 367
rect 518 335 548 367
rect 626 335 656 367
rect 260 319 548 335
rect 102 289 177 305
rect 260 299 287 319
rect 102 255 127 289
rect 161 255 177 289
rect 102 239 177 255
rect 253 285 287 299
rect 321 285 355 319
rect 389 285 423 319
rect 457 285 491 319
rect 525 285 548 319
rect 253 269 548 285
rect 590 319 656 335
rect 590 285 606 319
rect 640 285 656 319
rect 590 269 656 285
rect 698 335 728 367
rect 806 335 836 367
rect 698 319 764 335
rect 698 285 714 319
rect 748 285 764 319
rect 698 269 764 285
rect 806 319 872 335
rect 806 285 822 319
rect 856 285 872 319
rect 806 269 872 285
rect 102 217 132 239
rect 253 217 283 269
rect 339 217 369 269
rect 425 217 455 269
rect 511 217 541 269
rect 613 217 643 269
rect 699 217 729 269
rect 806 217 836 269
rect 102 107 132 133
rect 253 23 283 49
rect 339 23 369 49
rect 425 23 455 49
rect 511 23 541 49
rect 613 23 643 49
rect 699 23 729 49
rect 806 23 836 49
<< polycont >>
rect 127 255 161 289
rect 287 285 321 319
rect 355 285 389 319
rect 423 285 457 319
rect 491 285 525 319
rect 606 285 640 319
rect 714 285 748 319
rect 822 285 856 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 199 573 265 649
rect 199 539 215 573
rect 249 539 265 573
rect 199 531 265 539
rect 371 573 437 649
rect 371 539 387 573
rect 421 539 437 573
rect 371 531 437 539
rect 554 573 620 649
rect 554 539 570 573
rect 604 539 620 573
rect 831 599 942 615
rect 831 565 847 599
rect 881 565 942 599
rect 831 552 942 565
rect 554 531 620 539
rect 852 503 942 552
rect 41 463 818 497
rect 41 426 91 463
rect 41 392 57 426
rect 41 192 91 392
rect 41 158 57 192
rect 41 142 91 158
rect 125 289 167 424
rect 125 255 127 289
rect 161 255 167 289
rect 125 94 167 255
rect 201 413 545 429
rect 201 379 301 413
rect 335 379 473 413
rect 507 379 545 413
rect 201 363 545 379
rect 201 249 237 363
rect 271 319 570 329
rect 271 285 287 319
rect 321 285 355 319
rect 389 285 423 319
rect 457 285 491 319
rect 525 285 570 319
rect 271 283 570 285
rect 201 215 502 249
rect 286 205 330 215
rect 201 165 252 181
rect 201 131 208 165
rect 242 131 252 165
rect 201 95 252 131
rect 201 61 208 95
rect 242 61 252 95
rect 201 17 252 61
rect 286 171 294 205
rect 328 171 330 205
rect 464 205 502 215
rect 286 101 330 171
rect 286 67 294 101
rect 328 67 330 101
rect 286 51 330 67
rect 364 147 380 181
rect 414 147 430 181
rect 364 95 430 147
rect 364 61 380 95
rect 414 61 430 95
rect 364 17 430 61
rect 464 171 466 205
rect 500 171 502 205
rect 536 235 570 283
rect 604 319 655 429
rect 604 285 606 319
rect 640 285 655 319
rect 604 269 655 285
rect 689 319 748 429
rect 689 285 714 319
rect 689 269 748 285
rect 784 329 818 463
rect 886 469 942 503
rect 852 413 942 469
rect 886 379 942 413
rect 852 363 942 379
rect 784 319 872 329
rect 784 285 822 319
rect 856 285 872 319
rect 784 269 872 285
rect 906 235 942 363
rect 536 205 942 235
rect 536 201 654 205
rect 464 101 502 171
rect 644 171 654 201
rect 688 201 847 205
rect 688 171 701 201
rect 464 67 466 101
rect 500 67 502 101
rect 464 51 502 67
rect 544 133 560 167
rect 594 133 610 167
rect 544 91 610 133
rect 544 57 560 91
rect 594 57 610 91
rect 544 17 610 57
rect 644 101 701 171
rect 835 171 847 201
rect 881 171 942 205
rect 644 67 654 101
rect 688 67 701 101
rect 644 51 701 67
rect 735 133 751 167
rect 785 133 801 167
rect 735 91 801 133
rect 735 57 751 91
rect 785 57 801 91
rect 735 17 801 57
rect 835 101 942 171
rect 835 67 847 101
rect 881 67 942 101
rect 835 51 942 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or3b_4
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1632100
string GDS_START 1623912
<< end >>
