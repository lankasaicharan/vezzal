magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 1 49 582 241
rect 0 0 672 49
<< scnmos >>
rect 80 131 110 215
rect 199 47 229 215
rect 294 47 324 215
rect 387 47 417 215
rect 473 47 503 215
<< scpmoshvt >>
rect 110 367 140 451
rect 215 367 245 619
rect 301 367 331 619
rect 387 367 417 619
rect 473 367 503 619
<< ndiff >>
rect 27 187 80 215
rect 27 153 35 187
rect 69 153 80 187
rect 27 131 80 153
rect 110 187 199 215
rect 110 153 121 187
rect 155 153 199 187
rect 110 131 199 153
rect 132 93 199 131
rect 132 59 154 93
rect 188 59 199 93
rect 132 47 199 59
rect 229 181 294 215
rect 229 147 240 181
rect 274 147 294 181
rect 229 93 294 147
rect 229 59 240 93
rect 274 59 294 93
rect 229 47 294 59
rect 324 175 387 215
rect 324 141 342 175
rect 376 141 387 175
rect 324 47 387 141
rect 417 93 473 215
rect 417 59 428 93
rect 462 59 473 93
rect 417 47 473 59
rect 503 95 556 215
rect 503 61 514 95
rect 548 61 556 95
rect 503 47 556 61
<< pdiff >>
rect 162 607 215 619
rect 162 573 170 607
rect 204 573 215 607
rect 162 526 215 573
rect 162 492 170 526
rect 204 492 215 526
rect 162 451 215 492
rect 53 426 110 451
rect 53 392 65 426
rect 99 392 110 426
rect 53 367 110 392
rect 140 441 215 451
rect 140 407 151 441
rect 185 407 215 441
rect 140 367 215 407
rect 245 599 301 619
rect 245 565 256 599
rect 290 565 301 599
rect 245 525 301 565
rect 245 491 256 525
rect 290 491 301 525
rect 245 457 301 491
rect 245 423 256 457
rect 290 423 301 457
rect 245 367 301 423
rect 331 607 387 619
rect 331 573 342 607
rect 376 573 387 607
rect 331 514 387 573
rect 331 480 342 514
rect 376 480 387 514
rect 331 367 387 480
rect 417 599 473 619
rect 417 565 428 599
rect 462 565 473 599
rect 417 506 473 565
rect 417 472 428 506
rect 462 472 473 506
rect 417 416 473 472
rect 417 382 428 416
rect 462 382 473 416
rect 417 367 473 382
rect 503 607 556 619
rect 503 573 514 607
rect 548 573 556 607
rect 503 499 556 573
rect 503 465 514 499
rect 548 465 556 499
rect 503 367 556 465
<< ndiffc >>
rect 35 153 69 187
rect 121 153 155 187
rect 154 59 188 93
rect 240 147 274 181
rect 240 59 274 93
rect 342 141 376 175
rect 428 59 462 93
rect 514 61 548 95
<< pdiffc >>
rect 170 573 204 607
rect 170 492 204 526
rect 65 392 99 426
rect 151 407 185 441
rect 256 565 290 599
rect 256 491 290 525
rect 256 423 290 457
rect 342 573 376 607
rect 342 480 376 514
rect 428 565 462 599
rect 428 472 462 506
rect 428 382 462 416
rect 514 573 548 607
rect 514 465 548 499
<< poly >>
rect 215 619 245 645
rect 301 619 331 645
rect 387 619 417 645
rect 473 619 503 645
rect 110 451 140 477
rect 110 303 140 367
rect 215 303 245 367
rect 301 335 331 367
rect 387 335 417 367
rect 294 319 428 335
rect 72 287 140 303
rect 72 253 88 287
rect 122 273 140 287
rect 186 287 252 303
rect 122 253 138 273
rect 72 237 138 253
rect 186 253 202 287
rect 236 253 252 287
rect 186 237 252 253
rect 294 285 310 319
rect 344 285 428 319
rect 294 269 428 285
rect 473 303 503 367
rect 473 287 539 303
rect 80 215 110 237
rect 199 215 229 237
rect 294 215 324 269
rect 387 215 417 269
rect 473 253 489 287
rect 523 253 539 287
rect 473 237 539 253
rect 473 215 503 237
rect 80 105 110 131
rect 199 21 229 47
rect 294 21 324 47
rect 387 21 417 47
rect 473 21 503 47
<< polycont >>
rect 88 253 122 287
rect 202 253 236 287
rect 310 285 344 319
rect 489 253 523 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 135 607 212 649
rect 135 573 170 607
rect 204 573 212 607
rect 135 526 212 573
rect 135 492 170 526
rect 204 492 212 526
rect 18 426 101 442
rect 18 392 65 426
rect 99 392 101 426
rect 135 441 212 492
rect 135 407 151 441
rect 185 407 212 441
rect 246 599 292 615
rect 246 565 256 599
rect 290 565 292 599
rect 246 525 292 565
rect 246 491 256 525
rect 290 491 292 525
rect 246 457 292 491
rect 326 607 392 649
rect 326 573 342 607
rect 376 573 392 607
rect 326 514 392 573
rect 326 480 342 514
rect 376 480 392 514
rect 326 475 392 480
rect 426 599 464 615
rect 426 565 428 599
rect 462 565 464 599
rect 426 506 464 565
rect 246 423 256 457
rect 290 441 292 457
rect 426 472 428 506
rect 462 472 464 506
rect 426 441 464 472
rect 498 607 564 649
rect 498 573 514 607
rect 548 573 564 607
rect 498 499 564 573
rect 498 465 514 499
rect 548 465 564 499
rect 498 458 564 465
rect 290 424 464 441
rect 290 423 655 424
rect 246 416 655 423
rect 246 407 428 416
rect 18 373 101 392
rect 394 382 428 407
rect 462 382 655 416
rect 18 339 360 373
rect 394 366 655 382
rect 18 203 52 339
rect 294 319 360 339
rect 88 287 168 303
rect 122 253 168 287
rect 88 237 168 253
rect 202 287 260 303
rect 236 253 260 287
rect 294 285 310 319
rect 344 285 360 319
rect 294 283 360 285
rect 473 287 539 303
rect 202 249 260 253
rect 473 253 489 287
rect 523 253 539 287
rect 473 249 539 253
rect 202 215 539 249
rect 18 187 71 203
rect 18 153 35 187
rect 69 153 71 187
rect 18 137 71 153
rect 105 187 171 199
rect 105 153 121 187
rect 155 181 171 187
rect 575 181 655 366
rect 155 153 190 181
rect 105 93 190 153
rect 105 59 154 93
rect 188 59 190 93
rect 105 17 190 59
rect 224 147 240 181
rect 274 147 290 181
rect 224 97 290 147
rect 326 175 655 181
rect 326 141 342 175
rect 376 145 655 175
rect 376 141 392 145
rect 326 131 392 141
rect 224 93 478 97
rect 224 59 240 93
rect 274 59 428 93
rect 462 59 478 93
rect 224 51 478 59
rect 512 95 564 111
rect 512 61 514 95
rect 548 61 564 95
rect 512 17 564 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2b_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4430716
string GDS_START 4424710
<< end >>
