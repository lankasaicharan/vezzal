magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 1 49 577 157
rect 0 0 672 49
<< scnmos >>
rect 80 47 110 131
rect 152 47 182 131
rect 238 47 268 131
rect 310 47 340 131
rect 396 47 426 131
rect 468 47 498 131
<< scpmoshvt >>
rect 119 417 169 617
rect 225 417 275 617
rect 331 417 381 617
<< ndiff >>
rect 27 105 80 131
rect 27 71 35 105
rect 69 71 80 105
rect 27 47 80 71
rect 110 47 152 131
rect 182 105 238 131
rect 182 71 193 105
rect 227 71 238 105
rect 182 47 238 71
rect 268 47 310 131
rect 340 105 396 131
rect 340 71 351 105
rect 385 71 396 105
rect 340 47 396 71
rect 426 47 468 131
rect 498 105 551 131
rect 498 71 509 105
rect 543 71 551 105
rect 498 47 551 71
<< pdiff >>
rect 66 599 119 617
rect 66 565 74 599
rect 108 565 119 599
rect 66 531 119 565
rect 66 497 74 531
rect 108 497 119 531
rect 66 463 119 497
rect 66 429 74 463
rect 108 429 119 463
rect 66 417 119 429
rect 169 599 225 617
rect 169 565 180 599
rect 214 565 225 599
rect 169 531 225 565
rect 169 497 180 531
rect 214 497 225 531
rect 169 463 225 497
rect 169 429 180 463
rect 214 429 225 463
rect 169 417 225 429
rect 275 599 331 617
rect 275 565 286 599
rect 320 565 331 599
rect 275 531 331 565
rect 275 497 286 531
rect 320 497 331 531
rect 275 463 331 497
rect 275 429 286 463
rect 320 429 331 463
rect 275 417 331 429
rect 381 599 434 617
rect 381 565 392 599
rect 426 565 434 599
rect 381 531 434 565
rect 381 497 392 531
rect 426 497 434 531
rect 381 463 434 497
rect 381 429 392 463
rect 426 429 434 463
rect 381 417 434 429
<< ndiffc >>
rect 35 71 69 105
rect 193 71 227 105
rect 351 71 385 105
rect 509 71 543 105
<< pdiffc >>
rect 74 565 108 599
rect 74 497 108 531
rect 74 429 108 463
rect 180 565 214 599
rect 180 497 214 531
rect 180 429 214 463
rect 286 565 320 599
rect 286 497 320 531
rect 286 429 320 463
rect 392 565 426 599
rect 392 497 426 531
rect 392 429 426 463
<< poly >>
rect 119 617 169 645
rect 225 617 275 645
rect 331 617 381 645
rect 119 221 169 417
rect 225 309 275 417
rect 331 309 381 417
rect 211 293 500 309
rect 211 259 227 293
rect 261 259 500 293
rect 211 241 500 259
rect 80 210 169 221
rect 80 205 182 210
rect 80 171 119 205
rect 153 171 182 205
rect 80 155 182 171
rect 80 131 110 155
rect 152 131 182 155
rect 238 131 268 241
rect 310 131 340 241
rect 396 131 426 241
rect 468 131 498 241
rect 80 21 110 47
rect 152 21 182 47
rect 238 21 268 47
rect 310 21 340 47
rect 396 21 426 47
rect 468 21 498 47
<< polycont >>
rect 227 259 261 293
rect 119 171 153 205
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 58 599 124 615
rect 58 565 74 599
rect 108 565 124 599
rect 58 531 124 565
rect 58 497 74 531
rect 108 497 124 531
rect 58 463 124 497
rect 58 429 74 463
rect 108 429 124 463
rect 58 364 124 429
rect 164 599 230 649
rect 164 565 180 599
rect 214 565 230 599
rect 164 531 230 565
rect 164 497 180 531
rect 214 497 230 531
rect 164 463 230 497
rect 164 429 180 463
rect 214 429 230 463
rect 164 413 230 429
rect 264 599 336 615
rect 264 565 286 599
rect 320 565 336 599
rect 264 531 336 565
rect 264 497 286 531
rect 320 497 336 531
rect 264 463 336 497
rect 264 429 286 463
rect 320 429 336 463
rect 19 307 124 364
rect 264 375 336 429
rect 376 599 442 649
rect 376 565 392 599
rect 426 565 442 599
rect 376 531 442 565
rect 376 497 392 531
rect 426 497 442 531
rect 376 463 442 497
rect 376 429 392 463
rect 426 429 442 463
rect 376 417 442 429
rect 264 341 454 375
rect 19 293 277 307
rect 19 259 227 293
rect 261 259 277 293
rect 19 255 277 259
rect 19 105 75 255
rect 111 205 265 221
rect 111 171 119 205
rect 153 171 265 205
rect 111 155 265 171
rect 19 71 35 105
rect 69 71 75 105
rect 19 53 75 71
rect 177 105 243 121
rect 177 71 193 105
rect 227 71 243 105
rect 177 17 243 71
rect 311 105 454 341
rect 311 71 351 105
rect 385 71 454 105
rect 311 53 454 71
rect 493 105 559 121
rect 493 71 509 105
rect 543 71 559 105
rect 493 17 559 71
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkbuflp_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5393896
string GDS_START 5388348
<< end >>
