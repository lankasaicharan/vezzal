magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 103 49 830 165
rect 0 0 864 49
<< scnmos >>
rect 186 55 216 139
rect 272 55 302 139
rect 374 55 404 139
rect 615 55 645 139
rect 701 55 731 139
<< scpmoshvt >>
rect 170 419 220 619
rect 297 419 347 619
rect 395 419 445 619
rect 509 419 559 619
rect 607 419 657 619
<< ndiff >>
rect 129 115 186 139
rect 129 81 141 115
rect 175 81 186 115
rect 129 55 186 81
rect 216 115 272 139
rect 216 81 227 115
rect 261 81 272 115
rect 216 55 272 81
rect 302 115 374 139
rect 302 81 329 115
rect 363 81 374 115
rect 302 55 374 81
rect 404 101 615 139
rect 404 67 431 101
rect 465 67 615 101
rect 404 55 615 67
rect 645 115 701 139
rect 645 81 656 115
rect 690 81 701 115
rect 645 55 701 81
rect 731 115 804 139
rect 731 81 758 115
rect 792 81 804 115
rect 731 55 804 81
<< pdiff >>
rect 113 597 170 619
rect 113 563 125 597
rect 159 563 170 597
rect 113 465 170 563
rect 113 431 125 465
rect 159 431 170 465
rect 113 419 170 431
rect 220 602 297 619
rect 220 568 231 602
rect 265 568 297 602
rect 220 419 297 568
rect 347 419 395 619
rect 445 570 509 619
rect 445 536 456 570
rect 490 536 509 570
rect 445 419 509 536
rect 559 419 607 619
rect 657 575 714 619
rect 657 541 668 575
rect 702 541 714 575
rect 657 419 714 541
<< ndiffc >>
rect 141 81 175 115
rect 227 81 261 115
rect 329 81 363 115
rect 431 67 465 101
rect 656 81 690 115
rect 758 81 792 115
<< pdiffc >>
rect 125 563 159 597
rect 125 431 159 465
rect 231 568 265 602
rect 456 536 490 570
rect 668 541 702 575
<< poly >>
rect 170 619 220 645
rect 297 619 347 645
rect 395 619 445 645
rect 509 619 559 645
rect 607 619 657 645
rect 170 344 220 419
rect 297 370 347 419
rect 109 328 220 344
rect 109 294 125 328
rect 159 314 220 328
rect 272 354 347 370
rect 272 320 297 354
rect 331 320 347 354
rect 395 387 445 419
rect 395 371 461 387
rect 395 337 411 371
rect 445 337 461 371
rect 395 321 461 337
rect 509 365 559 419
rect 159 294 216 314
rect 109 260 216 294
rect 109 226 125 260
rect 159 226 216 260
rect 109 210 216 226
rect 186 139 216 210
rect 272 286 347 320
rect 272 252 297 286
rect 331 252 347 286
rect 509 273 539 365
rect 607 361 657 419
rect 607 317 637 361
rect 272 236 347 252
rect 404 257 539 273
rect 272 139 302 236
rect 404 223 420 257
rect 454 243 539 257
rect 587 301 653 317
rect 587 267 603 301
rect 637 267 653 301
rect 454 223 470 243
rect 404 188 470 223
rect 374 158 470 188
rect 587 233 653 267
rect 587 199 603 233
rect 637 199 653 233
rect 587 183 653 199
rect 701 297 767 313
rect 701 263 717 297
rect 751 263 767 297
rect 701 229 767 263
rect 701 195 717 229
rect 751 195 767 229
rect 374 139 404 158
rect 615 139 645 183
rect 701 179 767 195
rect 701 139 731 179
rect 186 29 216 55
rect 272 29 302 55
rect 374 29 404 55
rect 615 29 645 55
rect 701 29 731 55
<< polycont >>
rect 125 294 159 328
rect 297 320 331 354
rect 411 337 445 371
rect 125 226 159 260
rect 297 252 331 286
rect 420 223 454 257
rect 603 267 637 301
rect 603 199 637 233
rect 717 263 751 297
rect 717 195 751 229
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 25 597 175 613
rect 25 563 125 597
rect 159 563 175 597
rect 215 602 281 649
rect 215 568 231 602
rect 265 568 281 602
rect 215 563 281 568
rect 440 570 506 613
rect 25 527 175 563
rect 440 536 456 570
rect 490 536 506 570
rect 440 527 506 536
rect 25 493 506 527
rect 652 575 718 649
rect 652 541 668 575
rect 702 541 718 575
rect 652 493 718 541
rect 25 465 175 493
rect 25 431 125 465
rect 159 431 175 465
rect 25 384 175 431
rect 211 423 837 457
rect 25 143 59 384
rect 109 328 175 344
rect 109 294 125 328
rect 159 294 175 328
rect 109 260 175 294
rect 109 226 125 260
rect 159 226 175 260
rect 109 210 175 226
rect 211 179 245 423
rect 395 371 767 387
rect 281 354 359 370
rect 281 320 297 354
rect 331 320 359 354
rect 395 337 411 371
rect 445 353 767 371
rect 445 337 461 353
rect 395 321 461 337
rect 281 286 359 320
rect 281 252 297 286
rect 331 252 359 286
rect 587 301 653 317
rect 281 236 359 252
rect 404 257 551 282
rect 404 223 420 257
rect 454 223 551 257
rect 404 207 551 223
rect 587 267 603 301
rect 637 267 653 301
rect 587 233 653 267
rect 587 199 603 233
rect 637 199 653 233
rect 587 183 653 199
rect 697 297 767 353
rect 697 263 717 297
rect 751 263 767 297
rect 697 229 767 263
rect 697 195 717 229
rect 751 195 767 229
rect 697 179 767 195
rect 25 115 175 143
rect 25 81 141 115
rect 25 53 175 81
rect 211 115 277 179
rect 211 81 227 115
rect 261 81 277 115
rect 211 53 277 81
rect 313 143 551 171
rect 803 143 837 423
rect 313 137 706 143
rect 313 115 379 137
rect 313 81 329 115
rect 363 81 379 115
rect 517 115 706 137
rect 517 109 656 115
rect 313 53 379 81
rect 415 67 431 101
rect 465 67 481 101
rect 415 17 481 67
rect 640 81 656 109
rect 690 81 706 115
rect 640 53 706 81
rect 742 115 837 143
rect 742 81 758 115
rect 792 81 837 115
rect 742 53 837 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221ai_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5814792
string GDS_START 5807584
<< end >>
