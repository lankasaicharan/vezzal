magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 1 228 383 248
rect 585 228 860 248
rect 1 49 860 228
rect 0 0 864 49
<< scnmos >>
rect 84 74 114 222
rect 170 74 200 222
rect 270 74 300 222
rect 470 74 500 202
rect 548 74 578 202
rect 661 74 691 222
rect 747 74 777 222
<< scpmoshvt >>
rect 87 392 117 592
rect 171 392 201 592
rect 273 392 303 592
rect 402 393 432 561
rect 510 393 540 561
rect 658 368 688 592
rect 748 368 778 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 188 170 222
rect 114 154 125 188
rect 159 154 170 188
rect 114 116 170 154
rect 114 82 125 116
rect 159 82 170 116
rect 114 74 170 82
rect 200 210 270 222
rect 200 176 211 210
rect 245 176 270 210
rect 200 120 270 176
rect 200 86 211 120
rect 245 86 270 120
rect 200 74 270 86
rect 300 193 357 222
rect 611 202 661 222
rect 300 159 311 193
rect 345 159 357 193
rect 300 116 357 159
rect 300 82 311 116
rect 345 82 357 116
rect 300 74 357 82
rect 413 179 470 202
rect 413 145 425 179
rect 459 145 470 179
rect 413 74 470 145
rect 500 74 548 202
rect 578 193 661 202
rect 578 159 593 193
rect 627 159 661 193
rect 578 116 661 159
rect 578 82 593 116
rect 627 82 661 116
rect 578 74 661 82
rect 691 210 747 222
rect 691 176 702 210
rect 736 176 747 210
rect 691 120 747 176
rect 691 86 702 120
rect 736 86 747 120
rect 691 74 747 86
rect 777 210 834 222
rect 777 176 788 210
rect 822 176 834 210
rect 777 120 834 176
rect 777 86 788 120
rect 822 86 834 120
rect 777 74 834 86
<< pdiff >>
rect 321 597 384 609
rect 321 592 335 597
rect 28 580 87 592
rect 28 546 40 580
rect 74 546 87 580
rect 28 510 87 546
rect 28 476 40 510
rect 74 476 87 510
rect 28 440 87 476
rect 28 406 40 440
rect 74 406 87 440
rect 28 392 87 406
rect 117 392 171 592
rect 201 580 273 592
rect 201 546 226 580
rect 260 546 273 580
rect 201 510 273 546
rect 201 476 226 510
rect 260 476 273 510
rect 201 440 273 476
rect 201 406 226 440
rect 260 406 273 440
rect 201 392 273 406
rect 303 563 335 592
rect 369 563 384 597
rect 558 597 640 609
rect 303 561 384 563
rect 558 563 582 597
rect 616 592 640 597
rect 616 563 658 592
rect 558 561 658 563
rect 303 393 402 561
rect 432 445 510 561
rect 432 411 454 445
rect 488 411 510 445
rect 432 393 510 411
rect 540 393 658 561
rect 303 392 356 393
rect 605 368 658 393
rect 688 580 748 592
rect 688 546 701 580
rect 735 546 748 580
rect 688 497 748 546
rect 688 463 701 497
rect 735 463 748 497
rect 688 414 748 463
rect 688 380 701 414
rect 735 380 748 414
rect 688 368 748 380
rect 778 580 837 592
rect 778 546 791 580
rect 825 546 837 580
rect 778 497 837 546
rect 778 463 791 497
rect 825 463 837 497
rect 778 414 837 463
rect 778 380 791 414
rect 825 380 837 414
rect 778 368 837 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 154 159 188
rect 125 82 159 116
rect 211 176 245 210
rect 211 86 245 120
rect 311 159 345 193
rect 311 82 345 116
rect 425 145 459 179
rect 593 159 627 193
rect 593 82 627 116
rect 702 176 736 210
rect 702 86 736 120
rect 788 176 822 210
rect 788 86 822 120
<< pdiffc >>
rect 40 546 74 580
rect 40 476 74 510
rect 40 406 74 440
rect 226 546 260 580
rect 226 476 260 510
rect 226 406 260 440
rect 335 563 369 597
rect 582 563 616 597
rect 454 411 488 445
rect 701 546 735 580
rect 701 463 735 497
rect 701 380 735 414
rect 791 546 825 580
rect 791 463 825 497
rect 791 380 825 414
<< poly >>
rect 87 592 117 618
rect 171 592 201 618
rect 273 592 303 618
rect 402 561 432 587
rect 510 561 540 587
rect 658 592 688 618
rect 748 592 778 618
rect 87 377 117 392
rect 171 377 201 392
rect 273 377 303 392
rect 402 378 432 393
rect 510 378 540 393
rect 84 356 120 377
rect 168 356 204 377
rect 270 356 306 377
rect 399 361 435 378
rect 507 361 543 378
rect 48 340 120 356
rect 48 306 64 340
rect 98 326 120 340
rect 162 340 228 356
rect 98 306 114 326
rect 48 290 114 306
rect 162 306 178 340
rect 212 306 228 340
rect 162 290 228 306
rect 270 340 357 356
rect 270 306 307 340
rect 341 306 357 340
rect 270 290 357 306
rect 399 345 465 361
rect 399 311 415 345
rect 449 311 465 345
rect 399 295 465 311
rect 507 345 578 361
rect 658 353 688 368
rect 748 353 778 368
rect 507 311 523 345
rect 557 311 578 345
rect 655 327 691 353
rect 745 327 781 353
rect 507 295 578 311
rect 84 222 114 290
rect 170 222 200 290
rect 270 222 300 290
rect 435 247 465 295
rect 435 217 500 247
rect 470 202 500 217
rect 548 202 578 295
rect 620 311 781 327
rect 620 277 636 311
rect 670 277 781 311
rect 620 261 781 277
rect 661 222 691 261
rect 747 222 777 261
rect 84 48 114 74
rect 170 48 200 74
rect 270 48 300 74
rect 470 48 500 74
rect 548 48 578 74
rect 661 48 691 74
rect 747 48 777 74
<< polycont >>
rect 64 306 98 340
rect 178 306 212 340
rect 307 306 341 340
rect 415 311 449 345
rect 523 311 557 345
rect 636 277 670 311
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 24 580 90 649
rect 317 597 388 649
rect 24 546 40 580
rect 74 546 90 580
rect 24 510 90 546
rect 24 476 40 510
rect 74 476 90 510
rect 24 440 90 476
rect 24 406 40 440
rect 74 406 90 440
rect 24 390 90 406
rect 210 580 276 596
rect 210 546 226 580
rect 260 546 276 580
rect 317 563 335 597
rect 369 563 388 597
rect 317 547 388 563
rect 554 597 644 649
rect 554 563 582 597
rect 616 563 644 597
rect 554 547 644 563
rect 685 580 754 596
rect 210 513 276 546
rect 685 546 701 580
rect 735 546 754 580
rect 210 510 651 513
rect 210 476 226 510
rect 260 479 651 510
rect 260 476 276 479
rect 210 440 276 476
rect 210 406 226 440
rect 260 406 276 440
rect 210 390 276 406
rect 323 411 454 445
rect 488 411 513 445
rect 323 395 513 411
rect 323 356 357 395
rect 25 340 114 356
rect 25 306 64 340
rect 98 306 114 340
rect 25 290 114 306
rect 162 340 257 356
rect 162 306 178 340
rect 212 306 257 340
rect 162 290 257 306
rect 291 340 357 356
rect 291 306 307 340
rect 341 306 357 340
rect 291 290 357 306
rect 399 345 465 361
rect 399 311 415 345
rect 449 311 465 345
rect 399 295 465 311
rect 505 345 573 361
rect 505 311 523 345
rect 557 311 573 345
rect 505 295 573 311
rect 617 327 651 479
rect 685 497 754 546
rect 685 463 701 497
rect 735 463 754 497
rect 685 414 754 463
rect 685 380 701 414
rect 735 380 754 414
rect 685 364 754 380
rect 791 580 841 649
rect 825 546 841 580
rect 791 497 841 546
rect 825 463 841 497
rect 791 414 841 463
rect 825 380 841 414
rect 791 364 841 380
rect 617 311 686 327
rect 323 261 357 290
rect 617 277 636 311
rect 670 277 686 311
rect 617 261 686 277
rect 23 222 261 256
rect 323 227 475 261
rect 23 210 73 222
rect 23 176 39 210
rect 211 210 261 222
rect 23 120 73 176
rect 23 86 39 120
rect 23 70 73 86
rect 109 154 125 188
rect 159 154 175 188
rect 109 116 175 154
rect 109 82 125 116
rect 159 82 175 116
rect 109 17 175 82
rect 245 176 261 210
rect 211 120 261 176
rect 245 86 261 120
rect 211 70 261 86
rect 295 159 311 193
rect 345 159 361 193
rect 295 116 361 159
rect 409 179 475 227
rect 409 145 425 179
rect 459 145 475 179
rect 409 119 475 145
rect 509 227 651 261
rect 295 82 311 116
rect 345 85 361 116
rect 509 85 543 227
rect 720 226 754 364
rect 686 210 754 226
rect 345 82 543 85
rect 295 51 543 82
rect 577 159 593 193
rect 627 159 643 193
rect 577 116 643 159
rect 577 82 593 116
rect 627 82 643 116
rect 577 17 643 82
rect 686 176 702 210
rect 736 176 754 210
rect 686 120 754 176
rect 686 86 702 120
rect 736 86 754 120
rect 686 70 754 86
rect 788 210 838 226
rect 822 176 838 210
rect 788 120 838 176
rect 822 86 838 120
rect 788 17 838 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o2bb2a_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 2214212
string GDS_START 2206160
<< end >>
