magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3506 1852
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 1 21 2200 203
rect 29 -17 63 21
<< scnmos >>
rect 82 47 112 177
rect 176 47 206 177
rect 270 47 300 177
rect 374 47 404 177
rect 458 47 488 177
rect 552 47 582 177
rect 646 47 676 177
rect 740 47 770 177
rect 938 47 968 177
rect 1032 47 1062 177
rect 1126 47 1156 177
rect 1230 47 1260 177
rect 1314 47 1344 177
rect 1408 47 1438 177
rect 1502 47 1532 177
rect 1606 47 1636 177
rect 1796 47 1826 177
rect 1890 47 1920 177
rect 1984 47 2014 177
rect 2088 47 2118 177
<< scpmoshvt >>
rect 84 297 120 497
rect 178 297 214 497
rect 272 297 308 497
rect 366 297 402 497
rect 460 297 496 497
rect 554 297 590 497
rect 648 297 684 497
rect 742 297 778 497
rect 940 297 976 497
rect 1034 297 1070 497
rect 1128 297 1164 497
rect 1222 297 1258 497
rect 1316 297 1352 497
rect 1410 297 1446 497
rect 1504 297 1540 497
rect 1598 297 1634 497
rect 1798 297 1834 497
rect 1892 297 1928 497
rect 1986 297 2022 497
rect 2080 297 2116 497
<< ndiff >>
rect 27 95 82 177
rect 27 61 38 95
rect 72 61 82 95
rect 27 47 82 61
rect 112 163 176 177
rect 112 129 132 163
rect 166 129 176 163
rect 112 95 176 129
rect 112 61 132 95
rect 166 61 176 95
rect 112 47 176 61
rect 206 95 270 177
rect 206 61 226 95
rect 260 61 270 95
rect 206 47 270 61
rect 300 163 374 177
rect 300 129 320 163
rect 354 129 374 163
rect 300 95 374 129
rect 300 61 320 95
rect 354 61 374 95
rect 300 47 374 61
rect 404 95 458 177
rect 404 61 414 95
rect 448 61 458 95
rect 404 47 458 61
rect 488 163 552 177
rect 488 129 508 163
rect 542 129 552 163
rect 488 95 552 129
rect 488 61 508 95
rect 542 61 552 95
rect 488 47 552 61
rect 582 95 646 177
rect 582 61 602 95
rect 636 61 646 95
rect 582 47 646 61
rect 676 163 740 177
rect 676 129 696 163
rect 730 129 740 163
rect 676 95 740 129
rect 676 61 696 95
rect 730 61 740 95
rect 676 47 740 61
rect 770 163 832 177
rect 770 129 790 163
rect 824 129 832 163
rect 770 95 832 129
rect 770 61 790 95
rect 824 61 832 95
rect 770 47 832 61
rect 886 95 938 177
rect 886 61 894 95
rect 928 61 938 95
rect 886 47 938 61
rect 968 163 1032 177
rect 968 129 988 163
rect 1022 129 1032 163
rect 968 47 1032 129
rect 1062 95 1126 177
rect 1062 61 1082 95
rect 1116 61 1126 95
rect 1062 47 1126 61
rect 1156 163 1230 177
rect 1156 129 1176 163
rect 1210 129 1230 163
rect 1156 47 1230 129
rect 1260 163 1314 177
rect 1260 129 1270 163
rect 1304 129 1314 163
rect 1260 95 1314 129
rect 1260 61 1270 95
rect 1304 61 1314 95
rect 1260 47 1314 61
rect 1344 95 1408 177
rect 1344 61 1364 95
rect 1398 61 1408 95
rect 1344 47 1408 61
rect 1438 163 1502 177
rect 1438 129 1458 163
rect 1492 129 1502 163
rect 1438 95 1502 129
rect 1438 61 1458 95
rect 1492 61 1502 95
rect 1438 47 1502 61
rect 1532 95 1606 177
rect 1532 61 1552 95
rect 1586 61 1606 95
rect 1532 47 1606 61
rect 1636 163 1688 177
rect 1636 129 1646 163
rect 1680 129 1688 163
rect 1636 95 1688 129
rect 1636 61 1646 95
rect 1680 61 1688 95
rect 1636 47 1688 61
rect 1744 95 1796 177
rect 1744 61 1752 95
rect 1786 61 1796 95
rect 1744 47 1796 61
rect 1826 163 1890 177
rect 1826 129 1846 163
rect 1880 129 1890 163
rect 1826 95 1890 129
rect 1826 61 1846 95
rect 1880 61 1890 95
rect 1826 47 1890 61
rect 1920 95 1984 177
rect 1920 61 1940 95
rect 1974 61 1984 95
rect 1920 47 1984 61
rect 2014 163 2088 177
rect 2014 129 2034 163
rect 2068 129 2088 163
rect 2014 95 2088 129
rect 2014 61 2034 95
rect 2068 61 2088 95
rect 2014 47 2088 61
rect 2118 95 2174 177
rect 2118 61 2128 95
rect 2162 61 2174 95
rect 2118 47 2174 61
<< pdiff >>
rect 27 477 84 497
rect 27 443 38 477
rect 72 443 84 477
rect 27 409 84 443
rect 27 375 38 409
rect 72 375 84 409
rect 27 297 84 375
rect 120 485 178 497
rect 120 451 132 485
rect 166 451 178 485
rect 120 297 178 451
rect 214 477 272 497
rect 214 443 226 477
rect 260 443 272 477
rect 214 409 272 443
rect 214 375 226 409
rect 260 375 272 409
rect 214 297 272 375
rect 308 485 366 497
rect 308 451 320 485
rect 354 451 366 485
rect 308 297 366 451
rect 402 477 460 497
rect 402 443 414 477
rect 448 443 460 477
rect 402 409 460 443
rect 402 375 414 409
rect 448 375 460 409
rect 402 297 460 375
rect 496 409 554 497
rect 496 375 508 409
rect 542 375 554 409
rect 496 297 554 375
rect 590 477 648 497
rect 590 443 602 477
rect 636 443 648 477
rect 590 297 648 443
rect 684 409 742 497
rect 684 375 696 409
rect 730 375 742 409
rect 684 297 742 375
rect 778 477 832 497
rect 778 443 790 477
rect 824 443 832 477
rect 778 409 832 443
rect 778 375 790 409
rect 824 375 832 409
rect 778 297 832 375
rect 886 477 940 497
rect 886 443 894 477
rect 928 443 940 477
rect 886 409 940 443
rect 886 375 894 409
rect 928 375 940 409
rect 886 297 940 375
rect 976 485 1034 497
rect 976 451 988 485
rect 1022 451 1034 485
rect 976 297 1034 451
rect 1070 477 1128 497
rect 1070 443 1082 477
rect 1116 443 1128 477
rect 1070 409 1128 443
rect 1070 375 1082 409
rect 1116 375 1128 409
rect 1070 297 1128 375
rect 1164 485 1222 497
rect 1164 451 1176 485
rect 1210 451 1222 485
rect 1164 297 1222 451
rect 1258 477 1316 497
rect 1258 443 1270 477
rect 1304 443 1316 477
rect 1258 409 1316 443
rect 1258 375 1270 409
rect 1304 375 1316 409
rect 1258 297 1316 375
rect 1352 485 1410 497
rect 1352 451 1364 485
rect 1398 451 1410 485
rect 1352 297 1410 451
rect 1446 477 1504 497
rect 1446 443 1458 477
rect 1492 443 1504 477
rect 1446 409 1504 443
rect 1446 375 1458 409
rect 1492 375 1504 409
rect 1446 341 1504 375
rect 1446 307 1458 341
rect 1492 307 1504 341
rect 1446 297 1504 307
rect 1540 485 1598 497
rect 1540 451 1552 485
rect 1586 451 1598 485
rect 1540 297 1598 451
rect 1634 477 1688 497
rect 1634 443 1646 477
rect 1680 443 1688 477
rect 1634 409 1688 443
rect 1634 375 1646 409
rect 1680 375 1688 409
rect 1634 361 1688 375
rect 1742 409 1798 497
rect 1742 375 1752 409
rect 1786 375 1798 409
rect 1634 297 1686 361
rect 1742 346 1798 375
rect 1740 339 1798 346
rect 1740 305 1752 339
rect 1786 305 1798 339
rect 1740 297 1798 305
rect 1834 485 1892 497
rect 1834 451 1846 485
rect 1880 451 1892 485
rect 1834 417 1892 451
rect 1834 383 1846 417
rect 1880 383 1892 417
rect 1834 297 1892 383
rect 1928 409 1986 497
rect 1928 375 1940 409
rect 1974 375 1986 409
rect 1928 341 1986 375
rect 1928 307 1940 341
rect 1974 307 1986 341
rect 1928 297 1986 307
rect 2022 477 2080 497
rect 2022 443 2034 477
rect 2068 443 2080 477
rect 2022 409 2080 443
rect 2022 375 2034 409
rect 2068 375 2080 409
rect 2022 297 2080 375
rect 2116 477 2174 497
rect 2116 443 2128 477
rect 2162 443 2174 477
rect 2116 409 2174 443
rect 2116 375 2128 409
rect 2162 375 2174 409
rect 2116 341 2174 375
rect 2116 307 2128 341
rect 2162 307 2174 341
rect 2116 297 2174 307
<< ndiffc >>
rect 38 61 72 95
rect 132 129 166 163
rect 132 61 166 95
rect 226 61 260 95
rect 320 129 354 163
rect 320 61 354 95
rect 414 61 448 95
rect 508 129 542 163
rect 508 61 542 95
rect 602 61 636 95
rect 696 129 730 163
rect 696 61 730 95
rect 790 129 824 163
rect 790 61 824 95
rect 894 61 928 95
rect 988 129 1022 163
rect 1082 61 1116 95
rect 1176 129 1210 163
rect 1270 129 1304 163
rect 1270 61 1304 95
rect 1364 61 1398 95
rect 1458 129 1492 163
rect 1458 61 1492 95
rect 1552 61 1586 95
rect 1646 129 1680 163
rect 1646 61 1680 95
rect 1752 61 1786 95
rect 1846 129 1880 163
rect 1846 61 1880 95
rect 1940 61 1974 95
rect 2034 129 2068 163
rect 2034 61 2068 95
rect 2128 61 2162 95
<< pdiffc >>
rect 38 443 72 477
rect 38 375 72 409
rect 132 451 166 485
rect 226 443 260 477
rect 226 375 260 409
rect 320 451 354 485
rect 414 443 448 477
rect 414 375 448 409
rect 508 375 542 409
rect 602 443 636 477
rect 696 375 730 409
rect 790 443 824 477
rect 790 375 824 409
rect 894 443 928 477
rect 894 375 928 409
rect 988 451 1022 485
rect 1082 443 1116 477
rect 1082 375 1116 409
rect 1176 451 1210 485
rect 1270 443 1304 477
rect 1270 375 1304 409
rect 1364 451 1398 485
rect 1458 443 1492 477
rect 1458 375 1492 409
rect 1458 307 1492 341
rect 1552 451 1586 485
rect 1646 443 1680 477
rect 1646 375 1680 409
rect 1752 375 1786 409
rect 1752 305 1786 339
rect 1846 451 1880 485
rect 1846 383 1880 417
rect 1940 375 1974 409
rect 1940 307 1974 341
rect 2034 443 2068 477
rect 2034 375 2068 409
rect 2128 443 2162 477
rect 2128 375 2162 409
rect 2128 307 2162 341
<< poly >>
rect 84 497 120 523
rect 178 497 214 523
rect 272 497 308 523
rect 366 497 402 523
rect 460 497 496 523
rect 554 497 590 523
rect 648 497 684 523
rect 742 497 778 523
rect 940 497 976 523
rect 1034 497 1070 523
rect 1128 497 1164 523
rect 1222 497 1258 523
rect 1316 497 1352 523
rect 1410 497 1446 523
rect 1504 497 1540 523
rect 1598 497 1634 523
rect 1798 497 1834 523
rect 1892 497 1928 523
rect 1986 497 2022 523
rect 2080 497 2116 523
rect 84 282 120 297
rect 178 282 214 297
rect 272 282 308 297
rect 366 282 402 297
rect 460 282 496 297
rect 554 282 590 297
rect 648 282 684 297
rect 742 282 778 297
rect 940 282 976 297
rect 1034 282 1070 297
rect 1128 282 1164 297
rect 1222 282 1258 297
rect 1316 282 1352 297
rect 1410 282 1446 297
rect 1504 282 1540 297
rect 1598 282 1634 297
rect 1798 282 1834 297
rect 1892 282 1928 297
rect 1986 282 2022 297
rect 2080 282 2116 297
rect 82 265 122 282
rect 176 265 216 282
rect 270 265 310 282
rect 364 265 404 282
rect 82 249 404 265
rect 82 215 102 249
rect 136 215 180 249
rect 214 215 258 249
rect 292 215 336 249
rect 370 215 404 249
rect 82 199 404 215
rect 82 177 112 199
rect 176 177 206 199
rect 270 177 300 199
rect 374 177 404 199
rect 458 265 498 282
rect 552 265 592 282
rect 646 265 686 282
rect 740 265 780 282
rect 938 265 978 282
rect 1032 265 1072 282
rect 1126 265 1166 282
rect 1220 265 1260 282
rect 458 249 1260 265
rect 458 215 670 249
rect 704 215 748 249
rect 782 215 826 249
rect 860 215 894 249
rect 928 215 962 249
rect 996 215 1040 249
rect 1074 215 1260 249
rect 458 199 1260 215
rect 458 177 488 199
rect 552 177 582 199
rect 646 177 676 199
rect 740 177 770 199
rect 938 177 968 199
rect 1032 177 1062 199
rect 1126 177 1156 199
rect 1230 177 1260 199
rect 1314 265 1354 282
rect 1408 265 1448 282
rect 1502 265 1542 282
rect 1596 265 1636 282
rect 1314 249 1636 265
rect 1314 215 1337 249
rect 1371 215 1415 249
rect 1449 215 1493 249
rect 1527 215 1571 249
rect 1605 215 1636 249
rect 1314 199 1636 215
rect 1314 177 1344 199
rect 1408 177 1438 199
rect 1502 177 1532 199
rect 1606 177 1636 199
rect 1796 265 1836 282
rect 1890 265 1930 282
rect 1984 265 2024 282
rect 2078 265 2118 282
rect 1796 249 2118 265
rect 1796 215 1812 249
rect 1846 215 1894 249
rect 1928 215 1972 249
rect 2006 215 2118 249
rect 1796 199 2118 215
rect 1796 177 1826 199
rect 1890 177 1920 199
rect 1984 177 2014 199
rect 2088 177 2118 199
rect 82 21 112 47
rect 176 21 206 47
rect 270 21 300 47
rect 374 21 404 47
rect 458 21 488 47
rect 552 21 582 47
rect 646 21 676 47
rect 740 21 770 47
rect 938 21 968 47
rect 1032 21 1062 47
rect 1126 21 1156 47
rect 1230 21 1260 47
rect 1314 21 1344 47
rect 1408 21 1438 47
rect 1502 21 1532 47
rect 1606 21 1636 47
rect 1796 21 1826 47
rect 1890 21 1920 47
rect 1984 21 2014 47
rect 2088 21 2118 47
<< polycont >>
rect 102 215 136 249
rect 180 215 214 249
rect 258 215 292 249
rect 336 215 370 249
rect 670 215 704 249
rect 748 215 782 249
rect 826 215 860 249
rect 894 215 928 249
rect 962 215 996 249
rect 1040 215 1074 249
rect 1337 215 1371 249
rect 1415 215 1449 249
rect 1493 215 1527 249
rect 1571 215 1605 249
rect 1812 215 1846 249
rect 1894 215 1928 249
rect 1972 215 2006 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 17 477 80 493
rect 17 443 38 477
rect 72 443 80 477
rect 17 409 80 443
rect 124 485 174 527
rect 124 451 132 485
rect 166 451 174 485
rect 124 435 174 451
rect 218 477 268 493
rect 218 443 226 477
rect 260 443 268 477
rect 17 375 38 409
rect 72 401 80 409
rect 218 409 268 443
rect 312 485 362 527
rect 312 451 320 485
rect 354 451 362 485
rect 312 435 362 451
rect 406 477 832 493
rect 406 443 414 477
rect 448 459 602 477
rect 448 443 456 459
rect 218 401 226 409
rect 72 375 226 401
rect 260 401 268 409
rect 406 409 456 443
rect 594 443 602 459
rect 636 459 790 477
rect 636 443 644 459
rect 594 425 644 443
rect 782 443 790 459
rect 824 443 832 477
rect 406 401 414 409
rect 260 375 414 401
rect 448 375 456 409
rect 17 357 456 375
rect 500 409 550 425
rect 500 375 508 409
rect 542 391 550 409
rect 688 409 738 425
rect 688 391 696 409
rect 542 375 696 391
rect 730 375 738 409
rect 500 357 738 375
rect 782 409 832 443
rect 782 375 790 409
rect 824 375 832 409
rect 782 359 832 375
rect 886 477 936 493
rect 886 443 894 477
rect 928 443 936 477
rect 886 409 936 443
rect 980 485 1030 527
rect 980 451 988 485
rect 1022 451 1030 485
rect 980 435 1030 451
rect 1074 477 1124 493
rect 1074 443 1082 477
rect 1116 443 1124 477
rect 886 375 894 409
rect 928 401 936 409
rect 1074 409 1124 443
rect 1168 485 1218 527
rect 1168 451 1176 485
rect 1210 451 1218 485
rect 1168 435 1218 451
rect 1262 477 1312 493
rect 1262 443 1270 477
rect 1304 443 1312 477
rect 1074 401 1082 409
rect 928 375 1082 401
rect 1116 401 1124 409
rect 1262 409 1312 443
rect 1356 485 1406 527
rect 1356 451 1364 485
rect 1398 451 1406 485
rect 1356 435 1406 451
rect 1450 477 1500 493
rect 1450 443 1458 477
rect 1492 443 1500 477
rect 1262 401 1270 409
rect 1116 375 1270 401
rect 1304 401 1312 409
rect 1450 409 1500 443
rect 1544 485 1594 527
rect 1544 451 1552 485
rect 1586 451 1594 485
rect 1544 435 1594 451
rect 1638 485 2076 493
rect 1638 477 1846 485
rect 1638 443 1646 477
rect 1680 459 1846 477
rect 1680 443 1688 459
rect 1450 401 1458 409
rect 1304 375 1458 401
rect 1492 401 1500 409
rect 1638 409 1688 443
rect 1838 451 1846 459
rect 1880 477 2076 485
rect 1880 459 2034 477
rect 1880 451 1888 459
rect 1638 401 1646 409
rect 1492 375 1646 401
rect 1680 375 1688 409
rect 886 357 1688 375
rect 1736 409 1794 425
rect 1736 375 1752 409
rect 1786 375 1794 409
rect 500 323 534 357
rect 1450 341 1500 357
rect 17 289 437 323
rect 471 289 534 323
rect 576 289 1363 323
rect 1450 307 1458 341
rect 1492 307 1500 341
rect 1736 339 1794 375
rect 1838 417 1888 451
rect 2026 443 2034 459
rect 2068 443 2076 477
rect 1838 383 1846 417
rect 1880 383 1888 417
rect 1838 367 1888 383
rect 1932 409 1982 425
rect 1932 375 1940 409
rect 1974 375 1982 409
rect 1450 291 1500 307
rect 1602 289 1661 323
rect 1695 289 1702 323
rect 1736 305 1752 339
rect 1786 333 1794 339
rect 1932 341 1982 375
rect 2026 409 2076 443
rect 2026 375 2034 409
rect 2068 375 2076 409
rect 2026 359 2076 375
rect 2110 477 2191 493
rect 2110 443 2128 477
rect 2162 443 2191 477
rect 2110 409 2191 443
rect 2110 375 2128 409
rect 2162 375 2191 409
rect 1932 333 1940 341
rect 1786 307 1940 333
rect 1974 325 1982 341
rect 2110 341 2191 375
rect 2110 325 2128 341
rect 1974 307 2128 325
rect 2162 307 2191 341
rect 1786 305 2191 307
rect 1736 289 2191 305
rect 17 181 51 289
rect 576 255 620 289
rect 1319 255 1363 289
rect 1668 255 1702 289
rect 85 249 620 255
rect 85 215 102 249
rect 136 215 180 249
rect 214 215 258 249
rect 292 215 336 249
rect 370 215 620 249
rect 654 249 1268 255
rect 654 215 670 249
rect 704 215 748 249
rect 782 215 826 249
rect 860 215 894 249
rect 928 215 962 249
rect 996 215 1040 249
rect 1074 221 1268 249
rect 1319 249 1624 255
rect 1074 215 1100 221
rect 1319 215 1337 249
rect 1371 215 1415 249
rect 1449 215 1493 249
rect 1527 215 1571 249
rect 1605 215 1624 249
rect 1668 249 2026 255
rect 1668 215 1812 249
rect 1846 215 1894 249
rect 1928 215 1972 249
rect 2006 215 2026 249
rect 1130 181 1226 187
rect 2127 181 2191 289
rect 17 163 746 181
rect 913 179 1226 181
rect 17 147 132 163
rect 106 129 132 147
rect 166 145 320 163
rect 166 129 182 145
rect 17 95 72 113
rect 17 61 38 95
rect 17 17 72 61
rect 106 95 182 129
rect 294 129 320 145
rect 354 145 508 163
rect 354 129 370 145
rect 106 61 132 95
rect 166 61 182 95
rect 106 51 182 61
rect 226 95 260 111
rect 226 17 260 61
rect 294 95 370 129
rect 482 129 508 145
rect 542 145 696 163
rect 542 129 558 145
rect 294 61 320 95
rect 354 61 370 95
rect 294 51 370 61
rect 414 95 448 111
rect 414 17 448 61
rect 482 95 558 129
rect 670 129 696 145
rect 730 129 746 163
rect 482 61 508 95
rect 542 61 558 95
rect 482 51 558 61
rect 602 95 636 111
rect 602 17 636 61
rect 670 95 746 129
rect 670 61 696 95
rect 730 61 746 95
rect 670 51 746 61
rect 790 163 844 179
rect 824 129 844 163
rect 913 163 1141 179
rect 913 129 988 163
rect 1022 145 1141 163
rect 1175 163 1226 179
rect 1175 145 1176 163
rect 1022 129 1176 145
rect 1210 129 1226 163
rect 1270 163 1696 181
rect 1304 145 1458 163
rect 1304 129 1320 145
rect 790 95 844 129
rect 1270 95 1320 129
rect 1432 129 1458 145
rect 1492 145 1646 163
rect 1492 129 1508 145
rect 824 61 844 95
rect 790 17 844 61
rect 878 61 894 95
rect 928 61 1082 95
rect 1116 61 1270 95
rect 1304 61 1320 95
rect 878 51 1320 61
rect 1364 95 1398 111
rect 1364 17 1398 61
rect 1432 95 1508 129
rect 1620 129 1646 145
rect 1680 129 1696 163
rect 1730 179 2191 181
rect 1730 145 1753 179
rect 1787 163 2191 179
rect 1787 145 1846 163
rect 1432 61 1458 95
rect 1492 61 1508 95
rect 1432 51 1508 61
rect 1552 95 1586 111
rect 1552 17 1586 61
rect 1620 95 1696 129
rect 1820 129 1846 145
rect 1880 147 2034 163
rect 1880 129 1896 147
rect 1620 61 1646 95
rect 1680 61 1696 95
rect 1620 51 1696 61
rect 1752 95 1786 111
rect 1752 17 1786 61
rect 1820 95 1896 129
rect 2008 129 2034 147
rect 2068 147 2191 163
rect 2068 129 2084 147
rect 1820 61 1846 95
rect 1880 61 1896 95
rect 1820 51 1896 61
rect 1940 95 1974 111
rect 1940 17 1974 61
rect 2008 95 2084 129
rect 2008 61 2034 95
rect 2068 61 2084 95
rect 2008 51 2084 61
rect 2128 95 2162 111
rect 2128 17 2162 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 437 289 471 323
rect 1661 289 1695 323
rect 1141 145 1175 179
rect 1753 145 1787 179
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 425 323 483 329
rect 425 289 437 323
rect 471 320 483 323
rect 1649 323 1707 329
rect 1649 320 1661 323
rect 471 292 1661 320
rect 471 289 483 292
rect 425 283 483 289
rect 1649 289 1661 292
rect 1695 289 1707 323
rect 1649 283 1707 289
rect 1129 179 1799 185
rect 1129 145 1141 179
rect 1175 156 1753 179
rect 1175 145 1187 156
rect 1129 139 1187 145
rect 1741 145 1753 156
rect 1787 145 1799 179
rect 1741 139 1799 145
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel locali s 2143 357 2177 391 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel locali s 853 221 887 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xor2_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2208 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 27654
string GDS_START 12384
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
