magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 253 204 731 235
rect 42 49 731 204
rect 0 0 768 49
<< scnmos >>
rect 125 94 155 178
rect 227 94 257 178
rect 329 125 359 209
rect 437 125 467 209
rect 509 125 539 209
rect 621 125 651 209
<< scpmoshvt >>
rect 89 491 119 619
rect 197 491 227 575
rect 269 491 299 575
rect 393 515 423 599
rect 523 515 553 599
rect 644 515 674 599
<< ndiff >>
rect 279 178 329 209
rect 68 136 125 178
rect 68 102 80 136
rect 114 102 125 136
rect 68 94 125 102
rect 155 136 227 178
rect 155 102 182 136
rect 216 102 227 136
rect 155 94 227 102
rect 257 125 329 178
rect 359 184 437 209
rect 359 150 385 184
rect 419 150 437 184
rect 359 125 437 150
rect 467 125 509 209
rect 539 181 621 209
rect 539 147 563 181
rect 597 147 621 181
rect 539 125 621 147
rect 651 197 705 209
rect 651 163 663 197
rect 697 163 705 197
rect 651 125 705 163
rect 257 94 307 125
<< pdiff >>
rect 36 605 89 619
rect 36 571 44 605
rect 78 571 89 605
rect 36 537 89 571
rect 36 503 44 537
rect 78 503 89 537
rect 36 491 89 503
rect 119 607 172 619
rect 119 573 130 607
rect 164 575 172 607
rect 321 575 393 599
rect 164 573 197 575
rect 119 539 197 573
rect 119 505 152 539
rect 186 505 197 539
rect 119 491 197 505
rect 227 491 269 575
rect 299 542 393 575
rect 299 508 329 542
rect 363 515 393 542
rect 423 515 523 599
rect 553 582 644 599
rect 553 548 599 582
rect 633 548 644 582
rect 553 515 644 548
rect 674 572 727 599
rect 674 538 685 572
rect 719 538 727 572
rect 674 515 727 538
rect 363 508 371 515
rect 299 491 371 508
<< ndiffc >>
rect 80 102 114 136
rect 182 102 216 136
rect 385 150 419 184
rect 563 147 597 181
rect 663 163 697 197
<< pdiffc >>
rect 44 571 78 605
rect 44 503 78 537
rect 130 573 164 607
rect 152 505 186 539
rect 329 508 363 542
rect 599 548 633 582
rect 685 538 719 572
<< poly >>
rect 89 619 119 645
rect 197 575 227 601
rect 269 575 299 601
rect 393 599 423 625
rect 523 599 553 625
rect 644 599 674 625
rect 89 334 119 491
rect 197 459 227 491
rect 161 443 227 459
rect 161 409 177 443
rect 211 409 227 443
rect 161 393 227 409
rect 89 318 155 334
rect 89 284 105 318
rect 139 284 155 318
rect 89 250 155 284
rect 89 216 105 250
rect 139 216 155 250
rect 89 200 155 216
rect 197 230 227 393
rect 269 412 299 491
rect 393 483 423 515
rect 393 467 481 483
rect 393 433 431 467
rect 465 433 481 467
rect 393 417 481 433
rect 269 382 317 412
rect 287 343 317 382
rect 523 369 553 515
rect 644 450 674 515
rect 627 434 693 450
rect 627 400 643 434
rect 677 400 693 434
rect 509 353 579 369
rect 287 327 353 343
rect 287 293 303 327
rect 337 313 353 327
rect 509 319 529 353
rect 563 319 579 353
rect 627 366 693 400
rect 627 346 643 366
rect 337 293 467 313
rect 287 283 467 293
rect 287 277 353 283
rect 197 200 257 230
rect 329 209 359 235
rect 437 209 467 283
rect 509 285 579 319
rect 509 251 529 285
rect 563 251 579 285
rect 509 235 579 251
rect 621 332 643 346
rect 677 332 693 366
rect 621 316 693 332
rect 509 209 539 235
rect 621 209 651 316
rect 125 178 155 200
rect 227 178 257 200
rect 329 103 359 125
rect 125 68 155 94
rect 227 68 257 94
rect 329 87 395 103
rect 437 99 467 125
rect 509 99 539 125
rect 621 99 651 125
rect 329 53 345 87
rect 379 53 395 87
rect 329 37 395 53
<< polycont >>
rect 177 409 211 443
rect 105 284 139 318
rect 105 216 139 250
rect 431 433 465 467
rect 643 400 677 434
rect 303 293 337 327
rect 529 319 563 353
rect 529 251 563 285
rect 643 332 677 366
rect 345 53 379 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 605 94 609
rect 17 571 44 605
rect 78 571 94 605
rect 17 537 94 571
rect 17 503 44 537
rect 78 503 94 537
rect 17 487 94 503
rect 128 607 198 649
rect 128 573 130 607
rect 164 573 198 607
rect 128 539 198 573
rect 128 505 152 539
rect 186 505 198 539
rect 128 487 198 505
rect 232 581 561 615
rect 17 140 71 487
rect 232 453 266 581
rect 161 443 266 453
rect 161 409 177 443
rect 211 409 266 443
rect 313 542 379 547
rect 313 508 329 542
rect 363 508 379 542
rect 313 397 379 508
rect 413 467 493 541
rect 413 433 431 467
rect 465 433 493 467
rect 527 498 561 581
rect 595 582 635 649
rect 595 548 599 582
rect 633 548 635 582
rect 595 532 635 548
rect 669 572 747 588
rect 669 538 685 572
rect 719 538 747 572
rect 669 532 747 538
rect 527 464 677 498
rect 413 431 493 433
rect 313 363 423 397
rect 105 318 156 334
rect 139 284 156 318
rect 105 250 156 284
rect 139 216 156 250
rect 200 327 355 329
rect 200 293 303 327
rect 337 293 355 327
rect 200 242 355 293
rect 105 208 156 216
rect 389 208 423 363
rect 105 184 423 208
rect 105 174 385 184
rect 369 150 385 174
rect 419 150 423 184
rect 17 136 130 140
rect 17 102 80 136
rect 114 102 130 136
rect 17 94 130 102
rect 166 136 232 140
rect 166 102 182 136
rect 216 102 232 136
rect 369 134 423 150
rect 166 17 232 102
rect 459 100 493 431
rect 597 434 677 464
rect 597 400 643 434
rect 527 353 563 369
rect 527 319 529 353
rect 527 285 563 319
rect 597 366 677 400
rect 597 332 643 366
rect 597 303 677 332
rect 527 251 529 285
rect 713 269 747 532
rect 563 251 747 269
rect 527 235 747 251
rect 647 207 747 235
rect 647 197 713 207
rect 329 87 493 100
rect 329 53 345 87
rect 379 53 493 87
rect 547 181 613 197
rect 547 147 563 181
rect 597 147 613 181
rect 647 163 663 197
rect 697 163 713 197
rect 647 159 713 163
rect 547 17 613 147
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2_0
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1700566
string GDS_START 1693028
<< end >>
