magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 32 49 920 259
rect 0 0 960 49
<< scnmos >>
rect 111 65 141 233
rect 197 65 227 233
rect 283 65 313 233
rect 453 65 483 233
rect 539 65 569 233
rect 625 65 655 233
rect 725 65 755 233
rect 811 65 841 233
<< scpmoshvt >>
rect 97 367 127 619
rect 183 367 213 619
rect 269 367 299 619
rect 355 367 385 619
rect 545 367 575 619
rect 647 367 677 619
rect 764 367 794 619
rect 850 367 880 619
<< ndiff >>
rect 58 208 111 233
rect 58 174 66 208
rect 100 174 111 208
rect 58 113 111 174
rect 58 79 66 113
rect 100 79 111 113
rect 58 65 111 79
rect 141 132 197 233
rect 141 98 152 132
rect 186 98 197 132
rect 141 65 197 98
rect 227 208 283 233
rect 227 174 238 208
rect 272 174 283 208
rect 227 113 283 174
rect 227 79 238 113
rect 272 79 283 113
rect 227 65 283 79
rect 313 124 453 233
rect 313 90 324 124
rect 358 90 401 124
rect 435 90 453 124
rect 313 65 453 90
rect 483 181 539 233
rect 483 147 494 181
rect 528 147 539 181
rect 483 107 539 147
rect 483 73 494 107
rect 528 73 539 107
rect 483 65 539 73
rect 569 107 625 233
rect 569 73 580 107
rect 614 73 625 107
rect 569 65 625 73
rect 655 181 725 233
rect 655 147 666 181
rect 700 147 725 181
rect 655 107 725 147
rect 655 73 666 107
rect 700 73 725 107
rect 655 65 725 73
rect 755 225 811 233
rect 755 191 766 225
rect 800 191 811 225
rect 755 153 811 191
rect 755 119 766 153
rect 800 119 811 153
rect 755 65 811 119
rect 841 192 894 233
rect 841 158 852 192
rect 886 158 894 192
rect 841 111 894 158
rect 841 77 852 111
rect 886 77 894 111
rect 841 65 894 77
<< pdiff >>
rect 44 599 97 619
rect 44 565 52 599
rect 86 565 97 599
rect 44 505 97 565
rect 44 471 52 505
rect 86 471 97 505
rect 44 413 97 471
rect 44 379 52 413
rect 86 379 97 413
rect 44 367 97 379
rect 127 607 183 619
rect 127 573 138 607
rect 172 573 183 607
rect 127 539 183 573
rect 127 505 138 539
rect 172 505 183 539
rect 127 457 183 505
rect 127 423 138 457
rect 172 423 183 457
rect 127 367 183 423
rect 213 599 269 619
rect 213 565 224 599
rect 258 565 269 599
rect 213 505 269 565
rect 213 471 224 505
rect 258 471 269 505
rect 213 413 269 471
rect 213 379 224 413
rect 258 379 269 413
rect 213 367 269 379
rect 299 599 355 619
rect 299 565 310 599
rect 344 565 355 599
rect 299 529 355 565
rect 299 495 310 529
rect 344 495 355 529
rect 299 457 355 495
rect 299 423 310 457
rect 344 423 355 457
rect 299 367 355 423
rect 385 539 438 619
rect 385 505 396 539
rect 430 505 438 539
rect 385 413 438 505
rect 385 379 396 413
rect 430 379 438 413
rect 385 367 438 379
rect 492 539 545 619
rect 492 505 500 539
rect 534 505 545 539
rect 492 413 545 505
rect 492 379 500 413
rect 534 379 545 413
rect 492 367 545 379
rect 575 597 647 619
rect 575 563 586 597
rect 620 563 647 597
rect 575 508 647 563
rect 575 474 586 508
rect 620 474 647 508
rect 575 367 647 474
rect 677 599 764 619
rect 677 565 699 599
rect 733 565 764 599
rect 677 509 764 565
rect 677 475 699 509
rect 733 475 764 509
rect 677 419 764 475
rect 677 385 699 419
rect 733 385 764 419
rect 677 367 764 385
rect 794 607 850 619
rect 794 573 805 607
rect 839 573 850 607
rect 794 530 850 573
rect 794 496 805 530
rect 839 496 850 530
rect 794 453 850 496
rect 794 419 805 453
rect 839 419 850 453
rect 794 367 850 419
rect 880 599 933 619
rect 880 565 891 599
rect 925 565 933 599
rect 880 507 933 565
rect 880 473 891 507
rect 925 473 933 507
rect 880 413 933 473
rect 880 379 891 413
rect 925 379 933 413
rect 880 367 933 379
<< ndiffc >>
rect 66 174 100 208
rect 66 79 100 113
rect 152 98 186 132
rect 238 174 272 208
rect 238 79 272 113
rect 324 90 358 124
rect 401 90 435 124
rect 494 147 528 181
rect 494 73 528 107
rect 580 73 614 107
rect 666 147 700 181
rect 666 73 700 107
rect 766 191 800 225
rect 766 119 800 153
rect 852 158 886 192
rect 852 77 886 111
<< pdiffc >>
rect 52 565 86 599
rect 52 471 86 505
rect 52 379 86 413
rect 138 573 172 607
rect 138 505 172 539
rect 138 423 172 457
rect 224 565 258 599
rect 224 471 258 505
rect 224 379 258 413
rect 310 565 344 599
rect 310 495 344 529
rect 310 423 344 457
rect 396 505 430 539
rect 396 379 430 413
rect 500 505 534 539
rect 500 379 534 413
rect 586 563 620 597
rect 586 474 620 508
rect 699 565 733 599
rect 699 475 733 509
rect 699 385 733 419
rect 805 573 839 607
rect 805 496 839 530
rect 805 419 839 453
rect 891 565 925 599
rect 891 473 925 507
rect 891 379 925 413
<< poly >>
rect 97 619 127 645
rect 183 619 213 645
rect 269 619 299 645
rect 355 619 385 645
rect 545 619 575 645
rect 647 619 677 645
rect 764 619 794 645
rect 850 619 880 645
rect 97 321 127 367
rect 183 321 213 367
rect 269 321 299 367
rect 355 321 385 367
rect 545 335 575 367
rect 647 335 677 367
rect 75 305 227 321
rect 75 271 91 305
rect 125 271 177 305
rect 211 271 227 305
rect 75 255 227 271
rect 269 305 483 321
rect 269 271 307 305
rect 341 271 405 305
rect 439 271 483 305
rect 545 319 683 335
rect 764 333 794 367
rect 850 333 880 367
rect 545 299 633 319
rect 269 255 483 271
rect 111 233 141 255
rect 197 233 227 255
rect 283 233 313 255
rect 453 233 483 255
rect 539 285 633 299
rect 667 285 683 319
rect 539 269 683 285
rect 725 321 880 333
rect 725 317 918 321
rect 725 283 745 317
rect 779 305 918 317
rect 779 283 868 305
rect 725 271 868 283
rect 902 271 918 305
rect 539 233 569 269
rect 625 233 655 269
rect 725 255 918 271
rect 725 233 755 255
rect 811 233 841 255
rect 111 39 141 65
rect 197 39 227 65
rect 283 39 313 65
rect 453 39 483 65
rect 539 39 569 65
rect 625 39 655 65
rect 725 39 755 65
rect 811 39 841 65
<< polycont >>
rect 91 271 125 305
rect 177 271 211 305
rect 307 271 341 305
rect 405 271 439 305
rect 633 285 667 319
rect 745 283 779 317
rect 868 271 902 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 36 599 102 615
rect 36 565 52 599
rect 86 565 102 599
rect 36 505 102 565
rect 36 471 52 505
rect 86 471 102 505
rect 36 413 102 471
rect 36 379 52 413
rect 86 379 102 413
rect 136 607 174 649
rect 136 573 138 607
rect 172 573 174 607
rect 136 539 174 573
rect 136 505 138 539
rect 172 505 174 539
rect 136 457 174 505
rect 136 423 138 457
rect 172 423 174 457
rect 136 407 174 423
rect 208 599 274 615
rect 208 565 224 599
rect 258 565 274 599
rect 208 505 274 565
rect 208 471 224 505
rect 258 471 274 505
rect 208 413 274 471
rect 36 373 102 379
rect 208 379 224 413
rect 258 379 274 413
rect 308 599 636 615
rect 308 565 310 599
rect 344 597 636 599
rect 344 581 586 597
rect 344 565 346 581
rect 308 529 346 565
rect 584 563 586 581
rect 620 563 636 597
rect 308 495 310 529
rect 344 495 346 529
rect 308 457 346 495
rect 308 423 310 457
rect 344 423 346 457
rect 308 407 346 423
rect 380 539 446 547
rect 380 505 396 539
rect 430 505 446 539
rect 380 413 446 505
rect 208 373 274 379
rect 380 379 396 413
rect 430 379 446 413
rect 380 373 446 379
rect 36 339 446 373
rect 484 539 550 547
rect 484 505 500 539
rect 534 505 550 539
rect 484 424 550 505
rect 584 508 636 563
rect 584 474 586 508
rect 620 474 636 508
rect 584 458 636 474
rect 683 599 755 615
rect 683 565 699 599
rect 733 565 755 599
rect 683 509 755 565
rect 683 475 699 509
rect 733 475 755 509
rect 683 424 755 475
rect 484 419 755 424
rect 789 607 855 649
rect 789 573 805 607
rect 839 573 855 607
rect 789 530 855 573
rect 789 496 805 530
rect 839 496 855 530
rect 789 453 855 496
rect 789 419 805 453
rect 839 419 855 453
rect 889 599 941 615
rect 889 565 891 599
rect 925 565 941 599
rect 889 507 941 565
rect 889 473 891 507
rect 925 473 941 507
rect 484 413 699 419
rect 484 379 500 413
rect 534 385 699 413
rect 733 385 755 419
rect 889 413 941 473
rect 889 385 891 413
rect 534 379 571 385
rect 484 363 571 379
rect 31 271 91 305
rect 125 271 177 305
rect 211 271 257 305
rect 31 242 257 271
rect 291 271 307 305
rect 341 271 405 305
rect 439 271 455 305
rect 291 242 455 271
rect 537 249 571 363
rect 719 379 891 385
rect 925 379 941 413
rect 719 351 941 379
rect 607 319 683 351
rect 607 285 633 319
rect 667 285 683 319
rect 729 283 745 317
rect 779 305 943 317
rect 779 283 868 305
rect 852 271 868 283
rect 902 271 943 305
rect 537 225 816 249
rect 852 242 943 271
rect 537 215 766 225
rect 50 174 66 208
rect 100 174 238 208
rect 272 181 503 208
rect 750 191 766 215
rect 800 191 816 225
rect 272 174 494 181
rect 50 113 102 174
rect 50 79 66 113
rect 100 79 102 113
rect 50 63 102 79
rect 136 132 202 140
rect 136 98 152 132
rect 186 98 202 132
rect 136 17 202 98
rect 236 113 282 174
rect 469 147 494 174
rect 528 147 666 181
rect 700 147 716 181
rect 236 79 238 113
rect 272 79 282 113
rect 236 63 282 79
rect 316 124 435 140
rect 316 90 324 124
rect 358 90 401 124
rect 316 17 435 90
rect 469 107 530 147
rect 469 73 494 107
rect 528 73 530 107
rect 469 57 530 73
rect 564 107 630 113
rect 564 73 580 107
rect 614 73 630 107
rect 564 17 630 73
rect 664 107 716 147
rect 750 153 816 191
rect 750 119 766 153
rect 800 119 816 153
rect 850 192 902 208
rect 850 158 852 192
rect 886 158 902 192
rect 664 73 666 107
rect 700 85 716 107
rect 850 111 902 158
rect 850 85 852 111
rect 700 77 852 85
rect 886 77 902 111
rect 700 73 902 77
rect 664 51 902 73
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o31ai_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 353152
string GDS_START 344134
<< end >>
