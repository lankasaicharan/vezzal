magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 16 49 633 195
rect 0 0 768 49
<< scpmos >>
rect 82 392 282 592
rect 337 392 537 592
<< nmoslvt >>
rect 95 85 295 169
rect 350 85 550 169
<< ndiff >>
rect 42 145 95 169
rect 42 111 50 145
rect 84 111 95 145
rect 42 85 95 111
rect 295 145 350 169
rect 295 111 306 145
rect 340 111 350 145
rect 295 85 350 111
rect 550 145 607 169
rect 550 111 561 145
rect 595 111 607 145
rect 550 85 607 111
<< pdiff >>
rect 27 580 82 592
rect 27 546 35 580
rect 69 546 82 580
rect 27 509 82 546
rect 27 475 35 509
rect 69 475 82 509
rect 27 438 82 475
rect 27 404 35 438
rect 69 404 82 438
rect 27 392 82 404
rect 282 580 337 592
rect 282 546 293 580
rect 327 546 337 580
rect 282 509 337 546
rect 282 475 293 509
rect 327 475 337 509
rect 282 438 337 475
rect 282 404 293 438
rect 327 404 337 438
rect 282 392 337 404
rect 537 580 594 592
rect 537 546 548 580
rect 582 546 594 580
rect 537 509 594 546
rect 537 475 548 509
rect 582 475 594 509
rect 537 438 594 475
rect 537 404 548 438
rect 582 404 594 438
rect 537 392 594 404
<< ndiffc >>
rect 50 111 84 145
rect 306 111 340 145
rect 561 111 595 145
<< pdiffc >>
rect 35 546 69 580
rect 35 475 69 509
rect 35 404 69 438
rect 293 546 327 580
rect 293 475 327 509
rect 293 404 327 438
rect 548 546 582 580
rect 548 475 582 509
rect 548 404 582 438
<< poly >>
rect 82 592 282 618
rect 337 592 537 618
rect 82 366 282 392
rect 337 366 537 392
rect 82 301 148 366
rect 82 267 98 301
rect 132 267 148 301
rect 82 251 148 267
rect 229 300 416 316
rect 229 266 245 300
rect 279 266 366 300
rect 400 266 416 300
rect 229 238 416 266
rect 471 301 537 366
rect 471 267 487 301
rect 521 267 537 301
rect 471 251 537 267
rect 229 209 295 238
rect 95 169 295 209
rect 350 209 416 238
rect 350 169 550 209
rect 95 47 295 85
rect 350 47 550 85
<< polycont >>
rect 98 267 132 301
rect 245 266 279 300
rect 366 266 400 300
rect 487 267 521 301
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 19 580 85 649
rect 19 546 35 580
rect 69 546 85 580
rect 19 509 85 546
rect 19 475 35 509
rect 69 475 85 509
rect 19 438 85 475
rect 19 404 35 438
rect 69 404 85 438
rect 19 386 85 404
rect 229 580 416 649
rect 229 546 293 580
rect 327 546 416 580
rect 229 509 416 546
rect 229 475 293 509
rect 327 475 416 509
rect 229 438 416 475
rect 229 404 293 438
rect 327 404 416 438
rect 34 301 148 317
rect 34 267 98 301
rect 132 267 148 301
rect 34 145 148 267
rect 229 300 416 404
rect 532 580 598 649
rect 532 546 548 580
rect 582 546 598 580
rect 532 509 598 546
rect 532 475 548 509
rect 582 475 598 509
rect 532 438 598 475
rect 532 404 548 438
rect 582 404 598 438
rect 532 388 598 404
rect 229 266 245 300
rect 279 266 366 300
rect 400 266 416 300
rect 229 250 416 266
rect 471 301 611 316
rect 471 267 487 301
rect 521 267 611 301
rect 34 111 50 145
rect 84 111 148 145
rect 34 17 148 111
rect 290 145 356 161
rect 290 111 306 145
rect 340 111 356 145
rect 290 17 356 111
rect 471 145 611 267
rect 471 111 561 145
rect 595 111 611 145
rect 471 17 611 111
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 decap_8
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 3141892
string GDS_START 3137942
<< end >>
