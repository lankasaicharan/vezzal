magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 4242 1852
<< nwell >>
rect -38 261 2982 582
<< pwell >>
rect 1538 157 1919 201
rect 2408 157 2907 203
rect 1 21 2907 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 169 47 199 131
rect 265 47 295 131
rect 349 47 379 131
rect 557 47 587 131
rect 761 47 791 131
rect 849 47 879 131
rect 1053 47 1083 131
rect 1147 47 1177 131
rect 1219 47 1249 131
rect 1437 47 1467 131
rect 1509 47 1539 131
rect 1625 47 1655 175
rect 1803 47 1833 175
rect 1947 47 1977 131
rect 2019 47 2049 131
rect 2177 47 2207 131
rect 2298 47 2328 131
rect 2486 47 2516 177
rect 2694 47 2724 131
rect 2799 47 2829 177
<< scpmoshvt >>
rect 81 369 117 497
rect 175 369 211 497
rect 257 369 293 497
rect 351 369 387 497
rect 549 369 585 497
rect 747 369 783 497
rect 841 369 877 497
rect 1039 413 1075 497
rect 1133 413 1169 497
rect 1245 413 1281 497
rect 1373 413 1409 497
rect 1490 413 1526 497
rect 1616 329 1652 497
rect 1699 329 1735 497
rect 1834 413 1870 497
rect 1932 413 1968 497
rect 2081 413 2117 497
rect 2289 413 2325 497
rect 2488 297 2524 497
rect 2686 355 2722 483
rect 2791 297 2827 497
<< ndiff >>
rect 1564 131 1625 175
rect 27 103 79 131
rect 27 69 35 103
rect 69 69 79 103
rect 27 47 79 69
rect 109 47 169 131
rect 199 98 265 131
rect 199 64 221 98
rect 255 64 265 98
rect 199 47 265 64
rect 295 47 349 131
rect 379 93 447 131
rect 379 59 405 93
rect 439 59 447 93
rect 379 47 447 59
rect 501 105 557 131
rect 501 71 509 105
rect 543 71 557 105
rect 501 47 557 71
rect 587 93 645 131
rect 587 59 603 93
rect 637 59 645 93
rect 587 47 645 59
rect 699 105 761 131
rect 699 71 707 105
rect 741 71 761 105
rect 699 47 761 71
rect 791 89 849 131
rect 791 55 801 89
rect 835 55 849 89
rect 791 47 849 55
rect 879 101 937 131
rect 879 67 895 101
rect 929 67 937 101
rect 879 47 937 67
rect 991 101 1053 131
rect 991 67 999 101
rect 1033 67 1053 101
rect 991 47 1053 67
rect 1083 101 1147 131
rect 1083 67 1093 101
rect 1127 67 1147 101
rect 1083 47 1147 67
rect 1177 47 1219 131
rect 1249 93 1311 131
rect 1249 59 1269 93
rect 1303 59 1311 93
rect 1249 47 1311 59
rect 1365 119 1437 131
rect 1365 85 1373 119
rect 1407 85 1437 119
rect 1365 47 1437 85
rect 1467 47 1509 131
rect 1539 89 1625 131
rect 1539 55 1559 89
rect 1593 55 1625 89
rect 1539 47 1625 55
rect 1655 47 1803 175
rect 1833 131 1893 175
rect 2434 161 2486 177
rect 1833 89 1947 131
rect 1833 55 1858 89
rect 1892 55 1947 89
rect 1833 47 1947 55
rect 1977 47 2019 131
rect 2049 47 2177 131
rect 2207 89 2298 131
rect 2207 55 2244 89
rect 2278 55 2298 89
rect 2207 47 2298 55
rect 2328 101 2380 131
rect 2328 67 2338 101
rect 2372 67 2380 101
rect 2328 47 2380 67
rect 2434 127 2442 161
rect 2476 127 2486 161
rect 2434 93 2486 127
rect 2434 59 2442 93
rect 2476 59 2486 93
rect 2434 47 2486 59
rect 2516 161 2578 177
rect 2516 127 2536 161
rect 2570 127 2578 161
rect 2739 131 2799 177
rect 2516 93 2578 127
rect 2516 59 2536 93
rect 2570 59 2578 93
rect 2516 47 2578 59
rect 2632 105 2694 131
rect 2632 71 2640 105
rect 2674 71 2694 105
rect 2632 47 2694 71
rect 2724 103 2799 131
rect 2724 69 2745 103
rect 2779 69 2799 103
rect 2724 47 2799 69
rect 2829 165 2881 177
rect 2829 131 2839 165
rect 2873 131 2881 165
rect 2829 97 2881 131
rect 2829 63 2839 97
rect 2873 63 2881 97
rect 2829 47 2881 63
<< pdiff >>
rect 27 431 81 497
rect 27 397 35 431
rect 69 397 81 431
rect 27 369 81 397
rect 117 489 175 497
rect 117 455 129 489
rect 163 455 175 489
rect 117 369 175 455
rect 211 369 257 497
rect 293 411 351 497
rect 293 377 305 411
rect 339 377 351 411
rect 293 369 351 377
rect 387 485 441 497
rect 387 451 399 485
rect 433 451 441 485
rect 387 369 441 451
rect 495 415 549 497
rect 495 381 503 415
rect 537 381 549 415
rect 495 369 549 381
rect 585 485 639 497
rect 585 451 597 485
rect 631 451 639 485
rect 585 369 639 451
rect 693 449 747 497
rect 693 415 701 449
rect 735 415 747 449
rect 693 369 747 415
rect 783 489 841 497
rect 783 455 795 489
rect 829 455 841 489
rect 783 369 841 455
rect 877 477 931 497
rect 877 443 889 477
rect 923 443 931 477
rect 877 369 931 443
rect 985 477 1039 497
rect 985 443 993 477
rect 1027 443 1039 477
rect 985 413 1039 443
rect 1075 477 1133 497
rect 1075 443 1087 477
rect 1121 443 1133 477
rect 1075 413 1133 443
rect 1169 413 1245 497
rect 1281 489 1373 497
rect 1281 455 1305 489
rect 1339 455 1373 489
rect 1281 413 1373 455
rect 1409 474 1490 497
rect 1409 440 1425 474
rect 1459 440 1490 474
rect 1409 413 1490 440
rect 1526 489 1616 497
rect 1526 455 1547 489
rect 1581 455 1616 489
rect 1526 413 1616 455
rect 1564 329 1616 413
rect 1652 329 1699 497
rect 1735 475 1834 497
rect 1735 441 1776 475
rect 1810 441 1834 475
rect 1735 413 1834 441
rect 1870 413 1932 497
rect 1968 489 2081 497
rect 1968 455 2025 489
rect 2059 455 2081 489
rect 1968 413 2081 455
rect 2117 474 2171 497
rect 2117 440 2129 474
rect 2163 440 2171 474
rect 2117 413 2171 440
rect 2235 485 2289 497
rect 2235 451 2243 485
rect 2277 451 2289 485
rect 2235 413 2289 451
rect 2325 474 2379 497
rect 2325 440 2337 474
rect 2371 440 2379 474
rect 2325 413 2379 440
rect 2434 485 2488 497
rect 2434 451 2442 485
rect 2476 451 2488 485
rect 2434 417 2488 451
rect 1735 329 1787 413
rect 2434 383 2442 417
rect 2476 383 2488 417
rect 2434 349 2488 383
rect 2434 315 2442 349
rect 2476 315 2488 349
rect 2434 297 2488 315
rect 2524 484 2578 497
rect 2524 450 2536 484
rect 2570 450 2578 484
rect 2739 483 2791 497
rect 2524 416 2578 450
rect 2524 382 2536 416
rect 2570 382 2578 416
rect 2524 348 2578 382
rect 2632 471 2686 483
rect 2632 437 2640 471
rect 2674 437 2686 471
rect 2632 403 2686 437
rect 2632 369 2640 403
rect 2674 369 2686 403
rect 2632 355 2686 369
rect 2722 465 2791 483
rect 2722 431 2745 465
rect 2779 431 2791 465
rect 2722 397 2791 431
rect 2722 363 2745 397
rect 2779 363 2791 397
rect 2722 355 2791 363
rect 2524 314 2536 348
rect 2570 314 2578 348
rect 2524 297 2578 314
rect 2739 297 2791 355
rect 2827 485 2881 497
rect 2827 451 2839 485
rect 2873 451 2881 485
rect 2827 417 2881 451
rect 2827 383 2839 417
rect 2873 383 2881 417
rect 2827 349 2881 383
rect 2827 315 2839 349
rect 2873 315 2881 349
rect 2827 297 2881 315
<< ndiffc >>
rect 35 69 69 103
rect 221 64 255 98
rect 405 59 439 93
rect 509 71 543 105
rect 603 59 637 93
rect 707 71 741 105
rect 801 55 835 89
rect 895 67 929 101
rect 999 67 1033 101
rect 1093 67 1127 101
rect 1269 59 1303 93
rect 1373 85 1407 119
rect 1559 55 1593 89
rect 1858 55 1892 89
rect 2244 55 2278 89
rect 2338 67 2372 101
rect 2442 127 2476 161
rect 2442 59 2476 93
rect 2536 127 2570 161
rect 2536 59 2570 93
rect 2640 71 2674 105
rect 2745 69 2779 103
rect 2839 131 2873 165
rect 2839 63 2873 97
<< pdiffc >>
rect 35 397 69 431
rect 129 455 163 489
rect 305 377 339 411
rect 399 451 433 485
rect 503 381 537 415
rect 597 451 631 485
rect 701 415 735 449
rect 795 455 829 489
rect 889 443 923 477
rect 993 443 1027 477
rect 1087 443 1121 477
rect 1305 455 1339 489
rect 1425 440 1459 474
rect 1547 455 1581 489
rect 1776 441 1810 475
rect 2025 455 2059 489
rect 2129 440 2163 474
rect 2243 451 2277 485
rect 2337 440 2371 474
rect 2442 451 2476 485
rect 2442 383 2476 417
rect 2442 315 2476 349
rect 2536 450 2570 484
rect 2536 382 2570 416
rect 2640 437 2674 471
rect 2640 369 2674 403
rect 2745 431 2779 465
rect 2745 363 2779 397
rect 2536 314 2570 348
rect 2839 451 2873 485
rect 2839 383 2873 417
rect 2839 315 2873 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 257 497 293 523
rect 351 497 387 523
rect 549 497 585 523
rect 747 497 783 523
rect 841 497 877 523
rect 1039 497 1075 523
rect 1133 497 1169 523
rect 1245 497 1281 523
rect 1373 497 1409 523
rect 1490 497 1526 523
rect 1616 497 1652 523
rect 1699 497 1735 523
rect 1834 497 1870 523
rect 1932 497 1968 523
rect 2081 497 2117 523
rect 2289 497 2325 523
rect 2488 497 2524 523
rect 1039 398 1075 413
rect 1133 398 1169 413
rect 1245 398 1281 413
rect 1373 398 1409 413
rect 1490 398 1526 413
rect 81 354 117 369
rect 175 354 211 369
rect 257 354 293 369
rect 351 354 387 369
rect 549 354 585 369
rect 747 354 783 369
rect 841 354 877 369
rect 978 368 1077 398
rect 1131 381 1171 398
rect 1243 381 1283 398
rect 49 324 119 354
rect 49 265 79 324
rect 173 282 213 354
rect 22 249 79 265
rect 22 215 35 249
rect 69 215 79 249
rect 128 266 213 282
rect 128 232 138 266
rect 172 253 213 266
rect 172 232 199 253
rect 128 216 199 232
rect 255 219 295 354
rect 22 199 79 215
rect 49 176 79 199
rect 49 146 109 176
rect 79 131 109 146
rect 169 131 199 216
rect 241 203 295 219
rect 241 169 251 203
rect 285 169 295 203
rect 241 153 295 169
rect 265 131 295 153
rect 349 265 389 354
rect 547 265 587 354
rect 733 324 785 354
rect 733 284 763 324
rect 839 284 879 354
rect 978 284 1008 368
rect 1119 365 1183 381
rect 1119 331 1129 365
rect 1163 331 1183 365
rect 1119 315 1183 331
rect 1243 365 1329 381
rect 1243 331 1285 365
rect 1319 331 1329 365
rect 1243 315 1329 331
rect 349 249 469 265
rect 349 215 413 249
rect 447 215 469 249
rect 349 199 469 215
rect 520 249 587 265
rect 520 215 530 249
rect 564 215 587 249
rect 709 268 763 284
rect 709 234 719 268
rect 753 234 763 268
rect 709 218 763 234
rect 815 268 879 284
rect 815 234 825 268
rect 859 234 879 268
rect 815 218 879 234
rect 924 268 1008 284
rect 924 234 934 268
rect 968 248 1008 268
rect 968 234 1177 248
rect 924 218 1177 234
rect 520 199 587 215
rect 349 131 379 199
rect 557 131 587 199
rect 733 176 763 218
rect 849 176 879 218
rect 733 146 791 176
rect 761 131 791 146
rect 849 146 1083 176
rect 849 131 879 146
rect 1053 131 1083 146
rect 1147 131 1177 218
rect 1243 213 1283 315
rect 1371 273 1411 398
rect 1488 369 1528 398
rect 1453 353 1528 369
rect 1453 319 1473 353
rect 1507 319 1528 353
rect 1834 398 1870 413
rect 1932 398 1968 413
rect 2081 398 2117 413
rect 2289 398 2325 413
rect 1832 381 1872 398
rect 1824 365 1888 381
rect 1824 345 1844 365
rect 1803 331 1844 345
rect 1878 331 1888 365
rect 1453 303 1528 319
rect 1616 314 1652 329
rect 1699 314 1735 329
rect 1803 315 1888 331
rect 1930 325 1970 398
rect 2079 397 2119 398
rect 2079 367 2207 397
rect 2287 375 2327 398
rect 2143 339 2207 367
rect 1337 263 1411 273
rect 1337 229 1353 263
rect 1387 229 1411 263
rect 1488 273 1528 303
rect 1488 232 1539 273
rect 1614 265 1654 314
rect 1697 265 1737 314
rect 1337 219 1411 229
rect 1219 203 1295 213
rect 1219 169 1235 203
rect 1269 169 1295 203
rect 1219 159 1295 169
rect 1373 176 1411 219
rect 1219 131 1249 159
rect 1373 146 1467 176
rect 1437 131 1467 146
rect 1509 131 1539 232
rect 1591 249 1655 265
rect 1591 215 1601 249
rect 1635 215 1655 249
rect 1591 199 1655 215
rect 1697 249 1761 265
rect 1697 215 1707 249
rect 1741 215 1761 249
rect 1697 199 1761 215
rect 1625 175 1655 199
rect 1803 175 1833 315
rect 1930 295 2059 325
rect 1912 233 1977 249
rect 1912 199 1923 233
rect 1957 199 1977 233
rect 1912 183 1977 199
rect 1947 131 1977 183
rect 2019 237 2059 295
rect 2143 305 2153 339
rect 2187 305 2207 339
rect 2143 289 2207 305
rect 2019 221 2083 237
rect 2019 187 2029 221
rect 2063 187 2083 221
rect 2019 171 2083 187
rect 2019 131 2049 171
rect 2177 131 2207 289
rect 2249 355 2327 375
rect 2249 321 2259 355
rect 2293 321 2327 355
rect 2249 265 2327 321
rect 2686 483 2722 523
rect 2791 497 2827 523
rect 2686 340 2722 355
rect 2488 282 2524 297
rect 2486 265 2526 282
rect 2684 265 2724 340
rect 2791 282 2827 297
rect 2789 265 2829 282
rect 2249 203 2724 265
rect 2249 169 2259 203
rect 2293 199 2724 203
rect 2766 249 2829 265
rect 2766 215 2776 249
rect 2810 215 2829 249
rect 2766 199 2829 215
rect 2293 169 2328 199
rect 2486 177 2516 199
rect 2249 153 2328 169
rect 2298 131 2328 153
rect 2694 131 2724 199
rect 2799 177 2829 199
rect 79 21 109 47
rect 169 21 199 47
rect 265 21 295 47
rect 349 21 379 47
rect 557 21 587 47
rect 761 21 791 47
rect 849 21 879 47
rect 1053 21 1083 47
rect 1147 21 1177 47
rect 1219 21 1249 47
rect 1437 21 1467 47
rect 1509 21 1539 47
rect 1625 21 1655 47
rect 1803 21 1833 47
rect 1947 21 1977 47
rect 2019 21 2049 47
rect 2177 21 2207 47
rect 2298 21 2328 47
rect 2486 21 2516 47
rect 2694 21 2724 47
rect 2799 21 2829 47
<< polycont >>
rect 35 215 69 249
rect 138 232 172 266
rect 251 169 285 203
rect 1129 331 1163 365
rect 1285 331 1319 365
rect 413 215 447 249
rect 530 215 564 249
rect 719 234 753 268
rect 825 234 859 268
rect 934 234 968 268
rect 1473 319 1507 353
rect 1844 331 1878 365
rect 1353 229 1387 263
rect 1235 169 1269 203
rect 1601 215 1635 249
rect 1707 215 1741 249
rect 1923 199 1957 233
rect 2153 305 2187 339
rect 2029 187 2063 221
rect 2259 321 2293 355
rect 2259 169 2293 203
rect 2776 215 2810 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2944 561
rect 17 431 69 493
rect 103 489 163 527
rect 103 455 129 489
rect 103 439 163 455
rect 207 485 449 493
rect 207 451 399 485
rect 433 451 449 485
rect 17 397 35 431
rect 207 405 241 451
rect 494 417 537 493
rect 588 485 656 527
rect 588 451 597 485
rect 631 451 656 485
rect 769 489 845 527
rect 588 428 656 451
rect 701 449 735 465
rect 769 455 795 489
rect 829 455 845 489
rect 889 477 958 493
rect 413 415 537 417
rect 69 397 241 405
rect 17 369 241 397
rect 279 411 369 415
rect 279 377 305 411
rect 339 377 369 411
rect 279 374 369 377
rect 17 249 73 335
rect 17 215 35 249
rect 69 215 73 249
rect 17 153 73 215
rect 110 266 172 335
rect 110 255 138 266
rect 110 221 126 255
rect 160 221 172 232
rect 110 153 172 221
rect 206 203 285 335
rect 206 169 251 203
rect 206 153 285 169
rect 331 323 369 374
rect 331 289 335 323
rect 17 103 86 119
rect 331 112 369 289
rect 413 381 503 415
rect 923 443 958 477
rect 889 427 958 443
rect 413 354 537 381
rect 413 249 480 354
rect 571 344 667 394
rect 701 391 735 415
rect 701 357 825 391
rect 701 355 859 357
rect 631 318 667 344
rect 447 215 480 249
rect 514 255 590 310
rect 514 221 529 255
rect 563 249 590 255
rect 514 215 530 221
rect 564 215 590 249
rect 631 268 763 318
rect 631 234 719 268
rect 753 234 763 268
rect 413 181 480 215
rect 631 211 763 234
rect 807 268 859 355
rect 807 234 825 268
rect 413 143 543 181
rect 807 177 859 234
rect 17 69 35 103
rect 69 69 86 103
rect 17 17 86 69
rect 195 98 369 112
rect 195 64 221 98
rect 255 64 369 98
rect 195 56 369 64
rect 405 93 441 109
rect 439 59 441 93
rect 405 17 441 59
rect 492 105 543 143
rect 704 143 859 177
rect 903 284 958 427
rect 992 477 1036 493
rect 992 443 993 477
rect 1027 443 1036 477
rect 992 323 1036 443
rect 1086 477 1241 493
rect 1086 443 1087 477
rect 1121 443 1241 477
rect 1289 489 1355 527
rect 1289 455 1305 489
rect 1339 455 1355 489
rect 1420 474 1473 490
rect 1086 427 1241 443
rect 992 318 1002 323
rect 1155 365 1173 391
rect 1121 331 1129 357
rect 1163 331 1173 365
rect 1121 315 1173 331
rect 903 268 968 284
rect 903 255 934 268
rect 903 221 917 255
rect 951 221 968 234
rect 903 218 968 221
rect 492 71 509 105
rect 492 51 543 71
rect 588 93 656 111
rect 588 59 603 93
rect 637 59 656 93
rect 588 17 656 59
rect 704 105 741 143
rect 903 117 937 218
rect 1002 184 1036 289
rect 1207 279 1241 427
rect 1420 440 1425 474
rect 1459 440 1473 474
rect 1420 421 1473 440
rect 1531 489 1742 527
rect 1531 455 1547 489
rect 1581 455 1742 489
rect 1531 425 1742 455
rect 1776 475 1947 492
rect 1810 441 1947 475
rect 2009 489 2085 527
rect 2009 455 2025 489
rect 2059 455 2085 489
rect 2009 447 2085 455
rect 2129 474 2172 490
rect 1776 425 1947 441
rect 1285 387 1473 421
rect 1913 413 1947 425
rect 2163 440 2172 474
rect 2227 485 2293 527
rect 2227 451 2243 485
rect 2277 451 2293 485
rect 2227 447 2293 451
rect 2337 474 2389 493
rect 2129 413 2172 440
rect 2371 440 2389 474
rect 1285 365 1319 387
rect 1582 357 1641 391
rect 1675 357 1751 391
rect 1285 315 1319 331
rect 1438 319 1473 353
rect 1507 323 1545 353
rect 1438 289 1489 319
rect 1523 289 1545 323
rect 1582 299 1751 357
rect 1097 263 1387 279
rect 1097 255 1353 263
rect 704 71 707 105
rect 704 51 741 71
rect 786 89 848 109
rect 786 55 801 89
rect 835 55 848 89
rect 786 17 848 55
rect 892 101 937 117
rect 892 67 895 101
rect 929 67 937 101
rect 892 51 937 67
rect 971 101 1036 184
rect 971 67 999 101
rect 1033 67 1036 101
rect 971 51 1036 67
rect 1080 245 1353 255
rect 1080 101 1178 245
rect 1350 229 1353 245
rect 1590 255 1672 265
rect 1387 249 1672 255
rect 1387 229 1601 249
rect 1350 215 1601 229
rect 1635 215 1672 249
rect 1212 169 1235 203
rect 1269 169 1295 203
rect 1350 195 1672 215
rect 1707 249 1751 299
rect 1741 215 1751 249
rect 1823 365 1879 381
rect 1913 379 2293 413
rect 1823 331 1844 365
rect 1878 331 1879 365
rect 2249 355 2293 379
rect 1823 255 1879 331
rect 1937 339 2215 345
rect 1937 323 2153 339
rect 1937 289 1947 323
rect 1981 305 2153 323
rect 2187 305 2215 339
rect 2249 321 2259 355
rect 2249 305 2293 321
rect 1981 289 1992 305
rect 1937 283 1992 289
rect 2337 271 2389 440
rect 2434 485 2476 527
rect 2434 451 2442 485
rect 2434 417 2476 451
rect 2434 383 2442 417
rect 2434 349 2476 383
rect 2434 315 2442 349
rect 2434 297 2476 315
rect 2510 484 2586 493
rect 2510 450 2536 484
rect 2570 450 2586 484
rect 2510 416 2586 450
rect 2510 382 2536 416
rect 2570 382 2586 416
rect 2510 348 2586 382
rect 2510 314 2536 348
rect 2570 314 2586 348
rect 1823 221 1845 255
rect 1823 215 1879 221
rect 1922 233 1978 249
rect 1212 161 1295 169
rect 1707 179 1751 215
rect 1922 199 1923 233
rect 1957 199 1978 233
rect 1922 179 1978 199
rect 1212 127 1417 161
rect 1707 139 1978 179
rect 2028 237 2389 271
rect 2028 221 2073 237
rect 2028 187 2029 221
rect 2063 187 2073 221
rect 2028 171 2073 187
rect 2121 169 2259 203
rect 2293 169 2309 203
rect 1080 67 1093 101
rect 1127 67 1178 101
rect 1355 119 1417 127
rect 1080 51 1178 67
rect 1212 59 1269 93
rect 1303 59 1319 93
rect 1212 17 1319 59
rect 1355 85 1373 119
rect 1407 85 1417 119
rect 1355 51 1417 85
rect 1508 89 1655 138
rect 2121 89 2155 169
rect 1508 55 1559 89
rect 1593 55 1655 89
rect 1832 55 1858 89
rect 1892 55 2155 89
rect 2244 89 2278 109
rect 2353 108 2389 237
rect 1508 17 1655 55
rect 2244 17 2278 55
rect 2312 101 2389 108
rect 2312 67 2338 101
rect 2372 67 2389 101
rect 2312 51 2389 67
rect 2434 161 2476 177
rect 2434 127 2442 161
rect 2434 93 2476 127
rect 2434 59 2442 93
rect 2434 17 2476 59
rect 2510 161 2586 314
rect 2510 127 2536 161
rect 2570 127 2586 161
rect 2510 93 2586 127
rect 2510 59 2536 93
rect 2570 59 2586 93
rect 2510 51 2586 59
rect 2632 471 2674 493
rect 2632 437 2640 471
rect 2632 403 2674 437
rect 2632 369 2640 403
rect 2632 265 2674 369
rect 2745 465 2779 527
rect 2745 397 2779 431
rect 2745 315 2779 363
rect 2813 485 2925 490
rect 2813 451 2839 485
rect 2873 451 2925 485
rect 2813 417 2925 451
rect 2813 383 2839 417
rect 2873 383 2925 417
rect 2813 349 2925 383
rect 2813 315 2839 349
rect 2873 315 2925 349
rect 2813 299 2925 315
rect 2632 249 2810 265
rect 2632 215 2776 249
rect 2632 199 2810 215
rect 2632 105 2674 199
rect 2854 165 2925 299
rect 2632 71 2640 105
rect 2632 51 2674 71
rect 2738 103 2779 165
rect 2738 69 2745 103
rect 2738 17 2779 69
rect 2813 131 2839 165
rect 2873 131 2925 165
rect 2813 97 2925 131
rect 2813 63 2839 97
rect 2873 63 2925 97
rect 2813 55 2925 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2944 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 126 232 138 255
rect 138 232 160 255
rect 126 221 160 232
rect 335 289 369 323
rect 825 357 859 391
rect 529 249 563 255
rect 529 221 530 249
rect 530 221 563 249
rect 1002 289 1036 323
rect 1121 365 1155 391
rect 1121 357 1129 365
rect 1129 357 1155 365
rect 917 234 934 255
rect 934 234 951 255
rect 917 221 951 234
rect 1641 357 1675 391
rect 1489 319 1507 323
rect 1507 319 1523 323
rect 1489 289 1523 319
rect 1947 289 1981 323
rect 1845 221 1879 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
<< metal1 >>
rect 0 561 2944 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2944 561
rect 0 496 2944 527
rect 813 391 881 397
rect 813 357 825 391
rect 859 388 881 391
rect 1109 391 1177 397
rect 1109 388 1121 391
rect 859 360 1121 388
rect 859 357 881 360
rect 813 351 881 357
rect 1109 357 1121 360
rect 1155 388 1177 391
rect 1629 391 1687 397
rect 1629 388 1641 391
rect 1155 360 1641 388
rect 1155 357 1177 360
rect 1109 351 1177 357
rect 1629 357 1641 360
rect 1675 357 1687 391
rect 1629 351 1687 357
rect 323 323 391 329
rect 323 289 335 323
rect 369 320 391 323
rect 990 323 1048 329
rect 990 320 1002 323
rect 369 292 1002 320
rect 369 289 391 292
rect 323 283 391 289
rect 990 289 1002 292
rect 1036 289 1048 323
rect 990 283 1048 289
rect 1477 323 1545 329
rect 1477 289 1489 323
rect 1523 320 1545 323
rect 1935 323 1993 329
rect 1935 320 1947 323
rect 1523 292 1947 320
rect 1523 289 1545 292
rect 1477 283 1545 289
rect 1935 289 1947 292
rect 1981 289 1993 323
rect 1935 283 1993 289
rect 114 255 172 261
rect 114 221 126 255
rect 160 252 172 255
rect 517 255 575 261
rect 517 252 529 255
rect 160 224 529 252
rect 160 221 172 224
rect 114 215 172 221
rect 517 221 529 224
rect 563 221 575 255
rect 517 215 575 221
rect 905 255 963 261
rect 905 221 917 255
rect 951 252 963 255
rect 1823 255 1891 261
rect 1823 252 1845 255
rect 951 224 1845 252
rect 951 221 963 224
rect 905 215 963 221
rect 1823 221 1845 224
rect 1879 221 1891 255
rect 1823 215 1891 221
rect 0 17 2944 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2944 17
rect 0 -48 2944 -17
<< labels >>
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 SCD
port 3 nsew signal input
flabel locali s 581 357 615 391 0 FreeSans 200 0 0 0 CLK
port 1 nsew signal input
flabel locali s 2513 357 2547 391 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 213 289 247 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 2513 425 2547 459 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 SCD
port 3 nsew signal input
flabel locali s 2513 289 2547 323 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2513 221 2547 255 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2513 153 2547 187 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2513 85 2547 119 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 213 153 247 187 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew signal input
flabel locali s 2881 357 2915 391 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2881 425 2915 459 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2881 221 2915 255 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2881 153 2915 187 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2881 85 2915 119 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2881 289 2915 323 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 1501 289 1535 323 0 FreeSans 200 0 0 0 SET_B
port 5 nsew signal input
flabel metal1 s 121 221 155 255 0 FreeSans 200 0 0 0 SCE
port 4 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel comment s 2441 225 2441 225 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfsbp_1
flabel comment s 1260 297 1260 297 0 FreeSans 200 0 0 0 no_jumper_check
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2944 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2775766
string GDS_START 2753694
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
