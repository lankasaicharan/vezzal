magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 471 167 1055 184
rect 37 49 1055 167
rect 0 0 1056 49
<< scnmos >>
rect 120 57 150 141
rect 198 57 228 141
rect 284 57 314 141
rect 356 57 386 141
rect 554 74 584 158
rect 626 74 656 158
rect 712 74 742 158
rect 784 74 814 158
rect 870 74 900 158
rect 942 74 972 158
<< scpmoshvt >>
rect 100 408 150 608
rect 206 408 256 608
rect 317 408 367 608
rect 606 409 656 609
rect 744 409 794 609
rect 842 409 892 609
<< ndiff >>
rect 63 116 120 141
rect 63 82 75 116
rect 109 82 120 116
rect 63 57 120 82
rect 150 57 198 141
rect 228 107 284 141
rect 228 73 239 107
rect 273 73 284 107
rect 228 57 284 73
rect 314 57 356 141
rect 386 116 443 141
rect 386 82 397 116
rect 431 82 443 116
rect 386 57 443 82
rect 497 133 554 158
rect 497 99 509 133
rect 543 99 554 133
rect 497 74 554 99
rect 584 74 626 158
rect 656 133 712 158
rect 656 99 667 133
rect 701 99 712 133
rect 656 74 712 99
rect 742 74 784 158
rect 814 133 870 158
rect 814 99 825 133
rect 859 99 870 133
rect 814 74 870 99
rect 900 74 942 158
rect 972 133 1029 158
rect 972 99 983 133
rect 1017 99 1029 133
rect 972 74 1029 99
<< pdiff >>
rect 43 596 100 608
rect 43 562 55 596
rect 89 562 100 596
rect 43 525 100 562
rect 43 491 55 525
rect 89 491 100 525
rect 43 454 100 491
rect 43 420 55 454
rect 89 420 100 454
rect 43 408 100 420
rect 150 596 206 608
rect 150 562 161 596
rect 195 562 206 596
rect 150 524 206 562
rect 150 490 161 524
rect 195 490 206 524
rect 150 408 206 490
rect 256 596 317 608
rect 256 562 267 596
rect 301 562 317 596
rect 256 525 317 562
rect 256 491 267 525
rect 301 491 317 525
rect 256 454 317 491
rect 256 420 267 454
rect 301 420 317 454
rect 256 408 317 420
rect 367 454 485 608
rect 367 420 439 454
rect 473 420 485 454
rect 367 408 485 420
rect 549 455 606 609
rect 549 421 561 455
rect 595 421 606 455
rect 549 409 606 421
rect 656 601 744 609
rect 656 567 683 601
rect 717 567 744 601
rect 656 409 744 567
rect 794 409 842 609
rect 892 597 949 609
rect 892 563 903 597
rect 937 563 949 597
rect 892 526 949 563
rect 892 492 903 526
rect 937 492 949 526
rect 892 455 949 492
rect 892 421 903 455
rect 937 421 949 455
rect 892 409 949 421
<< ndiffc >>
rect 75 82 109 116
rect 239 73 273 107
rect 397 82 431 116
rect 509 99 543 133
rect 667 99 701 133
rect 825 99 859 133
rect 983 99 1017 133
<< pdiffc >>
rect 55 562 89 596
rect 55 491 89 525
rect 55 420 89 454
rect 161 562 195 596
rect 161 490 195 524
rect 267 562 301 596
rect 267 491 301 525
rect 267 420 301 454
rect 439 420 473 454
rect 561 421 595 455
rect 683 567 717 601
rect 903 563 937 597
rect 903 492 937 526
rect 903 421 937 455
<< poly >>
rect 100 608 150 634
rect 206 608 256 634
rect 317 608 367 634
rect 606 609 656 635
rect 744 609 794 635
rect 842 609 892 635
rect 100 368 150 408
rect 206 368 256 408
rect 317 368 367 408
rect 84 352 150 368
rect 84 318 100 352
rect 134 318 150 352
rect 84 284 150 318
rect 84 250 100 284
rect 134 250 150 284
rect 84 234 150 250
rect 120 141 150 234
rect 198 352 269 368
rect 198 318 219 352
rect 253 318 269 352
rect 198 284 269 318
rect 198 250 219 284
rect 253 250 269 284
rect 198 234 269 250
rect 317 352 386 368
rect 317 318 336 352
rect 370 318 386 352
rect 317 284 386 318
rect 317 250 336 284
rect 370 250 386 284
rect 317 234 386 250
rect 198 141 228 234
rect 356 186 386 234
rect 434 316 500 332
rect 434 282 450 316
rect 484 282 500 316
rect 434 248 500 282
rect 434 214 450 248
rect 484 228 500 248
rect 606 228 656 409
rect 744 370 794 409
rect 484 214 656 228
rect 434 198 656 214
rect 284 156 386 186
rect 554 158 584 198
rect 626 158 656 198
rect 712 354 794 370
rect 712 320 728 354
rect 762 320 794 354
rect 712 286 794 320
rect 842 356 892 409
rect 842 340 972 356
rect 842 314 922 340
rect 712 252 728 286
rect 762 266 794 286
rect 862 306 922 314
rect 956 306 972 340
rect 862 272 972 306
rect 762 252 814 266
rect 712 236 814 252
rect 712 158 742 236
rect 784 158 814 236
rect 862 238 922 272
rect 956 238 972 272
rect 862 222 972 238
rect 870 158 900 222
rect 942 158 972 222
rect 284 141 314 156
rect 356 141 386 156
rect 120 31 150 57
rect 198 31 228 57
rect 284 31 314 57
rect 356 31 386 57
rect 554 48 584 74
rect 626 48 656 74
rect 712 48 742 74
rect 784 48 814 74
rect 870 48 900 74
rect 942 48 972 74
<< polycont >>
rect 100 318 134 352
rect 100 250 134 284
rect 219 318 253 352
rect 219 250 253 284
rect 336 318 370 352
rect 336 250 370 284
rect 450 282 484 316
rect 450 214 484 248
rect 728 320 762 354
rect 728 252 762 286
rect 922 306 956 340
rect 922 238 956 272
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 39 596 105 612
rect 39 562 55 596
rect 89 562 105 596
rect 39 525 105 562
rect 39 491 55 525
rect 89 491 105 525
rect 39 454 105 491
rect 145 596 211 649
rect 145 562 161 596
rect 195 562 211 596
rect 145 524 211 562
rect 145 490 161 524
rect 195 490 211 524
rect 145 474 211 490
rect 251 596 317 612
rect 251 562 267 596
rect 301 562 317 596
rect 667 601 733 649
rect 667 567 683 601
rect 717 567 733 601
rect 853 597 953 613
rect 251 525 317 562
rect 853 563 903 597
rect 937 563 953 597
rect 853 533 953 563
rect 251 491 267 525
rect 301 491 317 525
rect 39 420 55 454
rect 89 438 105 454
rect 251 454 317 491
rect 251 438 267 454
rect 89 420 267 438
rect 301 420 317 454
rect 39 404 317 420
rect 353 526 953 533
rect 353 499 903 526
rect 353 368 387 499
rect 819 492 903 499
rect 937 492 953 526
rect 25 352 167 368
rect 25 318 100 352
rect 134 318 167 352
rect 25 284 167 318
rect 25 250 100 284
rect 134 250 167 284
rect 25 234 167 250
rect 203 352 269 368
rect 203 318 219 352
rect 253 318 269 352
rect 203 284 269 318
rect 203 250 219 284
rect 253 250 269 284
rect 203 234 269 250
rect 320 352 387 368
rect 320 318 336 352
rect 370 318 387 352
rect 320 284 387 318
rect 320 250 336 284
rect 370 250 387 284
rect 320 234 387 250
rect 423 454 489 465
rect 423 420 439 454
rect 473 420 489 454
rect 423 332 489 420
rect 536 455 611 465
rect 536 421 561 455
rect 595 430 611 455
rect 819 455 953 492
rect 595 421 647 430
rect 536 384 647 421
rect 423 316 500 332
rect 423 282 450 316
rect 484 282 500 316
rect 423 248 500 282
rect 423 214 450 248
rect 484 214 500 248
rect 423 198 500 214
rect 59 164 457 198
rect 59 116 125 164
rect 59 82 75 116
rect 109 82 125 116
rect 59 53 125 82
rect 223 107 289 128
rect 223 73 239 107
rect 273 73 289 107
rect 223 17 289 73
rect 381 116 447 164
rect 536 162 570 384
rect 697 354 778 430
rect 697 320 728 354
rect 762 320 778 354
rect 697 286 778 320
rect 697 252 728 286
rect 762 252 778 286
rect 697 236 778 252
rect 819 421 903 455
rect 937 421 953 455
rect 819 405 953 421
rect 819 162 853 405
rect 889 340 1031 356
rect 889 306 922 340
rect 956 306 1031 340
rect 889 272 1031 306
rect 889 238 922 272
rect 956 238 1031 272
rect 889 222 1031 238
rect 381 82 397 116
rect 431 82 447 116
rect 381 53 447 82
rect 493 133 570 162
rect 493 99 509 133
rect 543 99 570 133
rect 493 70 570 99
rect 651 133 717 162
rect 651 99 667 133
rect 701 99 717 133
rect 651 17 717 99
rect 809 133 875 162
rect 809 99 825 133
rect 859 99 875 133
rect 809 70 875 99
rect 967 133 1033 162
rect 967 99 983 133
rect 1017 99 1033 133
rect 967 17 1033 99
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2bb2o_lp
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5869690
string GDS_START 5860744
<< end >>
