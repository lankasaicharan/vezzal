magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 149 228 1151 248
rect 28 49 1151 228
rect 0 0 1152 49
<< scpmos >>
rect 83 392 119 592
rect 285 368 321 592
rect 375 368 411 592
rect 465 368 501 592
rect 555 368 591 592
rect 757 368 793 592
rect 847 368 883 592
rect 937 368 973 592
rect 1029 368 1065 592
<< nmoslvt >>
rect 111 74 141 202
rect 225 74 255 222
rect 325 74 355 222
rect 463 74 493 222
rect 549 74 579 222
rect 659 74 689 222
rect 763 74 793 222
rect 938 74 968 222
rect 1035 74 1065 222
<< ndiff >>
rect 175 202 225 222
rect 54 190 111 202
rect 54 156 66 190
rect 100 156 111 190
rect 54 120 111 156
rect 54 86 66 120
rect 100 86 111 120
rect 54 74 111 86
rect 141 184 225 202
rect 141 150 166 184
rect 200 150 225 184
rect 141 116 225 150
rect 141 82 166 116
rect 200 82 225 116
rect 141 74 225 82
rect 255 184 325 222
rect 255 150 266 184
rect 300 150 325 184
rect 255 116 325 150
rect 255 82 266 116
rect 300 82 325 116
rect 255 74 325 82
rect 355 120 463 222
rect 355 86 385 120
rect 419 86 463 120
rect 355 74 463 86
rect 493 210 549 222
rect 493 176 504 210
rect 538 176 549 210
rect 493 120 549 176
rect 493 86 504 120
rect 538 86 549 120
rect 493 74 549 86
rect 579 152 659 222
rect 579 118 604 152
rect 638 118 659 152
rect 579 74 659 118
rect 689 210 763 222
rect 689 176 704 210
rect 738 176 763 210
rect 689 120 763 176
rect 689 86 704 120
rect 738 86 763 120
rect 689 74 763 86
rect 793 142 938 222
rect 793 108 804 142
rect 838 108 893 142
rect 927 108 938 142
rect 793 74 938 108
rect 968 210 1035 222
rect 968 176 979 210
rect 1013 176 1035 210
rect 968 120 1035 176
rect 968 86 979 120
rect 1013 86 1035 120
rect 968 74 1035 86
rect 1065 210 1125 222
rect 1065 176 1079 210
rect 1113 176 1125 210
rect 1065 120 1125 176
rect 1065 86 1079 120
rect 1113 86 1125 120
rect 1065 74 1125 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 509 83 546
rect 27 475 39 509
rect 73 475 83 509
rect 27 438 83 475
rect 27 404 39 438
rect 73 404 83 438
rect 27 392 83 404
rect 119 580 175 592
rect 119 546 129 580
rect 163 546 175 580
rect 119 512 175 546
rect 119 478 129 512
rect 163 478 175 512
rect 119 444 175 478
rect 119 410 129 444
rect 163 410 175 444
rect 119 392 175 410
rect 229 580 285 592
rect 229 546 241 580
rect 275 546 285 580
rect 229 497 285 546
rect 229 463 241 497
rect 275 463 285 497
rect 229 414 285 463
rect 229 380 241 414
rect 275 380 285 414
rect 229 368 285 380
rect 321 531 375 592
rect 321 497 331 531
rect 365 497 375 531
rect 321 414 375 497
rect 321 380 331 414
rect 365 380 375 414
rect 321 368 375 380
rect 411 580 465 592
rect 411 546 421 580
rect 455 546 465 580
rect 411 508 465 546
rect 411 474 421 508
rect 455 474 465 508
rect 411 368 465 474
rect 501 578 555 592
rect 501 544 511 578
rect 545 544 555 578
rect 501 368 555 544
rect 591 519 647 592
rect 591 485 601 519
rect 635 485 647 519
rect 591 368 647 485
rect 701 531 757 592
rect 701 497 713 531
rect 747 497 757 531
rect 701 424 757 497
rect 701 390 713 424
rect 747 390 757 424
rect 701 368 757 390
rect 793 580 847 592
rect 793 546 803 580
rect 837 546 847 580
rect 793 508 847 546
rect 793 474 803 508
rect 837 474 847 508
rect 793 368 847 474
rect 883 580 937 592
rect 883 546 893 580
rect 927 546 937 580
rect 883 502 937 546
rect 883 468 893 502
rect 927 468 937 502
rect 883 424 937 468
rect 883 390 893 424
rect 927 390 937 424
rect 883 368 937 390
rect 973 580 1029 592
rect 973 546 983 580
rect 1017 546 1029 580
rect 973 508 1029 546
rect 973 474 983 508
rect 1017 474 1029 508
rect 973 368 1029 474
rect 1065 580 1121 592
rect 1065 546 1075 580
rect 1109 546 1121 580
rect 1065 502 1121 546
rect 1065 468 1075 502
rect 1109 468 1121 502
rect 1065 424 1121 468
rect 1065 390 1075 424
rect 1109 390 1121 424
rect 1065 368 1121 390
<< ndiffc >>
rect 66 156 100 190
rect 66 86 100 120
rect 166 150 200 184
rect 166 82 200 116
rect 266 150 300 184
rect 266 82 300 116
rect 385 86 419 120
rect 504 176 538 210
rect 504 86 538 120
rect 604 118 638 152
rect 704 176 738 210
rect 704 86 738 120
rect 804 108 838 142
rect 893 108 927 142
rect 979 176 1013 210
rect 979 86 1013 120
rect 1079 176 1113 210
rect 1079 86 1113 120
<< pdiffc >>
rect 39 546 73 580
rect 39 475 73 509
rect 39 404 73 438
rect 129 546 163 580
rect 129 478 163 512
rect 129 410 163 444
rect 241 546 275 580
rect 241 463 275 497
rect 241 380 275 414
rect 331 497 365 531
rect 331 380 365 414
rect 421 546 455 580
rect 421 474 455 508
rect 511 544 545 578
rect 601 485 635 519
rect 713 497 747 531
rect 713 390 747 424
rect 803 546 837 580
rect 803 474 837 508
rect 893 546 927 580
rect 893 468 927 502
rect 893 390 927 424
rect 983 546 1017 580
rect 983 474 1017 508
rect 1075 546 1109 580
rect 1075 468 1109 502
rect 1075 390 1109 424
<< poly >>
rect 83 592 119 618
rect 285 592 321 618
rect 375 592 411 618
rect 465 592 501 618
rect 555 592 591 618
rect 757 592 793 618
rect 847 592 883 618
rect 937 592 973 618
rect 1029 592 1065 618
rect 83 360 119 392
rect 83 344 173 360
rect 83 310 123 344
rect 157 310 173 344
rect 285 310 321 368
rect 375 310 411 368
rect 465 336 501 368
rect 555 336 591 368
rect 757 336 793 368
rect 847 336 883 368
rect 937 336 973 368
rect 1029 336 1065 368
rect 83 294 173 310
rect 221 294 411 310
rect 111 202 141 294
rect 221 260 237 294
rect 271 260 305 294
rect 339 260 411 294
rect 221 244 411 260
rect 463 320 591 336
rect 463 286 479 320
rect 513 286 591 320
rect 463 270 591 286
rect 659 320 883 336
rect 659 286 675 320
rect 709 286 743 320
rect 777 306 883 320
rect 931 320 1065 336
rect 777 286 793 306
rect 659 270 793 286
rect 931 286 947 320
rect 981 286 1015 320
rect 1049 286 1065 320
rect 931 270 1065 286
rect 225 222 255 244
rect 325 222 355 244
rect 463 222 493 270
rect 549 222 579 270
rect 659 222 689 270
rect 763 222 793 270
rect 938 222 968 270
rect 1035 222 1065 270
rect 111 48 141 74
rect 225 48 255 74
rect 325 48 355 74
rect 463 48 493 74
rect 549 48 579 74
rect 659 48 689 74
rect 763 48 793 74
rect 938 48 968 74
rect 1035 48 1065 74
<< polycont >>
rect 123 310 157 344
rect 237 260 271 294
rect 305 260 339 294
rect 479 286 513 320
rect 675 286 709 320
rect 743 286 777 320
rect 947 286 981 320
rect 1015 286 1049 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 580 73 596
rect 23 546 39 580
rect 23 509 73 546
rect 23 475 39 509
rect 23 438 73 475
rect 23 404 39 438
rect 23 260 73 404
rect 113 580 179 649
rect 113 546 129 580
rect 163 546 179 580
rect 113 512 179 546
rect 113 478 129 512
rect 163 478 179 512
rect 113 444 179 478
rect 113 410 129 444
rect 163 410 179 444
rect 113 394 179 410
rect 225 581 455 615
rect 225 580 291 581
rect 225 546 241 580
rect 275 546 291 580
rect 405 580 455 581
rect 225 497 291 546
rect 225 463 241 497
rect 275 463 291 497
rect 225 414 291 463
rect 225 380 241 414
rect 275 380 291 414
rect 225 364 291 380
rect 331 531 365 547
rect 331 424 365 497
rect 405 546 421 580
rect 405 508 455 546
rect 495 581 853 615
rect 495 578 561 581
rect 495 544 511 578
rect 545 544 561 578
rect 787 580 853 581
rect 495 526 561 544
rect 405 474 421 508
rect 601 519 651 547
rect 455 485 601 492
rect 635 485 651 519
rect 455 474 651 485
rect 405 458 651 474
rect 697 531 747 547
rect 697 497 713 531
rect 697 424 747 497
rect 787 546 803 580
rect 837 546 853 580
rect 787 508 853 546
rect 787 474 803 508
rect 837 474 853 508
rect 787 458 853 474
rect 893 580 927 596
rect 893 502 927 546
rect 893 424 927 468
rect 967 580 1033 649
rect 967 546 983 580
rect 1017 546 1033 580
rect 967 508 1033 546
rect 967 474 983 508
rect 1017 474 1033 508
rect 967 458 1033 474
rect 1075 580 1125 596
rect 1109 546 1125 580
rect 1075 502 1125 546
rect 1109 468 1125 502
rect 1075 424 1125 468
rect 331 414 619 424
rect 365 390 619 414
rect 697 390 713 424
rect 747 390 893 424
rect 927 390 1075 424
rect 1109 390 1125 424
rect 331 364 365 380
rect 107 344 173 360
rect 107 310 123 344
rect 157 310 173 344
rect 409 320 551 356
rect 107 294 173 310
rect 221 294 355 310
rect 221 260 237 294
rect 271 260 305 294
rect 339 260 355 294
rect 409 286 479 320
rect 513 286 551 320
rect 409 270 551 286
rect 23 226 355 260
rect 585 236 619 390
rect 659 320 839 356
rect 659 286 675 320
rect 709 286 743 320
rect 777 286 839 320
rect 659 270 839 286
rect 889 320 1127 356
rect 889 286 947 320
rect 981 286 1015 320
rect 1049 286 1127 320
rect 889 270 1127 286
rect 23 190 116 226
rect 488 210 1029 236
rect 488 192 504 210
rect 23 156 66 190
rect 100 156 116 190
rect 23 120 116 156
rect 23 86 66 120
rect 100 86 116 120
rect 23 70 116 86
rect 150 184 216 192
rect 150 150 166 184
rect 200 150 216 184
rect 150 116 216 150
rect 150 82 166 116
rect 200 82 216 116
rect 150 17 216 82
rect 250 184 504 192
rect 250 150 266 184
rect 300 176 504 184
rect 538 202 704 210
rect 538 176 554 202
rect 300 158 554 176
rect 688 176 704 202
rect 738 202 979 210
rect 738 176 754 202
rect 300 150 316 158
rect 250 116 316 150
rect 488 120 554 158
rect 250 82 266 116
rect 300 82 316 116
rect 250 66 316 82
rect 350 86 385 120
rect 419 86 454 120
rect 350 17 454 86
rect 488 86 504 120
rect 538 86 554 120
rect 488 70 554 86
rect 588 152 654 168
rect 588 118 604 152
rect 638 118 654 152
rect 588 17 654 118
rect 688 120 754 176
rect 963 176 979 202
rect 1013 176 1029 210
rect 688 86 704 120
rect 738 86 754 120
rect 688 70 754 86
rect 788 142 929 158
rect 788 108 804 142
rect 838 108 893 142
rect 927 108 929 142
rect 788 17 929 108
rect 963 120 1029 176
rect 963 86 979 120
rect 1013 86 1029 120
rect 963 70 1029 86
rect 1063 210 1129 226
rect 1063 176 1079 210
rect 1113 176 1129 210
rect 1063 120 1129 176
rect 1063 86 1079 120
rect 1113 86 1129 120
rect 1063 17 1129 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4b_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 931758
string GDS_START 921826
<< end >>
