magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1778 1975
<< nwell >>
rect -38 331 518 704
<< pwell >>
rect 2 49 448 241
rect 0 0 480 49
<< scnmos >>
rect 81 47 111 215
rect 167 47 197 215
rect 253 47 283 215
rect 339 47 369 215
<< scpmoshvt >>
rect 81 367 111 619
rect 167 367 197 619
rect 253 367 283 619
rect 339 367 369 619
<< ndiff >>
rect 28 192 81 215
rect 28 158 36 192
rect 70 158 81 192
rect 28 93 81 158
rect 28 59 36 93
rect 70 59 81 93
rect 28 47 81 59
rect 111 192 167 215
rect 111 158 122 192
rect 156 158 167 192
rect 111 101 167 158
rect 111 67 122 101
rect 156 67 167 101
rect 111 47 167 67
rect 197 124 253 215
rect 197 90 208 124
rect 242 90 253 124
rect 197 47 253 90
rect 283 192 339 215
rect 283 158 294 192
rect 328 158 339 192
rect 283 101 339 158
rect 283 67 294 101
rect 328 67 339 101
rect 283 47 339 67
rect 369 118 422 215
rect 369 84 380 118
rect 414 84 422 118
rect 369 47 422 84
<< pdiff >>
rect 28 607 81 619
rect 28 573 36 607
rect 70 573 81 607
rect 28 507 81 573
rect 28 473 36 507
rect 70 473 81 507
rect 28 413 81 473
rect 28 379 36 413
rect 70 379 81 413
rect 28 367 81 379
rect 111 599 167 619
rect 111 565 122 599
rect 156 565 167 599
rect 111 509 167 565
rect 111 475 122 509
rect 156 475 167 509
rect 111 413 167 475
rect 111 379 122 413
rect 156 379 167 413
rect 111 367 167 379
rect 197 607 253 619
rect 197 573 208 607
rect 242 573 253 607
rect 197 539 253 573
rect 197 505 208 539
rect 242 505 253 539
rect 197 469 253 505
rect 197 435 208 469
rect 242 435 253 469
rect 197 367 253 435
rect 283 599 339 619
rect 283 565 294 599
rect 328 565 339 599
rect 283 509 339 565
rect 283 475 294 509
rect 328 475 339 509
rect 283 413 339 475
rect 283 379 294 413
rect 328 379 339 413
rect 283 367 339 379
rect 369 607 422 619
rect 369 573 380 607
rect 414 573 422 607
rect 369 539 422 573
rect 369 505 380 539
rect 414 505 422 539
rect 369 469 422 505
rect 369 435 380 469
rect 414 435 422 469
rect 369 367 422 435
<< ndiffc >>
rect 36 158 70 192
rect 36 59 70 93
rect 122 158 156 192
rect 122 67 156 101
rect 208 90 242 124
rect 294 158 328 192
rect 294 67 328 101
rect 380 84 414 118
<< pdiffc >>
rect 36 573 70 607
rect 36 473 70 507
rect 36 379 70 413
rect 122 565 156 599
rect 122 475 156 509
rect 122 379 156 413
rect 208 573 242 607
rect 208 505 242 539
rect 208 435 242 469
rect 294 565 328 599
rect 294 475 328 509
rect 294 379 328 413
rect 380 573 414 607
rect 380 505 414 539
rect 380 435 414 469
<< poly >>
rect 81 619 111 645
rect 167 619 197 645
rect 253 619 283 645
rect 339 619 369 645
rect 81 303 111 367
rect 167 303 197 367
rect 253 303 283 367
rect 339 303 369 367
rect 31 287 369 303
rect 31 253 47 287
rect 81 253 115 287
rect 149 253 183 287
rect 217 253 251 287
rect 285 253 319 287
rect 353 253 369 287
rect 31 237 369 253
rect 81 215 111 237
rect 167 215 197 237
rect 253 215 283 237
rect 339 215 369 237
rect 81 21 111 47
rect 167 21 197 47
rect 253 21 283 47
rect 339 21 369 47
<< polycont >>
rect 47 253 81 287
rect 115 253 149 287
rect 183 253 217 287
rect 251 253 285 287
rect 319 253 353 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 20 607 78 649
rect 20 573 36 607
rect 70 573 78 607
rect 20 507 78 573
rect 20 473 36 507
rect 70 473 78 507
rect 20 413 78 473
rect 20 379 36 413
rect 70 379 78 413
rect 20 363 78 379
rect 112 599 165 615
rect 112 565 122 599
rect 156 565 165 599
rect 112 509 165 565
rect 112 475 122 509
rect 156 475 165 509
rect 112 413 165 475
rect 199 607 250 649
rect 199 573 208 607
rect 242 573 250 607
rect 199 539 250 573
rect 199 505 208 539
rect 242 505 250 539
rect 199 469 250 505
rect 199 435 208 469
rect 242 435 250 469
rect 199 419 250 435
rect 284 599 337 615
rect 284 565 294 599
rect 328 565 337 599
rect 284 509 337 565
rect 284 475 294 509
rect 328 475 337 509
rect 112 379 122 413
rect 156 385 165 413
rect 284 413 337 475
rect 371 607 430 649
rect 371 573 380 607
rect 414 573 430 607
rect 371 539 430 573
rect 371 505 380 539
rect 414 505 430 539
rect 371 469 430 505
rect 371 435 380 469
rect 414 435 430 469
rect 371 419 430 435
rect 284 385 294 413
rect 156 379 294 385
rect 328 385 337 413
rect 328 379 460 385
rect 112 351 460 379
rect 20 287 369 303
rect 20 253 47 287
rect 81 253 115 287
rect 149 253 183 287
rect 217 253 251 287
rect 285 253 319 287
rect 353 253 369 287
rect 20 242 369 253
rect 405 208 460 351
rect 20 192 79 208
rect 20 158 36 192
rect 70 158 79 192
rect 20 93 79 158
rect 20 59 36 93
rect 70 59 79 93
rect 20 17 79 59
rect 113 192 460 208
rect 113 158 122 192
rect 156 174 294 192
rect 156 158 165 174
rect 113 101 165 158
rect 285 158 294 174
rect 328 168 460 192
rect 328 158 337 168
rect 113 67 122 101
rect 156 67 165 101
rect 113 51 165 67
rect 199 124 251 140
rect 199 90 208 124
rect 242 90 251 124
rect 199 17 251 90
rect 285 101 337 158
rect 285 67 294 101
rect 328 67 337 101
rect 285 51 337 67
rect 371 118 430 134
rect 371 84 380 118
rect 414 84 430 118
rect 371 17 430 84
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 inv_4
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5442026
string GDS_START 5436540
<< end >>
