magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 24 49 861 251
rect 0 0 864 49
<< scnmos >>
rect 107 141 137 225
rect 185 141 215 225
rect 299 141 329 225
rect 413 141 443 225
rect 527 141 557 225
rect 652 141 682 225
rect 730 141 760 225
<< scpmoshvt >>
rect 87 419 137 619
rect 193 419 243 619
rect 299 419 349 619
rect 421 419 471 619
rect 527 419 577 619
rect 730 419 780 619
<< ndiff >>
rect 50 191 107 225
rect 50 157 62 191
rect 96 157 107 191
rect 50 141 107 157
rect 137 141 185 225
rect 215 191 299 225
rect 215 157 254 191
rect 288 157 299 191
rect 215 141 299 157
rect 329 141 413 225
rect 443 141 527 225
rect 557 187 652 225
rect 557 153 585 187
rect 619 153 652 187
rect 557 141 652 153
rect 682 141 730 225
rect 760 200 835 225
rect 760 166 789 200
rect 823 166 835 200
rect 760 141 835 166
<< pdiff >>
rect 30 597 87 619
rect 30 563 42 597
rect 76 563 87 597
rect 30 467 87 563
rect 30 433 42 467
rect 76 433 87 467
rect 30 419 87 433
rect 137 497 193 619
rect 137 463 148 497
rect 182 463 193 497
rect 137 419 193 463
rect 243 567 299 619
rect 243 533 254 567
rect 288 533 299 567
rect 243 419 299 533
rect 349 607 421 619
rect 349 573 360 607
rect 394 573 421 607
rect 349 419 421 573
rect 471 567 527 619
rect 471 533 482 567
rect 516 533 527 567
rect 471 419 527 533
rect 577 607 730 619
rect 577 573 601 607
rect 635 573 730 607
rect 577 536 730 573
rect 577 502 601 536
rect 635 502 730 536
rect 577 465 730 502
rect 577 431 601 465
rect 635 431 730 465
rect 577 419 730 431
rect 780 597 837 619
rect 780 563 791 597
rect 825 563 837 597
rect 780 465 837 563
rect 780 431 791 465
rect 825 431 837 465
rect 780 419 837 431
<< ndiffc >>
rect 62 157 96 191
rect 254 157 288 191
rect 585 153 619 187
rect 789 166 823 200
<< pdiffc >>
rect 42 563 76 597
rect 42 433 76 467
rect 148 463 182 497
rect 254 533 288 567
rect 360 573 394 607
rect 482 533 516 567
rect 601 573 635 607
rect 601 502 635 536
rect 601 431 635 465
rect 791 563 825 597
rect 791 431 825 465
<< poly >>
rect 87 619 137 645
rect 193 619 243 645
rect 299 619 349 645
rect 421 619 471 645
rect 527 619 577 645
rect 730 619 780 645
rect 87 381 137 419
rect 193 381 243 419
rect 299 381 349 419
rect 421 381 471 419
rect 71 365 137 381
rect 71 331 87 365
rect 121 331 137 365
rect 71 297 137 331
rect 71 263 87 297
rect 121 263 137 297
rect 71 247 137 263
rect 107 225 137 247
rect 185 365 251 381
rect 185 331 201 365
rect 235 331 251 365
rect 185 297 251 331
rect 185 263 201 297
rect 235 263 251 297
rect 185 247 251 263
rect 299 365 365 381
rect 299 331 315 365
rect 349 331 365 365
rect 299 297 365 331
rect 299 263 315 297
rect 349 263 365 297
rect 299 247 365 263
rect 413 365 479 381
rect 413 331 429 365
rect 463 331 479 365
rect 413 297 479 331
rect 413 263 429 297
rect 463 263 479 297
rect 413 247 479 263
rect 527 376 577 419
rect 527 360 651 376
rect 527 326 601 360
rect 635 326 651 360
rect 527 310 651 326
rect 185 225 215 247
rect 299 225 329 247
rect 413 225 443 247
rect 527 225 557 310
rect 730 270 780 419
rect 652 225 682 251
rect 730 225 760 270
rect 107 115 137 141
rect 185 115 215 141
rect 299 115 329 141
rect 413 115 443 141
rect 527 115 557 141
rect 652 119 682 141
rect 730 119 760 141
rect 652 103 760 119
rect 652 69 687 103
rect 721 69 760 103
rect 652 53 760 69
<< polycont >>
rect 87 331 121 365
rect 87 263 121 297
rect 201 331 235 365
rect 201 263 235 297
rect 315 331 349 365
rect 315 263 349 297
rect 429 331 463 365
rect 429 263 463 297
rect 601 326 635 360
rect 687 69 721 103
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 26 597 304 613
rect 26 563 42 597
rect 76 579 304 597
rect 76 563 92 579
rect 26 467 92 563
rect 238 567 304 579
rect 26 433 42 467
rect 76 433 92 467
rect 26 417 92 433
rect 132 497 198 543
rect 132 463 148 497
rect 182 463 198 497
rect 238 533 254 567
rect 288 533 304 567
rect 344 607 410 649
rect 344 573 360 607
rect 394 573 410 607
rect 344 557 410 573
rect 466 567 532 613
rect 238 521 304 533
rect 466 533 482 567
rect 516 533 532 567
rect 466 521 532 533
rect 238 487 532 521
rect 585 607 651 649
rect 585 573 601 607
rect 635 573 651 607
rect 585 536 651 573
rect 585 502 601 536
rect 635 502 651 536
rect 132 451 198 463
rect 585 465 651 502
rect 132 417 549 451
rect 25 365 137 381
rect 25 331 87 365
rect 121 331 137 365
rect 25 297 137 331
rect 25 263 87 297
rect 121 263 137 297
rect 25 247 137 263
rect 185 365 263 381
rect 185 331 201 365
rect 235 331 263 365
rect 185 297 263 331
rect 185 263 201 297
rect 235 263 263 297
rect 185 247 263 263
rect 299 365 365 381
rect 299 331 315 365
rect 349 331 365 365
rect 299 297 365 331
rect 299 263 315 297
rect 349 263 365 297
rect 299 247 365 263
rect 409 365 479 381
rect 409 331 429 365
rect 463 331 479 365
rect 409 297 479 331
rect 409 263 429 297
rect 463 263 479 297
rect 46 191 112 211
rect 46 157 62 191
rect 96 157 112 191
rect 46 17 112 157
rect 238 191 304 211
rect 238 157 254 191
rect 288 157 304 191
rect 409 162 479 263
rect 515 274 549 417
rect 585 431 601 465
rect 635 431 651 465
rect 585 415 651 431
rect 773 597 841 613
rect 773 563 791 597
rect 825 563 841 597
rect 773 465 841 563
rect 773 431 791 465
rect 825 431 841 465
rect 585 360 651 376
rect 585 326 601 360
rect 635 326 651 360
rect 585 310 651 326
rect 515 240 737 274
rect 238 126 304 157
rect 515 126 549 240
rect 238 92 549 126
rect 585 187 635 204
rect 619 153 635 187
rect 585 17 635 153
rect 671 103 737 240
rect 671 69 687 103
rect 721 69 737 103
rect 773 200 841 431
rect 773 166 789 200
rect 823 166 841 200
rect 773 88 841 166
rect 671 53 737 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a32o_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2058004
string GDS_START 2050418
<< end >>
