magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2494 1852
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1193 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 196 47 226 177
rect 396 47 426 177
rect 500 47 530 177
rect 709 47 739 177
rect 803 47 833 177
rect 897 47 927 177
rect 991 47 1021 177
rect 1085 47 1115 177
<< scpmoshvt >>
rect 81 297 117 497
rect 186 297 222 497
rect 388 297 424 497
rect 492 297 528 497
rect 701 297 737 497
rect 795 297 831 497
rect 889 297 925 497
rect 983 297 1019 497
rect 1077 297 1113 497
<< ndiff >>
rect 27 109 89 177
rect 27 75 35 109
rect 69 75 89 109
rect 27 47 89 75
rect 119 93 196 177
rect 119 59 129 93
rect 163 59 196 93
rect 119 47 196 59
rect 226 47 396 177
rect 426 93 500 177
rect 426 59 441 93
rect 475 59 500 93
rect 426 47 500 59
rect 530 47 709 177
rect 739 93 803 177
rect 739 59 749 93
rect 783 59 803 93
rect 739 47 803 59
rect 833 101 897 177
rect 833 67 843 101
rect 877 67 897 101
rect 833 47 897 67
rect 927 93 991 177
rect 927 59 937 93
rect 971 59 991 93
rect 927 47 991 59
rect 1021 101 1085 177
rect 1021 67 1031 101
rect 1065 67 1085 101
rect 1021 47 1085 67
rect 1115 93 1167 177
rect 1115 59 1125 93
rect 1159 59 1167 93
rect 1115 47 1167 59
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 297 81 375
rect 117 485 186 497
rect 117 451 129 485
rect 163 451 186 485
rect 117 417 186 451
rect 117 383 129 417
rect 163 383 186 417
rect 117 297 186 383
rect 222 489 280 497
rect 222 455 234 489
rect 268 455 280 489
rect 222 421 280 455
rect 222 387 238 421
rect 272 387 280 421
rect 222 297 280 387
rect 334 421 388 497
rect 334 387 342 421
rect 376 387 388 421
rect 334 297 388 387
rect 424 353 492 497
rect 424 319 442 353
rect 476 319 492 353
rect 424 297 492 319
rect 528 489 590 497
rect 528 455 544 489
rect 578 455 590 489
rect 528 297 590 455
rect 647 477 701 497
rect 647 443 655 477
rect 689 443 701 477
rect 647 297 701 443
rect 737 485 795 497
rect 737 451 749 485
rect 783 451 795 485
rect 737 297 795 451
rect 831 477 889 497
rect 831 443 843 477
rect 877 443 889 477
rect 831 409 889 443
rect 831 375 843 409
rect 877 375 889 409
rect 831 297 889 375
rect 925 485 983 497
rect 925 451 937 485
rect 971 451 983 485
rect 925 417 983 451
rect 925 383 937 417
rect 971 383 983 417
rect 925 297 983 383
rect 1019 477 1077 497
rect 1019 443 1031 477
rect 1065 443 1077 477
rect 1019 409 1077 443
rect 1019 375 1031 409
rect 1065 375 1077 409
rect 1019 297 1077 375
rect 1113 485 1167 497
rect 1113 451 1125 485
rect 1159 451 1167 485
rect 1113 417 1167 451
rect 1113 383 1125 417
rect 1159 383 1167 417
rect 1113 297 1167 383
<< ndiffc >>
rect 35 75 69 109
rect 129 59 163 93
rect 441 59 475 93
rect 749 59 783 93
rect 843 67 877 101
rect 937 59 971 93
rect 1031 67 1065 101
rect 1125 59 1159 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 451 163 485
rect 129 383 163 417
rect 234 455 268 489
rect 238 387 272 421
rect 342 387 376 421
rect 442 319 476 353
rect 544 455 578 489
rect 655 443 689 477
rect 749 451 783 485
rect 843 443 877 477
rect 843 375 877 409
rect 937 451 971 485
rect 937 383 971 417
rect 1031 443 1065 477
rect 1031 375 1065 409
rect 1125 451 1159 485
rect 1125 383 1159 417
<< poly >>
rect 81 497 117 523
rect 186 497 222 523
rect 388 497 424 523
rect 492 497 528 523
rect 701 497 737 523
rect 795 497 831 523
rect 889 497 925 523
rect 983 497 1019 523
rect 1077 497 1113 523
rect 81 282 117 297
rect 186 282 222 297
rect 388 282 424 297
rect 492 282 528 297
rect 701 282 737 297
rect 795 282 831 297
rect 889 282 925 297
rect 983 282 1019 297
rect 1077 282 1113 297
rect 79 265 119 282
rect 184 265 224 282
rect 386 265 426 282
rect 490 265 530 282
rect 699 265 739 282
rect 76 249 140 265
rect 76 215 86 249
rect 120 215 140 249
rect 76 199 140 215
rect 182 249 246 265
rect 182 215 192 249
rect 226 215 246 249
rect 182 199 246 215
rect 315 249 426 265
rect 315 215 325 249
rect 359 215 426 249
rect 315 199 426 215
rect 473 249 537 265
rect 473 215 483 249
rect 517 215 537 249
rect 473 199 537 215
rect 607 249 739 265
rect 793 265 833 282
rect 887 265 927 282
rect 981 265 1021 282
rect 1075 265 1115 282
rect 793 259 1115 265
rect 607 215 617 249
rect 651 215 685 249
rect 719 215 739 249
rect 607 199 739 215
rect 786 249 1115 259
rect 786 215 802 249
rect 836 215 880 249
rect 914 215 958 249
rect 992 215 1036 249
rect 1070 215 1115 249
rect 786 205 1115 215
rect 89 177 119 199
rect 196 177 226 199
rect 396 177 426 199
rect 500 177 530 199
rect 709 177 739 199
rect 803 199 1115 205
rect 803 177 833 199
rect 897 177 927 199
rect 991 177 1021 199
rect 1085 177 1115 199
rect 89 21 119 47
rect 196 21 226 47
rect 396 21 426 47
rect 500 21 530 47
rect 709 21 739 47
rect 803 21 833 47
rect 897 21 927 47
rect 991 21 1021 47
rect 1085 21 1115 47
<< polycont >>
rect 86 215 120 249
rect 192 215 226 249
rect 325 215 359 249
rect 483 215 517 249
rect 617 215 651 249
rect 685 215 719 249
rect 802 215 836 249
rect 880 215 914 249
rect 958 215 992 249
rect 1036 215 1070 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 18 477 69 493
rect 18 443 35 477
rect 18 409 69 443
rect 18 375 35 409
rect 18 333 69 375
rect 103 485 174 527
rect 103 451 129 485
rect 163 451 174 485
rect 103 417 174 451
rect 103 383 129 417
rect 163 383 174 417
rect 208 455 234 489
rect 268 455 544 489
rect 578 455 594 489
rect 655 477 689 493
rect 208 421 288 455
rect 723 485 799 527
rect 723 451 749 485
rect 783 451 799 485
rect 843 477 877 493
rect 655 421 689 443
rect 208 387 238 421
rect 272 387 288 421
rect 326 387 342 421
rect 376 387 689 421
rect 843 409 877 443
rect 103 367 174 383
rect 911 485 987 527
rect 911 451 937 485
rect 971 451 987 485
rect 911 417 987 451
rect 911 383 937 417
rect 971 383 987 417
rect 1031 477 1065 493
rect 1031 409 1065 443
rect 18 299 236 333
rect 18 125 52 299
rect 86 249 158 265
rect 120 215 158 249
rect 86 199 158 215
rect 192 249 236 299
rect 226 215 236 249
rect 192 199 236 215
rect 290 249 359 323
rect 426 319 442 353
rect 476 319 797 353
rect 290 215 325 249
rect 290 199 359 215
rect 393 249 517 265
rect 393 215 483 249
rect 393 199 517 215
rect 576 249 719 265
rect 576 215 617 249
rect 651 215 685 249
rect 576 199 719 215
rect 763 249 797 319
rect 843 349 877 375
rect 1099 485 1175 527
rect 1099 451 1125 485
rect 1159 451 1175 485
rect 1099 417 1175 451
rect 1099 383 1125 417
rect 1159 383 1175 417
rect 1031 349 1065 375
rect 843 315 1176 349
rect 763 215 802 249
rect 836 215 880 249
rect 914 215 958 249
rect 992 215 1036 249
rect 1070 215 1086 249
rect 124 161 158 199
rect 576 161 610 199
rect 763 165 797 215
rect 124 127 610 161
rect 652 131 797 165
rect 1130 161 1176 315
rect 18 109 69 125
rect 18 75 35 109
rect 652 93 686 131
rect 843 127 1176 161
rect 843 101 877 127
rect 18 59 69 75
rect 103 59 129 93
rect 163 59 179 93
rect 415 59 441 93
rect 475 59 686 93
rect 723 59 749 93
rect 783 59 799 93
rect 103 17 179 59
rect 723 17 799 59
rect 1031 101 1065 127
rect 843 51 877 67
rect 911 59 937 93
rect 971 59 987 93
rect 911 17 987 59
rect 1031 51 1065 67
rect 1099 59 1125 93
rect 1159 59 1175 93
rect 1099 17 1175 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 1133 153 1167 187 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 1133 289 1167 323 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 305 289 339 323 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 mux2_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1066690
string GDS_START 1057924
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
