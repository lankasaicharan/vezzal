magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3026 1975
<< nwell >>
rect -38 331 1766 704
<< pwell >>
rect 801 229 993 273
rect 1447 229 1721 273
rect 233 172 1721 229
rect 1 49 1721 172
rect 0 0 1728 49
<< scnmos >>
rect 80 62 110 146
rect 316 119 346 203
rect 402 119 432 203
rect 521 119 551 203
rect 607 119 637 203
rect 679 119 709 203
rect 884 119 914 247
rect 989 119 1019 203
rect 1103 119 1133 203
rect 1175 119 1205 203
rect 1313 75 1343 203
rect 1526 79 1556 247
rect 1612 79 1642 247
<< scpmoshvt >>
rect 80 480 110 608
rect 293 443 323 571
rect 449 443 479 527
rect 535 443 565 527
rect 675 443 705 527
rect 747 443 777 527
rect 872 379 902 547
rect 974 379 1004 547
rect 1133 379 1163 463
rect 1205 379 1235 463
rect 1313 379 1343 547
rect 1526 367 1556 619
rect 1612 367 1642 619
<< ndiff >>
rect 827 203 884 247
rect 259 178 316 203
rect 27 121 80 146
rect 27 87 35 121
rect 69 87 80 121
rect 27 62 80 87
rect 110 116 163 146
rect 259 144 267 178
rect 301 144 316 178
rect 259 119 316 144
rect 346 178 402 203
rect 346 144 357 178
rect 391 144 402 178
rect 346 119 402 144
rect 432 178 521 203
rect 432 144 461 178
rect 495 144 521 178
rect 432 119 521 144
rect 551 178 607 203
rect 551 144 562 178
rect 596 144 607 178
rect 551 119 607 144
rect 637 119 679 203
rect 709 171 884 203
rect 709 137 720 171
rect 754 137 835 171
rect 869 137 884 171
rect 709 119 884 137
rect 914 235 967 247
rect 914 201 925 235
rect 959 203 967 235
rect 1473 235 1526 247
rect 959 201 989 203
rect 914 167 989 201
rect 914 133 925 167
rect 959 133 989 167
rect 914 119 989 133
rect 1019 179 1103 203
rect 1019 145 1045 179
rect 1079 145 1103 179
rect 1019 119 1103 145
rect 1133 119 1175 203
rect 1205 183 1313 203
rect 1205 149 1216 183
rect 1250 149 1313 183
rect 1205 119 1313 149
rect 110 82 121 116
rect 155 82 163 116
rect 110 62 163 82
rect 1240 117 1313 119
rect 1240 83 1268 117
rect 1302 83 1313 117
rect 1240 75 1313 83
rect 1343 189 1396 203
rect 1343 155 1354 189
rect 1388 155 1396 189
rect 1343 121 1396 155
rect 1343 87 1354 121
rect 1388 87 1396 121
rect 1343 75 1396 87
rect 1473 201 1481 235
rect 1515 201 1526 235
rect 1473 125 1526 201
rect 1473 91 1481 125
rect 1515 91 1526 125
rect 1473 79 1526 91
rect 1556 235 1612 247
rect 1556 201 1567 235
rect 1601 201 1612 235
rect 1556 125 1612 201
rect 1556 91 1567 125
rect 1601 91 1612 125
rect 1556 79 1612 91
rect 1642 235 1695 247
rect 1642 201 1653 235
rect 1687 201 1695 235
rect 1642 125 1695 201
rect 1642 91 1653 125
rect 1687 91 1695 125
rect 1642 79 1695 91
<< pdiff >>
rect 27 574 80 608
rect 27 540 35 574
rect 69 540 80 574
rect 27 480 80 540
rect 110 594 163 608
rect 110 560 121 594
rect 155 560 163 594
rect 110 526 163 560
rect 110 492 121 526
rect 155 492 163 526
rect 110 480 163 492
rect 240 557 293 571
rect 240 523 248 557
rect 282 523 293 557
rect 240 489 293 523
rect 240 455 248 489
rect 282 455 293 489
rect 240 443 293 455
rect 323 563 380 571
rect 323 529 334 563
rect 368 529 380 563
rect 323 527 380 529
rect 799 561 857 569
rect 799 527 811 561
rect 845 547 857 561
rect 1473 607 1526 619
rect 1473 573 1481 607
rect 1515 573 1526 607
rect 845 527 872 547
rect 323 495 449 527
rect 323 461 334 495
rect 368 461 449 495
rect 323 443 449 461
rect 479 502 535 527
rect 479 468 490 502
rect 524 468 535 502
rect 479 443 535 468
rect 565 502 675 527
rect 565 468 630 502
rect 664 468 675 502
rect 565 443 675 468
rect 705 443 747 527
rect 777 443 872 527
rect 799 379 872 443
rect 902 421 974 547
rect 902 387 913 421
rect 947 387 974 421
rect 902 379 974 387
rect 1004 535 1111 547
rect 1004 501 1069 535
rect 1103 501 1111 535
rect 1004 463 1111 501
rect 1260 535 1313 547
rect 1260 501 1268 535
rect 1302 501 1313 535
rect 1260 463 1313 501
rect 1004 425 1133 463
rect 1004 391 1069 425
rect 1103 391 1133 425
rect 1004 379 1133 391
rect 1163 379 1205 463
rect 1235 438 1313 463
rect 1235 404 1246 438
rect 1280 404 1313 438
rect 1235 379 1313 404
rect 1343 535 1396 547
rect 1343 501 1354 535
rect 1388 501 1396 535
rect 1343 425 1396 501
rect 1343 391 1354 425
rect 1388 391 1396 425
rect 1343 379 1396 391
rect 1473 510 1526 573
rect 1473 476 1481 510
rect 1515 476 1526 510
rect 1473 413 1526 476
rect 1473 379 1481 413
rect 1515 379 1526 413
rect 1473 367 1526 379
rect 1556 599 1612 619
rect 1556 565 1567 599
rect 1601 565 1612 599
rect 1556 501 1612 565
rect 1556 467 1567 501
rect 1601 467 1612 501
rect 1556 420 1612 467
rect 1556 386 1567 420
rect 1601 386 1612 420
rect 1556 367 1612 386
rect 1642 607 1695 619
rect 1642 573 1653 607
rect 1687 573 1695 607
rect 1642 510 1695 573
rect 1642 476 1653 510
rect 1687 476 1695 510
rect 1642 413 1695 476
rect 1642 379 1653 413
rect 1687 379 1695 413
rect 1642 367 1695 379
<< ndiffc >>
rect 35 87 69 121
rect 267 144 301 178
rect 357 144 391 178
rect 461 144 495 178
rect 562 144 596 178
rect 720 137 754 171
rect 835 137 869 171
rect 925 201 959 235
rect 925 133 959 167
rect 1045 145 1079 179
rect 1216 149 1250 183
rect 121 82 155 116
rect 1268 83 1302 117
rect 1354 155 1388 189
rect 1354 87 1388 121
rect 1481 201 1515 235
rect 1481 91 1515 125
rect 1567 201 1601 235
rect 1567 91 1601 125
rect 1653 201 1687 235
rect 1653 91 1687 125
<< pdiffc >>
rect 35 540 69 574
rect 121 560 155 594
rect 121 492 155 526
rect 248 523 282 557
rect 248 455 282 489
rect 334 529 368 563
rect 811 527 845 561
rect 1481 573 1515 607
rect 334 461 368 495
rect 490 468 524 502
rect 630 468 664 502
rect 913 387 947 421
rect 1069 501 1103 535
rect 1268 501 1302 535
rect 1069 391 1103 425
rect 1246 404 1280 438
rect 1354 501 1388 535
rect 1354 391 1388 425
rect 1481 476 1515 510
rect 1481 379 1515 413
rect 1567 565 1601 599
rect 1567 467 1601 501
rect 1567 386 1601 420
rect 1653 573 1687 607
rect 1653 476 1687 510
rect 1653 379 1687 413
<< poly >>
rect 80 608 110 634
rect 293 615 1004 645
rect 1526 619 1556 645
rect 1612 619 1642 645
rect 293 571 323 615
rect 80 302 110 480
rect 449 527 479 553
rect 535 527 565 553
rect 675 527 705 615
rect 747 527 777 553
rect 872 547 902 573
rect 974 547 1004 615
rect 1313 547 1343 573
rect 31 286 110 302
rect 31 252 47 286
rect 81 252 110 286
rect 31 218 110 252
rect 158 364 224 380
rect 158 330 174 364
rect 208 330 224 364
rect 158 296 224 330
rect 158 262 174 296
rect 208 276 224 296
rect 293 276 323 443
rect 449 360 479 443
rect 388 344 479 360
rect 388 310 404 344
rect 438 310 479 344
rect 388 276 479 310
rect 535 411 565 443
rect 675 417 705 443
rect 535 395 610 411
rect 535 361 560 395
rect 594 361 610 395
rect 535 327 610 361
rect 747 347 777 443
rect 1133 463 1163 489
rect 1205 463 1235 489
rect 535 293 560 327
rect 594 307 610 327
rect 679 331 787 347
rect 872 335 902 379
rect 974 353 1004 379
rect 1133 357 1163 379
rect 594 293 637 307
rect 535 277 637 293
rect 208 262 346 276
rect 158 246 346 262
rect 31 184 47 218
rect 81 184 110 218
rect 316 203 346 246
rect 388 242 404 276
rect 438 242 479 276
rect 388 226 479 242
rect 402 203 432 226
rect 521 203 551 229
rect 607 203 637 277
rect 679 297 737 331
rect 771 297 787 331
rect 679 281 787 297
rect 835 319 914 335
rect 835 285 851 319
rect 885 285 914 319
rect 1052 327 1163 357
rect 1205 345 1235 379
rect 1205 329 1271 345
rect 1052 311 1082 327
rect 679 203 709 281
rect 835 269 914 285
rect 884 247 914 269
rect 989 295 1082 311
rect 989 261 1011 295
rect 1045 281 1082 295
rect 1205 295 1221 329
rect 1255 295 1271 329
rect 1045 261 1061 281
rect 1205 279 1271 295
rect 31 168 110 184
rect 80 146 110 168
rect 989 245 1061 261
rect 1175 249 1271 279
rect 1313 291 1343 379
rect 1526 335 1556 367
rect 1421 319 1556 335
rect 1313 275 1379 291
rect 989 203 1019 245
rect 1103 203 1133 229
rect 1175 203 1205 249
rect 1313 241 1329 275
rect 1363 241 1379 275
rect 1421 285 1437 319
rect 1471 299 1556 319
rect 1612 299 1642 367
rect 1471 285 1642 299
rect 1421 269 1642 285
rect 1526 247 1556 269
rect 1612 247 1642 269
rect 1313 225 1379 241
rect 1313 203 1343 225
rect 80 36 110 62
rect 316 51 346 119
rect 402 93 432 119
rect 521 51 551 119
rect 607 93 637 119
rect 679 93 709 119
rect 884 93 914 119
rect 989 93 1019 119
rect 1103 51 1133 119
rect 1175 93 1205 119
rect 316 21 1133 51
rect 1313 49 1343 75
rect 1526 53 1556 79
rect 1612 53 1642 79
<< polycont >>
rect 47 252 81 286
rect 174 330 208 364
rect 174 262 208 296
rect 404 310 438 344
rect 560 361 594 395
rect 560 293 594 327
rect 47 184 81 218
rect 404 242 438 276
rect 737 297 771 331
rect 851 285 885 319
rect 1011 261 1045 295
rect 1221 295 1255 329
rect 1329 241 1363 275
rect 1437 285 1471 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 19 574 85 649
rect 19 540 35 574
rect 69 540 85 574
rect 19 532 85 540
rect 119 594 208 610
rect 119 560 121 594
rect 155 560 208 594
rect 119 526 208 560
rect 17 286 85 498
rect 17 252 47 286
rect 81 252 85 286
rect 17 218 85 252
rect 17 184 47 218
rect 81 184 85 218
rect 17 168 85 184
rect 119 492 121 526
rect 155 492 208 526
rect 119 364 208 492
rect 119 330 174 364
rect 119 296 208 330
rect 119 262 174 296
rect 19 121 85 134
rect 19 87 35 121
rect 69 87 85 121
rect 19 17 85 87
rect 119 116 208 262
rect 242 557 284 573
rect 242 523 248 557
rect 282 523 284 557
rect 242 489 284 523
rect 242 455 248 489
rect 282 455 284 489
rect 318 563 384 649
rect 318 529 334 563
rect 368 529 384 563
rect 318 495 384 529
rect 318 461 334 495
rect 368 461 384 495
rect 318 457 384 461
rect 418 552 738 588
rect 242 421 284 455
rect 418 421 454 552
rect 242 387 454 421
rect 488 502 526 518
rect 488 468 490 502
rect 524 468 526 502
rect 242 178 317 387
rect 388 344 454 353
rect 388 310 404 344
rect 438 310 454 344
rect 388 276 454 310
rect 388 242 404 276
rect 438 242 454 276
rect 388 228 454 242
rect 488 244 526 468
rect 560 395 594 552
rect 560 327 594 361
rect 560 277 594 293
rect 628 502 670 518
rect 628 468 630 502
rect 664 468 670 502
rect 628 245 670 468
rect 704 491 738 552
rect 795 561 861 649
rect 795 527 811 561
rect 845 527 861 561
rect 795 525 861 527
rect 1067 535 1131 551
rect 1067 501 1069 535
rect 1103 501 1131 535
rect 704 457 1033 491
rect 721 421 963 423
rect 721 387 913 421
rect 947 387 963 421
rect 721 383 963 387
rect 721 331 787 383
rect 721 297 737 331
rect 771 297 787 331
rect 721 281 787 297
rect 835 319 885 335
rect 835 285 851 319
rect 835 245 885 285
rect 488 194 524 244
rect 628 211 885 245
rect 919 235 961 383
rect 997 311 1033 457
rect 1067 425 1131 501
rect 1067 391 1069 425
rect 1103 391 1131 425
rect 1230 535 1306 649
rect 1467 607 1523 649
rect 1467 573 1481 607
rect 1515 573 1523 607
rect 1230 501 1268 535
rect 1302 501 1306 535
rect 1230 438 1306 501
rect 1230 404 1246 438
rect 1280 404 1306 438
rect 1230 395 1306 404
rect 1350 535 1433 551
rect 1350 501 1354 535
rect 1388 501 1433 535
rect 1350 425 1433 501
rect 1067 375 1131 391
rect 997 295 1061 311
rect 995 261 1011 295
rect 1045 261 1061 295
rect 995 259 1061 261
rect 1097 259 1131 375
rect 1350 391 1354 425
rect 1388 391 1433 425
rect 1350 361 1433 391
rect 1467 510 1523 573
rect 1467 476 1481 510
rect 1515 476 1523 510
rect 1467 413 1523 476
rect 1467 379 1481 413
rect 1515 379 1523 413
rect 1467 363 1523 379
rect 1557 599 1610 615
rect 1557 565 1567 599
rect 1601 565 1610 599
rect 1557 501 1610 565
rect 1557 467 1567 501
rect 1601 467 1610 501
rect 1557 420 1610 467
rect 1557 386 1567 420
rect 1601 386 1610 420
rect 1205 329 1433 361
rect 1205 295 1221 329
rect 1255 327 1487 329
rect 1255 295 1271 327
rect 1205 293 1271 295
rect 1399 319 1487 327
rect 1313 275 1365 291
rect 1313 259 1329 275
rect 628 207 668 211
rect 242 144 267 178
rect 301 144 317 178
rect 242 128 317 144
rect 351 178 407 194
rect 351 144 357 178
rect 391 144 407 178
rect 119 82 121 116
rect 155 82 208 116
rect 119 66 208 82
rect 351 17 407 144
rect 445 178 524 194
rect 445 144 461 178
rect 495 144 524 178
rect 445 128 524 144
rect 558 178 668 207
rect 558 144 562 178
rect 596 173 668 178
rect 919 201 925 235
rect 959 201 961 235
rect 1097 241 1329 259
rect 1363 241 1365 275
rect 1097 225 1365 241
rect 1399 285 1437 319
rect 1471 285 1487 319
rect 596 144 612 173
rect 558 128 612 144
rect 704 171 885 177
rect 704 137 720 171
rect 754 137 835 171
rect 869 137 885 171
rect 704 17 885 137
rect 919 167 961 201
rect 919 133 925 167
rect 959 133 961 167
rect 919 117 961 133
rect 1029 179 1131 225
rect 1399 189 1433 285
rect 1029 145 1045 179
rect 1079 145 1131 179
rect 1029 129 1131 145
rect 1200 183 1304 189
rect 1200 149 1216 183
rect 1250 149 1304 183
rect 1200 117 1304 149
rect 1200 83 1268 117
rect 1302 83 1304 117
rect 1338 155 1354 189
rect 1388 155 1433 189
rect 1338 121 1433 155
rect 1338 87 1354 121
rect 1388 87 1433 121
rect 1338 83 1433 87
rect 1467 235 1523 251
rect 1467 201 1481 235
rect 1515 201 1523 235
rect 1467 125 1523 201
rect 1467 91 1481 125
rect 1515 91 1523 125
rect 1200 17 1304 83
rect 1467 17 1523 91
rect 1557 235 1610 386
rect 1644 607 1691 649
rect 1644 573 1653 607
rect 1687 573 1691 607
rect 1644 510 1691 573
rect 1644 476 1653 510
rect 1687 476 1691 510
rect 1644 413 1691 476
rect 1644 379 1653 413
rect 1687 379 1691 413
rect 1644 363 1691 379
rect 1557 201 1567 235
rect 1601 201 1610 235
rect 1557 125 1610 201
rect 1557 91 1567 125
rect 1601 91 1610 125
rect 1557 75 1610 91
rect 1644 235 1691 251
rect 1644 201 1653 235
rect 1687 201 1691 235
rect 1644 125 1691 201
rect 1644 91 1653 125
rect 1687 91 1691 125
rect 1644 17 1691 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfxtp_2
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1003074
string GDS_START 989846
<< end >>
