magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2218 1852
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 108 157 900 203
rect 1 21 900 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 198 47 228 177
rect 302 47 332 177
rect 510 47 540 177
rect 604 47 634 177
rect 688 47 718 177
rect 792 47 822 177
<< scpmoshvt >>
rect 81 413 117 497
rect 200 297 236 497
rect 294 297 330 497
rect 388 297 424 497
rect 482 297 518 497
rect 690 297 726 497
rect 784 297 820 497
<< ndiff >>
rect 134 161 198 177
rect 134 131 142 161
rect 27 101 79 131
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 127 142 131
rect 176 127 198 161
rect 109 93 198 127
rect 109 59 142 93
rect 176 59 198 93
rect 109 47 198 59
rect 228 161 302 177
rect 228 127 248 161
rect 282 127 302 161
rect 228 93 302 127
rect 228 59 248 93
rect 282 59 302 93
rect 228 47 302 59
rect 332 93 384 177
rect 332 59 342 93
rect 376 59 384 93
rect 332 47 384 59
rect 448 93 510 177
rect 448 59 456 93
rect 490 59 510 93
rect 448 47 510 59
rect 540 161 604 177
rect 540 127 550 161
rect 584 127 604 161
rect 540 47 604 127
rect 634 161 688 177
rect 634 127 644 161
rect 678 127 688 161
rect 634 93 688 127
rect 634 59 644 93
rect 678 59 688 93
rect 634 47 688 59
rect 718 169 792 177
rect 718 135 738 169
rect 772 135 792 169
rect 718 47 792 135
rect 822 93 874 177
rect 822 59 832 93
rect 866 59 874 93
rect 822 47 874 59
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 413 81 443
rect 117 485 200 497
rect 117 451 142 485
rect 176 451 200 485
rect 117 417 200 451
rect 117 413 142 417
rect 134 383 142 413
rect 176 383 200 417
rect 134 297 200 383
rect 236 485 294 497
rect 236 451 248 485
rect 282 451 294 485
rect 236 417 294 451
rect 236 383 248 417
rect 282 383 294 417
rect 236 297 294 383
rect 330 485 388 497
rect 330 451 342 485
rect 376 451 388 485
rect 330 297 388 451
rect 424 485 482 497
rect 424 451 436 485
rect 470 451 482 485
rect 424 417 482 451
rect 424 383 436 417
rect 470 383 482 417
rect 424 297 482 383
rect 518 485 572 497
rect 518 451 530 485
rect 564 451 572 485
rect 518 297 572 451
rect 636 485 690 497
rect 636 451 644 485
rect 678 451 690 485
rect 636 297 690 451
rect 726 477 784 497
rect 726 443 738 477
rect 772 443 784 477
rect 726 409 784 443
rect 726 375 738 409
rect 772 375 784 409
rect 726 297 784 375
rect 820 485 874 497
rect 820 451 832 485
rect 866 451 874 485
rect 820 297 874 451
<< ndiffc >>
rect 35 67 69 101
rect 142 127 176 161
rect 142 59 176 93
rect 248 127 282 161
rect 248 59 282 93
rect 342 59 376 93
rect 456 59 490 93
rect 550 127 584 161
rect 644 127 678 161
rect 644 59 678 93
rect 738 135 772 169
rect 832 59 866 93
<< pdiffc >>
rect 35 443 69 477
rect 142 451 176 485
rect 142 383 176 417
rect 248 451 282 485
rect 248 383 282 417
rect 342 451 376 485
rect 436 451 470 485
rect 436 383 470 417
rect 530 451 564 485
rect 644 451 678 485
rect 738 443 772 477
rect 738 375 772 409
rect 832 451 866 485
<< poly >>
rect 81 497 117 523
rect 200 497 236 523
rect 294 497 330 523
rect 388 497 424 523
rect 482 497 518 523
rect 690 497 726 523
rect 784 497 820 523
rect 81 398 117 413
rect 79 265 119 398
rect 200 282 236 297
rect 294 282 330 297
rect 388 282 424 297
rect 482 282 518 297
rect 690 282 726 297
rect 784 282 820 297
rect 79 249 156 265
rect 79 215 102 249
rect 136 215 156 249
rect 79 199 156 215
rect 198 259 238 282
rect 292 259 332 282
rect 198 249 332 259
rect 198 215 248 249
rect 282 215 332 249
rect 198 205 332 215
rect 386 259 426 282
rect 480 259 520 282
rect 688 259 728 282
rect 782 259 822 282
rect 386 249 634 259
rect 386 215 446 249
rect 480 215 528 249
rect 562 215 634 249
rect 386 205 634 215
rect 79 131 109 199
rect 198 177 228 205
rect 302 177 332 205
rect 510 177 540 205
rect 604 177 634 205
rect 688 249 822 259
rect 688 215 750 249
rect 784 215 822 249
rect 688 205 822 215
rect 688 177 718 205
rect 792 177 822 205
rect 79 21 109 47
rect 198 21 228 47
rect 302 21 332 47
rect 510 21 540 47
rect 604 21 634 47
rect 688 21 718 47
rect 792 21 822 47
<< polycont >>
rect 102 215 136 249
rect 248 215 282 249
rect 446 215 480 249
rect 528 215 562 249
rect 750 215 784 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 477 82 493
rect 18 443 35 477
rect 69 443 82 477
rect 18 413 82 443
rect 126 485 188 527
rect 126 451 142 485
rect 176 451 188 485
rect 126 417 188 451
rect 18 323 52 413
rect 126 383 142 417
rect 176 383 188 417
rect 126 367 188 383
rect 222 485 298 493
rect 222 451 248 485
rect 282 451 298 485
rect 222 417 298 451
rect 342 485 376 527
rect 342 435 376 451
rect 410 485 486 493
rect 410 451 436 485
rect 470 451 486 485
rect 222 383 248 417
rect 282 401 298 417
rect 410 417 486 451
rect 530 485 580 527
rect 564 451 580 485
rect 530 435 580 451
rect 618 485 678 527
rect 618 451 644 485
rect 618 435 678 451
rect 712 477 772 493
rect 712 443 738 477
rect 410 401 436 417
rect 282 383 436 401
rect 470 391 486 417
rect 712 409 772 443
rect 832 485 890 527
rect 866 451 890 485
rect 832 435 890 451
rect 712 391 738 409
rect 470 383 738 391
rect 222 375 738 383
rect 772 375 898 401
rect 222 357 898 375
rect 18 289 800 323
rect 18 131 52 289
rect 86 249 166 255
rect 86 215 102 249
rect 136 215 166 249
rect 213 249 378 255
rect 213 215 248 249
rect 282 215 378 249
rect 430 249 688 255
rect 430 215 446 249
rect 480 215 528 249
rect 562 215 688 249
rect 734 249 800 289
rect 734 215 750 249
rect 784 215 800 249
rect 850 181 898 357
rect 126 161 188 181
rect 18 101 82 131
rect 18 67 35 101
rect 69 67 82 101
rect 18 51 82 67
rect 126 127 142 161
rect 176 127 188 161
rect 126 93 188 127
rect 126 59 142 93
rect 176 59 188 93
rect 126 17 188 59
rect 222 161 600 181
rect 222 127 248 161
rect 282 143 550 161
rect 282 127 298 143
rect 440 127 550 143
rect 584 127 600 161
rect 644 161 678 181
rect 712 169 898 181
rect 712 135 738 169
rect 772 135 898 169
rect 712 127 898 135
rect 222 93 298 127
rect 222 59 248 93
rect 282 59 298 93
rect 222 51 298 59
rect 342 93 392 109
rect 644 93 678 127
rect 376 59 392 93
rect 342 17 392 59
rect 440 59 456 93
rect 490 59 644 93
rect 678 59 832 93
rect 866 59 890 93
rect 440 51 890 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 850 221 884 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 224 221 258 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 132 221 166 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 438 221 472 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 850 289 884 323 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 454 238 454 238 0 FreeSans 200 0 0 0 B
port 2 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand3b_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2236236
string GDS_START 2228904
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
