magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1265 -1309 2705 2641
<< nwell >>
rect -5 997 1445 1370
rect -5 -38 1445 335
<< pwell >>
rect 5 912 91 921
rect 1349 912 1435 921
rect 5 776 786 912
rect 5 420 630 776
rect 1078 692 1435 912
rect 5 411 91 420
rect 1349 411 1435 692
<< scnmos >>
rect 176 718 206 886
rect 248 718 278 886
rect 334 718 364 886
rect 406 718 436 886
rect 601 802 631 886
rect 673 802 703 886
rect 1161 718 1191 886
rect 1233 718 1263 886
rect 176 446 206 530
rect 248 446 278 530
rect 517 446 547 614
<< scpmoshvt >>
rect 176 1085 206 1285
rect 248 1085 278 1285
rect 334 1085 364 1285
rect 406 1085 436 1285
rect 601 1085 631 1285
rect 687 1085 717 1285
rect 759 1085 789 1285
rect 1003 1085 1033 1285
rect 1075 1085 1105 1285
rect 1161 1085 1191 1285
rect 1233 1085 1263 1285
rect 176 47 206 247
rect 248 47 278 247
<< ndiff >>
rect 123 874 176 886
rect 123 840 131 874
rect 165 840 176 874
rect 123 767 176 840
rect 123 733 131 767
rect 165 733 176 767
rect 123 718 176 733
rect 206 718 248 886
rect 278 878 334 886
rect 278 844 289 878
rect 323 844 334 878
rect 278 767 334 844
rect 278 733 289 767
rect 323 733 334 767
rect 278 718 334 733
rect 364 718 406 886
rect 436 864 493 886
rect 436 830 447 864
rect 481 830 493 864
rect 436 718 493 830
rect 548 848 601 886
rect 548 814 556 848
rect 590 814 601 848
rect 548 802 601 814
rect 631 802 673 886
rect 703 848 760 886
rect 703 814 714 848
rect 748 814 760 848
rect 703 802 760 814
rect 1104 846 1161 886
rect 1104 812 1116 846
rect 1150 812 1161 846
rect 1104 760 1161 812
rect 1104 726 1116 760
rect 1150 726 1161 760
rect 1104 718 1161 726
rect 1191 718 1233 886
rect 1263 874 1316 886
rect 1263 840 1274 874
rect 1308 840 1316 874
rect 1263 764 1316 840
rect 1263 730 1274 764
rect 1308 730 1316 764
rect 1263 718 1316 730
rect 464 602 517 614
rect 464 568 472 602
rect 506 568 517 602
rect 123 505 176 530
rect 123 471 131 505
rect 165 471 176 505
rect 123 446 176 471
rect 206 446 248 530
rect 278 505 331 530
rect 278 471 289 505
rect 323 471 331 505
rect 278 446 331 471
rect 464 516 517 568
rect 464 482 472 516
rect 506 482 517 516
rect 464 446 517 482
rect 547 606 604 614
rect 547 572 558 606
rect 592 572 604 606
rect 547 520 604 572
rect 547 486 558 520
rect 592 486 604 520
rect 547 446 604 486
<< pdiff >>
rect 123 1273 176 1285
rect 123 1239 131 1273
rect 165 1239 176 1273
rect 123 1199 176 1239
rect 123 1165 131 1199
rect 165 1165 176 1199
rect 123 1131 176 1165
rect 123 1097 131 1131
rect 165 1097 176 1131
rect 123 1085 176 1097
rect 206 1085 248 1285
rect 278 1277 334 1285
rect 278 1243 289 1277
rect 323 1243 334 1277
rect 278 1173 334 1243
rect 278 1139 289 1173
rect 323 1139 334 1173
rect 278 1085 334 1139
rect 364 1085 406 1285
rect 436 1195 493 1285
rect 436 1161 447 1195
rect 481 1161 493 1195
rect 436 1127 493 1161
rect 436 1093 447 1127
rect 481 1093 493 1127
rect 436 1085 493 1093
rect 547 1273 601 1285
rect 547 1239 556 1273
rect 590 1239 601 1273
rect 547 1205 601 1239
rect 547 1171 556 1205
rect 590 1171 601 1205
rect 547 1137 601 1171
rect 547 1103 556 1137
rect 590 1103 601 1137
rect 547 1085 601 1103
rect 631 1277 687 1285
rect 631 1243 642 1277
rect 676 1243 687 1277
rect 631 1209 687 1243
rect 631 1175 642 1209
rect 676 1175 687 1209
rect 631 1141 687 1175
rect 631 1107 642 1141
rect 676 1107 687 1141
rect 631 1085 687 1107
rect 717 1085 759 1285
rect 789 1195 846 1285
rect 789 1161 800 1195
rect 834 1161 846 1195
rect 789 1127 846 1161
rect 789 1093 800 1127
rect 834 1093 846 1127
rect 789 1085 846 1093
rect 946 1277 1003 1285
rect 946 1243 958 1277
rect 992 1243 1003 1277
rect 946 1202 1003 1243
rect 946 1168 958 1202
rect 992 1168 1003 1202
rect 946 1134 1003 1168
rect 946 1100 958 1134
rect 992 1100 1003 1134
rect 946 1085 1003 1100
rect 1033 1085 1075 1285
rect 1105 1277 1161 1285
rect 1105 1243 1116 1277
rect 1150 1243 1161 1277
rect 1105 1202 1161 1243
rect 1105 1168 1116 1202
rect 1150 1168 1161 1202
rect 1105 1085 1161 1168
rect 1191 1085 1233 1285
rect 1263 1273 1316 1285
rect 1263 1239 1274 1273
rect 1308 1239 1316 1273
rect 1263 1202 1316 1239
rect 1263 1168 1274 1202
rect 1308 1168 1316 1202
rect 1263 1131 1316 1168
rect 1263 1097 1274 1131
rect 1308 1097 1316 1131
rect 1263 1085 1316 1097
rect 123 235 176 247
rect 123 201 131 235
rect 165 201 176 235
rect 123 164 176 201
rect 123 130 131 164
rect 165 130 176 164
rect 123 93 176 130
rect 123 59 131 93
rect 165 59 176 93
rect 123 47 176 59
rect 206 47 248 247
rect 278 235 331 247
rect 278 201 289 235
rect 323 201 331 235
rect 278 164 331 201
rect 278 130 289 164
rect 323 130 331 164
rect 278 93 331 130
rect 278 59 289 93
rect 323 59 331 93
rect 278 47 331 59
<< ndiffc >>
rect 131 840 165 874
rect 131 733 165 767
rect 289 844 323 878
rect 289 733 323 767
rect 447 830 481 864
rect 556 814 590 848
rect 714 814 748 848
rect 1116 812 1150 846
rect 1116 726 1150 760
rect 1274 840 1308 874
rect 1274 730 1308 764
rect 472 568 506 602
rect 131 471 165 505
rect 289 471 323 505
rect 472 482 506 516
rect 558 572 592 606
rect 558 486 592 520
<< pdiffc >>
rect 131 1239 165 1273
rect 131 1165 165 1199
rect 131 1097 165 1131
rect 289 1243 323 1277
rect 289 1139 323 1173
rect 447 1161 481 1195
rect 447 1093 481 1127
rect 556 1239 590 1273
rect 556 1171 590 1205
rect 556 1103 590 1137
rect 642 1243 676 1277
rect 642 1175 676 1209
rect 642 1107 676 1141
rect 800 1161 834 1195
rect 800 1093 834 1127
rect 958 1243 992 1277
rect 958 1168 992 1202
rect 958 1100 992 1134
rect 1116 1243 1150 1277
rect 1116 1168 1150 1202
rect 1274 1239 1308 1273
rect 1274 1168 1308 1202
rect 1274 1097 1308 1131
rect 131 201 165 235
rect 131 130 165 164
rect 131 59 165 93
rect 289 201 323 235
rect 289 130 323 164
rect 289 59 323 93
<< psubdiff >>
rect 31 871 65 895
rect 31 788 65 837
rect 31 730 65 754
rect 1375 871 1409 895
rect 1375 788 1409 837
rect 1375 730 1409 754
rect 31 578 65 602
rect 31 495 65 544
rect 31 437 65 461
rect 1375 578 1409 602
rect 1375 495 1409 544
rect 1375 437 1409 461
<< nsubdiff >>
rect 31 1244 65 1268
rect 31 1157 65 1210
rect 31 1099 65 1123
rect 1375 1244 1409 1268
rect 1375 1157 1409 1210
rect 1375 1099 1409 1123
rect 31 209 65 233
rect 31 122 65 175
rect 31 64 65 88
rect 1375 209 1409 233
rect 1375 122 1409 175
rect 1375 64 1409 88
<< psubdiffcont >>
rect 31 837 65 871
rect 31 754 65 788
rect 1375 837 1409 871
rect 1375 754 1409 788
rect 31 544 65 578
rect 31 461 65 495
rect 1375 544 1409 578
rect 1375 461 1409 495
<< nsubdiffcont >>
rect 31 1210 65 1244
rect 31 1123 65 1157
rect 1375 1210 1409 1244
rect 1375 1123 1409 1157
rect 31 175 65 209
rect 31 88 65 122
rect 1375 175 1409 209
rect 1375 88 1409 122
<< poly >>
rect 176 1285 206 1311
rect 248 1285 278 1311
rect 334 1285 364 1311
rect 406 1285 436 1311
rect 601 1285 631 1311
rect 687 1285 717 1311
rect 759 1285 789 1311
rect 1003 1285 1033 1311
rect 1075 1285 1105 1311
rect 1161 1285 1191 1311
rect 1233 1285 1263 1311
rect 176 1053 206 1085
rect 248 1053 278 1085
rect 334 1070 364 1085
rect 406 1070 436 1085
rect 334 1053 549 1070
rect 176 1037 278 1053
rect 176 1003 216 1037
rect 250 1003 278 1037
rect 176 987 278 1003
rect 320 1040 549 1053
rect 320 1037 386 1040
rect 320 1003 336 1037
rect 370 1003 386 1037
rect 320 987 386 1003
rect 483 1037 549 1040
rect 483 1003 499 1037
rect 533 1003 549 1037
rect 483 987 549 1003
rect 601 974 631 1085
rect 687 974 717 1085
rect 601 958 717 974
rect 601 931 634 958
rect 600 924 634 931
rect 668 931 717 958
rect 759 931 789 1085
rect 1003 931 1033 1085
rect 1075 931 1105 1085
rect 1161 1039 1191 1085
rect 1233 1039 1263 1085
rect 1161 1023 1263 1039
rect 1161 989 1177 1023
rect 1211 989 1263 1023
rect 1161 973 1263 989
rect 668 924 789 931
rect 176 886 206 912
rect 248 886 278 912
rect 334 886 364 912
rect 406 886 436 912
rect 600 901 789 924
rect 904 901 1191 931
rect 601 886 631 901
rect 673 886 703 901
rect 601 776 631 802
rect 673 776 703 802
rect 904 783 934 901
rect 1161 886 1191 901
rect 1233 886 1263 973
rect 766 767 934 783
rect 766 733 782 767
rect 816 753 934 767
rect 816 733 832 753
rect 176 628 206 718
rect 248 628 278 718
rect 334 703 364 718
rect 406 703 436 718
rect 334 673 436 703
rect 766 717 832 733
rect 176 618 278 628
rect 399 618 429 673
rect 766 659 796 717
rect 1161 692 1191 718
rect 1233 692 1263 718
rect 176 602 314 618
rect 176 598 264 602
rect 248 568 264 598
rect 298 568 314 602
rect 176 530 206 556
rect 248 552 314 568
rect 363 602 429 618
rect 517 629 796 659
rect 517 614 547 629
rect 363 568 379 602
rect 413 568 429 602
rect 363 552 429 568
rect 248 530 278 552
rect 176 426 206 446
rect 248 426 278 446
rect 117 408 278 426
rect 517 420 547 446
rect 117 374 133 408
rect 167 374 201 408
rect 235 374 278 408
rect 117 358 278 374
rect 176 247 206 358
rect 248 247 278 358
rect 176 21 206 47
rect 248 21 278 47
<< polycont >>
rect 216 1003 250 1037
rect 336 1003 370 1037
rect 499 1003 533 1037
rect 634 924 668 958
rect 1177 989 1211 1023
rect 782 733 816 767
rect 264 568 298 602
rect 379 568 413 602
rect 133 374 167 408
rect 201 374 235 408
<< locali >>
rect 0 1315 31 1349
rect 65 1315 127 1349
rect 161 1315 223 1349
rect 257 1315 319 1349
rect 353 1315 415 1349
rect 449 1315 511 1349
rect 545 1315 607 1349
rect 641 1315 703 1349
rect 737 1315 799 1349
rect 833 1315 895 1349
rect 929 1315 991 1349
rect 1025 1315 1087 1349
rect 1121 1315 1183 1349
rect 1217 1315 1279 1349
rect 1313 1315 1375 1349
rect 1409 1315 1440 1349
rect 18 1244 78 1279
rect 18 1210 31 1244
rect 65 1210 78 1244
rect 18 1157 78 1210
rect 18 1123 31 1157
rect 65 1123 78 1157
rect 18 1044 78 1123
rect 115 1273 185 1281
rect 115 1239 131 1273
rect 165 1239 185 1273
rect 115 1199 185 1239
rect 115 1165 131 1199
rect 165 1165 185 1199
rect 115 1131 185 1165
rect 273 1277 606 1281
rect 273 1243 289 1277
rect 323 1273 606 1277
rect 323 1247 556 1273
rect 323 1243 339 1247
rect 273 1173 339 1243
rect 540 1239 556 1247
rect 590 1239 606 1273
rect 273 1139 289 1173
rect 323 1139 339 1173
rect 431 1195 497 1211
rect 431 1161 447 1195
rect 481 1161 497 1195
rect 115 1097 131 1131
rect 165 1097 185 1131
rect 431 1127 497 1161
rect 431 1105 447 1127
rect 115 1087 185 1097
rect 232 1093 447 1105
rect 481 1093 497 1127
rect 540 1205 606 1239
rect 540 1171 556 1205
rect 590 1171 606 1205
rect 540 1137 606 1171
rect 540 1103 556 1137
rect 590 1103 606 1137
rect 540 1093 606 1103
rect 642 1277 676 1315
rect 642 1209 676 1243
rect 642 1141 676 1175
rect 115 964 166 1087
rect 232 1071 465 1093
rect 642 1091 676 1107
rect 726 1247 903 1281
rect 232 1053 266 1071
rect 200 1037 266 1053
rect 200 1003 216 1037
rect 250 1003 266 1037
rect 200 998 266 1003
rect 304 1003 336 1037
rect 370 1003 386 1037
rect 304 1002 386 1003
rect 304 964 338 1002
rect 18 871 78 954
rect 18 837 31 871
rect 65 837 78 871
rect 18 788 78 837
rect 18 754 31 788
rect 65 754 78 788
rect 18 683 78 754
rect 115 930 338 964
rect 115 874 171 930
rect 115 840 131 874
rect 165 840 171 874
rect 115 767 171 840
rect 115 733 131 767
rect 165 733 171 767
rect 115 717 171 733
rect 273 878 329 896
rect 273 844 289 878
rect 323 844 329 878
rect 273 767 329 844
rect 431 880 465 1071
rect 726 1057 760 1247
rect 499 1037 760 1057
rect 533 1016 760 1037
rect 794 1195 834 1211
rect 794 1161 800 1195
rect 794 1127 834 1161
rect 794 1093 800 1127
rect 499 987 533 1003
rect 794 982 834 1093
rect 567 958 684 982
rect 567 924 634 958
rect 668 924 684 958
rect 567 901 684 924
rect 718 948 834 982
rect 868 1039 903 1247
rect 942 1277 1008 1281
rect 942 1243 958 1277
rect 992 1243 1008 1277
rect 942 1202 1008 1243
rect 942 1168 958 1202
rect 992 1168 1008 1202
rect 942 1134 1008 1168
rect 1100 1277 1166 1315
rect 1100 1243 1116 1277
rect 1150 1243 1166 1277
rect 1100 1202 1166 1243
rect 1100 1168 1116 1202
rect 1150 1168 1166 1202
rect 1100 1152 1166 1168
rect 1258 1273 1324 1281
rect 1258 1239 1274 1273
rect 1308 1239 1324 1273
rect 1258 1202 1324 1239
rect 1258 1168 1274 1202
rect 1308 1168 1324 1202
rect 942 1100 958 1134
rect 992 1118 1008 1134
rect 1258 1131 1324 1168
rect 1258 1118 1274 1131
rect 992 1100 1274 1118
rect 942 1097 1274 1100
rect 1308 1097 1324 1131
rect 942 1084 1324 1097
rect 868 1023 1211 1039
rect 868 989 1177 1023
rect 868 973 1211 989
rect 431 864 497 880
rect 431 830 447 864
rect 481 830 497 864
rect 718 848 763 948
rect 1258 874 1324 1084
rect 1362 1244 1422 1279
rect 1362 1210 1375 1244
rect 1409 1210 1422 1244
rect 1362 1157 1422 1210
rect 1362 1123 1375 1157
rect 1409 1123 1422 1157
rect 1362 1044 1422 1123
rect 431 814 497 830
rect 540 814 556 848
rect 590 814 606 848
rect 273 733 289 767
rect 323 751 329 767
rect 323 733 497 751
rect 273 717 497 733
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 429 683
rect 18 578 78 649
rect 18 544 31 578
rect 65 544 78 578
rect 18 495 78 544
rect 18 461 31 495
rect 65 461 78 495
rect 115 505 181 649
rect 463 618 497 717
rect 540 683 606 814
rect 698 814 714 848
rect 748 814 764 848
rect 698 783 764 814
rect 1100 812 1116 846
rect 1150 812 1166 846
rect 698 767 816 783
rect 698 733 782 767
rect 698 717 816 733
rect 1100 760 1166 812
rect 1100 726 1116 760
rect 1150 726 1166 760
rect 1100 683 1166 726
rect 1258 840 1274 874
rect 1308 840 1324 874
rect 1258 764 1324 840
rect 1258 730 1274 764
rect 1308 730 1324 764
rect 1258 717 1324 730
rect 1362 871 1422 954
rect 1362 837 1375 871
rect 1409 837 1422 871
rect 1362 788 1422 837
rect 1362 754 1375 788
rect 1409 754 1422 788
rect 1362 683 1422 754
rect 540 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1374 683
rect 1408 649 1440 683
rect 115 471 131 505
rect 165 471 181 505
rect 115 461 181 471
rect 215 602 329 615
rect 215 568 264 602
rect 298 568 329 602
rect 215 555 329 568
rect 363 602 429 615
rect 363 568 379 602
rect 413 568 429 602
rect 18 378 78 461
rect 215 427 249 555
rect 363 521 429 568
rect 117 408 249 427
rect 117 374 133 408
rect 167 374 201 408
rect 235 374 249 408
rect 117 306 249 374
rect 283 505 429 521
rect 283 471 289 505
rect 323 487 429 505
rect 463 602 506 618
rect 463 568 472 602
rect 463 516 506 568
rect 323 471 343 487
rect 18 209 78 288
rect 283 272 343 471
rect 463 482 472 516
rect 540 606 608 649
rect 540 572 558 606
rect 592 572 608 606
rect 540 520 608 572
rect 540 486 558 520
rect 592 486 608 520
rect 1362 578 1422 649
rect 1362 544 1375 578
rect 1409 544 1422 578
rect 1362 495 1422 544
rect 463 466 506 482
rect 1362 461 1375 495
rect 1409 461 1422 495
rect 1362 378 1422 461
rect 273 235 343 272
rect 18 175 31 209
rect 65 175 78 209
rect 18 122 78 175
rect 18 88 31 122
rect 65 88 78 122
rect 18 53 78 88
rect 115 201 131 235
rect 165 201 181 235
rect 115 164 181 201
rect 115 130 131 164
rect 165 130 181 164
rect 115 93 181 130
rect 115 59 131 93
rect 165 59 181 93
rect 115 17 181 59
rect 273 201 289 235
rect 323 201 343 235
rect 273 164 343 201
rect 273 130 289 164
rect 323 130 343 164
rect 273 93 343 130
rect 273 59 289 93
rect 323 59 343 93
rect 273 53 343 59
rect 1362 209 1422 288
rect 1362 175 1375 209
rect 1409 175 1422 209
rect 1362 122 1422 175
rect 1362 88 1375 122
rect 1409 88 1422 122
rect 1362 53 1422 88
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 1315 65 1349
rect 127 1315 161 1349
rect 223 1315 257 1349
rect 319 1315 353 1349
rect 415 1315 449 1349
rect 511 1315 545 1349
rect 607 1315 641 1349
rect 703 1315 737 1349
rect 799 1315 833 1349
rect 895 1315 929 1349
rect 991 1315 1025 1349
rect 1087 1315 1121 1349
rect 1183 1315 1217 1349
rect 1279 1315 1313 1349
rect 1375 1315 1409 1349
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1374 649 1408 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 1349 1440 1381
rect 0 1315 31 1349
rect 65 1315 127 1349
rect 161 1315 223 1349
rect 257 1315 319 1349
rect 353 1315 415 1349
rect 449 1315 511 1349
rect 545 1315 607 1349
rect 641 1315 703 1349
rect 737 1315 799 1349
rect 833 1315 895 1349
rect 929 1315 991 1349
rect 1025 1315 1087 1349
rect 1121 1315 1183 1349
rect 1217 1315 1279 1349
rect 1313 1315 1375 1349
rect 1409 1315 1440 1349
rect 0 1283 1440 1315
rect 0 683 1440 713
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1374 683
rect 1408 649 1440 683
rect 0 615 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel locali s 1279 1204 1313 1238 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 128 383 162 417 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1279 760 1313 794 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 1279 908 1313 942 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 1279 834 1313 868 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 1279 1056 1313 1090 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 1279 982 1313 1016 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 128 316 162 350 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1279 1130 1313 1164 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 607 908 641 942 0 FreeSans 200 0 0 0 SLEEP
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 31 1204 65 1238 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
flabel locali s 31 1130 65 1164 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
flabel locali s 1375 94 1409 128 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 1375 168 1409 202 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 1375 1204 1409 1238 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
flabel locali s 1375 1130 1409 1164 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
flabel locali s 1375 1056 1409 1090 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
flabel locali s 31 1056 65 1090 0 FreeSans 150 0 0 0 DESTVPB
port 3 nsew power bidirectional
rlabel comment s 0 0 0 0 4 lsbuf_lp
flabel comment s 441 1056 441 1056 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 0 1440 49 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 1283 1440 1332 0 FreeSans 200 0 0 0 DESTPWR
port 2 nsew power bidirectional
flabel metal1 s 0 615 1440 713 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 1332
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1297896
string GDS_START 1281058
<< end >>
