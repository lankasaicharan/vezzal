magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2065 1975
<< nwell >>
rect -38 331 805 704
<< pwell >>
rect 1 49 753 203
rect 0 0 768 49
<< scnmos >>
rect 82 93 112 177
rect 154 93 184 177
rect 310 93 340 177
rect 382 93 412 177
rect 572 93 602 177
rect 644 93 674 177
<< scpmoshvt >>
rect 82 489 112 573
rect 154 489 184 573
rect 240 489 270 573
rect 312 489 342 573
rect 402 489 432 573
rect 474 489 504 573
rect 572 367 602 619
rect 644 367 674 619
<< ndiff >>
rect 27 161 82 177
rect 27 127 37 161
rect 71 127 82 161
rect 27 93 82 127
rect 112 93 154 177
rect 184 152 310 177
rect 184 118 195 152
rect 229 118 265 152
rect 299 118 310 152
rect 184 93 310 118
rect 340 93 382 177
rect 412 161 465 177
rect 412 127 423 161
rect 457 127 465 161
rect 412 93 465 127
rect 519 161 572 177
rect 519 127 527 161
rect 561 127 572 161
rect 519 93 572 127
rect 602 93 644 177
rect 674 161 727 177
rect 674 127 685 161
rect 719 127 727 161
rect 674 93 727 127
<< pdiff >>
rect 519 581 572 619
rect 519 573 527 581
rect 27 539 82 573
rect 27 505 37 539
rect 71 505 82 539
rect 27 489 82 505
rect 112 489 154 573
rect 184 539 240 573
rect 184 505 195 539
rect 229 505 240 539
rect 184 489 240 505
rect 270 489 312 573
rect 342 539 402 573
rect 342 505 357 539
rect 391 505 402 539
rect 342 489 402 505
rect 432 489 474 573
rect 504 547 527 573
rect 561 547 572 581
rect 504 493 572 547
rect 504 489 527 493
rect 519 459 527 489
rect 561 459 572 493
rect 519 367 572 459
rect 602 367 644 619
rect 674 597 727 619
rect 674 563 685 597
rect 719 563 727 597
rect 674 514 727 563
rect 674 480 685 514
rect 719 480 727 514
rect 674 442 727 480
rect 674 408 685 442
rect 719 408 727 442
rect 674 367 727 408
<< ndiffc >>
rect 37 127 71 161
rect 195 118 229 152
rect 265 118 299 152
rect 423 127 457 161
rect 527 127 561 161
rect 685 127 719 161
<< pdiffc >>
rect 37 505 71 539
rect 195 505 229 539
rect 357 505 391 539
rect 527 547 561 581
rect 527 459 561 493
rect 685 563 719 597
rect 685 480 719 514
rect 685 408 719 442
<< poly >>
rect 572 619 602 645
rect 644 619 674 645
rect 82 573 112 599
rect 154 573 184 599
rect 240 573 270 599
rect 312 573 342 599
rect 402 573 432 599
rect 474 573 504 599
rect 82 397 112 489
rect 154 397 184 489
rect 82 379 184 397
rect 82 345 125 379
rect 159 345 184 379
rect 82 310 184 345
rect 82 276 125 310
rect 159 276 184 310
rect 82 260 184 276
rect 240 397 270 489
rect 312 397 342 489
rect 240 380 342 397
rect 240 346 269 380
rect 303 346 342 380
rect 240 312 342 346
rect 402 329 432 489
rect 474 329 504 489
rect 572 337 602 367
rect 644 337 674 367
rect 240 278 269 312
rect 303 278 342 312
rect 240 265 342 278
rect 396 313 530 329
rect 396 279 412 313
rect 446 279 480 313
rect 514 279 530 313
rect 240 262 340 265
rect 82 177 112 260
rect 154 177 184 260
rect 310 177 340 262
rect 396 263 530 279
rect 572 319 674 337
rect 572 285 595 319
rect 629 285 674 319
rect 396 229 426 263
rect 382 199 426 229
rect 572 251 674 285
rect 572 217 595 251
rect 629 217 674 251
rect 572 201 674 217
rect 382 177 412 199
rect 572 177 602 201
rect 644 177 674 201
rect 82 67 112 93
rect 154 67 184 93
rect 310 67 340 93
rect 382 67 412 93
rect 572 67 602 93
rect 644 67 674 93
<< polycont >>
rect 125 345 159 379
rect 125 276 159 310
rect 269 346 303 380
rect 269 278 303 312
rect 412 279 446 313
rect 480 279 514 313
rect 595 285 629 319
rect 595 217 629 251
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 179 572 245 584
rect 31 539 75 571
rect 31 505 37 539
rect 71 505 75 539
rect 31 447 75 505
rect 179 505 195 572
rect 229 505 245 572
rect 505 581 582 615
rect 505 572 527 581
rect 179 489 245 505
rect 353 539 395 571
rect 353 505 357 539
rect 391 505 395 539
rect 31 413 319 447
rect 31 161 75 413
rect 240 380 319 413
rect 353 425 395 505
rect 505 538 523 572
rect 561 547 582 581
rect 557 538 582 547
rect 505 493 582 538
rect 505 459 527 493
rect 561 459 582 493
rect 680 597 751 615
rect 680 563 685 597
rect 719 563 751 597
rect 680 514 751 563
rect 680 480 685 514
rect 719 480 751 514
rect 680 442 751 480
rect 353 391 646 425
rect 109 345 125 379
rect 159 345 184 379
rect 109 310 184 345
rect 109 276 125 310
rect 159 276 184 310
rect 240 346 269 380
rect 303 346 319 380
rect 240 312 319 346
rect 240 278 269 312
rect 303 278 319 312
rect 396 313 530 350
rect 396 279 412 313
rect 446 279 480 313
rect 514 279 530 313
rect 564 319 646 391
rect 564 285 595 319
rect 629 285 646 319
rect 109 232 184 276
rect 564 251 646 285
rect 564 245 595 251
rect 419 217 595 245
rect 629 217 646 251
rect 419 201 646 217
rect 680 408 685 442
rect 719 408 751 442
rect 31 127 37 161
rect 71 127 75 161
rect 31 86 75 127
rect 179 152 315 168
rect 179 118 195 152
rect 229 118 265 152
rect 299 118 315 152
rect 179 17 315 118
rect 419 161 461 201
rect 419 127 423 161
rect 457 127 461 161
rect 419 86 461 127
rect 510 161 577 167
rect 510 127 527 161
rect 561 127 577 161
rect 510 17 577 127
rect 680 161 751 408
rect 680 127 685 161
rect 719 127 751 161
rect 680 93 751 127
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 195 539 229 572
rect 195 538 229 539
rect 523 547 527 572
rect 527 547 557 572
rect 523 538 557 547
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 14 572 754 578
rect 14 538 195 572
rect 229 538 523 572
rect 557 538 754 572
rect 14 532 754 538
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel locali s 703 390 737 424 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 200 0 0 0 SLEEP
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 200 0 0 0 SLEEP
port 3 nsew signal input
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 iso0p_lp
flabel metal1 s 14 532 754 578 0 FreeSans 340 0 0 0 KAPWR
port 2 nsew power bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5925670
string GDS_START 5919166
<< end >>
