magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 4466 1975
<< nwell >>
rect -38 332 3206 704
<< pwell >>
rect 590 207 886 248
rect 2554 242 3146 248
rect 590 191 998 207
rect 590 184 1330 191
rect 1545 184 2130 228
rect 2554 184 3167 242
rect 1 49 3167 184
rect 0 0 3168 49
<< scpmos >>
rect 84 464 114 592
rect 174 464 204 592
rect 258 464 288 592
rect 384 464 414 592
rect 468 464 498 592
rect 687 368 717 592
rect 777 368 807 592
rect 1003 457 1033 541
rect 1110 495 1140 579
rect 1211 457 1241 541
rect 1358 457 1388 541
rect 1454 457 1484 541
rect 1590 373 1620 541
rect 1680 373 1710 541
rect 1882 424 1912 592
rect 1972 424 2002 592
rect 2073 508 2103 592
rect 2198 508 2228 592
rect 2288 508 2318 592
rect 2490 508 2520 592
rect 2591 424 2621 592
rect 2681 424 2711 592
rect 2782 368 2812 592
rect 2872 368 2902 592
rect 2962 368 2992 592
rect 3052 368 3082 592
<< nmoslvt >>
rect 84 74 114 158
rect 192 74 222 158
rect 270 74 300 158
rect 387 74 417 158
rect 465 74 495 158
rect 673 74 703 222
rect 773 74 803 222
rect 987 81 1017 165
rect 1123 81 1153 165
rect 1201 81 1231 165
rect 1415 74 1445 158
rect 1493 74 1523 158
rect 1647 74 1677 202
rect 1733 74 1763 202
rect 1931 74 1961 202
rect 2017 74 2047 202
rect 2119 74 2149 158
rect 2197 74 2227 158
rect 2305 74 2335 158
rect 2439 74 2469 158
rect 2637 74 2667 222
rect 2737 74 2767 222
rect 2854 74 2884 222
rect 2954 74 2984 222
rect 3040 74 3070 222
<< ndiff >>
rect 616 202 673 222
rect 616 168 628 202
rect 662 168 673 202
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 126 192 158
rect 114 92 139 126
rect 173 92 192 126
rect 114 74 192 92
rect 222 74 270 158
rect 300 132 387 158
rect 300 98 326 132
rect 360 98 387 132
rect 300 74 387 98
rect 417 74 465 158
rect 495 126 552 158
rect 495 92 506 126
rect 540 92 552 126
rect 495 74 552 92
rect 616 120 673 168
rect 616 86 628 120
rect 662 86 673 120
rect 616 74 673 86
rect 703 202 773 222
rect 703 168 728 202
rect 762 168 773 202
rect 703 120 773 168
rect 703 86 728 120
rect 762 86 773 120
rect 703 74 773 86
rect 803 210 860 222
rect 803 176 814 210
rect 848 176 860 210
rect 803 120 860 176
rect 803 86 814 120
rect 848 86 860 120
rect 803 74 860 86
rect 914 169 972 181
rect 914 135 926 169
rect 960 165 972 169
rect 960 135 987 165
rect 914 81 987 135
rect 1017 140 1123 165
rect 1017 106 1078 140
rect 1112 106 1123 140
rect 1017 81 1123 106
rect 1153 81 1201 165
rect 1231 96 1304 165
rect 1571 184 1647 202
rect 1571 158 1602 184
rect 1231 81 1258 96
rect 1246 62 1258 81
rect 1292 62 1304 96
rect 1358 133 1415 158
rect 1358 99 1370 133
rect 1404 99 1415 133
rect 1358 74 1415 99
rect 1445 74 1493 158
rect 1523 150 1602 158
rect 1636 150 1647 184
rect 1523 133 1647 150
rect 1523 99 1534 133
rect 1568 116 1647 133
rect 1568 99 1602 116
rect 1523 82 1602 99
rect 1636 82 1647 116
rect 1523 74 1647 82
rect 1677 190 1733 202
rect 1677 156 1688 190
rect 1722 156 1733 190
rect 1677 120 1733 156
rect 1677 86 1688 120
rect 1722 86 1733 120
rect 1677 74 1733 86
rect 1763 188 1820 202
rect 1763 154 1774 188
rect 1808 154 1820 188
rect 1763 120 1820 154
rect 1763 86 1774 120
rect 1808 86 1820 120
rect 1763 74 1820 86
rect 1874 188 1931 202
rect 1874 154 1886 188
rect 1920 154 1931 188
rect 1874 120 1931 154
rect 1874 86 1886 120
rect 1920 86 1931 120
rect 1874 74 1931 86
rect 1961 179 2017 202
rect 1961 145 1972 179
rect 2006 145 2017 179
rect 1961 74 2017 145
rect 2047 190 2104 202
rect 2047 156 2058 190
rect 2092 158 2104 190
rect 2580 210 2637 222
rect 2580 176 2592 210
rect 2626 176 2637 210
rect 2092 156 2119 158
rect 2047 120 2119 156
rect 2047 86 2058 120
rect 2092 86 2119 120
rect 2047 74 2119 86
rect 2149 74 2197 158
rect 2227 74 2305 158
rect 2335 120 2439 158
rect 2335 86 2363 120
rect 2397 86 2439 120
rect 2335 74 2439 86
rect 2469 133 2526 158
rect 2469 99 2480 133
rect 2514 99 2526 133
rect 2469 74 2526 99
rect 2580 120 2637 176
rect 2580 86 2592 120
rect 2626 86 2637 120
rect 2580 74 2637 86
rect 2667 210 2737 222
rect 2667 176 2692 210
rect 2726 176 2737 210
rect 2667 120 2737 176
rect 2667 86 2692 120
rect 2726 86 2737 120
rect 2667 74 2737 86
rect 2767 210 2854 222
rect 2767 176 2795 210
rect 2829 176 2854 210
rect 2767 120 2854 176
rect 2767 86 2795 120
rect 2829 86 2854 120
rect 2767 74 2854 86
rect 2884 146 2954 222
rect 2884 112 2895 146
rect 2929 112 2954 146
rect 2884 74 2954 112
rect 2984 210 3040 222
rect 2984 176 2995 210
rect 3029 176 3040 210
rect 2984 120 3040 176
rect 2984 86 2995 120
rect 3029 86 3040 120
rect 2984 74 3040 86
rect 3070 216 3120 222
rect 3070 204 3141 216
rect 3070 170 3095 204
rect 3129 170 3141 204
rect 3070 120 3141 170
rect 3070 86 3095 120
rect 3129 86 3141 120
rect 3070 74 3141 86
rect 1246 43 1304 62
<< pdiff >>
rect 516 616 574 628
rect 516 592 528 616
rect 27 580 84 592
rect 27 546 37 580
rect 71 546 84 580
rect 27 510 84 546
rect 27 476 37 510
rect 71 476 84 510
rect 27 464 84 476
rect 114 573 174 592
rect 114 539 127 573
rect 161 539 174 573
rect 114 464 174 539
rect 204 464 258 592
rect 288 566 384 592
rect 288 532 319 566
rect 353 532 384 566
rect 288 464 384 532
rect 414 464 468 592
rect 498 582 528 592
rect 562 582 574 616
rect 498 464 574 582
rect 628 414 687 592
rect 628 380 640 414
rect 674 380 687 414
rect 628 368 687 380
rect 717 573 777 592
rect 717 539 730 573
rect 764 539 777 573
rect 717 368 777 539
rect 807 573 876 592
rect 807 539 830 573
rect 864 539 876 573
rect 807 520 876 539
rect 807 368 860 520
rect 1057 541 1110 579
rect 944 516 1003 541
rect 944 482 956 516
rect 990 482 1003 516
rect 944 457 1003 482
rect 1033 517 1110 541
rect 1033 483 1046 517
rect 1080 495 1110 517
rect 1140 541 1193 579
rect 1259 576 1317 588
rect 1259 542 1271 576
rect 1305 542 1317 576
rect 1823 575 1882 592
rect 1259 541 1317 542
rect 1823 541 1835 575
rect 1869 541 1882 575
rect 1140 495 1211 541
rect 1080 483 1092 495
rect 1033 457 1092 483
rect 1158 457 1211 495
rect 1241 457 1358 541
rect 1388 516 1454 541
rect 1388 482 1407 516
rect 1441 482 1454 516
rect 1388 457 1454 482
rect 1484 518 1590 541
rect 1484 484 1543 518
rect 1577 484 1590 518
rect 1484 457 1590 484
rect 1537 373 1590 457
rect 1620 527 1680 541
rect 1620 493 1633 527
rect 1667 493 1680 527
rect 1620 458 1680 493
rect 1620 424 1633 458
rect 1667 424 1680 458
rect 1620 373 1680 424
rect 1710 527 1769 541
rect 1710 493 1723 527
rect 1757 493 1769 527
rect 1823 524 1882 541
rect 1710 480 1769 493
rect 1710 373 1763 480
rect 1829 424 1882 524
rect 1912 538 1972 592
rect 1912 504 1925 538
rect 1959 504 1972 538
rect 1912 470 1972 504
rect 1912 436 1925 470
rect 1959 436 1972 470
rect 1912 424 1972 436
rect 2002 566 2073 592
rect 2002 532 2025 566
rect 2059 532 2073 566
rect 2002 508 2073 532
rect 2103 580 2198 592
rect 2103 546 2133 580
rect 2167 546 2198 580
rect 2103 508 2198 546
rect 2228 580 2288 592
rect 2228 546 2241 580
rect 2275 546 2288 580
rect 2228 508 2288 546
rect 2318 567 2377 592
rect 2318 533 2331 567
rect 2365 533 2377 567
rect 2318 508 2377 533
rect 2431 580 2490 592
rect 2431 546 2443 580
rect 2477 546 2490 580
rect 2431 508 2490 546
rect 2520 567 2591 592
rect 2520 533 2544 567
rect 2578 533 2591 567
rect 2520 508 2591 533
rect 2002 424 2055 508
rect 2538 424 2591 508
rect 2621 580 2681 592
rect 2621 546 2634 580
rect 2668 546 2681 580
rect 2621 470 2681 546
rect 2621 436 2634 470
rect 2668 436 2681 470
rect 2621 424 2681 436
rect 2711 580 2782 592
rect 2711 546 2724 580
rect 2758 546 2782 580
rect 2711 470 2782 546
rect 2711 436 2724 470
rect 2758 436 2782 470
rect 2711 424 2782 436
rect 2729 368 2782 424
rect 2812 580 2872 592
rect 2812 546 2825 580
rect 2859 546 2872 580
rect 2812 497 2872 546
rect 2812 463 2825 497
rect 2859 463 2872 497
rect 2812 414 2872 463
rect 2812 380 2825 414
rect 2859 380 2872 414
rect 2812 368 2872 380
rect 2902 580 2962 592
rect 2902 546 2915 580
rect 2949 546 2962 580
rect 2902 498 2962 546
rect 2902 464 2915 498
rect 2949 464 2962 498
rect 2902 368 2962 464
rect 2992 580 3052 592
rect 2992 546 3005 580
rect 3039 546 3052 580
rect 2992 497 3052 546
rect 2992 463 3005 497
rect 3039 463 3052 497
rect 2992 414 3052 463
rect 2992 380 3005 414
rect 3039 380 3052 414
rect 2992 368 3052 380
rect 3082 580 3141 592
rect 3082 546 3095 580
rect 3129 546 3141 580
rect 3082 510 3141 546
rect 3082 476 3095 510
rect 3129 476 3141 510
rect 3082 440 3141 476
rect 3082 406 3095 440
rect 3129 406 3141 440
rect 3082 368 3141 406
<< ndiffc >>
rect 628 168 662 202
rect 39 99 73 133
rect 139 92 173 126
rect 326 98 360 132
rect 506 92 540 126
rect 628 86 662 120
rect 728 168 762 202
rect 728 86 762 120
rect 814 176 848 210
rect 814 86 848 120
rect 926 135 960 169
rect 1078 106 1112 140
rect 1258 62 1292 96
rect 1370 99 1404 133
rect 1602 150 1636 184
rect 1534 99 1568 133
rect 1602 82 1636 116
rect 1688 156 1722 190
rect 1688 86 1722 120
rect 1774 154 1808 188
rect 1774 86 1808 120
rect 1886 154 1920 188
rect 1886 86 1920 120
rect 1972 145 2006 179
rect 2058 156 2092 190
rect 2592 176 2626 210
rect 2058 86 2092 120
rect 2363 86 2397 120
rect 2480 99 2514 133
rect 2592 86 2626 120
rect 2692 176 2726 210
rect 2692 86 2726 120
rect 2795 176 2829 210
rect 2795 86 2829 120
rect 2895 112 2929 146
rect 2995 176 3029 210
rect 2995 86 3029 120
rect 3095 170 3129 204
rect 3095 86 3129 120
<< pdiffc >>
rect 37 546 71 580
rect 37 476 71 510
rect 127 539 161 573
rect 319 532 353 566
rect 528 582 562 616
rect 640 380 674 414
rect 730 539 764 573
rect 830 539 864 573
rect 956 482 990 516
rect 1046 483 1080 517
rect 1271 542 1305 576
rect 1835 541 1869 575
rect 1407 482 1441 516
rect 1543 484 1577 518
rect 1633 493 1667 527
rect 1633 424 1667 458
rect 1723 493 1757 527
rect 1925 504 1959 538
rect 1925 436 1959 470
rect 2025 532 2059 566
rect 2133 546 2167 580
rect 2241 546 2275 580
rect 2331 533 2365 567
rect 2443 546 2477 580
rect 2544 533 2578 567
rect 2634 546 2668 580
rect 2634 436 2668 470
rect 2724 546 2758 580
rect 2724 436 2758 470
rect 2825 546 2859 580
rect 2825 463 2859 497
rect 2825 380 2859 414
rect 2915 546 2949 580
rect 2915 464 2949 498
rect 3005 546 3039 580
rect 3005 463 3039 497
rect 3005 380 3039 414
rect 3095 546 3129 580
rect 3095 476 3129 510
rect 3095 406 3129 440
<< poly >>
rect 84 592 114 618
rect 174 592 204 618
rect 258 592 288 618
rect 384 592 414 618
rect 468 592 498 618
rect 687 592 717 618
rect 777 592 807 618
rect 891 615 2005 645
rect 84 449 114 464
rect 174 449 204 464
rect 258 449 288 464
rect 384 449 414 464
rect 468 449 498 464
rect 81 430 117 449
rect 171 430 207 449
rect 255 430 291 449
rect 381 432 417 449
rect 81 414 207 430
rect 81 380 121 414
rect 155 400 207 414
rect 249 414 315 430
rect 155 380 201 400
rect 81 346 201 380
rect 249 380 265 414
rect 299 380 315 414
rect 249 364 315 380
rect 357 416 423 432
rect 357 382 373 416
rect 407 382 423 416
rect 357 366 423 382
rect 465 422 501 449
rect 465 406 572 422
rect 465 372 522 406
rect 556 372 572 406
rect 81 312 121 346
rect 155 312 201 346
rect 81 296 201 312
rect 84 158 114 296
rect 162 232 228 248
rect 162 198 178 232
rect 212 198 228 232
rect 162 182 228 198
rect 192 158 222 182
rect 270 158 300 364
rect 465 338 572 372
rect 891 424 921 615
rect 1107 594 1143 615
rect 1879 607 1915 615
rect 1969 607 2005 615
rect 1110 579 1140 594
rect 1882 592 1912 607
rect 1972 592 2002 607
rect 2073 592 2103 618
rect 2198 592 2228 618
rect 2288 592 2318 618
rect 2490 592 2520 618
rect 2591 592 2621 618
rect 2681 592 2711 618
rect 2782 592 2812 618
rect 2872 592 2902 618
rect 2962 592 2992 618
rect 3052 592 3082 618
rect 1003 541 1033 567
rect 1211 541 1241 567
rect 1358 541 1388 567
rect 1454 541 1484 567
rect 1590 541 1620 567
rect 1680 541 1710 567
rect 1110 469 1140 495
rect 1003 442 1033 457
rect 1211 442 1241 457
rect 1358 442 1388 457
rect 1454 442 1484 457
rect 875 394 921 424
rect 687 353 717 368
rect 777 353 807 368
rect 343 300 417 316
rect 343 266 359 300
rect 393 266 417 300
rect 343 250 417 266
rect 387 158 417 250
rect 465 304 522 338
rect 556 304 572 338
rect 684 310 720 353
rect 774 336 810 353
rect 875 336 905 394
rect 1000 346 1036 442
rect 1208 422 1244 442
rect 1100 405 1166 421
rect 1100 371 1116 405
rect 1150 371 1166 405
rect 1100 346 1166 371
rect 1208 406 1274 422
rect 1208 372 1224 406
rect 1258 372 1274 406
rect 1208 356 1274 372
rect 1355 356 1391 442
rect 1451 356 1487 442
rect 2073 493 2103 508
rect 2198 493 2228 508
rect 2288 493 2318 508
rect 2490 493 2520 508
rect 2070 427 2106 493
rect 1882 398 1912 424
rect 1972 409 2002 424
rect 2070 411 2153 427
rect 1590 358 1620 373
rect 1680 358 1710 373
rect 773 320 905 336
rect 465 270 572 304
rect 465 236 522 270
rect 556 236 572 270
rect 665 294 731 310
rect 665 260 681 294
rect 715 260 731 294
rect 665 244 731 260
rect 773 286 793 320
rect 827 286 905 320
rect 773 270 905 286
rect 947 330 1166 346
rect 947 296 963 330
rect 997 316 1166 330
rect 997 296 1036 316
rect 947 280 1036 296
rect 465 220 572 236
rect 673 222 703 244
rect 773 222 803 270
rect 875 238 905 270
rect 465 158 495 220
rect 875 208 1017 238
rect 987 165 1017 208
rect 1123 165 1153 316
rect 1237 253 1267 356
rect 1201 237 1267 253
rect 1201 203 1217 237
rect 1251 203 1267 237
rect 1325 340 1391 356
rect 1325 306 1341 340
rect 1375 306 1391 340
rect 1325 272 1391 306
rect 1439 340 1523 356
rect 1439 306 1455 340
rect 1489 306 1523 340
rect 1439 290 1523 306
rect 1325 238 1341 272
rect 1375 238 1391 272
rect 1325 222 1391 238
rect 1201 187 1267 203
rect 1361 203 1391 222
rect 1201 165 1231 187
rect 1361 173 1445 203
rect 1415 158 1445 173
rect 1493 158 1523 290
rect 1587 290 1623 358
rect 1677 290 1713 358
rect 1809 340 1875 356
rect 1809 306 1825 340
rect 1859 306 1875 340
rect 1969 319 2005 409
rect 2070 377 2103 411
rect 2137 377 2153 411
rect 2070 361 2153 377
rect 1809 290 1875 306
rect 1587 274 1713 290
rect 1587 240 1603 274
rect 1637 247 1713 274
rect 1845 247 1875 290
rect 1975 289 2149 319
rect 1637 240 1763 247
rect 1587 224 1763 240
rect 1647 217 1763 224
rect 1845 217 2047 247
rect 1647 202 1677 217
rect 1733 202 1763 217
rect 1931 202 1961 217
rect 2017 202 2047 217
rect 84 48 114 74
rect 192 48 222 74
rect 270 48 300 74
rect 387 48 417 74
rect 465 48 495 74
rect 673 48 703 74
rect 773 48 803 74
rect 987 55 1017 81
rect 1123 55 1153 81
rect 1201 55 1231 81
rect 2119 158 2149 289
rect 2195 246 2231 493
rect 2285 428 2321 493
rect 2285 412 2360 428
rect 2285 378 2310 412
rect 2344 378 2360 412
rect 2487 408 2523 493
rect 2591 409 2621 424
rect 2681 409 2711 424
rect 2588 408 2624 409
rect 2678 408 2714 409
rect 2285 344 2360 378
rect 2285 310 2310 344
rect 2344 310 2360 344
rect 2285 294 2360 310
rect 2408 386 2714 408
rect 2408 352 2424 386
rect 2458 378 2714 386
rect 2458 352 2523 378
rect 2408 318 2523 352
rect 2191 230 2257 246
rect 2191 196 2207 230
rect 2241 196 2257 230
rect 2191 180 2257 196
rect 2197 158 2227 180
rect 2305 158 2335 294
rect 2408 284 2424 318
rect 2458 284 2523 318
rect 2408 268 2523 284
rect 2439 158 2469 268
rect 2637 222 2667 378
rect 2782 353 2812 368
rect 2872 353 2902 368
rect 2962 353 2992 368
rect 3052 353 3082 368
rect 2779 330 2815 353
rect 2869 330 2905 353
rect 2959 330 2995 353
rect 2737 314 2995 330
rect 2737 280 2753 314
rect 2787 280 2821 314
rect 2855 280 2889 314
rect 2923 294 2995 314
rect 3049 294 3085 353
rect 2923 280 3085 294
rect 2737 264 3085 280
rect 2737 222 2767 264
rect 2854 222 2884 264
rect 2954 222 2984 264
rect 3040 222 3070 264
rect 1415 48 1445 74
rect 1493 48 1523 74
rect 1647 48 1677 74
rect 1733 48 1763 74
rect 1931 48 1961 74
rect 2017 48 2047 74
rect 2119 48 2149 74
rect 2197 48 2227 74
rect 2305 48 2335 74
rect 2439 48 2469 74
rect 2637 48 2667 74
rect 2737 48 2767 74
rect 2854 48 2884 74
rect 2954 48 2984 74
rect 3040 48 3070 74
<< polycont >>
rect 121 380 155 414
rect 265 380 299 414
rect 373 382 407 416
rect 522 372 556 406
rect 121 312 155 346
rect 178 198 212 232
rect 359 266 393 300
rect 522 304 556 338
rect 1116 371 1150 405
rect 1224 372 1258 406
rect 522 236 556 270
rect 681 260 715 294
rect 793 286 827 320
rect 963 296 997 330
rect 1217 203 1251 237
rect 1341 306 1375 340
rect 1455 306 1489 340
rect 1341 238 1375 272
rect 1825 306 1859 340
rect 2103 377 2137 411
rect 1603 240 1637 274
rect 2310 378 2344 412
rect 2310 310 2344 344
rect 2424 352 2458 386
rect 2207 196 2241 230
rect 2424 284 2458 318
rect 2753 280 2787 314
rect 2821 280 2855 314
rect 2889 280 2923 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 21 580 71 596
rect 21 546 37 580
rect 21 510 71 546
rect 111 573 177 649
rect 512 616 578 649
rect 512 582 528 616
rect 562 582 578 616
rect 111 539 127 573
rect 161 539 177 573
rect 111 532 177 539
rect 285 566 477 582
rect 512 566 578 582
rect 714 573 780 649
rect 285 532 319 566
rect 353 532 477 566
rect 714 539 730 573
rect 764 539 780 573
rect 21 476 37 510
rect 443 498 635 532
rect 714 516 780 539
rect 814 579 1166 613
rect 814 573 880 579
rect 814 539 830 573
rect 864 539 880 573
rect 814 516 880 539
rect 940 516 1006 545
rect 71 476 409 498
rect 21 464 409 476
rect 21 248 71 464
rect 105 414 171 430
rect 105 380 121 414
rect 155 380 171 414
rect 105 346 171 380
rect 221 414 315 430
rect 221 380 265 414
rect 299 380 315 414
rect 221 364 315 380
rect 357 416 409 464
rect 357 382 373 416
rect 407 382 409 416
rect 357 366 409 382
rect 105 312 121 346
rect 155 316 171 346
rect 155 312 409 316
rect 105 300 409 312
rect 105 282 359 300
rect 343 266 359 282
rect 393 266 409 300
rect 343 250 409 266
rect 21 232 228 248
rect 21 198 178 232
rect 212 198 228 232
rect 443 216 477 498
rect 601 482 635 498
rect 940 482 956 516
rect 990 482 1006 516
rect 601 448 1006 482
rect 511 406 567 430
rect 511 372 522 406
rect 556 372 567 406
rect 511 338 567 372
rect 511 304 522 338
rect 556 304 567 338
rect 511 270 567 304
rect 511 236 522 270
rect 556 236 567 270
rect 511 220 567 236
rect 601 380 640 414
rect 674 380 843 414
rect 601 364 843 380
rect 21 182 228 198
rect 358 182 477 216
rect 601 202 635 364
rect 777 320 843 364
rect 669 294 743 310
rect 669 260 681 294
rect 715 260 743 294
rect 777 286 793 320
rect 827 286 843 320
rect 777 270 843 286
rect 882 380 1006 448
rect 1040 517 1096 545
rect 1040 483 1046 517
rect 1080 483 1096 517
rect 1040 455 1096 483
rect 1132 492 1166 579
rect 1255 576 1305 649
rect 1255 542 1271 576
rect 1255 526 1305 542
rect 1339 579 1509 613
rect 1339 492 1373 579
rect 1132 458 1373 492
rect 1407 516 1441 545
rect 669 236 743 260
rect 814 210 848 226
rect 21 133 89 182
rect 358 148 392 182
rect 601 168 628 202
rect 662 168 678 202
rect 21 99 39 133
rect 73 99 89 133
rect 21 70 89 99
rect 123 126 189 148
rect 123 92 139 126
rect 173 92 189 126
rect 123 17 189 92
rect 295 132 392 148
rect 295 98 326 132
rect 360 98 392 132
rect 295 82 392 98
rect 490 126 556 148
rect 490 92 506 126
rect 540 92 556 126
rect 490 17 556 92
rect 601 120 678 168
rect 601 86 628 120
rect 662 86 678 120
rect 601 70 678 86
rect 712 168 728 202
rect 762 168 778 202
rect 712 120 778 168
rect 712 86 728 120
rect 762 86 778 120
rect 712 17 778 86
rect 814 120 848 176
rect 882 185 916 380
rect 950 330 1006 346
rect 950 296 963 330
rect 997 296 1006 330
rect 950 253 1006 296
rect 1040 321 1074 455
rect 1132 421 1166 458
rect 1407 424 1441 482
rect 1108 405 1166 421
rect 1108 371 1116 405
rect 1150 371 1166 405
rect 1108 355 1166 371
rect 1208 406 1441 424
rect 1208 372 1224 406
rect 1258 390 1441 406
rect 1475 424 1509 579
rect 1543 518 1577 649
rect 1543 458 1577 484
rect 1617 527 1673 543
rect 1617 493 1633 527
rect 1667 493 1673 527
rect 1617 458 1673 493
rect 1707 527 1773 649
rect 1707 493 1723 527
rect 1757 493 1773 527
rect 1819 575 2075 615
rect 1819 541 1835 575
rect 1869 572 2075 575
rect 1869 541 1875 572
rect 1819 520 1875 541
rect 2009 566 2075 572
rect 1707 492 1773 493
rect 1909 504 1925 538
rect 1959 504 1975 538
rect 1909 470 1975 504
rect 1909 458 1925 470
rect 1617 424 1633 458
rect 1667 436 1925 458
rect 1959 436 1975 470
rect 2009 532 2025 566
rect 2059 532 2075 566
rect 2009 496 2075 532
rect 2109 580 2191 596
rect 2109 546 2133 580
rect 2167 546 2191 580
rect 2109 530 2191 546
rect 2225 580 2275 649
rect 2225 546 2241 580
rect 2225 530 2275 546
rect 2315 567 2381 596
rect 2315 533 2331 567
rect 2365 533 2381 567
rect 2315 496 2381 533
rect 2427 580 2510 596
rect 2427 546 2443 580
rect 2477 546 2510 580
rect 2427 530 2510 546
rect 2009 462 2442 496
rect 1667 424 1975 436
rect 1475 390 1579 424
rect 1909 420 1975 424
rect 2087 411 2153 427
rect 1258 372 1274 390
rect 1208 356 1274 372
rect 1545 386 1875 390
rect 2087 386 2103 411
rect 1545 377 2103 386
rect 2137 377 2153 411
rect 1545 356 2153 377
rect 1325 340 1391 356
rect 1325 321 1341 340
rect 1040 306 1341 321
rect 1375 306 1391 340
rect 1040 287 1391 306
rect 1439 350 1511 356
rect 1439 340 1471 350
rect 1439 306 1455 340
rect 1505 316 1511 350
rect 1489 306 1511 316
rect 1439 290 1511 306
rect 1809 352 2153 356
rect 1809 340 1875 352
rect 1809 306 1825 340
rect 1859 306 1875 340
rect 2187 314 2221 462
rect 1809 290 1875 306
rect 950 219 1028 253
rect 882 169 960 185
rect 882 135 926 169
rect 882 119 960 135
rect 814 85 848 86
rect 994 85 1028 219
rect 814 51 1028 85
rect 1062 140 1128 287
rect 1325 272 1391 287
rect 1201 237 1267 253
rect 1201 203 1217 237
rect 1251 203 1267 237
rect 1325 238 1341 272
rect 1375 256 1391 272
rect 1587 274 1653 290
rect 1587 256 1603 274
rect 1375 240 1603 256
rect 1637 240 1653 274
rect 2042 280 2221 314
rect 2294 412 2374 428
rect 2294 378 2310 412
rect 2344 378 2374 412
rect 2294 350 2374 378
rect 2294 344 2335 350
rect 2294 310 2310 344
rect 2369 316 2374 350
rect 2344 310 2374 316
rect 2294 294 2374 310
rect 2408 402 2442 462
rect 2476 470 2510 530
rect 2544 567 2594 649
rect 2578 533 2594 567
rect 2544 504 2594 533
rect 2634 580 2668 596
rect 2634 470 2668 546
rect 2476 436 2542 470
rect 2408 386 2474 402
rect 2408 352 2424 386
rect 2458 352 2474 386
rect 2408 318 2474 352
rect 2408 284 2424 318
rect 2458 284 2474 318
rect 1375 238 1653 240
rect 1325 222 1653 238
rect 1688 222 2006 256
rect 1201 188 1267 203
rect 1688 190 1722 222
rect 1201 154 1420 188
rect 1062 106 1078 140
rect 1112 106 1128 140
rect 1354 133 1420 154
rect 1062 77 1128 106
rect 1242 96 1308 120
rect 1242 62 1258 96
rect 1292 62 1308 96
rect 1354 99 1370 133
rect 1404 99 1420 133
rect 1354 70 1420 99
rect 1518 184 1652 186
rect 1518 150 1602 184
rect 1636 150 1652 184
rect 1518 133 1652 150
rect 1518 99 1534 133
rect 1568 116 1652 133
rect 1568 99 1602 116
rect 1518 82 1602 99
rect 1636 82 1652 116
rect 1242 17 1308 62
rect 1518 17 1652 82
rect 1688 120 1722 156
rect 1688 70 1722 86
rect 1758 154 1774 188
rect 1808 154 1824 188
rect 1758 120 1824 154
rect 1758 86 1774 120
rect 1808 86 1824 120
rect 1758 17 1824 86
rect 1870 154 1886 188
rect 1920 154 1936 188
rect 1870 120 1936 154
rect 1870 86 1886 120
rect 1920 86 1936 120
rect 1972 179 2006 222
rect 1972 119 2006 145
rect 2042 190 2108 280
rect 2408 268 2474 284
rect 2042 156 2058 190
rect 2092 156 2108 190
rect 2191 230 2257 246
rect 2191 196 2207 230
rect 2241 214 2257 230
rect 2508 214 2542 436
rect 2634 330 2668 436
rect 2708 580 2774 649
rect 2708 546 2724 580
rect 2758 546 2774 580
rect 2708 470 2774 546
rect 2708 436 2724 470
rect 2758 436 2774 470
rect 2708 420 2774 436
rect 2809 580 2865 596
rect 2809 546 2825 580
rect 2859 546 2865 580
rect 2809 497 2865 546
rect 2809 463 2825 497
rect 2859 463 2865 497
rect 2899 580 2965 649
rect 2899 546 2915 580
rect 2949 546 2965 580
rect 2899 498 2965 546
rect 2899 464 2915 498
rect 2949 464 2965 498
rect 3005 580 3039 596
rect 3005 497 3039 546
rect 2809 430 2865 463
rect 3005 430 3039 463
rect 2809 414 3039 430
rect 2809 380 2825 414
rect 2859 380 3005 414
rect 3079 580 3145 649
rect 3079 546 3095 580
rect 3129 546 3145 580
rect 3079 510 3145 546
rect 3079 476 3095 510
rect 3129 476 3145 510
rect 3079 440 3145 476
rect 3079 406 3095 440
rect 3129 406 3145 440
rect 3079 390 3145 406
rect 2809 364 3039 380
rect 3005 356 3039 364
rect 2634 314 2939 330
rect 3005 322 3143 356
rect 2634 298 2753 314
rect 2241 196 2542 214
rect 2191 180 2542 196
rect 2042 120 2108 156
rect 1870 85 1936 86
rect 2042 86 2058 120
rect 2092 86 2108 120
rect 2042 85 2108 86
rect 1870 51 2108 85
rect 2330 120 2430 136
rect 2330 86 2363 120
rect 2397 86 2430 120
rect 2330 17 2430 86
rect 2464 133 2542 180
rect 2464 99 2480 133
rect 2514 99 2542 133
rect 2464 70 2542 99
rect 2576 280 2753 298
rect 2787 280 2821 314
rect 2855 280 2889 314
rect 2923 280 2939 314
rect 3097 288 3143 322
rect 2576 264 2939 280
rect 2576 210 2642 264
rect 2979 254 3143 288
rect 2979 230 3045 254
rect 2576 176 2592 210
rect 2626 176 2642 210
rect 2576 120 2642 176
rect 2576 86 2592 120
rect 2626 86 2642 120
rect 2576 70 2642 86
rect 2676 210 2742 226
rect 2676 176 2692 210
rect 2726 176 2742 210
rect 2676 120 2742 176
rect 2676 86 2692 120
rect 2726 86 2742 120
rect 2676 17 2742 86
rect 2779 210 3045 230
rect 2779 176 2795 210
rect 2829 196 2995 210
rect 2829 176 2845 196
rect 2779 120 2845 176
rect 2979 176 2995 196
rect 3029 176 3045 210
rect 2779 86 2795 120
rect 2829 86 2845 120
rect 2779 70 2845 86
rect 2879 146 2945 162
rect 2879 112 2895 146
rect 2929 112 2945 146
rect 2879 17 2945 112
rect 2979 120 3045 176
rect 2979 86 2995 120
rect 3029 86 3045 120
rect 2979 70 3045 86
rect 3079 204 3145 220
rect 3079 170 3095 204
rect 3129 170 3145 204
rect 3079 120 3145 170
rect 3079 86 3095 120
rect 3129 86 3145 120
rect 3079 17 3145 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 1471 340 1505 350
rect 1471 316 1489 340
rect 1489 316 1505 340
rect 2335 344 2369 350
rect 2335 316 2344 344
rect 2344 316 2369 344
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
<< metal1 >>
rect 0 683 3168 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 0 617 3168 649
rect 1459 350 1517 356
rect 1459 316 1471 350
rect 1505 347 1517 350
rect 2323 350 2381 356
rect 2323 347 2335 350
rect 1505 319 2335 347
rect 1505 316 1517 319
rect 1459 310 1517 316
rect 2323 316 2335 319
rect 2369 316 2381 350
rect 2323 310 2381 316
rect 0 17 3168 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
rect 0 -49 3168 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfstp_4
flabel comment s 1252 275 1252 275 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 1100 328 1100 328 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 3168 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 3168 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 2335 316 2369 350 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel metal1 s 0 617 3168 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 3168 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 3103 316 3137 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3168 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 177418
string GDS_START 154454
<< end >>
