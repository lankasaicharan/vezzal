magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 331 1958 704
rect 331 299 973 331
<< pwell >>
rect 337 229 923 241
rect 1 49 1917 229
rect 0 0 1920 49
<< scnmos >>
rect 84 119 114 203
rect 170 119 200 203
rect 420 131 450 215
rect 556 47 586 215
rect 642 47 672 215
rect 728 47 758 215
rect 814 47 844 215
rect 922 119 952 203
rect 994 119 1024 203
rect 1080 119 1110 203
rect 1152 119 1182 203
rect 1337 119 1367 203
rect 1409 119 1439 203
rect 1495 119 1525 203
rect 1589 119 1619 203
rect 1804 119 1834 203
<< scpmoshvt >>
rect 84 402 114 530
rect 170 402 200 530
rect 417 335 447 463
rect 526 335 556 587
rect 612 335 642 587
rect 698 335 728 587
rect 784 335 814 587
rect 969 431 999 559
rect 1041 431 1071 559
rect 1127 431 1157 559
rect 1229 419 1259 547
rect 1373 419 1403 547
rect 1445 419 1475 547
rect 1559 431 1589 559
rect 1661 419 1691 547
rect 1747 419 1777 547
<< ndiff >>
rect 27 165 84 203
rect 27 131 35 165
rect 69 131 84 165
rect 27 119 84 131
rect 114 165 170 203
rect 114 131 125 165
rect 159 131 170 165
rect 114 119 170 131
rect 200 178 253 203
rect 200 144 211 178
rect 245 144 253 178
rect 200 119 253 144
rect 363 178 420 215
rect 363 144 371 178
rect 405 144 420 178
rect 363 131 420 144
rect 450 131 556 215
rect 503 93 556 131
rect 503 59 511 93
rect 545 59 556 93
rect 503 47 556 59
rect 586 190 642 215
rect 586 156 597 190
rect 631 156 642 190
rect 586 122 642 156
rect 586 88 597 122
rect 631 88 642 122
rect 586 47 642 88
rect 672 93 728 215
rect 672 59 683 93
rect 717 59 728 93
rect 672 47 728 59
rect 758 190 814 215
rect 758 156 769 190
rect 803 156 814 190
rect 758 122 814 156
rect 758 88 769 122
rect 803 88 814 122
rect 758 47 814 88
rect 844 203 897 215
rect 844 161 922 203
rect 844 127 855 161
rect 889 127 922 161
rect 844 119 922 127
rect 952 119 994 203
rect 1024 175 1080 203
rect 1024 141 1035 175
rect 1069 141 1080 175
rect 1024 119 1080 141
rect 1110 119 1152 203
rect 1182 140 1337 203
rect 1182 119 1209 140
rect 844 93 897 119
rect 844 59 855 93
rect 889 59 897 93
rect 844 47 897 59
rect 1197 106 1209 119
rect 1243 119 1337 140
rect 1367 119 1409 203
rect 1439 165 1495 203
rect 1439 131 1450 165
rect 1484 131 1495 165
rect 1439 119 1495 131
rect 1525 119 1589 203
rect 1619 165 1804 203
rect 1619 131 1630 165
rect 1664 131 1804 165
rect 1619 119 1804 131
rect 1834 191 1891 203
rect 1834 157 1849 191
rect 1883 157 1891 191
rect 1834 119 1891 157
rect 1243 106 1255 119
rect 1197 98 1255 106
<< pdiff >>
rect 27 516 84 530
rect 27 482 35 516
rect 69 482 84 516
rect 27 448 84 482
rect 27 414 35 448
rect 69 414 84 448
rect 27 402 84 414
rect 114 516 170 530
rect 114 482 125 516
rect 159 482 170 516
rect 114 448 170 482
rect 114 414 125 448
rect 159 414 170 448
rect 114 402 170 414
rect 200 518 253 530
rect 200 484 211 518
rect 245 484 253 518
rect 200 450 253 484
rect 469 579 526 587
rect 469 545 481 579
rect 515 545 526 579
rect 469 463 526 545
rect 200 416 211 450
rect 245 416 253 450
rect 200 402 253 416
rect 317 438 417 463
rect 317 404 329 438
rect 363 404 417 438
rect 317 396 417 404
rect 367 335 417 396
rect 447 335 526 463
rect 556 381 612 587
rect 556 347 567 381
rect 601 347 612 381
rect 556 335 612 347
rect 642 579 698 587
rect 642 545 653 579
rect 687 545 698 579
rect 642 335 698 545
rect 728 381 784 587
rect 728 347 739 381
rect 773 347 784 381
rect 728 335 784 347
rect 814 575 937 587
rect 814 541 895 575
rect 929 559 937 575
rect 929 541 969 559
rect 814 507 969 541
rect 814 473 895 507
rect 929 473 969 507
rect 814 431 969 473
rect 999 431 1041 559
rect 1071 538 1127 559
rect 1071 504 1082 538
rect 1116 504 1127 538
rect 1071 431 1127 504
rect 1157 547 1207 559
rect 1509 547 1559 559
rect 1157 431 1229 547
rect 814 335 937 431
rect 1179 419 1229 431
rect 1259 535 1373 547
rect 1259 501 1270 535
rect 1304 501 1373 535
rect 1259 419 1373 501
rect 1403 419 1445 547
rect 1475 536 1559 547
rect 1475 502 1486 536
rect 1520 502 1559 536
rect 1475 468 1559 502
rect 1475 434 1486 468
rect 1520 434 1559 468
rect 1475 431 1559 434
rect 1589 547 1639 559
rect 1589 431 1661 547
rect 1475 419 1532 431
rect 1611 419 1661 431
rect 1691 535 1747 547
rect 1691 501 1702 535
rect 1736 501 1747 535
rect 1691 419 1747 501
rect 1777 533 1830 547
rect 1777 499 1788 533
rect 1822 499 1830 533
rect 1777 465 1830 499
rect 1777 431 1788 465
rect 1822 431 1830 465
rect 1777 419 1830 431
<< ndiffc >>
rect 35 131 69 165
rect 125 131 159 165
rect 211 144 245 178
rect 371 144 405 178
rect 511 59 545 93
rect 597 156 631 190
rect 597 88 631 122
rect 683 59 717 93
rect 769 156 803 190
rect 769 88 803 122
rect 855 127 889 161
rect 1035 141 1069 175
rect 855 59 889 93
rect 1209 106 1243 140
rect 1450 131 1484 165
rect 1630 131 1664 165
rect 1849 157 1883 191
<< pdiffc >>
rect 35 482 69 516
rect 35 414 69 448
rect 125 482 159 516
rect 125 414 159 448
rect 211 484 245 518
rect 481 545 515 579
rect 211 416 245 450
rect 329 404 363 438
rect 567 347 601 381
rect 653 545 687 579
rect 739 347 773 381
rect 895 541 929 575
rect 895 473 929 507
rect 1082 504 1116 538
rect 1270 501 1304 535
rect 1486 502 1520 536
rect 1486 434 1520 468
rect 1702 501 1736 535
rect 1788 499 1822 533
rect 1788 431 1822 465
<< poly >>
rect 1127 615 1777 645
rect 526 587 556 613
rect 612 587 642 613
rect 698 587 728 613
rect 784 587 814 613
rect 84 530 114 556
rect 170 552 447 582
rect 170 530 200 552
rect 417 463 447 552
rect 84 307 114 402
rect 170 376 200 402
rect 269 348 335 364
rect 269 314 285 348
rect 319 314 335 348
rect 969 559 999 585
rect 1041 559 1071 585
rect 1127 559 1157 615
rect 1229 547 1259 573
rect 1373 547 1403 573
rect 1445 547 1475 573
rect 1559 559 1589 615
rect 269 307 335 314
rect 84 280 335 307
rect 417 303 447 335
rect 526 303 556 335
rect 612 303 642 335
rect 698 303 728 335
rect 784 303 814 335
rect 969 307 999 431
rect 1041 363 1071 431
rect 1127 405 1157 431
rect 1661 547 1691 573
rect 1747 547 1777 615
rect 1229 382 1259 419
rect 1373 382 1403 419
rect 1229 366 1295 382
rect 1041 347 1171 363
rect 1041 333 1121 347
rect 84 277 285 280
rect 84 203 114 229
rect 170 203 200 277
rect 269 246 285 277
rect 319 246 335 280
rect 269 230 335 246
rect 399 287 465 303
rect 399 253 415 287
rect 449 253 465 287
rect 399 237 465 253
rect 526 287 814 303
rect 526 253 542 287
rect 576 253 610 287
rect 644 253 678 287
rect 712 267 814 287
rect 886 287 999 307
rect 712 253 844 267
rect 526 237 844 253
rect 886 253 902 287
rect 936 277 999 287
rect 1080 313 1121 333
rect 1155 313 1171 347
rect 1080 297 1171 313
rect 1229 332 1245 366
rect 1279 332 1295 366
rect 1229 316 1295 332
rect 1337 366 1403 382
rect 1337 332 1353 366
rect 1387 332 1403 366
rect 1337 316 1403 332
rect 1445 359 1475 419
rect 1559 405 1589 431
rect 1661 363 1691 419
rect 1445 343 1547 359
rect 1445 329 1497 343
rect 936 253 952 277
rect 886 237 952 253
rect 420 215 450 237
rect 556 215 586 237
rect 642 215 672 237
rect 728 215 758 237
rect 814 215 844 237
rect 84 51 114 119
rect 170 93 200 119
rect 420 51 450 131
rect 84 21 450 51
rect 922 203 952 237
rect 994 203 1024 229
rect 1080 203 1110 297
rect 1229 255 1259 316
rect 1152 225 1259 255
rect 1152 203 1182 225
rect 1337 203 1367 316
rect 1481 309 1497 329
rect 1531 309 1547 343
rect 1603 347 1691 363
rect 1603 327 1619 347
rect 1481 275 1547 309
rect 1481 241 1497 275
rect 1531 241 1547 275
rect 1409 203 1439 229
rect 1481 225 1547 241
rect 1589 313 1619 327
rect 1653 313 1691 347
rect 1589 297 1691 313
rect 1747 359 1777 419
rect 1747 343 1834 359
rect 1747 309 1763 343
rect 1797 309 1834 343
rect 1495 203 1525 225
rect 1589 203 1619 297
rect 1747 275 1834 309
rect 1747 241 1763 275
rect 1797 241 1834 275
rect 1747 225 1834 241
rect 1804 203 1834 225
rect 922 93 952 119
rect 994 51 1024 119
rect 1080 93 1110 119
rect 1152 93 1182 119
rect 1337 93 1367 119
rect 1409 51 1439 119
rect 1495 93 1525 119
rect 1589 93 1619 119
rect 1804 51 1834 119
rect 556 21 586 47
rect 642 21 672 47
rect 728 21 758 47
rect 814 21 844 47
rect 994 21 1834 51
<< polycont >>
rect 285 314 319 348
rect 285 246 319 280
rect 415 253 449 287
rect 542 253 576 287
rect 610 253 644 287
rect 678 253 712 287
rect 902 253 936 287
rect 1121 313 1155 347
rect 1245 332 1279 366
rect 1353 332 1387 366
rect 1497 309 1531 343
rect 1497 241 1531 275
rect 1619 313 1653 347
rect 1763 309 1797 343
rect 1763 241 1797 275
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 465 579 531 649
rect 465 545 481 579
rect 515 545 531 579
rect 637 579 703 649
rect 637 545 653 579
rect 687 545 703 579
rect 879 575 945 649
rect 879 541 895 575
rect 929 541 945 575
rect 31 516 73 532
rect 31 482 35 516
rect 69 482 73 516
rect 31 448 73 482
rect 31 414 35 448
rect 69 414 73 448
rect 31 165 73 414
rect 31 131 35 165
rect 69 131 73 165
rect 31 128 73 131
rect 65 94 73 128
rect 121 516 159 532
rect 121 482 125 516
rect 121 448 159 482
rect 121 414 125 448
rect 121 165 159 414
rect 121 131 125 165
rect 121 92 159 131
rect 207 518 249 534
rect 207 484 211 518
rect 245 508 249 518
rect 245 484 843 508
rect 207 474 843 484
rect 207 450 249 474
rect 207 416 211 450
rect 245 416 249 450
rect 207 178 249 416
rect 313 404 329 438
rect 363 404 379 438
rect 809 433 843 474
rect 879 507 945 541
rect 879 473 895 507
rect 929 473 945 507
rect 879 469 945 473
rect 981 538 1120 554
rect 981 504 1082 538
rect 1116 504 1120 538
rect 981 488 1120 504
rect 1254 535 1320 649
rect 1254 501 1270 535
rect 1304 501 1320 535
rect 1254 497 1320 501
rect 1482 536 1524 552
rect 1482 502 1486 536
rect 1520 502 1524 536
rect 981 433 1015 488
rect 1482 468 1524 502
rect 1482 452 1486 468
rect 313 364 379 404
rect 285 348 379 364
rect 319 314 379 348
rect 285 280 379 314
rect 319 246 379 280
rect 285 230 379 246
rect 415 287 449 424
rect 809 399 1015 433
rect 563 381 773 397
rect 563 347 567 381
rect 601 347 739 381
rect 773 347 833 363
rect 563 329 833 347
rect 415 237 449 253
rect 523 253 542 287
rect 576 253 610 287
rect 644 253 678 287
rect 712 253 728 287
rect 207 144 211 178
rect 245 144 249 178
rect 207 128 249 144
rect 345 194 379 230
rect 523 201 557 253
rect 773 242 833 329
rect 895 287 936 350
rect 895 253 902 287
rect 773 206 807 242
rect 895 237 936 253
rect 345 178 405 194
rect 345 144 371 178
rect 345 128 405 144
rect 441 167 557 201
rect 593 190 807 206
rect 441 92 475 167
rect 593 156 597 190
rect 631 172 769 190
rect 631 156 635 172
rect 593 122 635 156
rect 121 58 475 92
rect 511 93 549 109
rect 545 59 549 93
rect 593 88 597 122
rect 631 88 635 122
rect 765 156 769 172
rect 803 156 807 190
rect 981 191 1015 399
rect 1051 434 1486 452
rect 1520 434 1524 468
rect 1051 418 1524 434
rect 1051 261 1085 418
rect 1245 366 1313 382
rect 1121 347 1209 363
rect 1155 313 1209 347
rect 1279 332 1313 366
rect 1245 316 1313 332
rect 1353 366 1409 382
rect 1387 332 1409 366
rect 1353 316 1409 332
rect 1497 343 1531 359
rect 1121 297 1209 313
rect 1175 280 1209 297
rect 1497 280 1531 309
rect 1567 347 1653 572
rect 1698 535 1740 649
rect 1698 501 1702 535
rect 1736 501 1740 535
rect 1698 485 1740 501
rect 1784 533 1826 549
rect 1784 499 1788 533
rect 1822 499 1826 533
rect 1784 465 1826 499
rect 1784 431 1788 465
rect 1822 431 1826 465
rect 1784 429 1826 431
rect 1567 313 1619 347
rect 1567 297 1653 313
rect 1689 395 1899 429
rect 1175 275 1531 280
rect 1051 227 1139 261
rect 1175 246 1497 275
rect 1105 210 1139 227
rect 1689 259 1723 395
rect 1531 241 1723 259
rect 1497 225 1723 241
rect 1759 343 1797 359
rect 1759 309 1763 343
rect 1759 275 1797 309
rect 1759 241 1763 275
rect 765 122 807 156
rect 593 72 635 88
rect 679 93 721 109
rect 511 17 549 59
rect 679 59 683 93
rect 717 59 721 93
rect 765 88 769 122
rect 803 88 807 122
rect 765 72 807 88
rect 851 161 893 177
rect 851 127 855 161
rect 889 127 893 161
rect 851 93 893 127
rect 981 175 1069 191
rect 1105 181 1329 210
rect 1105 176 1505 181
rect 981 141 1035 175
rect 1295 165 1505 176
rect 1295 147 1450 165
rect 981 125 1069 141
rect 679 17 721 59
rect 851 59 855 93
rect 889 59 893 93
rect 851 17 893 59
rect 1193 106 1209 140
rect 1243 106 1259 140
rect 1193 17 1259 106
rect 1446 131 1450 147
rect 1484 131 1505 165
rect 1446 128 1505 131
rect 1446 94 1471 128
rect 1614 165 1680 169
rect 1614 131 1630 165
rect 1664 131 1680 165
rect 1614 17 1680 131
rect 1759 94 1797 241
rect 1833 191 1899 395
rect 1833 157 1849 191
rect 1883 157 1899 191
rect 1833 153 1899 157
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 94 65 128
rect 1471 94 1505 128
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 19 128 77 134
rect 19 94 31 128
rect 65 125 77 128
rect 1459 128 1517 134
rect 1459 125 1471 128
rect 65 97 1471 125
rect 65 94 77 97
rect 19 88 77 94
rect 1459 94 1471 97
rect 1505 94 1517 128
rect 1459 88 1517 94
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux4_4
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 1759 94 1793 128 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 1759 168 1793 202 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 1759 316 1793 350 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1536282
string GDS_START 1522208
<< end >>
