magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
rect 296 325 1760 331
rect 296 273 494 325
<< pwell >>
rect 1747 241 2015 247
rect 1 157 433 221
rect 1020 157 2015 241
rect 1 49 2015 157
rect 0 0 2016 49
<< scnmos >>
rect 84 111 114 195
rect 156 111 186 195
rect 242 111 272 195
rect 320 111 350 195
rect 526 47 556 131
rect 604 47 634 131
rect 690 47 720 131
rect 768 47 798 131
rect 870 47 900 131
rect 978 47 1008 131
rect 1103 47 1133 215
rect 1175 47 1205 215
rect 1373 47 1403 215
rect 1445 47 1475 215
rect 1554 131 1584 215
rect 1632 131 1662 215
rect 1830 53 1860 221
rect 1902 53 1932 221
<< scpmoshvt >>
rect 82 481 112 609
rect 154 481 184 609
rect 248 481 278 609
rect 320 481 350 609
rect 537 475 567 603
rect 609 475 639 603
rect 711 475 741 603
rect 789 475 819 603
rect 897 519 927 603
rect 975 519 1005 603
rect 1122 361 1152 613
rect 1194 361 1224 613
rect 1388 361 1418 613
rect 1460 361 1490 613
rect 1567 361 1597 489
rect 1639 361 1669 489
rect 1833 367 1863 619
rect 1905 367 1935 619
<< ndiff >>
rect 27 170 84 195
rect 27 136 39 170
rect 73 136 84 170
rect 27 111 84 136
rect 114 111 156 195
rect 186 170 242 195
rect 186 136 197 170
rect 231 136 242 170
rect 186 111 242 136
rect 272 111 320 195
rect 350 170 407 195
rect 350 136 361 170
rect 395 136 407 170
rect 350 111 407 136
rect 1046 203 1103 215
rect 1046 169 1058 203
rect 1092 169 1103 203
rect 1046 131 1103 169
rect 469 111 526 131
rect 469 77 481 111
rect 515 77 526 111
rect 469 47 526 77
rect 556 47 604 131
rect 634 103 690 131
rect 634 69 645 103
rect 679 69 690 103
rect 634 47 690 69
rect 720 47 768 131
rect 798 103 870 131
rect 798 69 825 103
rect 859 69 870 103
rect 798 47 870 69
rect 900 47 978 131
rect 1008 93 1103 131
rect 1008 59 1058 93
rect 1092 59 1103 93
rect 1008 47 1103 59
rect 1133 47 1175 215
rect 1205 203 1262 215
rect 1205 169 1216 203
rect 1250 169 1262 203
rect 1205 103 1262 169
rect 1205 69 1216 103
rect 1250 69 1262 103
rect 1205 47 1262 69
rect 1316 203 1373 215
rect 1316 169 1328 203
rect 1362 169 1373 203
rect 1316 103 1373 169
rect 1316 69 1328 103
rect 1362 69 1373 103
rect 1316 47 1373 69
rect 1403 47 1445 215
rect 1475 131 1554 215
rect 1584 131 1632 215
rect 1662 190 1719 215
rect 1662 156 1673 190
rect 1707 156 1719 190
rect 1662 131 1719 156
rect 1773 209 1830 221
rect 1773 175 1785 209
rect 1819 175 1830 209
rect 1475 113 1532 131
rect 1475 79 1486 113
rect 1520 79 1532 113
rect 1475 47 1532 79
rect 1773 99 1830 175
rect 1773 65 1785 99
rect 1819 65 1830 99
rect 1773 53 1830 65
rect 1860 53 1902 221
rect 1932 209 1989 221
rect 1932 175 1943 209
rect 1977 175 1989 209
rect 1932 103 1989 175
rect 1932 69 1943 103
rect 1977 69 1989 103
rect 1932 53 1989 69
<< pdiff >>
rect 27 597 82 609
rect 27 563 37 597
rect 71 563 82 597
rect 27 527 82 563
rect 27 493 37 527
rect 71 493 82 527
rect 27 481 82 493
rect 112 481 154 609
rect 184 597 248 609
rect 184 563 195 597
rect 229 563 248 597
rect 184 481 248 563
rect 278 481 320 609
rect 350 481 428 609
rect 1067 603 1122 613
rect 372 355 428 481
rect 482 524 537 603
rect 482 490 492 524
rect 526 490 537 524
rect 482 475 537 490
rect 567 475 609 603
rect 639 558 711 603
rect 639 524 666 558
rect 700 524 711 558
rect 639 475 711 524
rect 741 475 789 603
rect 819 578 897 603
rect 819 544 830 578
rect 864 544 897 578
rect 819 519 897 544
rect 927 519 975 603
rect 1005 580 1122 603
rect 1005 546 1077 580
rect 1111 546 1122 580
rect 1005 519 1122 546
rect 819 475 875 519
rect 372 321 384 355
rect 418 321 428 355
rect 372 309 428 321
rect 1067 361 1122 519
rect 1152 361 1194 613
rect 1224 597 1279 613
rect 1224 563 1235 597
rect 1269 563 1279 597
rect 1224 502 1279 563
rect 1224 468 1235 502
rect 1269 468 1279 502
rect 1224 407 1279 468
rect 1224 373 1235 407
rect 1269 373 1279 407
rect 1224 361 1279 373
rect 1333 597 1388 613
rect 1333 563 1343 597
rect 1377 563 1388 597
rect 1333 502 1388 563
rect 1333 468 1343 502
rect 1377 468 1388 502
rect 1333 407 1388 468
rect 1333 373 1343 407
rect 1377 373 1388 407
rect 1333 361 1388 373
rect 1418 361 1460 613
rect 1490 601 1545 613
rect 1490 567 1501 601
rect 1535 567 1545 601
rect 1490 489 1545 567
rect 1778 607 1833 619
rect 1778 573 1788 607
rect 1822 573 1833 607
rect 1778 510 1833 573
rect 1490 477 1567 489
rect 1490 443 1501 477
rect 1535 443 1567 477
rect 1490 361 1567 443
rect 1597 361 1639 489
rect 1669 477 1724 489
rect 1669 443 1680 477
rect 1714 443 1724 477
rect 1669 407 1724 443
rect 1669 373 1680 407
rect 1714 373 1724 407
rect 1669 361 1724 373
rect 1778 476 1788 510
rect 1822 476 1833 510
rect 1778 413 1833 476
rect 1778 379 1788 413
rect 1822 379 1833 413
rect 1778 367 1833 379
rect 1863 367 1905 619
rect 1935 597 1989 619
rect 1935 563 1946 597
rect 1980 563 1989 597
rect 1935 505 1989 563
rect 1935 471 1946 505
rect 1980 471 1989 505
rect 1935 413 1989 471
rect 1935 379 1946 413
rect 1980 379 1989 413
rect 1935 367 1989 379
<< ndiffc >>
rect 39 136 73 170
rect 197 136 231 170
rect 361 136 395 170
rect 1058 169 1092 203
rect 481 77 515 111
rect 645 69 679 103
rect 825 69 859 103
rect 1058 59 1092 93
rect 1216 169 1250 203
rect 1216 69 1250 103
rect 1328 169 1362 203
rect 1328 69 1362 103
rect 1673 156 1707 190
rect 1785 175 1819 209
rect 1486 79 1520 113
rect 1785 65 1819 99
rect 1943 175 1977 209
rect 1943 69 1977 103
<< pdiffc >>
rect 37 563 71 597
rect 37 493 71 527
rect 195 563 229 597
rect 492 490 526 524
rect 666 524 700 558
rect 830 544 864 578
rect 1077 546 1111 580
rect 384 321 418 355
rect 1235 563 1269 597
rect 1235 468 1269 502
rect 1235 373 1269 407
rect 1343 563 1377 597
rect 1343 468 1377 502
rect 1343 373 1377 407
rect 1501 567 1535 601
rect 1788 573 1822 607
rect 1501 443 1535 477
rect 1680 443 1714 477
rect 1680 373 1714 407
rect 1788 476 1822 510
rect 1788 379 1822 413
rect 1946 563 1980 597
rect 1946 471 1980 505
rect 1946 379 1980 413
<< poly >>
rect 82 609 112 635
rect 154 609 184 635
rect 248 609 278 635
rect 320 609 350 635
rect 537 603 567 629
rect 609 603 639 629
rect 711 603 741 629
rect 789 603 819 629
rect 897 603 927 629
rect 975 603 1005 629
rect 1122 613 1152 639
rect 1194 613 1224 639
rect 1388 613 1418 639
rect 1460 613 1490 639
rect 1833 619 1863 645
rect 1905 619 1935 645
rect 82 370 112 481
rect 154 370 184 481
rect 248 439 278 481
rect 320 439 350 481
rect 82 354 184 370
rect 82 340 130 354
rect 84 320 130 340
rect 164 320 184 354
rect 84 286 184 320
rect 226 423 350 439
rect 226 389 242 423
rect 276 389 350 423
rect 226 355 350 389
rect 226 321 242 355
rect 276 321 350 355
rect 226 305 350 321
rect 537 447 567 475
rect 526 417 567 447
rect 526 369 556 417
rect 609 369 639 475
rect 711 439 741 475
rect 681 423 747 439
rect 681 389 697 423
rect 731 389 747 423
rect 681 373 747 389
rect 789 433 819 475
rect 789 417 855 433
rect 789 383 805 417
rect 839 383 855 417
rect 526 353 639 369
rect 526 319 542 353
rect 576 319 639 353
rect 84 252 130 286
rect 164 257 184 286
rect 164 252 186 257
rect 84 227 186 252
rect 84 195 114 227
rect 156 195 186 227
rect 242 195 272 305
rect 320 195 350 305
rect 526 285 639 319
rect 684 319 714 373
rect 789 367 855 383
rect 684 289 720 319
rect 897 309 927 519
rect 975 473 1005 519
rect 969 457 1035 473
rect 969 423 985 457
rect 1019 423 1035 457
rect 969 407 1035 423
rect 526 251 542 285
rect 576 251 639 285
rect 526 235 639 251
rect 526 131 556 235
rect 604 131 634 235
rect 690 131 720 289
rect 762 279 927 309
rect 762 215 828 279
rect 762 181 778 215
rect 812 181 828 215
rect 762 165 828 181
rect 870 215 936 231
rect 870 181 886 215
rect 920 181 936 215
rect 870 165 936 181
rect 768 131 798 165
rect 870 131 900 165
rect 978 131 1008 407
rect 1567 489 1597 515
rect 1639 489 1669 515
rect 1122 321 1152 361
rect 1194 321 1224 361
rect 1388 321 1418 361
rect 1460 321 1490 361
rect 1567 321 1597 361
rect 1122 305 1224 321
rect 1122 285 1144 305
rect 1103 271 1144 285
rect 1178 285 1224 305
rect 1323 305 1597 321
rect 1178 271 1275 285
rect 1103 255 1275 271
rect 1323 271 1339 305
rect 1373 271 1407 305
rect 1441 271 1475 305
rect 1509 291 1597 305
rect 1639 291 1669 361
rect 1833 327 1863 367
rect 1905 327 1935 367
rect 1509 271 1669 291
rect 1323 261 1669 271
rect 1825 311 1935 327
rect 1825 277 1841 311
rect 1875 277 1935 311
rect 1825 261 1935 277
rect 1323 255 1584 261
rect 1103 215 1133 255
rect 1175 215 1205 255
rect 1373 215 1403 255
rect 1445 215 1475 255
rect 1554 215 1584 255
rect 1632 215 1662 261
rect 1830 221 1860 261
rect 1902 221 1932 261
rect 84 85 114 111
rect 156 85 186 111
rect 242 85 272 111
rect 320 85 350 111
rect 1554 105 1584 131
rect 1632 105 1662 131
rect 526 21 556 47
rect 604 21 634 47
rect 690 21 720 47
rect 768 21 798 47
rect 870 21 900 47
rect 978 21 1008 47
rect 1103 21 1133 47
rect 1175 21 1205 47
rect 1373 21 1403 47
rect 1445 21 1475 47
rect 1830 27 1860 53
rect 1902 27 1932 53
<< polycont >>
rect 130 320 164 354
rect 242 389 276 423
rect 242 321 276 355
rect 697 389 731 423
rect 805 383 839 417
rect 542 319 576 353
rect 130 252 164 286
rect 985 423 1019 457
rect 542 251 576 285
rect 778 181 812 215
rect 886 181 920 215
rect 1144 271 1178 305
rect 1339 271 1373 305
rect 1407 271 1441 305
rect 1475 271 1509 305
rect 1841 277 1875 311
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 21 597 87 613
rect 21 563 37 597
rect 71 563 87 597
rect 21 527 87 563
rect 179 597 245 649
rect 179 563 195 597
rect 229 563 245 597
rect 179 547 245 563
rect 281 579 614 613
rect 21 493 37 527
rect 71 511 87 527
rect 281 511 315 579
rect 71 493 315 511
rect 21 477 315 493
rect 476 524 542 543
rect 476 490 492 524
rect 526 490 542 524
rect 21 199 55 477
rect 476 441 542 490
rect 114 354 180 430
rect 114 320 130 354
rect 164 320 180 354
rect 114 286 180 320
rect 217 423 278 439
rect 217 389 242 423
rect 276 389 278 423
rect 217 355 278 389
rect 217 321 242 355
rect 276 321 278 355
rect 217 305 278 321
rect 314 407 542 441
rect 580 439 614 579
rect 650 558 716 649
rect 650 524 666 558
rect 700 524 716 558
rect 650 475 716 524
rect 814 578 880 607
rect 814 544 830 578
rect 864 549 880 578
rect 1061 580 1127 649
rect 864 544 925 549
rect 814 515 925 544
rect 580 423 747 439
rect 114 252 130 286
rect 164 252 180 286
rect 314 269 348 407
rect 580 405 697 423
rect 681 389 697 405
rect 731 389 747 423
rect 681 373 747 389
rect 789 417 855 433
rect 789 383 805 417
rect 839 383 855 417
rect 114 236 180 252
rect 275 235 348 269
rect 384 369 434 371
rect 384 355 592 369
rect 418 353 592 355
rect 418 321 542 353
rect 384 319 542 321
rect 576 319 592 353
rect 384 305 592 319
rect 21 170 89 199
rect 21 136 39 170
rect 73 136 89 170
rect 21 107 89 136
rect 181 170 231 199
rect 181 136 197 170
rect 181 17 231 136
rect 275 87 309 235
rect 384 199 418 305
rect 526 301 592 305
rect 789 301 855 383
rect 891 371 925 515
rect 1061 546 1077 580
rect 1111 546 1127 580
rect 1061 509 1127 546
rect 1219 597 1285 613
rect 1219 563 1235 597
rect 1269 563 1285 597
rect 1219 502 1285 563
rect 1219 473 1235 502
rect 969 468 1235 473
rect 1269 468 1285 502
rect 969 457 1285 468
rect 969 423 985 457
rect 1019 423 1285 457
rect 969 407 1285 423
rect 1219 373 1235 407
rect 1269 373 1285 407
rect 891 337 1006 371
rect 1219 357 1285 373
rect 1327 597 1393 613
rect 1327 563 1343 597
rect 1377 563 1393 597
rect 1327 502 1393 563
rect 1327 468 1343 502
rect 1377 468 1393 502
rect 1327 407 1393 468
rect 1485 601 1551 649
rect 1485 567 1501 601
rect 1535 567 1551 601
rect 1485 477 1551 567
rect 1772 607 1838 649
rect 1772 573 1788 607
rect 1822 573 1838 607
rect 1772 510 1838 573
rect 1485 443 1501 477
rect 1535 443 1551 477
rect 1485 427 1551 443
rect 1657 477 1730 493
rect 1657 443 1680 477
rect 1714 443 1730 477
rect 1327 373 1343 407
rect 1377 391 1393 407
rect 1657 407 1730 443
rect 1377 373 1607 391
rect 1327 357 1607 373
rect 972 321 1006 337
rect 1232 321 1285 357
rect 972 305 1194 321
rect 526 285 904 301
rect 526 251 542 285
rect 576 267 904 285
rect 576 251 592 267
rect 526 235 592 251
rect 870 231 904 267
rect 972 271 1144 305
rect 1178 271 1194 305
rect 972 255 1194 271
rect 1232 305 1525 321
rect 1232 271 1339 305
rect 1373 271 1407 305
rect 1441 271 1475 305
rect 1509 271 1525 305
rect 1232 255 1525 271
rect 762 215 828 231
rect 762 199 778 215
rect 345 170 418 199
rect 345 136 361 170
rect 395 136 418 170
rect 345 123 418 136
rect 465 181 778 199
rect 812 181 828 215
rect 465 165 828 181
rect 870 215 936 231
rect 870 181 886 215
rect 920 181 936 215
rect 870 165 936 181
rect 465 111 531 165
rect 972 129 1006 255
rect 1232 219 1266 255
rect 1561 219 1607 357
rect 465 87 481 111
rect 275 77 481 87
rect 515 77 531 111
rect 275 53 531 77
rect 629 103 695 129
rect 629 69 645 103
rect 679 69 695 103
rect 629 17 695 69
rect 809 103 1006 129
rect 809 69 825 103
rect 859 69 1006 103
rect 809 59 1006 69
rect 1042 203 1108 219
rect 1042 169 1058 203
rect 1092 169 1108 203
rect 1042 93 1108 169
rect 1042 59 1058 93
rect 1092 59 1108 93
rect 1042 17 1108 59
rect 1200 203 1266 219
rect 1200 169 1216 203
rect 1250 169 1266 203
rect 1200 103 1266 169
rect 1200 69 1216 103
rect 1250 69 1266 103
rect 1200 53 1266 69
rect 1312 203 1607 219
rect 1312 169 1328 203
rect 1362 185 1607 203
rect 1657 373 1680 407
rect 1714 373 1730 407
rect 1657 327 1730 373
rect 1772 476 1788 510
rect 1822 476 1838 510
rect 1772 413 1838 476
rect 1772 379 1788 413
rect 1822 379 1838 413
rect 1772 363 1838 379
rect 1927 597 1996 613
rect 1927 563 1946 597
rect 1980 563 1996 597
rect 1927 505 1996 563
rect 1927 471 1946 505
rect 1980 471 1996 505
rect 1927 413 1996 471
rect 1927 379 1946 413
rect 1980 379 1996 413
rect 1657 311 1891 327
rect 1657 277 1841 311
rect 1875 277 1891 311
rect 1657 261 1891 277
rect 1657 190 1723 261
rect 1362 169 1378 185
rect 1312 103 1378 169
rect 1657 156 1673 190
rect 1707 156 1723 190
rect 1312 69 1328 103
rect 1362 69 1378 103
rect 1312 53 1378 69
rect 1470 113 1536 149
rect 1657 127 1723 156
rect 1769 209 1835 225
rect 1769 175 1785 209
rect 1819 175 1835 209
rect 1470 79 1486 113
rect 1520 79 1536 113
rect 1470 17 1536 79
rect 1769 99 1835 175
rect 1769 65 1785 99
rect 1819 65 1835 99
rect 1769 17 1835 65
rect 1927 209 1996 379
rect 1927 175 1943 209
rect 1977 175 1996 209
rect 1927 103 1996 175
rect 1927 69 1943 103
rect 1977 69 1996 103
rect 1927 53 1996 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlxbp_lp
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1951 94 1985 128 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 168 1985 202 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 390 1985 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 464 1985 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 538 1985 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2307856
string GDS_START 2293500
<< end >>
