magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 18 243 1177 259
rect 18 49 1625 243
rect 0 0 1632 49
<< scnmos >>
rect 97 65 127 233
rect 251 65 281 233
rect 337 65 367 233
rect 423 65 453 233
rect 517 65 547 233
rect 607 65 637 233
rect 780 65 810 233
rect 880 65 910 233
rect 966 65 996 233
rect 1053 65 1083 233
rect 1258 49 1288 217
rect 1344 49 1374 217
rect 1430 49 1460 217
rect 1516 49 1546 217
<< scpmoshvt >>
rect 165 367 195 619
rect 251 367 281 619
rect 337 367 367 619
rect 431 367 461 619
rect 517 367 547 619
rect 603 367 633 619
rect 793 367 823 619
rect 880 367 910 619
rect 966 367 996 619
rect 1052 367 1082 619
rect 1258 367 1288 619
rect 1344 367 1374 619
rect 1430 367 1460 619
rect 1516 367 1546 619
<< ndiff >>
rect 44 221 97 233
rect 44 187 52 221
rect 86 187 97 221
rect 44 111 97 187
rect 44 77 52 111
rect 86 77 97 111
rect 44 65 97 77
rect 127 183 251 233
rect 127 149 138 183
rect 172 149 251 183
rect 127 124 251 149
rect 127 107 206 124
rect 127 73 138 107
rect 172 90 206 107
rect 240 90 251 124
rect 172 73 251 90
rect 127 65 251 73
rect 281 175 337 233
rect 281 141 292 175
rect 326 141 337 175
rect 281 107 337 141
rect 281 73 292 107
rect 326 73 337 107
rect 281 65 337 73
rect 367 136 423 233
rect 367 102 378 136
rect 412 102 423 136
rect 367 65 423 102
rect 453 179 517 233
rect 453 145 470 179
rect 504 145 517 179
rect 453 111 517 145
rect 453 77 470 111
rect 504 77 517 111
rect 453 65 517 77
rect 547 136 607 233
rect 547 102 562 136
rect 596 102 607 136
rect 547 65 607 102
rect 637 192 780 233
rect 637 158 662 192
rect 696 158 735 192
rect 769 158 780 192
rect 637 111 780 158
rect 637 77 662 111
rect 696 77 735 111
rect 769 77 780 111
rect 637 65 780 77
rect 810 221 880 233
rect 810 187 821 221
rect 855 187 880 221
rect 810 153 880 187
rect 810 119 821 153
rect 855 119 880 153
rect 810 65 880 119
rect 910 124 966 233
rect 910 90 921 124
rect 955 90 966 124
rect 910 65 966 90
rect 996 225 1053 233
rect 996 191 1007 225
rect 1041 191 1053 225
rect 996 157 1053 191
rect 996 123 1007 157
rect 1041 123 1053 157
rect 996 65 1053 123
rect 1083 179 1151 233
rect 1083 145 1109 179
rect 1143 145 1151 179
rect 1083 111 1151 145
rect 1083 77 1109 111
rect 1143 77 1151 111
rect 1083 65 1151 77
rect 1205 181 1258 217
rect 1205 147 1213 181
rect 1247 147 1258 181
rect 1205 95 1258 147
rect 1205 61 1213 95
rect 1247 61 1258 95
rect 1205 49 1258 61
rect 1288 205 1344 217
rect 1288 171 1299 205
rect 1333 171 1344 205
rect 1288 101 1344 171
rect 1288 67 1299 101
rect 1333 67 1344 101
rect 1288 49 1344 67
rect 1374 177 1430 217
rect 1374 143 1385 177
rect 1419 143 1430 177
rect 1374 91 1430 143
rect 1374 57 1385 91
rect 1419 57 1430 91
rect 1374 49 1430 57
rect 1460 205 1516 217
rect 1460 171 1471 205
rect 1505 171 1516 205
rect 1460 101 1516 171
rect 1460 67 1471 101
rect 1505 67 1516 101
rect 1460 49 1516 67
rect 1546 177 1599 217
rect 1546 143 1557 177
rect 1591 143 1599 177
rect 1546 95 1599 143
rect 1546 61 1557 95
rect 1591 61 1599 95
rect 1546 49 1599 61
<< pdiff >>
rect 112 597 165 619
rect 112 563 120 597
rect 154 563 165 597
rect 112 521 165 563
rect 112 487 120 521
rect 154 487 165 521
rect 112 441 165 487
rect 112 407 120 441
rect 154 407 165 441
rect 112 367 165 407
rect 195 599 251 619
rect 195 565 206 599
rect 240 565 251 599
rect 195 509 251 565
rect 195 475 206 509
rect 240 475 251 509
rect 195 367 251 475
rect 281 585 337 619
rect 281 551 292 585
rect 326 551 337 585
rect 281 367 337 551
rect 367 599 431 619
rect 367 565 386 599
rect 420 565 431 599
rect 367 509 431 565
rect 367 475 386 509
rect 420 475 431 509
rect 367 367 431 475
rect 461 599 517 619
rect 461 565 472 599
rect 506 565 517 599
rect 461 507 517 565
rect 461 473 472 507
rect 506 473 517 507
rect 461 413 517 473
rect 461 379 472 413
rect 506 379 517 413
rect 461 367 517 379
rect 547 599 603 619
rect 547 565 558 599
rect 592 565 603 599
rect 547 522 603 565
rect 547 488 558 522
rect 592 488 603 522
rect 547 443 603 488
rect 547 409 558 443
rect 592 409 603 443
rect 547 367 603 409
rect 633 531 686 619
rect 633 497 644 531
rect 678 497 686 531
rect 633 413 686 497
rect 633 379 644 413
rect 678 379 686 413
rect 633 367 686 379
rect 740 599 793 619
rect 740 565 748 599
rect 782 565 793 599
rect 740 521 793 565
rect 740 487 748 521
rect 782 487 793 521
rect 740 441 793 487
rect 740 407 748 441
rect 782 407 793 441
rect 740 367 793 407
rect 823 599 880 619
rect 823 565 834 599
rect 868 565 880 599
rect 823 509 880 565
rect 823 475 834 509
rect 868 475 880 509
rect 823 367 880 475
rect 910 584 966 619
rect 910 550 921 584
rect 955 550 966 584
rect 910 367 966 550
rect 996 599 1052 619
rect 996 565 1007 599
rect 1041 565 1052 599
rect 996 509 1052 565
rect 996 475 1007 509
rect 1041 475 1052 509
rect 996 367 1052 475
rect 1082 599 1135 619
rect 1082 565 1093 599
rect 1127 565 1135 599
rect 1082 520 1135 565
rect 1082 486 1093 520
rect 1127 486 1135 520
rect 1082 441 1135 486
rect 1082 407 1093 441
rect 1127 407 1135 441
rect 1082 367 1135 407
rect 1205 607 1258 619
rect 1205 573 1213 607
rect 1247 573 1258 607
rect 1205 512 1258 573
rect 1205 478 1213 512
rect 1247 478 1258 512
rect 1205 367 1258 478
rect 1288 599 1344 619
rect 1288 565 1299 599
rect 1333 565 1344 599
rect 1288 511 1344 565
rect 1288 477 1299 511
rect 1333 477 1344 511
rect 1288 413 1344 477
rect 1288 379 1299 413
rect 1333 379 1344 413
rect 1288 367 1344 379
rect 1374 607 1430 619
rect 1374 573 1385 607
rect 1419 573 1430 607
rect 1374 528 1430 573
rect 1374 494 1385 528
rect 1419 494 1430 528
rect 1374 453 1430 494
rect 1374 419 1385 453
rect 1419 419 1430 453
rect 1374 367 1430 419
rect 1460 599 1516 619
rect 1460 565 1471 599
rect 1505 565 1516 599
rect 1460 511 1516 565
rect 1460 477 1471 511
rect 1505 477 1516 511
rect 1460 413 1516 477
rect 1460 379 1471 413
rect 1505 379 1516 413
rect 1460 367 1516 379
rect 1546 607 1599 619
rect 1546 573 1557 607
rect 1591 573 1599 607
rect 1546 528 1599 573
rect 1546 494 1557 528
rect 1591 494 1599 528
rect 1546 453 1599 494
rect 1546 419 1557 453
rect 1591 419 1599 453
rect 1546 367 1599 419
<< ndiffc >>
rect 52 187 86 221
rect 52 77 86 111
rect 138 149 172 183
rect 138 73 172 107
rect 206 90 240 124
rect 292 141 326 175
rect 292 73 326 107
rect 378 102 412 136
rect 470 145 504 179
rect 470 77 504 111
rect 562 102 596 136
rect 662 158 696 192
rect 735 158 769 192
rect 662 77 696 111
rect 735 77 769 111
rect 821 187 855 221
rect 821 119 855 153
rect 921 90 955 124
rect 1007 191 1041 225
rect 1007 123 1041 157
rect 1109 145 1143 179
rect 1109 77 1143 111
rect 1213 147 1247 181
rect 1213 61 1247 95
rect 1299 171 1333 205
rect 1299 67 1333 101
rect 1385 143 1419 177
rect 1385 57 1419 91
rect 1471 171 1505 205
rect 1471 67 1505 101
rect 1557 143 1591 177
rect 1557 61 1591 95
<< pdiffc >>
rect 120 563 154 597
rect 120 487 154 521
rect 120 407 154 441
rect 206 565 240 599
rect 206 475 240 509
rect 292 551 326 585
rect 386 565 420 599
rect 386 475 420 509
rect 472 565 506 599
rect 472 473 506 507
rect 472 379 506 413
rect 558 565 592 599
rect 558 488 592 522
rect 558 409 592 443
rect 644 497 678 531
rect 644 379 678 413
rect 748 565 782 599
rect 748 487 782 521
rect 748 407 782 441
rect 834 565 868 599
rect 834 475 868 509
rect 921 550 955 584
rect 1007 565 1041 599
rect 1007 475 1041 509
rect 1093 565 1127 599
rect 1093 486 1127 520
rect 1093 407 1127 441
rect 1213 573 1247 607
rect 1213 478 1247 512
rect 1299 565 1333 599
rect 1299 477 1333 511
rect 1299 379 1333 413
rect 1385 573 1419 607
rect 1385 494 1419 528
rect 1385 419 1419 453
rect 1471 565 1505 599
rect 1471 477 1505 511
rect 1471 379 1505 413
rect 1557 573 1591 607
rect 1557 494 1591 528
rect 1557 419 1591 453
<< poly >>
rect 165 619 195 645
rect 251 619 281 645
rect 337 619 367 645
rect 431 619 461 645
rect 517 619 547 645
rect 603 619 633 645
rect 793 619 823 645
rect 880 619 910 645
rect 966 619 996 645
rect 1052 619 1082 645
rect 1258 619 1288 645
rect 1344 619 1374 645
rect 1430 619 1460 645
rect 1516 619 1546 645
rect 165 335 195 367
rect 97 319 195 335
rect 97 285 137 319
rect 171 285 195 319
rect 97 269 195 285
rect 251 321 281 367
rect 337 321 367 367
rect 431 321 461 367
rect 517 321 547 367
rect 603 321 633 367
rect 793 335 823 367
rect 251 305 367 321
rect 251 271 316 305
rect 350 271 367 305
rect 97 233 127 269
rect 251 255 367 271
rect 409 305 475 321
rect 409 271 425 305
rect 459 271 475 305
rect 409 255 475 271
rect 517 305 690 321
rect 517 271 551 305
rect 585 271 619 305
rect 653 271 690 305
rect 517 255 690 271
rect 772 319 838 335
rect 772 285 788 319
rect 822 285 838 319
rect 772 270 838 285
rect 251 233 281 255
rect 337 233 367 255
rect 423 233 453 255
rect 517 233 547 255
rect 607 251 690 255
rect 780 269 838 270
rect 880 321 910 367
rect 966 321 996 367
rect 880 305 996 321
rect 880 271 905 305
rect 939 271 996 305
rect 607 233 637 251
rect 780 233 810 269
rect 880 255 996 271
rect 1052 335 1082 367
rect 1052 319 1125 335
rect 1052 285 1075 319
rect 1109 285 1125 319
rect 1052 269 1125 285
rect 1258 331 1288 367
rect 1344 331 1374 367
rect 1430 331 1460 367
rect 1516 331 1546 367
rect 1258 315 1546 331
rect 1258 281 1274 315
rect 1308 281 1342 315
rect 1376 281 1410 315
rect 1444 281 1478 315
rect 1512 281 1546 315
rect 880 233 910 255
rect 966 233 996 255
rect 1053 233 1083 269
rect 1258 265 1546 281
rect 1258 217 1288 265
rect 1344 217 1374 265
rect 1430 217 1460 265
rect 1516 217 1546 265
rect 97 39 127 65
rect 251 39 281 65
rect 337 39 367 65
rect 423 39 453 65
rect 517 39 547 65
rect 607 39 637 65
rect 780 39 810 65
rect 880 39 910 65
rect 966 39 996 65
rect 1053 39 1083 65
rect 1258 23 1288 49
rect 1344 23 1374 49
rect 1430 23 1460 49
rect 1516 23 1546 49
<< polycont >>
rect 137 285 171 319
rect 316 271 350 305
rect 425 271 459 305
rect 551 271 585 305
rect 619 271 653 305
rect 788 285 822 319
rect 905 271 939 305
rect 1075 285 1109 319
rect 1274 281 1308 315
rect 1342 281 1376 315
rect 1410 281 1444 315
rect 1478 281 1512 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 104 597 156 613
rect 104 563 120 597
rect 154 563 156 597
rect 104 521 156 563
rect 104 487 120 521
rect 154 487 156 521
rect 104 441 156 487
rect 190 599 242 615
rect 190 565 206 599
rect 240 565 242 599
rect 190 509 242 565
rect 276 585 342 649
rect 276 551 292 585
rect 326 551 342 585
rect 276 543 342 551
rect 376 599 436 615
rect 376 565 386 599
rect 420 565 436 599
rect 376 509 436 565
rect 190 475 206 509
rect 240 475 386 509
rect 420 475 436 509
rect 470 599 508 615
rect 470 565 472 599
rect 506 565 508 599
rect 470 507 508 565
rect 470 473 472 507
rect 506 473 508 507
rect 470 441 508 473
rect 104 407 120 441
rect 154 413 508 441
rect 154 407 472 413
rect 470 379 472 407
rect 506 379 508 413
rect 542 599 784 615
rect 542 565 558 599
rect 592 581 748 599
rect 592 565 608 581
rect 542 522 608 565
rect 732 565 748 581
rect 782 565 784 599
rect 542 488 558 522
rect 592 488 608 522
rect 542 443 608 488
rect 542 409 558 443
rect 592 409 608 443
rect 642 531 694 547
rect 642 497 644 531
rect 678 497 694 531
rect 642 413 694 497
rect 470 375 508 379
rect 642 379 644 413
rect 678 379 694 413
rect 732 521 784 565
rect 732 487 748 521
rect 782 487 784 521
rect 732 441 784 487
rect 818 599 871 615
rect 818 565 834 599
rect 868 565 871 599
rect 818 509 871 565
rect 905 584 971 649
rect 905 550 921 584
rect 955 550 971 584
rect 905 543 971 550
rect 1005 599 1057 615
rect 1005 565 1007 599
rect 1041 565 1057 599
rect 1005 509 1057 565
rect 818 475 834 509
rect 868 475 1007 509
rect 1041 475 1057 509
rect 1091 599 1143 615
rect 1091 565 1093 599
rect 1127 565 1143 599
rect 1091 520 1143 565
rect 1091 486 1093 520
rect 1127 486 1143 520
rect 1091 441 1143 486
rect 1197 607 1263 649
rect 1197 573 1213 607
rect 1247 573 1263 607
rect 1197 512 1263 573
rect 1197 478 1213 512
rect 1247 478 1263 512
rect 1197 475 1263 478
rect 1297 599 1335 615
rect 1297 565 1299 599
rect 1333 565 1335 599
rect 1297 511 1335 565
rect 1297 477 1299 511
rect 1333 477 1335 511
rect 732 407 748 441
rect 782 407 1093 441
rect 1127 407 1260 441
rect 642 375 694 379
rect 17 339 436 373
rect 470 341 694 375
rect 17 319 266 339
rect 17 285 137 319
rect 171 285 266 319
rect 402 307 436 339
rect 772 339 1125 373
rect 772 319 839 339
rect 402 305 475 307
rect 300 271 316 305
rect 350 271 366 305
rect 36 221 266 251
rect 300 242 366 271
rect 402 271 425 305
rect 459 271 475 305
rect 402 254 475 271
rect 511 305 738 307
rect 511 271 551 305
rect 585 271 619 305
rect 653 271 738 305
rect 772 285 788 319
rect 822 285 839 319
rect 989 319 1125 339
rect 772 271 839 285
rect 889 271 905 305
rect 939 271 955 305
rect 989 285 1075 319
rect 1109 285 1125 319
rect 1159 317 1260 407
rect 1297 413 1335 477
rect 1369 607 1435 649
rect 1369 573 1385 607
rect 1419 573 1435 607
rect 1369 528 1435 573
rect 1369 494 1385 528
rect 1419 494 1435 528
rect 1369 453 1435 494
rect 1369 419 1385 453
rect 1419 419 1435 453
rect 1469 599 1507 615
rect 1469 565 1471 599
rect 1505 565 1507 599
rect 1469 511 1507 565
rect 1469 477 1471 511
rect 1505 477 1507 511
rect 1297 379 1299 413
rect 1333 385 1335 413
rect 1469 413 1507 477
rect 1541 607 1607 649
rect 1541 573 1557 607
rect 1591 573 1607 607
rect 1541 528 1607 573
rect 1541 494 1557 528
rect 1591 494 1607 528
rect 1541 453 1607 494
rect 1541 419 1557 453
rect 1591 419 1607 453
rect 1469 385 1471 413
rect 1333 379 1471 385
rect 1505 385 1507 413
rect 1505 379 1615 385
rect 1297 351 1615 379
rect 1159 315 1528 317
rect 511 242 738 271
rect 889 242 955 271
rect 1159 281 1274 315
rect 1308 281 1342 315
rect 1376 281 1410 315
rect 1444 281 1478 315
rect 1512 281 1528 315
rect 1159 279 1528 281
rect 1159 251 1260 279
rect 36 187 52 221
rect 86 217 266 221
rect 86 187 88 217
rect 36 111 88 187
rect 232 208 266 217
rect 805 221 855 237
rect 232 192 771 208
rect 36 77 52 111
rect 86 77 88 111
rect 36 61 88 77
rect 122 149 138 183
rect 172 149 188 183
rect 232 179 662 192
rect 232 175 470 179
rect 232 174 292 175
rect 122 140 188 149
rect 281 141 292 174
rect 326 174 470 175
rect 326 141 328 174
rect 122 124 247 140
rect 122 107 206 124
rect 122 73 138 107
rect 172 90 206 107
rect 240 90 247 124
rect 172 73 247 90
rect 122 17 247 73
rect 281 107 328 141
rect 462 145 470 174
rect 504 174 662 179
rect 504 145 512 174
rect 281 73 292 107
rect 326 73 328 107
rect 281 51 328 73
rect 362 136 428 140
rect 362 102 378 136
rect 412 102 428 136
rect 362 17 428 102
rect 462 111 512 145
rect 646 158 662 174
rect 696 158 735 192
rect 769 158 771 192
rect 462 77 470 111
rect 504 77 512 111
rect 462 61 512 77
rect 546 136 612 140
rect 546 102 562 136
rect 596 102 612 136
rect 546 17 612 102
rect 646 111 771 158
rect 805 187 821 221
rect 991 225 1260 251
rect 1562 245 1615 351
rect 991 208 1007 225
rect 855 191 1007 208
rect 1041 215 1260 225
rect 1041 191 1057 215
rect 855 187 1057 191
rect 805 174 1057 187
rect 1297 211 1615 245
rect 1297 205 1333 211
rect 805 153 871 174
rect 805 119 821 153
rect 855 119 871 153
rect 991 157 1057 174
rect 905 124 957 140
rect 646 77 662 111
rect 696 77 735 111
rect 769 85 771 111
rect 905 90 921 124
rect 955 90 957 124
rect 991 123 1007 157
rect 1041 123 1057 157
rect 1093 145 1109 179
rect 1143 145 1159 179
rect 905 87 957 90
rect 1093 111 1159 145
rect 1093 87 1109 111
rect 905 85 1109 87
rect 769 77 1109 85
rect 1143 77 1159 111
rect 646 51 1159 77
rect 1197 147 1213 181
rect 1247 147 1263 181
rect 1197 95 1263 147
rect 1197 61 1213 95
rect 1247 61 1263 95
rect 1197 17 1263 61
rect 1297 171 1299 205
rect 1469 205 1505 211
rect 1297 101 1333 171
rect 1297 67 1299 101
rect 1297 51 1333 67
rect 1369 143 1385 177
rect 1419 143 1435 177
rect 1369 91 1435 143
rect 1369 57 1385 91
rect 1419 57 1435 91
rect 1369 17 1435 57
rect 1469 171 1471 205
rect 1469 101 1505 171
rect 1469 67 1471 101
rect 1469 51 1505 67
rect 1541 143 1557 177
rect 1591 143 1607 177
rect 1541 95 1607 143
rect 1541 61 1557 95
rect 1591 61 1607 95
rect 1541 17 1607 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o32a_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1872074
string GDS_START 1858214
<< end >>
