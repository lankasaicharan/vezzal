magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 379 162 735 246
rect 1 49 735 162
rect 0 0 768 49
<< scnmos >>
rect 458 136 494 220
rect 80 52 110 136
rect 252 52 288 136
rect 626 52 656 220
<< scpmoshvt >>
rect 80 467 110 551
rect 252 467 288 551
rect 458 367 494 451
rect 626 367 656 619
<< ndiff >>
rect 405 192 458 220
rect 405 158 413 192
rect 447 158 458 192
rect 405 136 458 158
rect 494 168 626 220
rect 494 136 581 168
rect 27 111 80 136
rect 27 77 35 111
rect 69 77 80 111
rect 27 52 80 77
rect 110 111 252 136
rect 110 77 132 111
rect 166 77 252 111
rect 110 52 252 77
rect 288 111 341 136
rect 288 77 299 111
rect 333 77 341 111
rect 573 134 581 136
rect 615 134 626 168
rect 288 52 341 77
rect 573 100 626 134
rect 573 66 581 100
rect 615 66 626 100
rect 573 52 626 66
rect 656 208 709 220
rect 656 174 667 208
rect 701 174 709 208
rect 656 101 709 174
rect 656 67 667 101
rect 701 67 709 101
rect 656 52 709 67
<< pdiff >>
rect 573 607 626 619
rect 573 573 581 607
rect 615 573 626 607
rect 27 529 80 551
rect 27 495 35 529
rect 69 495 80 529
rect 27 467 80 495
rect 110 526 252 551
rect 110 492 130 526
rect 164 492 252 526
rect 110 467 252 492
rect 288 529 341 551
rect 288 495 299 529
rect 333 495 341 529
rect 288 467 341 495
rect 573 539 626 573
rect 573 505 581 539
rect 615 505 626 539
rect 573 471 626 505
rect 573 451 581 471
rect 405 422 458 451
rect 405 388 413 422
rect 447 388 458 422
rect 405 367 458 388
rect 494 437 581 451
rect 615 437 626 471
rect 494 367 626 437
rect 656 599 709 619
rect 656 565 667 599
rect 701 565 709 599
rect 656 510 709 565
rect 656 476 667 510
rect 701 476 709 510
rect 656 413 709 476
rect 656 379 667 413
rect 701 379 709 413
rect 656 367 709 379
<< ndiffc >>
rect 413 158 447 192
rect 35 77 69 111
rect 132 77 166 111
rect 299 77 333 111
rect 581 134 615 168
rect 581 66 615 100
rect 667 174 701 208
rect 667 67 701 101
<< pdiffc >>
rect 581 573 615 607
rect 35 495 69 529
rect 130 492 164 526
rect 299 495 333 529
rect 581 505 615 539
rect 413 388 447 422
rect 581 437 615 471
rect 667 565 701 599
rect 667 476 701 510
rect 667 379 701 413
<< poly >>
rect 626 619 656 645
rect 80 551 110 577
rect 252 551 288 577
rect 80 372 110 467
rect 252 386 288 467
rect 458 451 494 477
rect 80 356 146 372
rect 80 322 96 356
rect 130 322 146 356
rect 80 288 146 322
rect 80 254 96 288
rect 130 254 146 288
rect 80 238 146 254
rect 188 370 288 386
rect 188 336 211 370
rect 245 336 288 370
rect 188 302 288 336
rect 458 335 494 367
rect 188 268 211 302
rect 245 268 288 302
rect 414 319 558 335
rect 626 325 656 367
rect 414 285 430 319
rect 464 285 498 319
rect 532 285 558 319
rect 414 269 558 285
rect 600 309 666 325
rect 600 275 616 309
rect 650 275 666 309
rect 80 136 110 238
rect 188 234 288 268
rect 188 200 211 234
rect 245 200 288 234
rect 458 220 494 269
rect 600 259 666 275
rect 626 220 656 259
rect 188 184 288 200
rect 252 136 288 184
rect 458 110 494 136
rect 80 26 110 52
rect 252 26 288 52
rect 626 26 656 52
<< polycont >>
rect 96 322 130 356
rect 96 254 130 288
rect 211 336 245 370
rect 211 268 245 302
rect 430 285 464 319
rect 498 285 532 319
rect 616 275 650 309
rect 211 200 245 234
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 19 529 80 545
rect 19 495 35 529
rect 69 495 80 529
rect 19 441 80 495
rect 114 526 180 649
rect 565 607 631 649
rect 565 573 581 607
rect 615 573 631 607
rect 114 492 130 526
rect 164 492 180 526
rect 114 476 180 492
rect 283 529 344 545
rect 283 495 299 529
rect 333 495 344 529
rect 283 479 344 495
rect 19 406 261 441
rect 20 356 146 372
rect 20 322 96 356
rect 130 322 146 356
rect 20 288 146 322
rect 20 254 96 288
rect 130 254 146 288
rect 20 238 146 254
rect 195 370 261 406
rect 195 336 211 370
rect 245 336 261 370
rect 195 302 261 336
rect 195 268 211 302
rect 245 268 261 302
rect 195 234 261 268
rect 195 204 211 234
rect 19 200 211 204
rect 245 200 261 234
rect 19 164 261 200
rect 295 331 344 479
rect 565 539 631 573
rect 565 505 581 539
rect 615 505 631 539
rect 565 471 631 505
rect 397 422 469 438
rect 565 437 581 471
rect 615 437 631 471
rect 565 433 631 437
rect 665 599 748 615
rect 665 565 667 599
rect 701 565 748 599
rect 665 510 748 565
rect 665 476 667 510
rect 701 476 748 510
rect 397 388 413 422
rect 447 399 469 422
rect 665 413 748 476
rect 447 388 631 399
rect 397 365 631 388
rect 295 319 548 331
rect 295 285 430 319
rect 464 285 498 319
rect 532 285 548 319
rect 295 277 548 285
rect 582 325 631 365
rect 665 379 667 413
rect 701 379 748 413
rect 665 363 748 379
rect 582 309 656 325
rect 19 111 82 164
rect 19 77 35 111
rect 69 77 82 111
rect 19 61 82 77
rect 116 111 182 130
rect 295 127 344 277
rect 582 275 616 309
rect 650 275 656 309
rect 582 259 656 275
rect 582 243 631 259
rect 397 209 631 243
rect 690 224 748 363
rect 397 192 469 209
rect 397 158 413 192
rect 447 158 469 192
rect 665 208 748 224
rect 397 142 469 158
rect 565 168 631 175
rect 116 77 132 111
rect 166 77 182 111
rect 116 17 182 77
rect 283 111 344 127
rect 283 77 299 111
rect 333 77 344 111
rect 283 61 344 77
rect 565 134 581 168
rect 615 134 631 168
rect 565 100 631 134
rect 565 66 581 100
rect 615 66 631 100
rect 565 17 631 66
rect 665 174 667 208
rect 701 174 748 208
rect 665 101 748 174
rect 665 67 667 101
rect 701 67 748 101
rect 665 51 748 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlygate4s18_1
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 703 94 737 128 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6255696
string GDS_START 6249070
<< end >>
