magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2034 1852
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 410 157 735 203
rect 1 21 735 157
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 131
rect 297 47 327 131
rect 391 47 421 131
rect 499 47 529 177
rect 625 47 655 177
<< scpmoshvt >>
rect 81 413 117 497
rect 194 413 230 497
rect 292 413 328 497
rect 491 297 527 497
rect 617 297 653 497
<< ndiff >>
rect 436 131 499 177
rect 27 106 89 131
rect 27 72 35 106
rect 69 72 89 106
rect 27 47 89 72
rect 119 106 171 131
rect 119 72 129 106
rect 163 72 171 106
rect 119 47 171 72
rect 235 106 297 131
rect 235 72 243 106
rect 277 72 297 106
rect 235 47 297 72
rect 327 47 391 131
rect 421 111 499 131
rect 421 77 445 111
rect 479 77 499 111
rect 421 47 499 77
rect 529 127 625 177
rect 529 93 539 127
rect 573 93 625 127
rect 529 47 625 93
rect 655 127 709 177
rect 655 93 665 127
rect 699 93 709 127
rect 655 47 709 93
<< pdiff >>
rect 27 462 81 497
rect 27 428 35 462
rect 69 428 81 462
rect 27 413 81 428
rect 117 471 194 497
rect 117 437 129 471
rect 163 437 194 471
rect 117 413 194 437
rect 230 462 292 497
rect 230 428 244 462
rect 278 428 292 462
rect 230 413 292 428
rect 328 483 491 497
rect 328 449 350 483
rect 384 449 428 483
rect 462 449 491 483
rect 328 413 491 449
rect 439 297 491 413
rect 527 457 617 497
rect 527 423 539 457
rect 573 423 617 457
rect 527 384 617 423
rect 527 350 539 384
rect 573 350 617 384
rect 527 297 617 350
rect 653 457 707 497
rect 653 423 665 457
rect 699 423 707 457
rect 653 389 707 423
rect 653 355 665 389
rect 699 355 707 389
rect 653 297 707 355
<< ndiffc >>
rect 35 72 69 106
rect 129 72 163 106
rect 243 72 277 106
rect 445 77 479 111
rect 539 93 573 127
rect 665 93 699 127
<< pdiffc >>
rect 35 428 69 462
rect 129 437 163 471
rect 244 428 278 462
rect 350 449 384 483
rect 428 449 462 483
rect 539 423 573 457
rect 539 350 573 384
rect 665 423 699 457
rect 665 355 699 389
<< poly >>
rect 81 497 117 523
rect 194 497 230 523
rect 292 497 328 523
rect 491 497 527 523
rect 617 497 653 523
rect 81 398 117 413
rect 194 398 230 413
rect 292 398 328 413
rect 79 265 119 398
rect 40 249 119 265
rect 40 215 56 249
rect 90 215 119 249
rect 40 199 119 215
rect 89 131 119 199
rect 192 227 232 398
rect 290 379 330 398
rect 290 363 398 379
rect 290 329 347 363
rect 381 329 398 363
rect 290 305 398 329
rect 314 282 398 305
rect 491 282 527 297
rect 617 282 653 297
rect 314 233 421 282
rect 489 265 529 282
rect 615 265 655 282
rect 192 211 271 227
rect 192 177 211 211
rect 245 191 271 211
rect 245 177 327 191
rect 192 161 327 177
rect 297 131 327 161
rect 391 131 421 233
rect 463 249 655 265
rect 463 215 473 249
rect 507 215 655 249
rect 463 197 655 215
rect 499 177 529 197
rect 625 177 655 197
rect 89 21 119 47
rect 297 21 327 47
rect 391 21 421 47
rect 499 21 529 47
rect 625 21 655 47
<< polycont >>
rect 56 215 90 249
rect 347 329 381 363
rect 211 177 245 211
rect 473 215 507 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 35 462 69 489
rect 103 471 179 527
rect 103 437 129 471
rect 163 437 179 471
rect 219 462 286 484
rect 35 403 69 428
rect 219 428 244 462
rect 278 428 286 462
rect 332 483 479 527
rect 332 449 350 483
rect 384 449 428 483
rect 462 449 479 483
rect 332 433 479 449
rect 515 457 618 473
rect 35 357 181 403
rect 29 249 90 323
rect 29 215 56 249
rect 29 153 90 215
rect 134 227 181 357
rect 219 295 286 428
rect 515 423 539 457
rect 573 423 618 457
rect 331 363 480 391
rect 331 329 347 363
rect 381 329 480 363
rect 515 384 618 423
rect 515 350 539 384
rect 573 350 618 384
rect 515 316 618 350
rect 665 457 719 527
rect 699 423 719 457
rect 665 389 719 423
rect 699 355 719 389
rect 665 336 719 355
rect 219 265 421 295
rect 219 261 507 265
rect 289 249 507 261
rect 134 211 255 227
rect 134 177 211 211
rect 245 177 255 211
rect 134 161 255 177
rect 289 215 473 249
rect 289 189 507 215
rect 134 131 177 161
rect 19 106 85 118
rect 19 72 35 106
rect 69 72 85 106
rect 19 17 85 72
rect 129 106 177 131
rect 289 122 333 189
rect 551 155 618 316
rect 163 72 177 106
rect 129 56 177 72
rect 243 106 333 122
rect 539 127 618 155
rect 277 83 333 106
rect 421 111 495 116
rect 243 54 277 72
rect 421 77 445 111
rect 479 77 495 111
rect 421 17 495 77
rect 573 93 618 127
rect 539 51 618 93
rect 665 127 719 144
rect 699 93 719 127
rect 665 17 719 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 581 425 615 459 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 397 357 431 391 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 29 153 90 323 0 FreeSans 400 0 0 0 A_N
port 1 nsew signal input
flabel locali s 46 170 46 170 0 FreeSans 400 0 0 0 A_N
port 1 nsew
flabel locali s 29 289 63 323 0 FreeSans 400 0 0 0 A_N
port 1 nsew
flabel locali s 581 357 615 391 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
rlabel comment s 0 0 0 0 4 and2b_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1780836
string GDS_START 1774972
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
