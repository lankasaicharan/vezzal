magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 331 1958 704
rect 934 321 1150 331
<< pwell >>
rect 670 271 936 279
rect 33 241 936 271
rect 1196 247 1532 281
rect 1196 241 1896 247
rect 33 49 1896 241
rect 0 0 1920 49
<< scnmos >>
rect 116 117 146 245
rect 255 117 285 245
rect 395 117 425 245
rect 504 161 534 245
rect 644 117 674 245
rect 776 125 806 253
rect 1027 47 1057 215
rect 1333 127 1363 255
rect 1419 127 1449 255
rect 1658 137 1688 221
rect 1783 53 1813 221
<< scpmoshvt >>
rect 99 411 129 611
rect 263 411 293 611
rect 372 411 402 579
rect 474 411 504 539
rect 560 411 590 539
rect 669 377 699 545
rect 1027 357 1057 609
rect 1340 393 1370 561
rect 1426 393 1456 561
rect 1624 383 1654 511
rect 1797 367 1827 619
<< ndiff >>
rect 696 245 776 253
rect 59 233 116 245
rect 59 199 71 233
rect 105 199 116 233
rect 59 163 116 199
rect 59 129 71 163
rect 105 129 116 163
rect 59 117 116 129
rect 146 117 255 245
rect 285 233 395 245
rect 285 199 296 233
rect 330 199 395 233
rect 285 117 395 199
rect 425 233 504 245
rect 425 199 436 233
rect 470 199 504 233
rect 425 163 504 199
rect 425 129 436 163
rect 470 161 504 163
rect 534 203 644 245
rect 534 169 568 203
rect 602 169 644 203
rect 534 161 644 169
rect 470 129 482 161
rect 425 117 482 129
rect 556 117 644 161
rect 674 241 776 245
rect 674 207 708 241
rect 742 207 776 241
rect 674 163 776 207
rect 674 129 708 163
rect 742 129 776 163
rect 674 125 776 129
rect 806 227 910 253
rect 806 193 864 227
rect 898 193 910 227
rect 806 125 910 193
rect 674 117 754 125
rect 161 77 219 117
rect 161 43 173 77
rect 207 43 219 77
rect 161 31 219 43
rect 970 188 1027 215
rect 970 154 982 188
rect 1016 154 1027 188
rect 970 47 1027 154
rect 1057 98 1168 215
rect 1222 173 1333 255
rect 1222 139 1234 173
rect 1268 139 1333 173
rect 1222 127 1333 139
rect 1363 243 1419 255
rect 1363 209 1374 243
rect 1408 209 1419 243
rect 1363 127 1419 209
rect 1449 178 1506 255
rect 1449 144 1460 178
rect 1494 144 1506 178
rect 1449 127 1506 144
rect 1601 196 1658 221
rect 1601 162 1613 196
rect 1647 162 1658 196
rect 1601 137 1658 162
rect 1688 209 1783 221
rect 1688 175 1722 209
rect 1756 175 1783 209
rect 1688 137 1783 175
rect 1057 64 1122 98
rect 1156 64 1168 98
rect 1057 47 1168 64
rect 1710 99 1783 137
rect 1710 65 1722 99
rect 1756 65 1783 99
rect 1710 53 1783 65
rect 1813 209 1870 221
rect 1813 175 1824 209
rect 1858 175 1870 209
rect 1813 103 1870 175
rect 1813 69 1824 103
rect 1858 69 1870 103
rect 1813 53 1870 69
<< pdiff >>
rect 42 597 99 611
rect 42 563 54 597
rect 88 563 99 597
rect 42 527 99 563
rect 42 493 54 527
rect 88 493 99 527
rect 42 457 99 493
rect 42 423 54 457
rect 88 423 99 457
rect 42 411 99 423
rect 129 599 263 611
rect 129 565 140 599
rect 174 565 263 599
rect 129 489 263 565
rect 129 455 140 489
rect 174 455 263 489
rect 129 411 263 455
rect 293 597 350 611
rect 293 563 304 597
rect 338 579 350 597
rect 338 563 372 579
rect 293 527 372 563
rect 293 493 304 527
rect 338 493 372 527
rect 293 457 372 493
rect 293 423 304 457
rect 338 423 372 457
rect 293 411 372 423
rect 402 539 452 579
rect 619 539 669 545
rect 402 527 474 539
rect 402 493 413 527
rect 447 493 474 527
rect 402 457 474 493
rect 402 423 413 457
rect 447 423 474 457
rect 402 411 474 423
rect 504 457 560 539
rect 504 423 515 457
rect 549 423 560 457
rect 504 411 560 423
rect 590 440 669 539
rect 590 411 624 440
rect 612 406 624 411
rect 658 406 669 440
rect 612 377 669 406
rect 699 533 840 545
rect 699 499 794 533
rect 828 499 840 533
rect 699 431 840 499
rect 699 397 794 431
rect 828 397 840 431
rect 699 377 840 397
rect 970 597 1027 609
rect 970 563 982 597
rect 1016 563 1027 597
rect 970 500 1027 563
rect 970 466 982 500
rect 1016 466 1027 500
rect 970 403 1027 466
rect 970 369 982 403
rect 1016 369 1027 403
rect 970 357 1027 369
rect 1057 597 1114 609
rect 1057 563 1068 597
rect 1102 563 1114 597
rect 1676 607 1797 619
rect 1057 500 1114 563
rect 1676 573 1688 607
rect 1722 573 1797 607
rect 1057 466 1068 500
rect 1102 466 1114 500
rect 1057 403 1114 466
rect 1057 369 1068 403
rect 1102 369 1114 403
rect 1181 549 1340 561
rect 1181 515 1193 549
rect 1227 515 1340 549
rect 1181 439 1340 515
rect 1181 405 1193 439
rect 1227 405 1340 439
rect 1181 393 1340 405
rect 1370 527 1426 561
rect 1370 493 1381 527
rect 1415 493 1426 527
rect 1370 439 1426 493
rect 1370 405 1381 439
rect 1415 405 1426 439
rect 1370 393 1426 405
rect 1456 527 1513 561
rect 1456 493 1467 527
rect 1501 493 1513 527
rect 1676 511 1797 573
rect 1456 439 1513 493
rect 1456 405 1467 439
rect 1501 405 1513 439
rect 1456 393 1513 405
rect 1567 499 1624 511
rect 1567 465 1579 499
rect 1613 465 1624 499
rect 1057 357 1114 369
rect 1567 383 1624 465
rect 1654 510 1797 511
rect 1654 476 1688 510
rect 1722 476 1797 510
rect 1654 413 1797 476
rect 1654 383 1688 413
rect 1676 379 1688 383
rect 1722 379 1797 413
rect 1676 367 1797 379
rect 1827 597 1884 619
rect 1827 563 1838 597
rect 1872 563 1884 597
rect 1827 505 1884 563
rect 1827 471 1838 505
rect 1872 471 1884 505
rect 1827 413 1884 471
rect 1827 379 1838 413
rect 1872 379 1884 413
rect 1827 367 1884 379
<< ndiffc >>
rect 71 199 105 233
rect 71 129 105 163
rect 296 199 330 233
rect 436 199 470 233
rect 436 129 470 163
rect 568 169 602 203
rect 708 207 742 241
rect 708 129 742 163
rect 864 193 898 227
rect 173 43 207 77
rect 982 154 1016 188
rect 1234 139 1268 173
rect 1374 209 1408 243
rect 1460 144 1494 178
rect 1613 162 1647 196
rect 1722 175 1756 209
rect 1122 64 1156 98
rect 1722 65 1756 99
rect 1824 175 1858 209
rect 1824 69 1858 103
<< pdiffc >>
rect 54 563 88 597
rect 54 493 88 527
rect 54 423 88 457
rect 140 565 174 599
rect 140 455 174 489
rect 304 563 338 597
rect 304 493 338 527
rect 304 423 338 457
rect 413 493 447 527
rect 413 423 447 457
rect 515 423 549 457
rect 624 406 658 440
rect 794 499 828 533
rect 794 397 828 431
rect 982 563 1016 597
rect 982 466 1016 500
rect 982 369 1016 403
rect 1068 563 1102 597
rect 1688 573 1722 607
rect 1068 466 1102 500
rect 1068 369 1102 403
rect 1193 515 1227 549
rect 1193 405 1227 439
rect 1381 493 1415 527
rect 1381 405 1415 439
rect 1467 493 1501 527
rect 1467 405 1501 439
rect 1579 465 1613 499
rect 1688 476 1722 510
rect 1688 379 1722 413
rect 1838 563 1872 597
rect 1838 471 1872 505
rect 1838 379 1872 413
<< poly >>
rect 99 611 129 637
rect 263 611 293 637
rect 372 613 955 643
rect 372 579 402 613
rect 474 539 504 565
rect 560 539 590 613
rect 669 545 699 571
rect 99 371 129 411
rect 86 355 152 371
rect 86 321 102 355
rect 136 321 152 355
rect 263 333 293 411
rect 372 385 402 411
rect 86 305 152 321
rect 194 317 293 333
rect 116 245 146 305
rect 194 283 210 317
rect 244 283 293 317
rect 474 343 504 411
rect 560 385 590 411
rect 669 349 699 377
rect 669 343 838 349
rect 474 329 838 343
rect 474 313 788 329
rect 194 267 293 283
rect 255 245 285 267
rect 395 245 425 271
rect 504 245 534 313
rect 772 295 788 313
rect 822 295 838 329
rect 772 279 838 295
rect 644 245 674 271
rect 776 253 806 279
rect 925 267 955 613
rect 1027 609 1057 635
rect 1797 619 1827 645
rect 1340 561 1370 587
rect 1426 561 1456 587
rect 1624 511 1654 537
rect 1340 361 1370 393
rect 1027 303 1057 357
rect 1263 345 1370 361
rect 1263 311 1279 345
rect 1313 311 1370 345
rect 1027 287 1118 303
rect 1263 295 1370 311
rect 1426 343 1456 393
rect 1426 327 1508 343
rect 1426 307 1458 327
rect 1027 267 1068 287
rect 925 253 1068 267
rect 1102 253 1118 287
rect 1333 255 1363 295
rect 1419 293 1458 307
rect 1492 307 1508 327
rect 1624 307 1654 383
rect 1797 327 1827 367
rect 1736 311 1827 327
rect 1492 293 1688 307
rect 1419 277 1688 293
rect 1419 255 1449 277
rect 504 135 534 161
rect 925 237 1118 253
rect 116 91 146 117
rect 255 91 285 117
rect 395 51 425 117
rect 644 51 674 117
rect 776 99 806 125
rect 925 51 955 237
rect 1027 215 1057 237
rect 395 21 955 51
rect 1658 221 1688 277
rect 1736 277 1752 311
rect 1786 277 1827 311
rect 1736 261 1827 277
rect 1783 221 1813 261
rect 1333 101 1363 127
rect 1419 101 1449 127
rect 1658 111 1688 137
rect 1027 21 1057 47
rect 1783 27 1813 53
<< polycont >>
rect 102 321 136 355
rect 210 283 244 317
rect 788 295 822 329
rect 1279 311 1313 345
rect 1068 253 1102 287
rect 1458 293 1492 327
rect 1752 277 1786 311
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 18 597 88 613
rect 18 563 54 597
rect 18 527 88 563
rect 18 493 54 527
rect 18 457 88 493
rect 18 423 54 457
rect 124 599 190 649
rect 124 565 140 599
rect 174 565 190 599
rect 124 489 190 565
rect 124 455 140 489
rect 174 455 190 489
rect 124 439 190 455
rect 288 597 812 613
rect 288 563 304 597
rect 338 579 812 597
rect 338 563 354 579
rect 288 527 354 563
rect 778 549 812 579
rect 966 597 1016 613
rect 966 563 982 597
rect 288 493 304 527
rect 338 493 354 527
rect 288 457 354 493
rect 18 407 88 423
rect 288 423 304 457
rect 338 423 354 457
rect 18 249 52 407
rect 288 403 354 423
rect 397 527 742 543
rect 397 493 413 527
rect 447 509 742 527
rect 447 493 463 509
rect 397 457 463 493
rect 397 423 413 457
rect 447 423 463 457
rect 397 407 463 423
rect 499 457 565 473
rect 499 423 515 457
rect 549 423 565 457
rect 124 371 330 403
rect 88 369 330 371
rect 88 355 158 369
rect 88 321 102 355
rect 136 321 158 355
rect 88 305 158 321
rect 194 317 260 333
rect 194 283 210 317
rect 244 283 260 317
rect 18 233 121 249
rect 194 236 260 283
rect 18 199 71 233
rect 105 199 121 233
rect 18 163 121 199
rect 296 233 330 369
rect 499 319 565 423
rect 601 440 672 473
rect 601 424 624 440
rect 601 390 607 424
rect 658 406 672 440
rect 641 390 672 406
rect 601 373 672 390
rect 296 183 330 199
rect 366 285 565 319
rect 18 129 71 163
rect 105 147 121 163
rect 366 147 400 285
rect 531 249 565 285
rect 105 129 400 147
rect 18 113 400 129
rect 436 233 486 249
rect 470 199 486 233
rect 436 163 486 199
rect 470 129 486 163
rect 436 87 486 129
rect 531 203 602 249
rect 531 169 568 203
rect 531 123 602 169
rect 638 87 672 373
rect 157 43 173 77
rect 207 43 223 77
rect 436 53 672 87
rect 708 241 742 509
rect 778 533 914 549
rect 778 499 794 533
rect 828 499 914 533
rect 778 431 914 499
rect 778 397 794 431
rect 828 397 914 431
rect 778 381 914 397
rect 708 163 742 207
rect 708 87 742 129
rect 778 329 832 345
rect 778 295 788 329
rect 822 295 832 329
rect 778 279 832 295
rect 778 157 812 279
rect 880 243 914 381
rect 848 227 914 243
rect 848 193 864 227
rect 898 193 914 227
rect 966 500 1016 563
rect 966 466 982 500
rect 966 403 1016 466
rect 966 369 982 403
rect 966 188 1016 369
rect 1052 597 1118 649
rect 1052 563 1068 597
rect 1102 563 1118 597
rect 1263 579 1647 613
rect 1052 500 1118 563
rect 1052 466 1068 500
rect 1102 466 1118 500
rect 1052 403 1118 466
rect 1052 369 1068 403
rect 1102 369 1118 403
rect 1052 353 1118 369
rect 1177 549 1227 565
rect 1177 515 1193 549
rect 1177 439 1227 515
rect 1177 424 1193 439
rect 1177 390 1183 424
rect 1217 390 1227 405
rect 1052 287 1127 303
rect 1052 253 1068 287
rect 1102 253 1127 287
rect 1052 236 1127 253
rect 1177 259 1227 390
rect 1263 345 1329 579
rect 1365 527 1431 543
rect 1365 493 1381 527
rect 1415 493 1431 527
rect 1365 439 1431 493
rect 1365 424 1381 439
rect 1365 390 1375 424
rect 1415 405 1431 439
rect 1409 390 1431 405
rect 1365 384 1431 390
rect 1467 527 1543 543
rect 1501 493 1543 527
rect 1467 439 1543 493
rect 1579 499 1647 579
rect 1613 465 1647 499
rect 1579 449 1647 465
rect 1501 413 1543 439
rect 1501 405 1577 413
rect 1263 311 1279 345
rect 1313 311 1329 345
rect 1263 295 1329 311
rect 1177 225 1338 259
rect 966 157 982 188
rect 778 154 982 157
rect 778 123 1016 154
rect 1052 173 1268 189
rect 1052 155 1234 173
rect 1052 87 1086 155
rect 1218 139 1234 155
rect 708 53 1086 87
rect 1122 98 1172 119
rect 1156 64 1172 98
rect 157 17 223 43
rect 1122 17 1172 64
rect 1218 87 1268 139
rect 1304 157 1338 225
rect 1374 243 1408 384
rect 1467 379 1577 405
rect 1444 327 1507 343
rect 1444 293 1458 327
rect 1492 293 1507 327
rect 1444 236 1507 293
rect 1374 193 1408 209
rect 1444 178 1494 200
rect 1444 157 1460 178
rect 1304 144 1460 157
rect 1304 123 1494 144
rect 1543 87 1577 379
rect 1613 225 1647 449
rect 1688 607 1722 649
rect 1688 510 1722 573
rect 1688 413 1722 476
rect 1838 597 1895 613
rect 1872 563 1895 597
rect 1838 505 1895 563
rect 1872 471 1895 505
rect 1688 363 1722 379
rect 1758 424 1802 430
rect 1758 390 1759 424
rect 1793 390 1802 424
rect 1758 327 1802 390
rect 1736 311 1802 327
rect 1736 277 1752 311
rect 1786 277 1802 311
rect 1736 261 1802 277
rect 1838 413 1895 471
rect 1872 379 1895 413
rect 1838 225 1895 379
rect 1613 196 1663 225
rect 1647 162 1663 196
rect 1613 133 1663 162
rect 1706 209 1772 225
rect 1706 175 1722 209
rect 1756 175 1772 209
rect 1218 53 1577 87
rect 1706 99 1772 175
rect 1706 65 1722 99
rect 1756 65 1772 99
rect 1706 17 1772 65
rect 1808 209 1895 225
rect 1808 175 1824 209
rect 1858 175 1895 209
rect 1808 103 1895 175
rect 1808 69 1824 103
rect 1858 69 1895 103
rect 1808 53 1895 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 607 406 624 424
rect 624 406 641 424
rect 607 390 641 406
rect 1183 405 1193 424
rect 1193 405 1217 424
rect 1183 390 1217 405
rect 1375 405 1381 424
rect 1381 405 1409 424
rect 1375 390 1409 405
rect 1759 390 1793 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 595 424 653 430
rect 595 390 607 424
rect 641 421 653 424
rect 1171 424 1229 430
rect 1171 421 1183 424
rect 641 393 1183 421
rect 641 390 653 393
rect 595 384 653 390
rect 1171 390 1183 393
rect 1217 390 1229 424
rect 1171 384 1229 390
rect 1363 424 1421 430
rect 1363 390 1375 424
rect 1409 421 1421 424
rect 1747 424 1805 430
rect 1747 421 1759 424
rect 1409 393 1759 421
rect 1409 390 1421 393
rect 1363 384 1421 390
rect 1747 390 1759 393
rect 1793 390 1805 424
rect 1747 384 1805 390
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xor3_1
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1855 94 1889 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1855 168 1889 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1855 390 1889 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1855 464 1889 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1855 538 1889 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4783324
string GDS_START 4769684
<< end >>
