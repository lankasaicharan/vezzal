magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 49 49 919 176
rect 0 0 960 49
<< scnmos >>
rect 132 66 162 150
rect 204 66 234 150
rect 306 66 336 150
rect 384 66 414 150
rect 552 66 582 150
rect 630 66 660 150
rect 734 66 764 150
rect 806 66 836 150
<< scpmoshvt >>
rect 112 419 162 619
rect 272 419 322 619
rect 378 419 428 619
rect 602 400 652 600
rect 708 400 758 600
rect 814 400 864 600
<< ndiff >>
rect 75 121 132 150
rect 75 87 87 121
rect 121 87 132 121
rect 75 66 132 87
rect 162 66 204 150
rect 234 121 306 150
rect 234 87 261 121
rect 295 87 306 121
rect 234 66 306 87
rect 336 66 384 150
rect 414 125 552 150
rect 414 91 507 125
rect 541 91 552 125
rect 414 66 552 91
rect 582 66 630 150
rect 660 112 734 150
rect 660 78 671 112
rect 705 78 734 112
rect 660 66 734 78
rect 764 66 806 150
rect 836 125 893 150
rect 836 91 847 125
rect 881 91 893 125
rect 836 66 893 91
<< pdiff >>
rect 55 597 112 619
rect 55 563 67 597
rect 101 563 112 597
rect 55 465 112 563
rect 55 431 67 465
rect 101 431 112 465
rect 55 419 112 431
rect 162 607 272 619
rect 162 573 219 607
rect 253 573 272 607
rect 162 473 272 573
rect 162 439 219 473
rect 253 439 272 473
rect 162 419 272 439
rect 322 597 378 619
rect 322 563 333 597
rect 367 563 378 597
rect 322 465 378 563
rect 322 431 333 465
rect 367 431 378 465
rect 322 419 378 431
rect 428 607 485 619
rect 428 573 439 607
rect 473 573 485 607
rect 428 532 485 573
rect 428 498 439 532
rect 473 498 485 532
rect 428 419 485 498
rect 545 560 602 600
rect 545 526 557 560
rect 591 526 602 560
rect 545 400 602 526
rect 652 494 708 600
rect 652 460 663 494
rect 697 460 708 494
rect 652 400 708 460
rect 758 588 814 600
rect 758 554 769 588
rect 803 554 814 588
rect 758 454 814 554
rect 758 420 769 454
rect 803 420 814 454
rect 758 400 814 420
rect 864 588 921 600
rect 864 554 875 588
rect 909 554 921 588
rect 864 454 921 554
rect 864 420 875 454
rect 909 420 921 454
rect 864 400 921 420
<< ndiffc >>
rect 87 87 121 121
rect 261 87 295 121
rect 507 91 541 125
rect 671 78 705 112
rect 847 91 881 125
<< pdiffc >>
rect 67 563 101 597
rect 67 431 101 465
rect 219 573 253 607
rect 219 439 253 473
rect 333 563 367 597
rect 333 431 367 465
rect 439 573 473 607
rect 439 498 473 532
rect 557 526 591 560
rect 663 460 697 494
rect 769 554 803 588
rect 769 420 803 454
rect 875 554 909 588
rect 875 420 909 454
<< poly >>
rect 112 619 162 645
rect 272 619 322 645
rect 378 619 428 645
rect 500 615 652 645
rect 112 317 162 419
rect 272 387 322 419
rect 96 301 162 317
rect 96 267 112 301
rect 146 267 162 301
rect 96 233 162 267
rect 214 371 336 387
rect 214 337 230 371
rect 264 337 336 371
rect 214 303 336 337
rect 378 306 428 419
rect 214 269 230 303
rect 264 269 336 303
rect 214 253 336 269
rect 96 199 112 233
rect 146 199 162 233
rect 96 183 162 199
rect 132 150 162 183
rect 204 150 234 176
rect 306 150 336 253
rect 384 290 452 306
rect 384 256 402 290
rect 436 256 452 290
rect 384 222 452 256
rect 500 302 530 615
rect 602 600 652 615
rect 708 600 758 626
rect 814 600 864 626
rect 602 374 652 400
rect 708 309 758 400
rect 814 368 864 400
rect 500 286 582 302
rect 500 252 516 286
rect 550 252 582 286
rect 500 236 582 252
rect 384 188 402 222
rect 436 188 452 222
rect 384 172 452 188
rect 384 150 414 172
rect 552 150 582 236
rect 630 293 758 309
rect 630 259 693 293
rect 727 259 758 293
rect 630 243 758 259
rect 806 352 872 368
rect 806 318 822 352
rect 856 318 872 352
rect 806 284 872 318
rect 806 250 822 284
rect 856 250 872 284
rect 630 150 660 243
rect 806 234 872 250
rect 806 195 836 234
rect 734 165 836 195
rect 734 150 764 165
rect 806 150 836 165
rect 132 51 162 66
rect 204 51 234 66
rect 132 21 234 51
rect 306 40 336 66
rect 384 40 414 66
rect 552 40 582 66
rect 630 40 660 66
rect 734 40 764 66
rect 806 40 836 66
<< polycont >>
rect 112 267 146 301
rect 230 337 264 371
rect 230 269 264 303
rect 112 199 146 233
rect 402 256 436 290
rect 516 252 550 286
rect 402 188 436 222
rect 693 259 727 293
rect 822 318 856 352
rect 822 250 856 284
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 25 597 167 613
rect 25 563 67 597
rect 101 563 167 597
rect 25 465 167 563
rect 25 431 67 465
rect 101 431 167 465
rect 25 384 167 431
rect 203 607 269 649
rect 203 573 219 607
rect 253 573 269 607
rect 203 473 269 573
rect 203 439 219 473
rect 253 439 269 473
rect 203 423 269 439
rect 317 597 383 613
rect 317 563 333 597
rect 367 563 383 597
rect 317 465 383 563
rect 423 607 489 649
rect 423 573 439 607
rect 473 573 489 607
rect 423 532 489 573
rect 423 498 439 532
rect 473 498 489 532
rect 423 482 489 498
rect 541 588 819 613
rect 541 579 769 588
rect 541 560 607 579
rect 541 526 557 560
rect 591 526 607 560
rect 753 554 769 579
rect 803 554 819 588
rect 541 482 607 526
rect 647 494 713 543
rect 317 431 333 465
rect 367 446 383 465
rect 647 460 663 494
rect 697 460 713 494
rect 647 446 713 460
rect 367 431 713 446
rect 317 412 713 431
rect 753 454 819 554
rect 753 420 769 454
rect 803 420 819 454
rect 753 404 819 420
rect 859 588 942 604
rect 859 554 875 588
rect 909 554 942 588
rect 859 454 942 554
rect 859 420 875 454
rect 909 420 942 454
rect 859 404 942 420
rect 25 147 59 384
rect 214 371 280 387
rect 214 337 230 371
rect 264 337 280 371
rect 96 301 162 317
rect 96 267 112 301
rect 146 267 162 301
rect 96 233 162 267
rect 214 303 280 337
rect 214 269 230 303
rect 264 269 280 303
rect 214 253 280 269
rect 316 342 636 376
rect 96 199 112 233
rect 146 217 162 233
rect 316 217 350 342
rect 146 199 350 217
rect 96 183 350 199
rect 386 290 455 306
rect 386 256 402 290
rect 436 256 455 290
rect 386 222 455 256
rect 500 286 566 302
rect 500 252 516 286
rect 550 252 566 286
rect 500 236 566 252
rect 386 188 402 222
rect 436 188 455 222
rect 602 198 636 342
rect 677 293 743 356
rect 677 259 693 293
rect 727 259 743 293
rect 677 236 743 259
rect 793 352 872 368
rect 793 318 822 352
rect 856 318 872 352
rect 793 284 872 318
rect 793 250 822 284
rect 856 250 872 284
rect 793 234 872 250
rect 908 198 942 404
rect 25 121 137 147
rect 25 113 87 121
rect 71 87 87 113
rect 121 87 137 121
rect 71 62 137 87
rect 245 121 311 147
rect 245 87 261 121
rect 295 87 311 121
rect 386 88 455 188
rect 491 164 942 198
rect 491 125 557 164
rect 491 91 507 125
rect 541 91 557 125
rect 245 17 311 87
rect 491 62 557 91
rect 655 112 721 128
rect 655 78 671 112
rect 705 78 721 112
rect 655 17 721 78
rect 831 125 942 164
rect 831 91 847 125
rect 881 91 942 125
rect 831 62 942 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a221o_lp
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6112120
string GDS_START 6103656
<< end >>
