magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3122 1975
<< nwell >>
rect -38 331 1862 704
rect 824 303 1036 331
<< pwell >>
rect 525 241 1000 243
rect 525 180 1817 241
rect 23 49 1817 180
rect 0 0 1824 49
<< scnmos >>
rect 104 70 134 154
rect 197 70 227 154
rect 305 70 335 154
rect 604 133 634 217
rect 690 133 720 217
rect 762 133 792 217
rect 887 49 917 217
rect 1081 47 1111 131
rect 1186 47 1216 215
rect 1258 47 1288 215
rect 1450 47 1480 215
rect 1536 47 1566 215
rect 1622 47 1652 215
rect 1708 47 1738 215
<< scpmoshvt >>
rect 80 468 110 596
rect 152 468 182 596
rect 391 413 421 541
rect 604 463 634 547
rect 690 463 720 547
rect 762 463 792 547
rect 917 339 947 591
rect 1140 367 1170 495
rect 1245 367 1275 619
rect 1331 367 1361 619
rect 1438 367 1468 619
rect 1524 367 1554 619
rect 1610 367 1640 619
rect 1696 367 1726 619
<< ndiff >>
rect 49 124 104 154
rect 49 90 57 124
rect 91 90 104 124
rect 49 70 104 90
rect 134 129 197 154
rect 134 95 145 129
rect 179 95 197 129
rect 134 70 197 95
rect 227 129 305 154
rect 227 95 250 129
rect 284 95 305 129
rect 227 70 305 95
rect 335 129 388 154
rect 335 95 346 129
rect 380 95 388 129
rect 335 70 388 95
rect 551 192 604 217
rect 551 158 559 192
rect 593 158 604 192
rect 551 133 604 158
rect 634 192 690 217
rect 634 158 645 192
rect 679 158 690 192
rect 634 133 690 158
rect 720 133 762 217
rect 792 133 887 217
rect 814 69 887 133
rect 814 35 826 69
rect 860 49 887 69
rect 917 209 974 217
rect 917 175 928 209
rect 962 175 974 209
rect 917 49 974 175
rect 1133 203 1186 215
rect 1133 169 1141 203
rect 1175 169 1186 203
rect 1133 131 1186 169
rect 1028 106 1081 131
rect 1028 72 1036 106
rect 1070 72 1081 106
rect 860 35 872 49
rect 814 27 872 35
rect 1028 47 1081 72
rect 1111 93 1186 131
rect 1111 59 1141 93
rect 1175 59 1186 93
rect 1111 47 1186 59
rect 1216 47 1258 215
rect 1288 203 1341 215
rect 1288 169 1299 203
rect 1333 169 1341 203
rect 1288 101 1341 169
rect 1288 67 1299 101
rect 1333 67 1341 101
rect 1288 47 1341 67
rect 1397 165 1450 215
rect 1397 131 1405 165
rect 1439 131 1450 165
rect 1397 93 1450 131
rect 1397 59 1405 93
rect 1439 59 1450 93
rect 1397 47 1450 59
rect 1480 187 1536 215
rect 1480 153 1491 187
rect 1525 153 1536 187
rect 1480 101 1536 153
rect 1480 67 1491 101
rect 1525 67 1536 101
rect 1480 47 1536 67
rect 1566 125 1622 215
rect 1566 91 1577 125
rect 1611 91 1622 125
rect 1566 47 1622 91
rect 1652 203 1708 215
rect 1652 169 1663 203
rect 1697 169 1708 203
rect 1652 135 1708 169
rect 1652 101 1663 135
rect 1697 101 1708 135
rect 1652 47 1708 101
rect 1738 202 1791 215
rect 1738 168 1749 202
rect 1783 168 1791 202
rect 1738 93 1791 168
rect 1738 59 1749 93
rect 1783 59 1791 93
rect 1738 47 1791 59
<< pdiff >>
rect 27 582 80 596
rect 27 548 35 582
rect 69 548 80 582
rect 27 468 80 548
rect 110 468 152 596
rect 182 582 235 596
rect 182 548 193 582
rect 227 548 235 582
rect 182 514 235 548
rect 182 480 193 514
rect 227 480 235 514
rect 182 468 235 480
rect 1192 607 1245 619
rect 860 583 917 591
rect 860 549 872 583
rect 906 549 917 583
rect 860 547 917 549
rect 297 510 391 541
rect 297 476 305 510
rect 339 476 391 510
rect 297 413 391 476
rect 421 527 487 541
rect 421 493 445 527
rect 479 493 487 527
rect 421 459 487 493
rect 551 523 604 547
rect 551 489 559 523
rect 593 489 604 523
rect 551 463 604 489
rect 634 523 690 547
rect 634 489 645 523
rect 679 489 690 523
rect 634 463 690 489
rect 720 463 762 547
rect 792 522 917 547
rect 792 488 803 522
rect 837 515 917 522
rect 837 488 872 515
rect 792 481 872 488
rect 906 481 917 515
rect 792 463 917 481
rect 421 425 445 459
rect 479 425 487 459
rect 421 413 487 425
rect 860 447 917 463
rect 860 413 872 447
rect 906 413 917 447
rect 860 339 917 413
rect 947 570 1000 591
rect 947 536 958 570
rect 992 536 1000 570
rect 947 502 1000 536
rect 1192 573 1200 607
rect 1234 573 1245 607
rect 947 468 958 502
rect 992 468 1000 502
rect 1192 495 1245 573
rect 947 339 1000 468
rect 1087 424 1140 495
rect 1087 390 1095 424
rect 1129 390 1140 424
rect 1087 367 1140 390
rect 1170 367 1245 495
rect 1275 574 1331 619
rect 1275 540 1286 574
rect 1320 540 1331 574
rect 1275 506 1331 540
rect 1275 472 1286 506
rect 1320 472 1331 506
rect 1275 367 1331 472
rect 1361 611 1438 619
rect 1361 577 1393 611
rect 1427 577 1438 611
rect 1361 487 1438 577
rect 1361 453 1393 487
rect 1427 453 1438 487
rect 1361 367 1438 453
rect 1468 599 1524 619
rect 1468 565 1479 599
rect 1513 565 1524 599
rect 1468 504 1524 565
rect 1468 470 1479 504
rect 1513 470 1524 504
rect 1468 413 1524 470
rect 1468 379 1479 413
rect 1513 379 1524 413
rect 1468 367 1524 379
rect 1554 607 1610 619
rect 1554 573 1565 607
rect 1599 573 1610 607
rect 1554 520 1610 573
rect 1554 486 1565 520
rect 1599 486 1610 520
rect 1554 439 1610 486
rect 1554 405 1565 439
rect 1599 405 1610 439
rect 1554 367 1610 405
rect 1640 599 1696 619
rect 1640 565 1651 599
rect 1685 565 1696 599
rect 1640 504 1696 565
rect 1640 470 1651 504
rect 1685 470 1696 504
rect 1640 413 1696 470
rect 1640 379 1651 413
rect 1685 379 1696 413
rect 1640 367 1696 379
rect 1726 599 1779 619
rect 1726 565 1737 599
rect 1771 565 1779 599
rect 1726 504 1779 565
rect 1726 470 1737 504
rect 1771 470 1779 504
rect 1726 413 1779 470
rect 1726 379 1737 413
rect 1771 379 1779 413
rect 1726 367 1779 379
<< ndiffc >>
rect 57 90 91 124
rect 145 95 179 129
rect 250 95 284 129
rect 346 95 380 129
rect 559 158 593 192
rect 645 158 679 192
rect 826 35 860 69
rect 928 175 962 209
rect 1141 169 1175 203
rect 1036 72 1070 106
rect 1141 59 1175 93
rect 1299 169 1333 203
rect 1299 67 1333 101
rect 1405 131 1439 165
rect 1405 59 1439 93
rect 1491 153 1525 187
rect 1491 67 1525 101
rect 1577 91 1611 125
rect 1663 169 1697 203
rect 1663 101 1697 135
rect 1749 168 1783 202
rect 1749 59 1783 93
<< pdiffc >>
rect 35 548 69 582
rect 193 548 227 582
rect 193 480 227 514
rect 872 549 906 583
rect 305 476 339 510
rect 445 493 479 527
rect 559 489 593 523
rect 645 489 679 523
rect 803 488 837 522
rect 872 481 906 515
rect 445 425 479 459
rect 872 413 906 447
rect 958 536 992 570
rect 1200 573 1234 607
rect 958 468 992 502
rect 1095 390 1129 424
rect 1286 540 1320 574
rect 1286 472 1320 506
rect 1393 577 1427 611
rect 1393 453 1427 487
rect 1479 565 1513 599
rect 1479 470 1513 504
rect 1479 379 1513 413
rect 1565 573 1599 607
rect 1565 486 1599 520
rect 1565 405 1599 439
rect 1651 565 1685 599
rect 1651 470 1685 504
rect 1651 379 1685 413
rect 1737 565 1771 599
rect 1737 470 1771 504
rect 1737 379 1771 413
<< poly >>
rect 80 596 110 622
rect 152 596 182 622
rect 252 615 720 645
rect 1245 619 1275 645
rect 1331 619 1361 645
rect 1438 619 1468 645
rect 1524 619 1554 645
rect 1610 619 1640 645
rect 1696 619 1726 645
rect 80 325 110 468
rect 21 309 110 325
rect 21 275 37 309
rect 71 295 110 309
rect 152 319 182 468
rect 252 391 282 615
rect 391 541 421 567
rect 604 547 634 573
rect 690 547 720 615
rect 917 591 947 617
rect 762 547 792 573
rect 391 391 421 413
rect 252 361 421 391
rect 152 303 263 319
rect 71 275 104 295
rect 152 289 213 303
rect 21 241 104 275
rect 21 207 37 241
rect 71 221 104 241
rect 197 269 213 289
rect 247 269 263 303
rect 391 269 421 361
rect 469 365 535 381
rect 469 331 485 365
rect 519 347 535 365
rect 604 347 634 463
rect 690 437 720 463
rect 762 419 792 463
rect 762 403 828 419
rect 762 369 778 403
rect 812 369 828 403
rect 762 353 828 369
rect 519 331 712 347
rect 469 317 712 331
rect 469 315 535 317
rect 682 305 712 317
rect 682 275 720 305
rect 197 235 263 269
rect 71 207 134 221
rect 21 191 134 207
rect 104 154 134 191
rect 197 201 213 235
rect 247 201 263 235
rect 197 185 263 201
rect 305 239 634 269
rect 197 154 227 185
rect 305 154 335 239
rect 453 87 519 239
rect 604 217 634 239
rect 690 217 720 275
rect 762 217 792 353
rect 1140 495 1170 521
rect 1140 345 1170 367
rect 1245 345 1275 367
rect 917 305 947 339
rect 1140 335 1275 345
rect 1331 335 1361 367
rect 842 289 947 305
rect 842 255 858 289
rect 892 275 947 289
rect 1081 319 1275 335
rect 1081 285 1097 319
rect 1131 315 1275 319
rect 1317 319 1383 335
rect 1131 285 1216 315
rect 892 255 917 275
rect 842 239 917 255
rect 887 217 917 239
rect 1081 269 1216 285
rect 604 107 634 133
rect 690 107 720 133
rect 762 107 792 133
rect 104 44 134 70
rect 197 44 227 70
rect 305 44 335 70
rect 453 53 469 87
rect 503 53 519 87
rect 453 37 519 53
rect 1081 131 1111 269
rect 1186 215 1216 269
rect 1317 285 1333 319
rect 1367 285 1383 319
rect 1438 303 1468 367
rect 1524 303 1554 367
rect 1610 303 1640 367
rect 1696 303 1726 367
rect 1317 267 1383 285
rect 1258 237 1383 267
rect 1425 287 1738 303
rect 1425 253 1441 287
rect 1475 253 1509 287
rect 1543 253 1577 287
rect 1611 253 1738 287
rect 1425 237 1738 253
rect 1258 215 1288 237
rect 1450 215 1480 237
rect 1536 215 1566 237
rect 1622 215 1652 237
rect 1708 215 1738 237
rect 887 23 917 49
rect 1081 21 1111 47
rect 1186 21 1216 47
rect 1258 21 1288 47
rect 1450 21 1480 47
rect 1536 21 1566 47
rect 1622 21 1652 47
rect 1708 21 1738 47
<< polycont >>
rect 37 275 71 309
rect 37 207 71 241
rect 213 269 247 303
rect 485 331 519 365
rect 778 369 812 403
rect 213 201 247 235
rect 858 255 892 289
rect 1097 285 1131 319
rect 469 53 503 87
rect 1333 285 1367 319
rect 1441 253 1475 287
rect 1509 253 1543 287
rect 1577 253 1611 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 19 582 73 649
rect 19 548 35 582
rect 69 548 73 582
rect 19 532 73 548
rect 141 582 243 598
rect 141 548 193 582
rect 227 548 243 582
rect 141 514 243 548
rect 17 309 87 498
rect 17 275 37 309
rect 71 275 87 309
rect 17 241 87 275
rect 17 207 37 241
rect 71 207 87 241
rect 17 168 87 207
rect 141 480 193 514
rect 227 480 243 514
rect 141 426 243 480
rect 289 510 341 649
rect 289 476 305 510
rect 339 476 341 510
rect 289 460 341 476
rect 375 577 602 615
rect 375 426 409 577
rect 141 392 409 426
rect 445 527 521 543
rect 479 493 521 527
rect 445 459 521 493
rect 479 425 521 459
rect 445 409 521 425
rect 141 145 179 392
rect 485 365 521 409
rect 213 303 449 358
rect 247 269 449 303
rect 213 235 449 269
rect 247 209 449 235
rect 519 331 521 365
rect 247 201 263 209
rect 213 185 263 201
rect 485 157 521 331
rect 41 124 107 134
rect 41 90 57 124
rect 91 90 107 124
rect 41 17 107 90
rect 141 129 195 145
rect 141 95 145 129
rect 179 95 195 129
rect 141 79 195 95
rect 234 129 296 145
rect 234 95 250 129
rect 284 95 296 129
rect 234 17 296 95
rect 330 129 521 157
rect 555 523 602 577
rect 787 583 906 649
rect 1196 607 1238 649
rect 787 549 872 583
rect 555 489 559 523
rect 593 489 602 523
rect 555 192 602 489
rect 555 158 559 192
rect 593 158 602 192
rect 555 142 602 158
rect 636 523 695 539
rect 636 489 645 523
rect 679 489 695 523
rect 636 293 695 489
rect 787 522 906 549
rect 787 488 803 522
rect 837 515 906 522
rect 837 488 872 515
rect 787 481 872 488
rect 787 472 906 481
rect 868 447 906 472
rect 761 403 828 419
rect 761 369 778 403
rect 812 369 828 403
rect 868 413 872 447
rect 868 397 906 413
rect 942 570 1008 586
rect 942 536 958 570
rect 992 536 1008 570
rect 1196 573 1200 607
rect 1234 573 1238 607
rect 1391 611 1439 649
rect 1196 557 1238 573
rect 1282 574 1357 590
rect 942 502 1008 536
rect 942 468 958 502
rect 992 498 1008 502
rect 1282 540 1286 574
rect 1320 540 1357 574
rect 1282 506 1357 540
rect 992 468 1215 498
rect 942 462 1215 468
rect 761 361 828 369
rect 942 361 983 462
rect 761 327 983 361
rect 636 289 908 293
rect 636 255 858 289
rect 892 255 908 289
rect 636 250 908 255
rect 636 192 695 250
rect 944 216 983 327
rect 636 158 645 192
rect 679 158 695 192
rect 912 209 983 216
rect 912 175 928 209
rect 962 175 983 209
rect 912 173 983 175
rect 1017 424 1145 428
rect 1017 390 1095 424
rect 1129 390 1145 424
rect 1017 386 1145 390
rect 1181 420 1215 462
rect 1282 472 1286 506
rect 1320 472 1357 506
rect 1282 456 1357 472
rect 1181 386 1287 420
rect 636 142 695 158
rect 1017 139 1051 386
rect 1087 319 1217 352
rect 1087 285 1097 319
rect 1131 285 1217 319
rect 1087 242 1217 285
rect 1253 335 1287 386
rect 1323 403 1357 456
rect 1391 577 1393 611
rect 1427 577 1439 611
rect 1391 487 1439 577
rect 1391 453 1393 487
rect 1427 453 1439 487
rect 1391 437 1439 453
rect 1473 599 1522 615
rect 1473 565 1479 599
rect 1513 565 1522 599
rect 1473 504 1522 565
rect 1473 470 1479 504
rect 1513 470 1522 504
rect 1473 413 1522 470
rect 1323 369 1439 403
rect 1253 319 1371 335
rect 1253 285 1333 319
rect 1367 285 1371 319
rect 1253 269 1371 285
rect 1405 287 1439 369
rect 1473 379 1479 413
rect 1513 379 1522 413
rect 1556 607 1608 649
rect 1556 573 1565 607
rect 1599 573 1608 607
rect 1556 520 1608 573
rect 1556 486 1565 520
rect 1599 486 1608 520
rect 1556 439 1608 486
rect 1556 405 1565 439
rect 1599 405 1608 439
rect 1556 389 1608 405
rect 1642 599 1689 615
rect 1642 565 1651 599
rect 1685 565 1689 599
rect 1642 504 1689 565
rect 1642 470 1651 504
rect 1685 494 1689 504
rect 1735 599 1787 649
rect 1735 565 1737 599
rect 1771 565 1787 599
rect 1735 504 1787 565
rect 1685 470 1701 494
rect 1642 413 1701 470
rect 1473 355 1522 379
rect 1642 379 1651 413
rect 1685 379 1701 413
rect 1642 355 1701 379
rect 1735 470 1737 504
rect 1771 470 1787 504
rect 1735 413 1787 470
rect 1735 379 1737 413
rect 1771 379 1787 413
rect 1735 363 1787 379
rect 1473 321 1701 355
rect 1405 253 1441 287
rect 1475 253 1509 287
rect 1543 253 1577 287
rect 1611 253 1627 287
rect 1405 237 1627 253
rect 1405 235 1439 237
rect 1125 203 1191 208
rect 1125 169 1141 203
rect 1175 169 1191 203
rect 330 95 346 129
rect 380 123 521 129
rect 380 95 396 123
rect 330 79 396 95
rect 740 106 1086 139
rect 740 105 1036 106
rect 740 89 774 105
rect 453 87 774 89
rect 453 53 469 87
rect 503 53 774 87
rect 1017 72 1036 105
rect 1070 72 1086 106
rect 453 51 774 53
rect 810 69 876 71
rect 810 35 826 69
rect 860 35 876 69
rect 1017 54 1086 72
rect 1125 93 1191 169
rect 1125 59 1141 93
rect 1175 59 1191 93
rect 810 17 876 35
rect 1125 17 1191 59
rect 1283 203 1439 235
rect 1661 203 1701 321
rect 1283 169 1299 203
rect 1333 199 1439 203
rect 1333 169 1337 199
rect 1283 101 1337 169
rect 1489 187 1663 203
rect 1283 67 1299 101
rect 1333 67 1337 101
rect 1283 51 1337 67
rect 1389 131 1405 165
rect 1439 131 1455 165
rect 1389 93 1455 131
rect 1389 59 1405 93
rect 1439 59 1455 93
rect 1389 17 1455 59
rect 1489 153 1491 187
rect 1525 169 1663 187
rect 1697 169 1701 203
rect 1525 153 1527 169
rect 1489 101 1527 153
rect 1661 135 1701 169
rect 1489 67 1491 101
rect 1525 67 1527 101
rect 1489 51 1527 67
rect 1561 125 1627 135
rect 1561 91 1577 125
rect 1611 91 1627 125
rect 1561 17 1627 91
rect 1661 101 1663 135
rect 1697 101 1701 135
rect 1661 85 1701 101
rect 1735 202 1799 218
rect 1735 168 1749 202
rect 1783 168 1799 202
rect 1735 93 1799 168
rect 1735 59 1749 93
rect 1783 59 1799 93
rect 1735 17 1799 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdlclkp_4
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1663 94 1697 128 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1663 168 1697 202 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1663 390 1697 424 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1438542
string GDS_START 1423582
<< end >>
