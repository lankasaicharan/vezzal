magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 59 49 668 157
rect 0 0 672 49
<< scnmos >>
rect 142 47 172 131
rect 220 47 250 131
rect 306 47 336 131
rect 378 47 408 131
rect 483 47 513 131
rect 555 47 585 131
<< scpmoshvt >>
rect 86 409 136 609
rect 192 409 242 609
rect 298 409 348 609
rect 535 409 585 609
<< ndiff >>
rect 85 101 142 131
rect 85 67 97 101
rect 131 67 142 101
rect 85 47 142 67
rect 172 47 220 131
rect 250 111 306 131
rect 250 77 261 111
rect 295 77 306 111
rect 250 47 306 77
rect 336 47 378 131
rect 408 106 483 131
rect 408 72 419 106
rect 453 72 483 106
rect 408 47 483 72
rect 513 47 555 131
rect 585 108 642 131
rect 585 74 596 108
rect 630 74 642 108
rect 585 47 642 74
<< pdiff >>
rect 29 597 86 609
rect 29 563 41 597
rect 75 563 86 597
rect 29 526 86 563
rect 29 492 41 526
rect 75 492 86 526
rect 29 455 86 492
rect 29 421 41 455
rect 75 421 86 455
rect 29 409 86 421
rect 136 591 192 609
rect 136 557 147 591
rect 181 557 192 591
rect 136 409 192 557
rect 242 597 298 609
rect 242 563 253 597
rect 287 563 298 597
rect 242 516 298 563
rect 242 482 253 516
rect 287 482 298 516
rect 242 409 298 482
rect 348 597 405 609
rect 348 563 359 597
rect 393 563 405 597
rect 348 526 405 563
rect 348 492 359 526
rect 393 492 405 526
rect 348 455 405 492
rect 348 421 359 455
rect 393 421 405 455
rect 348 409 405 421
rect 478 597 535 609
rect 478 563 490 597
rect 524 563 535 597
rect 478 526 535 563
rect 478 492 490 526
rect 524 492 535 526
rect 478 455 535 492
rect 478 421 490 455
rect 524 421 535 455
rect 478 409 535 421
rect 585 597 642 609
rect 585 563 596 597
rect 630 563 642 597
rect 585 526 642 563
rect 585 492 596 526
rect 630 492 642 526
rect 585 455 642 492
rect 585 421 596 455
rect 630 421 642 455
rect 585 409 642 421
<< ndiffc >>
rect 97 67 131 101
rect 261 77 295 111
rect 419 72 453 106
rect 596 74 630 108
<< pdiffc >>
rect 41 563 75 597
rect 41 492 75 526
rect 41 421 75 455
rect 147 557 181 591
rect 253 563 287 597
rect 253 482 287 516
rect 359 563 393 597
rect 359 492 393 526
rect 359 421 393 455
rect 490 563 524 597
rect 490 492 524 526
rect 490 421 524 455
rect 596 563 630 597
rect 596 492 630 526
rect 596 421 630 455
<< poly >>
rect 86 609 136 635
rect 192 609 242 635
rect 298 609 348 635
rect 535 609 585 635
rect 86 228 136 409
rect 192 358 242 409
rect 184 342 250 358
rect 184 308 200 342
rect 234 308 250 342
rect 298 348 348 409
rect 298 332 435 348
rect 298 318 385 332
rect 184 292 250 308
rect 86 212 172 228
rect 86 178 102 212
rect 136 178 172 212
rect 86 162 172 178
rect 142 131 172 162
rect 220 131 250 292
rect 369 298 385 318
rect 419 298 435 332
rect 535 347 585 409
rect 535 299 565 347
rect 369 264 435 298
rect 369 244 385 264
rect 306 230 385 244
rect 419 230 435 264
rect 306 214 435 230
rect 483 283 585 299
rect 483 249 521 283
rect 555 249 585 283
rect 483 215 585 249
rect 306 131 336 214
rect 378 131 408 214
rect 483 181 521 215
rect 555 181 585 215
rect 483 165 585 181
rect 483 131 513 165
rect 555 131 585 165
rect 142 21 172 47
rect 220 21 250 47
rect 306 21 336 47
rect 378 21 408 47
rect 483 21 513 47
rect 555 21 585 47
<< polycont >>
rect 200 308 234 342
rect 102 178 136 212
rect 385 298 419 332
rect 385 230 419 264
rect 521 249 555 283
rect 521 181 555 215
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 25 597 91 613
rect 25 563 41 597
rect 75 563 91 597
rect 25 526 91 563
rect 131 591 197 649
rect 131 557 147 591
rect 181 557 197 591
rect 131 536 197 557
rect 237 597 303 613
rect 237 563 253 597
rect 287 563 303 597
rect 25 492 41 526
rect 75 500 91 526
rect 237 516 303 563
rect 237 500 253 516
rect 75 492 253 500
rect 25 482 253 492
rect 287 482 303 516
rect 25 466 303 482
rect 339 597 409 613
rect 339 563 359 597
rect 393 563 409 597
rect 339 526 409 563
rect 339 492 359 526
rect 393 492 409 526
rect 25 455 91 466
rect 25 421 41 455
rect 75 421 91 455
rect 339 455 409 492
rect 339 430 359 455
rect 25 405 91 421
rect 299 421 359 430
rect 393 421 409 455
rect 299 405 409 421
rect 474 597 540 649
rect 474 563 490 597
rect 524 563 540 597
rect 474 526 540 563
rect 474 492 490 526
rect 524 492 540 526
rect 474 455 540 492
rect 474 421 490 455
rect 524 421 540 455
rect 474 405 540 421
rect 580 597 646 613
rect 580 563 596 597
rect 630 563 646 597
rect 580 526 646 563
rect 580 492 596 526
rect 630 492 646 526
rect 580 455 646 492
rect 580 421 596 455
rect 630 421 646 455
rect 299 384 373 405
rect 25 342 263 358
rect 25 308 200 342
rect 234 308 263 342
rect 25 292 263 308
rect 25 212 167 228
rect 25 178 102 212
rect 136 178 167 212
rect 25 162 167 178
rect 299 135 333 384
rect 580 369 646 421
rect 409 348 646 369
rect 369 335 646 348
rect 369 332 443 335
rect 369 298 385 332
rect 419 298 443 332
rect 369 264 443 298
rect 369 230 385 264
rect 419 230 443 264
rect 369 214 443 230
rect 505 283 571 299
rect 505 249 521 283
rect 555 249 571 283
rect 505 215 571 249
rect 505 181 521 215
rect 555 181 571 215
rect 505 165 571 181
rect 81 101 147 126
rect 81 67 97 101
rect 131 67 147 101
rect 81 17 147 67
rect 245 111 333 135
rect 245 77 261 111
rect 295 77 333 111
rect 245 53 333 77
rect 403 106 469 135
rect 612 129 646 335
rect 403 72 419 106
rect 453 72 469 106
rect 403 17 469 72
rect 580 108 646 129
rect 580 74 596 108
rect 630 74 646 108
rect 580 53 646 74
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21boi_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5534528
string GDS_START 5528204
<< end >>
