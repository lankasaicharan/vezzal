magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 1 49 1949 241
rect 0 0 2016 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 252 47 282 215
rect 338 47 368 215
rect 424 47 454 215
rect 510 47 540 215
rect 596 47 626 215
rect 682 47 712 215
rect 782 47 812 215
rect 868 47 898 215
rect 954 47 984 215
rect 1040 47 1070 215
rect 1238 47 1268 215
rect 1324 47 1354 215
rect 1410 47 1440 215
rect 1496 47 1526 215
rect 1582 47 1612 215
rect 1668 47 1698 215
rect 1754 47 1784 215
rect 1840 47 1870 215
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 252 367 282 619
rect 338 367 368 619
rect 424 367 454 619
rect 510 367 540 619
rect 596 367 626 619
rect 688 367 718 619
rect 776 367 806 619
rect 862 367 892 619
rect 948 367 978 619
rect 1034 367 1064 619
rect 1252 367 1282 619
rect 1338 367 1368 619
rect 1424 367 1454 619
rect 1510 367 1540 619
rect 1596 367 1626 619
rect 1682 367 1712 619
rect 1768 367 1798 619
rect 1854 367 1884 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 93 80 169
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 203 166 215
rect 110 169 121 203
rect 155 169 166 203
rect 110 101 166 169
rect 110 67 121 101
rect 155 67 166 101
rect 110 47 166 67
rect 196 97 252 215
rect 196 63 207 97
rect 241 63 252 97
rect 196 47 252 63
rect 282 165 338 215
rect 282 131 293 165
rect 327 131 338 165
rect 282 97 338 131
rect 282 63 293 97
rect 327 63 338 97
rect 282 47 338 63
rect 368 177 424 215
rect 368 143 379 177
rect 413 143 424 177
rect 368 47 424 143
rect 454 93 510 215
rect 454 59 465 93
rect 499 59 510 93
rect 454 47 510 59
rect 540 177 596 215
rect 540 143 551 177
rect 585 143 596 177
rect 540 47 596 143
rect 626 93 682 215
rect 626 59 637 93
rect 671 59 682 93
rect 626 47 682 59
rect 712 97 782 215
rect 712 63 737 97
rect 771 63 782 97
rect 712 47 782 63
rect 812 203 868 215
rect 812 169 823 203
rect 857 169 868 203
rect 812 101 868 169
rect 812 67 823 101
rect 857 67 868 101
rect 812 47 868 67
rect 898 169 954 215
rect 898 135 909 169
rect 943 135 954 169
rect 898 93 954 135
rect 898 59 909 93
rect 943 59 954 93
rect 898 47 954 59
rect 984 203 1040 215
rect 984 169 995 203
rect 1029 169 1040 203
rect 984 101 1040 169
rect 984 67 995 101
rect 1029 67 1040 101
rect 984 47 1040 67
rect 1070 205 1238 215
rect 1070 171 1081 205
rect 1115 171 1238 205
rect 1070 130 1238 171
rect 1070 96 1193 130
rect 1227 96 1238 130
rect 1070 93 1238 96
rect 1070 59 1081 93
rect 1115 59 1238 93
rect 1070 47 1238 59
rect 1268 206 1324 215
rect 1268 172 1279 206
rect 1313 172 1324 206
rect 1268 101 1324 172
rect 1268 67 1279 101
rect 1313 67 1324 101
rect 1268 47 1324 67
rect 1354 130 1410 215
rect 1354 96 1365 130
rect 1399 96 1410 130
rect 1354 47 1410 96
rect 1440 206 1496 215
rect 1440 172 1451 206
rect 1485 172 1496 206
rect 1440 101 1496 172
rect 1440 67 1451 101
rect 1485 67 1496 101
rect 1440 47 1496 67
rect 1526 169 1582 215
rect 1526 135 1537 169
rect 1571 135 1582 169
rect 1526 93 1582 135
rect 1526 59 1537 93
rect 1571 59 1582 93
rect 1526 47 1582 59
rect 1612 203 1668 215
rect 1612 169 1623 203
rect 1657 169 1668 203
rect 1612 101 1668 169
rect 1612 67 1623 101
rect 1657 67 1668 101
rect 1612 47 1668 67
rect 1698 169 1754 215
rect 1698 135 1709 169
rect 1743 135 1754 169
rect 1698 93 1754 135
rect 1698 59 1709 93
rect 1743 59 1754 93
rect 1698 47 1754 59
rect 1784 203 1840 215
rect 1784 169 1795 203
rect 1829 169 1840 203
rect 1784 101 1840 169
rect 1784 67 1795 101
rect 1829 67 1840 101
rect 1784 47 1840 67
rect 1870 169 1923 215
rect 1870 135 1881 169
rect 1915 135 1923 169
rect 1870 93 1923 135
rect 1870 59 1881 93
rect 1915 59 1923 93
rect 1870 47 1923 59
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 505 80 565
rect 27 471 35 505
rect 69 471 80 505
rect 27 413 80 471
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 607 166 619
rect 110 573 121 607
rect 155 573 166 607
rect 110 525 166 573
rect 110 491 121 525
rect 155 491 166 525
rect 110 441 166 491
rect 110 407 121 441
rect 155 407 166 441
rect 110 367 166 407
rect 196 599 252 619
rect 196 565 207 599
rect 241 565 252 599
rect 196 505 252 565
rect 196 471 207 505
rect 241 471 252 505
rect 196 413 252 471
rect 196 379 207 413
rect 241 379 252 413
rect 196 367 252 379
rect 282 607 338 619
rect 282 573 293 607
rect 327 573 338 607
rect 282 495 338 573
rect 282 461 293 495
rect 327 461 338 495
rect 282 367 338 461
rect 368 599 424 619
rect 368 565 379 599
rect 413 565 424 599
rect 368 513 424 565
rect 368 479 379 513
rect 413 479 424 513
rect 368 423 424 479
rect 368 389 379 423
rect 413 389 424 423
rect 368 367 424 389
rect 454 607 510 619
rect 454 573 465 607
rect 499 573 510 607
rect 454 495 510 573
rect 454 461 465 495
rect 499 461 510 495
rect 454 367 510 461
rect 540 599 596 619
rect 540 565 551 599
rect 585 565 596 599
rect 540 513 596 565
rect 540 479 551 513
rect 585 479 596 513
rect 540 423 596 479
rect 540 389 551 423
rect 585 389 596 423
rect 540 367 596 389
rect 626 611 688 619
rect 626 577 640 611
rect 674 577 688 611
rect 626 495 688 577
rect 626 461 640 495
rect 674 461 688 495
rect 626 367 688 461
rect 718 599 776 619
rect 718 565 729 599
rect 763 565 776 599
rect 718 514 776 565
rect 718 480 729 514
rect 763 480 776 514
rect 718 439 776 480
rect 718 405 729 439
rect 763 405 776 439
rect 718 367 776 405
rect 806 505 862 619
rect 806 471 817 505
rect 851 471 862 505
rect 806 409 862 471
rect 806 375 817 409
rect 851 375 862 409
rect 806 367 862 375
rect 892 597 948 619
rect 892 563 903 597
rect 937 563 948 597
rect 892 367 948 563
rect 978 517 1034 619
rect 978 483 989 517
rect 1023 483 1034 517
rect 978 409 1034 483
rect 978 375 989 409
rect 1023 375 1034 409
rect 978 367 1034 375
rect 1064 607 1117 619
rect 1064 573 1075 607
rect 1109 573 1117 607
rect 1064 507 1117 573
rect 1064 473 1075 507
rect 1109 473 1117 507
rect 1064 413 1117 473
rect 1064 379 1075 413
rect 1109 379 1117 413
rect 1064 367 1117 379
rect 1199 599 1252 619
rect 1199 565 1207 599
rect 1241 565 1252 599
rect 1199 529 1252 565
rect 1199 495 1207 529
rect 1241 495 1252 529
rect 1199 461 1252 495
rect 1199 427 1207 461
rect 1241 427 1252 461
rect 1199 367 1252 427
rect 1282 607 1338 619
rect 1282 573 1293 607
rect 1327 573 1338 607
rect 1282 500 1338 573
rect 1282 466 1293 500
rect 1327 466 1338 500
rect 1282 367 1338 466
rect 1368 599 1424 619
rect 1368 565 1379 599
rect 1413 565 1424 599
rect 1368 521 1424 565
rect 1368 487 1379 521
rect 1413 487 1424 521
rect 1368 443 1424 487
rect 1368 409 1379 443
rect 1413 409 1424 443
rect 1368 367 1424 409
rect 1454 607 1510 619
rect 1454 573 1465 607
rect 1499 573 1510 607
rect 1454 500 1510 573
rect 1454 466 1465 500
rect 1499 466 1510 500
rect 1454 367 1510 466
rect 1540 599 1596 619
rect 1540 565 1551 599
rect 1585 565 1596 599
rect 1540 529 1596 565
rect 1540 495 1551 529
rect 1585 495 1596 529
rect 1540 459 1596 495
rect 1540 425 1551 459
rect 1585 425 1596 459
rect 1540 367 1596 425
rect 1626 531 1682 619
rect 1626 497 1637 531
rect 1671 497 1682 531
rect 1626 409 1682 497
rect 1626 375 1637 409
rect 1671 375 1682 409
rect 1626 367 1682 375
rect 1712 599 1768 619
rect 1712 565 1723 599
rect 1757 565 1768 599
rect 1712 529 1768 565
rect 1712 495 1723 529
rect 1757 495 1768 529
rect 1712 459 1768 495
rect 1712 425 1723 459
rect 1757 425 1768 459
rect 1712 367 1768 425
rect 1798 547 1854 619
rect 1798 513 1809 547
rect 1843 513 1854 547
rect 1798 477 1854 513
rect 1798 443 1809 477
rect 1843 443 1854 477
rect 1798 409 1854 443
rect 1798 375 1809 409
rect 1843 375 1854 409
rect 1798 367 1854 375
rect 1884 599 1937 619
rect 1884 565 1895 599
rect 1929 565 1937 599
rect 1884 529 1937 565
rect 1884 495 1895 529
rect 1929 495 1937 529
rect 1884 459 1937 495
rect 1884 425 1895 459
rect 1929 425 1937 459
rect 1884 367 1937 425
<< ndiffc >>
rect 35 169 69 203
rect 35 59 69 93
rect 121 169 155 203
rect 121 67 155 101
rect 207 63 241 97
rect 293 131 327 165
rect 293 63 327 97
rect 379 143 413 177
rect 465 59 499 93
rect 551 143 585 177
rect 637 59 671 93
rect 737 63 771 97
rect 823 169 857 203
rect 823 67 857 101
rect 909 135 943 169
rect 909 59 943 93
rect 995 169 1029 203
rect 995 67 1029 101
rect 1081 171 1115 205
rect 1193 96 1227 130
rect 1081 59 1115 93
rect 1279 172 1313 206
rect 1279 67 1313 101
rect 1365 96 1399 130
rect 1451 172 1485 206
rect 1451 67 1485 101
rect 1537 135 1571 169
rect 1537 59 1571 93
rect 1623 169 1657 203
rect 1623 67 1657 101
rect 1709 135 1743 169
rect 1709 59 1743 93
rect 1795 169 1829 203
rect 1795 67 1829 101
rect 1881 135 1915 169
rect 1881 59 1915 93
<< pdiffc >>
rect 35 565 69 599
rect 35 471 69 505
rect 35 379 69 413
rect 121 573 155 607
rect 121 491 155 525
rect 121 407 155 441
rect 207 565 241 599
rect 207 471 241 505
rect 207 379 241 413
rect 293 573 327 607
rect 293 461 327 495
rect 379 565 413 599
rect 379 479 413 513
rect 379 389 413 423
rect 465 573 499 607
rect 465 461 499 495
rect 551 565 585 599
rect 551 479 585 513
rect 551 389 585 423
rect 640 577 674 611
rect 640 461 674 495
rect 729 565 763 599
rect 729 480 763 514
rect 729 405 763 439
rect 817 471 851 505
rect 817 375 851 409
rect 903 563 937 597
rect 989 483 1023 517
rect 989 375 1023 409
rect 1075 573 1109 607
rect 1075 473 1109 507
rect 1075 379 1109 413
rect 1207 565 1241 599
rect 1207 495 1241 529
rect 1207 427 1241 461
rect 1293 573 1327 607
rect 1293 466 1327 500
rect 1379 565 1413 599
rect 1379 487 1413 521
rect 1379 409 1413 443
rect 1465 573 1499 607
rect 1465 466 1499 500
rect 1551 565 1585 599
rect 1551 495 1585 529
rect 1551 425 1585 459
rect 1637 497 1671 531
rect 1637 375 1671 409
rect 1723 565 1757 599
rect 1723 495 1757 529
rect 1723 425 1757 459
rect 1809 513 1843 547
rect 1809 443 1843 477
rect 1809 375 1843 409
rect 1895 565 1929 599
rect 1895 495 1929 529
rect 1895 425 1929 459
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 252 619 282 645
rect 338 619 368 645
rect 424 619 454 645
rect 510 619 540 645
rect 596 619 626 645
rect 688 619 718 645
rect 776 619 806 645
rect 862 619 892 645
rect 948 619 978 645
rect 1034 619 1064 645
rect 1252 619 1282 645
rect 1338 619 1368 645
rect 1424 619 1454 645
rect 1510 619 1540 645
rect 1596 619 1626 645
rect 1682 619 1712 645
rect 1768 619 1798 645
rect 1854 619 1884 645
rect 80 321 110 367
rect 166 321 196 367
rect 252 321 282 367
rect 80 305 282 321
rect 80 271 96 305
rect 130 271 164 305
rect 198 271 232 305
rect 266 271 282 305
rect 80 255 282 271
rect 80 215 110 255
rect 166 215 196 255
rect 252 215 282 255
rect 338 335 368 367
rect 424 335 454 367
rect 510 335 540 367
rect 596 335 626 367
rect 338 319 626 335
rect 338 285 363 319
rect 397 285 431 319
rect 465 285 499 319
rect 533 285 567 319
rect 601 285 626 319
rect 688 303 718 367
rect 776 321 806 367
rect 862 321 892 367
rect 948 321 978 367
rect 1034 321 1064 367
rect 1252 321 1282 367
rect 1338 321 1368 367
rect 1424 321 1454 367
rect 1510 321 1540 367
rect 1596 321 1626 367
rect 1682 321 1712 367
rect 1768 321 1798 367
rect 1854 321 1884 367
rect 776 305 1181 321
rect 338 269 626 285
rect 338 215 368 269
rect 424 215 454 269
rect 510 215 540 269
rect 596 215 626 269
rect 668 287 734 303
rect 668 253 684 287
rect 718 253 734 287
rect 776 271 905 305
rect 939 271 973 305
rect 1007 271 1063 305
rect 1097 271 1131 305
rect 1165 271 1181 305
rect 776 255 1181 271
rect 1238 305 1540 321
rect 1238 271 1277 305
rect 1311 271 1345 305
rect 1379 271 1413 305
rect 1447 271 1481 305
rect 1515 271 1540 305
rect 1238 255 1540 271
rect 1582 305 1920 321
rect 1582 271 1598 305
rect 1632 271 1666 305
rect 1700 271 1734 305
rect 1768 271 1802 305
rect 1836 271 1870 305
rect 1904 271 1920 305
rect 1582 255 1920 271
rect 668 237 734 253
rect 682 215 712 237
rect 782 215 812 255
rect 868 215 898 255
rect 954 215 984 255
rect 1040 215 1070 255
rect 1238 215 1268 255
rect 1324 215 1354 255
rect 1410 215 1440 255
rect 1496 215 1526 255
rect 1582 215 1612 255
rect 1668 215 1698 255
rect 1754 215 1784 255
rect 1840 215 1870 255
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 424 21 454 47
rect 510 21 540 47
rect 596 21 626 47
rect 682 21 712 47
rect 782 21 812 47
rect 868 21 898 47
rect 954 21 984 47
rect 1040 21 1070 47
rect 1238 21 1268 47
rect 1324 21 1354 47
rect 1410 21 1440 47
rect 1496 21 1526 47
rect 1582 21 1612 47
rect 1668 21 1698 47
rect 1754 21 1784 47
rect 1840 21 1870 47
<< polycont >>
rect 96 271 130 305
rect 164 271 198 305
rect 232 271 266 305
rect 363 285 397 319
rect 431 285 465 319
rect 499 285 533 319
rect 567 285 601 319
rect 684 253 718 287
rect 905 271 939 305
rect 973 271 1007 305
rect 1063 271 1097 305
rect 1131 271 1165 305
rect 1277 271 1311 305
rect 1345 271 1379 305
rect 1413 271 1447 305
rect 1481 271 1515 305
rect 1598 271 1632 305
rect 1666 271 1700 305
rect 1734 271 1768 305
rect 1802 271 1836 305
rect 1870 271 1904 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 19 599 71 615
rect 19 565 35 599
rect 69 565 71 599
rect 19 505 71 565
rect 19 471 35 505
rect 69 471 71 505
rect 19 413 71 471
rect 19 379 35 413
rect 69 379 71 413
rect 105 607 171 649
rect 105 573 121 607
rect 155 573 171 607
rect 105 525 171 573
rect 105 491 121 525
rect 155 491 171 525
rect 105 441 171 491
rect 105 407 121 441
rect 155 407 171 441
rect 205 599 243 615
rect 205 565 207 599
rect 241 565 243 599
rect 205 505 243 565
rect 205 471 207 505
rect 241 471 243 505
rect 205 423 243 471
rect 277 607 343 649
rect 277 573 293 607
rect 327 573 343 607
rect 277 495 343 573
rect 277 461 293 495
rect 327 461 343 495
rect 277 457 343 461
rect 377 599 415 615
rect 377 565 379 599
rect 413 565 415 599
rect 377 513 415 565
rect 377 479 379 513
rect 413 479 415 513
rect 377 423 415 479
rect 449 607 515 649
rect 449 573 465 607
rect 499 573 515 607
rect 449 495 515 573
rect 449 461 465 495
rect 499 461 515 495
rect 449 457 515 461
rect 549 599 590 615
rect 549 565 551 599
rect 585 565 590 599
rect 549 513 590 565
rect 549 479 551 513
rect 585 479 590 513
rect 549 423 590 479
rect 624 611 690 649
rect 624 577 640 611
rect 674 577 690 611
rect 624 495 690 577
rect 624 461 640 495
rect 674 461 690 495
rect 624 457 690 461
rect 725 607 1125 615
rect 725 599 1075 607
rect 725 565 729 599
rect 763 597 1075 599
rect 763 565 903 597
rect 725 563 903 565
rect 937 573 1075 597
rect 1109 573 1125 607
rect 937 563 1125 573
rect 725 555 1125 563
rect 725 514 765 555
rect 725 480 729 514
rect 763 480 765 514
rect 725 439 765 480
rect 725 423 729 439
rect 205 413 379 423
rect 19 373 71 379
rect 205 379 207 413
rect 241 389 379 413
rect 413 389 551 423
rect 585 405 729 423
rect 763 405 765 439
rect 585 389 765 405
rect 799 517 1039 521
rect 799 505 989 517
rect 799 471 817 505
rect 851 483 989 505
rect 1023 483 1039 517
rect 851 471 1039 483
rect 799 458 1039 471
rect 799 409 855 458
rect 241 379 245 389
rect 205 373 245 379
rect 19 339 245 373
rect 799 375 817 409
rect 851 375 855 409
rect 347 350 617 355
rect 347 319 511 350
rect 545 319 617 350
rect 80 271 96 305
rect 130 271 164 305
rect 198 271 232 305
rect 266 276 311 305
rect 347 285 363 319
rect 397 285 431 319
rect 465 285 499 319
rect 545 316 567 319
rect 533 285 567 316
rect 601 285 617 319
rect 347 283 617 285
rect 80 255 264 271
rect 252 242 264 255
rect 298 249 311 276
rect 668 253 684 287
rect 718 276 737 287
rect 668 249 703 253
rect 298 242 703 249
rect 19 203 85 219
rect 19 169 35 203
rect 69 169 85 203
rect 19 93 85 169
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 119 203 157 219
rect 252 215 737 242
rect 799 237 855 375
rect 973 409 1039 458
rect 973 375 989 409
rect 1023 375 1039 409
rect 973 369 1039 375
rect 1073 507 1125 555
rect 1073 473 1075 507
rect 1109 473 1125 507
rect 1073 413 1125 473
rect 1073 379 1075 413
rect 1109 379 1125 413
rect 1191 599 1243 615
rect 1191 565 1207 599
rect 1241 565 1243 599
rect 1191 529 1243 565
rect 1191 495 1207 529
rect 1241 495 1243 529
rect 1191 461 1243 495
rect 1277 607 1343 649
rect 1277 573 1293 607
rect 1327 573 1343 607
rect 1277 500 1343 573
rect 1277 466 1293 500
rect 1327 466 1343 500
rect 1277 462 1343 466
rect 1377 599 1415 615
rect 1377 565 1379 599
rect 1413 565 1415 599
rect 1377 521 1415 565
rect 1377 487 1379 521
rect 1413 487 1415 521
rect 1191 427 1207 461
rect 1241 428 1243 461
rect 1377 443 1415 487
rect 1449 607 1515 649
rect 1449 573 1465 607
rect 1499 573 1515 607
rect 1449 500 1515 573
rect 1449 466 1465 500
rect 1499 466 1515 500
rect 1449 462 1515 466
rect 1549 599 1945 615
rect 1549 565 1551 599
rect 1585 581 1723 599
rect 1585 565 1587 581
rect 1549 529 1587 565
rect 1721 565 1723 581
rect 1757 581 1895 599
rect 1757 565 1759 581
rect 1549 495 1551 529
rect 1585 495 1587 529
rect 1377 428 1379 443
rect 1241 427 1379 428
rect 1191 409 1379 427
rect 1413 428 1415 443
rect 1549 459 1587 495
rect 1549 428 1551 459
rect 1413 425 1551 428
rect 1585 425 1587 459
rect 1413 409 1587 425
rect 1191 394 1587 409
rect 1637 531 1687 547
rect 1671 497 1687 531
rect 1637 409 1687 497
rect 1721 529 1759 565
rect 1893 565 1895 581
rect 1929 565 1945 599
rect 1721 495 1723 529
rect 1757 495 1759 529
rect 1721 459 1759 495
rect 1721 425 1723 459
rect 1757 425 1759 459
rect 1721 409 1759 425
rect 1793 513 1809 547
rect 1843 513 1859 547
rect 1793 477 1859 513
rect 1793 443 1809 477
rect 1843 443 1859 477
rect 1793 409 1859 443
rect 1893 529 1945 565
rect 1893 495 1895 529
rect 1929 495 1945 529
rect 1893 459 1945 495
rect 1893 425 1895 459
rect 1929 425 1945 459
rect 1893 409 1945 425
rect 1073 363 1125 379
rect 1671 375 1687 409
rect 1793 375 1809 409
rect 1843 375 1859 409
rect 1565 350 1603 360
rect 1565 316 1567 350
rect 1601 316 1603 350
rect 1637 341 1999 375
rect 1565 307 1603 316
rect 889 305 1227 307
rect 889 271 905 305
rect 939 271 973 305
rect 1007 271 1063 305
rect 1097 271 1131 305
rect 119 169 121 203
rect 155 181 157 203
rect 799 203 1031 237
rect 799 181 823 203
rect 155 169 329 181
rect 119 165 329 169
rect 119 147 293 165
rect 119 101 163 147
rect 277 131 293 147
rect 327 131 329 165
rect 363 177 823 181
rect 363 143 379 177
rect 413 143 551 177
rect 585 169 823 177
rect 857 169 859 203
rect 993 169 995 203
rect 1029 169 1031 203
rect 585 143 859 169
rect 363 139 859 143
rect 119 67 121 101
rect 155 67 163 101
rect 119 51 163 67
rect 197 97 243 113
rect 197 63 207 97
rect 241 63 243 97
rect 197 17 243 63
rect 277 105 329 131
rect 277 97 687 105
rect 277 63 293 97
rect 327 93 687 97
rect 327 63 465 93
rect 277 59 465 63
rect 499 59 637 93
rect 671 59 687 93
rect 277 51 687 59
rect 721 97 787 105
rect 721 63 737 97
rect 771 63 787 97
rect 721 17 787 63
rect 821 101 859 139
rect 821 67 823 101
rect 857 67 859 101
rect 821 51 859 67
rect 893 135 909 169
rect 943 135 959 169
rect 893 93 959 135
rect 893 59 909 93
rect 943 59 959 93
rect 893 17 959 59
rect 993 101 1031 169
rect 993 67 995 101
rect 1029 67 1031 101
rect 993 51 1031 67
rect 1065 205 1131 221
rect 1065 171 1081 205
rect 1115 171 1131 205
rect 1165 206 1227 305
rect 1261 305 1531 307
rect 1261 271 1277 305
rect 1311 276 1345 305
rect 1313 271 1345 276
rect 1379 271 1413 305
rect 1447 271 1481 305
rect 1515 271 1531 305
rect 1565 305 1920 307
rect 1565 271 1598 305
rect 1632 271 1666 305
rect 1700 271 1734 305
rect 1768 271 1802 305
rect 1836 271 1870 305
rect 1904 271 1920 305
rect 1261 242 1279 271
rect 1313 242 1415 271
rect 1261 240 1415 242
rect 1954 237 1999 341
rect 1449 206 1999 237
rect 1165 172 1279 206
rect 1313 172 1451 206
rect 1485 203 1999 206
rect 1485 172 1487 203
rect 1065 138 1131 171
rect 1065 130 1243 138
rect 1065 96 1193 130
rect 1227 96 1243 130
rect 1065 93 1243 96
rect 1065 59 1081 93
rect 1115 59 1243 93
rect 1065 17 1243 59
rect 1277 101 1315 172
rect 1277 67 1279 101
rect 1313 67 1315 101
rect 1277 51 1315 67
rect 1349 130 1415 138
rect 1349 96 1365 130
rect 1399 96 1415 130
rect 1349 17 1415 96
rect 1449 101 1487 172
rect 1621 169 1623 203
rect 1657 169 1659 203
rect 1793 169 1795 203
rect 1829 169 1831 203
rect 1449 67 1451 101
rect 1485 67 1487 101
rect 1449 51 1487 67
rect 1521 135 1537 169
rect 1571 135 1587 169
rect 1521 93 1587 135
rect 1521 59 1537 93
rect 1571 59 1587 93
rect 1521 17 1587 59
rect 1621 101 1659 169
rect 1621 67 1623 101
rect 1657 67 1659 101
rect 1621 51 1659 67
rect 1693 135 1709 169
rect 1743 135 1759 169
rect 1693 93 1759 135
rect 1693 59 1709 93
rect 1743 59 1759 93
rect 1693 17 1759 59
rect 1793 101 1831 169
rect 1793 67 1795 101
rect 1829 67 1831 101
rect 1793 51 1831 67
rect 1865 135 1881 169
rect 1915 135 1931 169
rect 1865 93 1931 135
rect 1865 59 1881 93
rect 1915 59 1931 93
rect 1865 17 1931 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 511 319 545 350
rect 511 316 533 319
rect 533 316 545 319
rect 264 271 266 276
rect 266 271 298 276
rect 264 242 298 271
rect 703 253 718 276
rect 718 253 737 276
rect 703 242 737 253
rect 1567 316 1601 350
rect 1279 271 1311 276
rect 1311 271 1313 276
rect 1279 242 1313 271
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 499 350 557 356
rect 499 316 511 350
rect 545 347 557 350
rect 1555 350 1613 356
rect 1555 347 1567 350
rect 545 319 1567 347
rect 545 316 557 319
rect 499 310 557 316
rect 1555 316 1567 319
rect 1601 316 1613 350
rect 1555 310 1613 316
rect 252 276 310 282
rect 252 242 264 276
rect 298 273 310 276
rect 691 276 749 282
rect 691 273 703 276
rect 298 245 703 273
rect 298 242 310 245
rect 252 236 310 242
rect 691 242 703 245
rect 737 273 749 276
rect 1267 276 1325 282
rect 1267 273 1279 276
rect 737 245 1279 273
rect 737 242 749 245
rect 691 236 749 242
rect 1267 242 1279 245
rect 1313 242 1325 276
rect 1267 236 1325 242
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xor2_4
flabel metal1 s 1279 242 1313 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel metal1 s 1567 316 1601 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 895 464 929 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 991 464 1025 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2074158
string GDS_START 2058060
<< end >>
