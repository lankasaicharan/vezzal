magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 3506 1975
<< nwell >>
rect -38 332 2246 704
<< pwell >>
rect 1 49 2207 248
rect 0 0 2208 49
<< scpmos >>
rect 86 368 116 592
rect 221 368 251 592
rect 321 368 351 592
rect 411 368 441 592
rect 900 368 930 592
rect 1000 368 1030 592
rect 1104 368 1134 592
rect 1230 368 1260 592
rect 1320 368 1350 592
rect 1420 368 1450 592
rect 1530 368 1560 592
rect 1620 368 1650 592
rect 1822 368 1852 592
rect 1912 368 1942 592
rect 2002 368 2032 592
rect 2092 368 2122 592
<< nmoslvt >>
rect 84 74 114 222
rect 171 74 201 222
rect 257 74 287 222
rect 343 74 373 222
rect 429 74 459 222
rect 515 74 545 222
rect 601 74 631 222
rect 689 74 719 222
rect 943 74 973 222
rect 1029 74 1059 222
rect 1147 74 1177 222
rect 1233 74 1263 222
rect 1353 74 1383 222
rect 1439 74 1469 222
rect 1533 74 1563 222
rect 1634 74 1664 222
rect 1720 74 1750 222
rect 1806 74 1836 222
rect 2005 74 2035 222
rect 2094 74 2124 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 204 171 222
rect 114 170 125 204
rect 159 170 171 204
rect 114 74 171 170
rect 201 120 257 222
rect 201 86 212 120
rect 246 86 257 120
rect 201 74 257 86
rect 287 207 343 222
rect 287 173 298 207
rect 332 173 343 207
rect 287 74 343 173
rect 373 144 429 222
rect 373 110 384 144
rect 418 110 429 144
rect 373 74 429 110
rect 459 116 515 222
rect 459 82 470 116
rect 504 82 515 116
rect 459 74 515 82
rect 545 184 601 222
rect 545 150 556 184
rect 590 150 601 184
rect 545 74 601 150
rect 631 116 689 222
rect 631 82 643 116
rect 677 82 689 116
rect 631 74 689 82
rect 719 196 769 222
rect 719 184 776 196
rect 719 150 730 184
rect 764 150 776 184
rect 719 138 776 150
rect 719 74 769 138
rect 893 128 943 222
rect 886 116 943 128
rect 886 82 898 116
rect 932 82 943 116
rect 886 74 943 82
rect 973 144 1029 222
rect 973 110 984 144
rect 1018 110 1029 144
rect 973 74 1029 110
rect 1059 100 1147 222
rect 1059 74 1086 100
rect 1074 66 1086 74
rect 1120 74 1147 100
rect 1177 144 1233 222
rect 1177 110 1188 144
rect 1222 110 1233 144
rect 1177 74 1233 110
rect 1263 100 1353 222
rect 1263 74 1291 100
rect 1120 66 1132 74
rect 1074 54 1132 66
rect 1278 66 1291 74
rect 1325 74 1353 100
rect 1383 210 1439 222
rect 1383 176 1394 210
rect 1428 176 1439 210
rect 1383 120 1439 176
rect 1383 86 1394 120
rect 1428 86 1439 120
rect 1383 74 1439 86
rect 1469 149 1533 222
rect 1469 115 1480 149
rect 1514 115 1533 149
rect 1469 74 1533 115
rect 1563 210 1634 222
rect 1563 176 1589 210
rect 1623 176 1634 210
rect 1563 120 1634 176
rect 1563 86 1589 120
rect 1623 86 1634 120
rect 1563 74 1634 86
rect 1664 210 1720 222
rect 1664 176 1675 210
rect 1709 176 1720 210
rect 1664 120 1720 176
rect 1664 86 1675 120
rect 1709 86 1720 120
rect 1664 74 1720 86
rect 1750 210 1806 222
rect 1750 176 1761 210
rect 1795 176 1806 210
rect 1750 120 1806 176
rect 1750 86 1761 120
rect 1795 86 1806 120
rect 1750 74 1806 86
rect 1836 142 2005 222
rect 1836 108 1847 142
rect 1881 108 1960 142
rect 1994 108 2005 142
rect 1836 74 2005 108
rect 2035 210 2094 222
rect 2035 176 2049 210
rect 2083 176 2094 210
rect 2035 120 2094 176
rect 2035 86 2049 120
rect 2083 86 2094 120
rect 2035 74 2094 86
rect 2124 210 2181 222
rect 2124 176 2135 210
rect 2169 176 2181 210
rect 2124 120 2181 176
rect 2124 86 2135 120
rect 2169 86 2181 120
rect 2124 74 2181 86
rect 1325 66 1338 74
rect 1278 54 1338 66
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 440 86 476
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 580 221 592
rect 116 546 164 580
rect 198 546 221 580
rect 116 510 221 546
rect 116 476 164 510
rect 198 476 221 510
rect 116 440 221 476
rect 116 406 164 440
rect 198 406 221 440
rect 116 368 221 406
rect 251 580 321 592
rect 251 546 264 580
rect 298 546 321 580
rect 251 508 321 546
rect 251 474 264 508
rect 298 474 321 508
rect 251 368 321 474
rect 351 580 411 592
rect 351 546 364 580
rect 398 546 411 580
rect 351 497 411 546
rect 351 463 364 497
rect 398 463 411 497
rect 351 414 411 463
rect 351 380 364 414
rect 398 380 411 414
rect 351 368 411 380
rect 441 580 780 592
rect 441 546 454 580
rect 488 546 523 580
rect 557 546 592 580
rect 626 546 662 580
rect 696 546 731 580
rect 765 546 780 580
rect 441 508 780 546
rect 441 474 454 508
rect 488 474 523 508
rect 557 474 592 508
rect 626 474 662 508
rect 696 474 731 508
rect 765 474 780 508
rect 441 368 780 474
rect 841 580 900 592
rect 841 546 853 580
rect 887 546 900 580
rect 841 508 900 546
rect 841 474 853 508
rect 887 474 900 508
rect 841 368 900 474
rect 930 547 1000 592
rect 930 513 953 547
rect 987 513 1000 547
rect 930 479 1000 513
rect 930 445 953 479
rect 987 445 1000 479
rect 930 411 1000 445
rect 930 377 953 411
rect 987 377 1000 411
rect 930 368 1000 377
rect 1030 580 1104 592
rect 1030 546 1053 580
rect 1087 546 1104 580
rect 1030 508 1104 546
rect 1030 474 1053 508
rect 1087 474 1104 508
rect 1030 368 1104 474
rect 1134 531 1230 592
rect 1134 497 1153 531
rect 1187 497 1230 531
rect 1134 440 1230 497
rect 1134 406 1153 440
rect 1187 406 1230 440
rect 1134 368 1230 406
rect 1260 580 1320 592
rect 1260 546 1273 580
rect 1307 546 1320 580
rect 1260 508 1320 546
rect 1260 474 1273 508
rect 1307 474 1320 508
rect 1260 368 1320 474
rect 1350 531 1420 592
rect 1350 497 1373 531
rect 1407 497 1420 531
rect 1350 440 1420 497
rect 1350 406 1373 440
rect 1407 406 1420 440
rect 1350 368 1420 406
rect 1450 580 1530 592
rect 1450 546 1473 580
rect 1507 546 1530 580
rect 1450 508 1530 546
rect 1450 474 1473 508
rect 1507 474 1530 508
rect 1450 368 1530 474
rect 1560 531 1620 592
rect 1560 497 1573 531
rect 1607 497 1620 531
rect 1560 424 1620 497
rect 1560 390 1573 424
rect 1607 390 1620 424
rect 1560 368 1620 390
rect 1650 580 1709 592
rect 1650 546 1663 580
rect 1697 546 1709 580
rect 1650 500 1709 546
rect 1650 466 1663 500
rect 1697 466 1709 500
rect 1650 368 1709 466
rect 1763 580 1822 592
rect 1763 546 1775 580
rect 1809 546 1822 580
rect 1763 500 1822 546
rect 1763 466 1775 500
rect 1809 466 1822 500
rect 1763 368 1822 466
rect 1852 580 1912 592
rect 1852 546 1865 580
rect 1899 546 1912 580
rect 1852 508 1912 546
rect 1852 474 1865 508
rect 1899 474 1912 508
rect 1852 424 1912 474
rect 1852 390 1865 424
rect 1899 390 1912 424
rect 1852 368 1912 390
rect 1942 580 2002 592
rect 1942 546 1955 580
rect 1989 546 2002 580
rect 1942 500 2002 546
rect 1942 466 1955 500
rect 1989 466 2002 500
rect 1942 368 2002 466
rect 2032 580 2092 592
rect 2032 546 2045 580
rect 2079 546 2092 580
rect 2032 508 2092 546
rect 2032 474 2045 508
rect 2079 474 2092 508
rect 2032 424 2092 474
rect 2032 390 2045 424
rect 2079 390 2092 424
rect 2032 368 2092 390
rect 2122 580 2181 592
rect 2122 546 2135 580
rect 2169 546 2181 580
rect 2122 497 2181 546
rect 2122 463 2135 497
rect 2169 463 2181 497
rect 2122 414 2181 463
rect 2122 380 2135 414
rect 2169 380 2181 414
rect 2122 368 2181 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 170 159 204
rect 212 86 246 120
rect 298 173 332 207
rect 384 110 418 144
rect 470 82 504 116
rect 556 150 590 184
rect 643 82 677 116
rect 730 150 764 184
rect 898 82 932 116
rect 984 110 1018 144
rect 1086 66 1120 100
rect 1188 110 1222 144
rect 1291 66 1325 100
rect 1394 176 1428 210
rect 1394 86 1428 120
rect 1480 115 1514 149
rect 1589 176 1623 210
rect 1589 86 1623 120
rect 1675 176 1709 210
rect 1675 86 1709 120
rect 1761 176 1795 210
rect 1761 86 1795 120
rect 1847 108 1881 142
rect 1960 108 1994 142
rect 2049 176 2083 210
rect 2049 86 2083 120
rect 2135 176 2169 210
rect 2135 86 2169 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 164 546 198 580
rect 164 476 198 510
rect 164 406 198 440
rect 264 546 298 580
rect 264 474 298 508
rect 364 546 398 580
rect 364 463 398 497
rect 364 380 398 414
rect 454 546 488 580
rect 523 546 557 580
rect 592 546 626 580
rect 662 546 696 580
rect 731 546 765 580
rect 454 474 488 508
rect 523 474 557 508
rect 592 474 626 508
rect 662 474 696 508
rect 731 474 765 508
rect 853 546 887 580
rect 853 474 887 508
rect 953 513 987 547
rect 953 445 987 479
rect 953 377 987 411
rect 1053 546 1087 580
rect 1053 474 1087 508
rect 1153 497 1187 531
rect 1153 406 1187 440
rect 1273 546 1307 580
rect 1273 474 1307 508
rect 1373 497 1407 531
rect 1373 406 1407 440
rect 1473 546 1507 580
rect 1473 474 1507 508
rect 1573 497 1607 531
rect 1573 390 1607 424
rect 1663 546 1697 580
rect 1663 466 1697 500
rect 1775 546 1809 580
rect 1775 466 1809 500
rect 1865 546 1899 580
rect 1865 474 1899 508
rect 1865 390 1899 424
rect 1955 546 1989 580
rect 1955 466 1989 500
rect 2045 546 2079 580
rect 2045 474 2079 508
rect 2045 390 2079 424
rect 2135 546 2169 580
rect 2135 463 2169 497
rect 2135 380 2169 414
<< poly >>
rect 86 592 116 618
rect 221 592 251 618
rect 321 592 351 618
rect 411 592 441 618
rect 900 592 930 618
rect 1000 592 1030 618
rect 1104 592 1134 618
rect 1230 592 1260 618
rect 1320 592 1350 618
rect 1420 592 1450 618
rect 1530 592 1560 618
rect 1620 592 1650 618
rect 1822 592 1852 618
rect 1912 592 1942 618
rect 2002 592 2032 618
rect 2092 592 2122 618
rect 86 353 116 368
rect 221 353 251 368
rect 321 353 351 368
rect 411 353 441 368
rect 900 353 930 368
rect 1000 353 1030 368
rect 1104 353 1134 368
rect 1230 353 1260 368
rect 1320 353 1350 368
rect 1420 353 1450 368
rect 1530 353 1560 368
rect 1620 353 1650 368
rect 1822 353 1852 368
rect 1912 353 1942 368
rect 2002 353 2032 368
rect 2092 353 2122 368
rect 83 326 119 353
rect 218 326 254 353
rect 46 310 254 326
rect 318 345 354 353
rect 408 345 444 353
rect 318 320 719 345
rect 318 315 465 320
rect 46 276 62 310
rect 96 276 130 310
rect 164 276 198 310
rect 232 276 254 310
rect 46 267 254 276
rect 429 286 465 315
rect 499 286 533 320
rect 567 286 601 320
rect 635 286 669 320
rect 703 286 719 320
rect 429 270 719 286
rect 897 336 933 353
rect 997 336 1033 353
rect 1101 336 1137 353
rect 1227 336 1263 353
rect 897 320 1263 336
rect 897 286 917 320
rect 951 286 985 320
rect 1019 286 1053 320
rect 1087 286 1121 320
rect 1155 286 1189 320
rect 1223 286 1263 320
rect 897 270 1263 286
rect 1317 336 1353 353
rect 1417 336 1453 353
rect 1527 336 1563 353
rect 1317 328 1563 336
rect 1617 328 1653 353
rect 1819 336 1855 353
rect 1909 336 1945 353
rect 1999 336 2035 353
rect 2089 336 2125 353
rect 1317 320 1653 328
rect 1317 286 1369 320
rect 1403 286 1437 320
rect 1471 286 1505 320
rect 1539 286 1653 320
rect 1317 270 1653 286
rect 1720 320 2125 336
rect 1720 306 1849 320
rect 46 237 373 267
rect 84 222 114 237
rect 171 222 201 237
rect 257 222 287 237
rect 343 222 373 237
rect 429 222 459 270
rect 515 222 545 270
rect 601 222 631 270
rect 689 222 719 270
rect 943 222 973 270
rect 1029 222 1059 270
rect 1147 222 1177 270
rect 1233 222 1263 270
rect 1353 222 1383 270
rect 1439 222 1469 270
rect 1533 240 1664 270
rect 1533 222 1563 240
rect 1634 222 1664 240
rect 1720 222 1750 306
rect 1806 286 1849 306
rect 1883 286 1917 320
rect 1951 286 1985 320
rect 2019 286 2053 320
rect 2087 286 2125 320
rect 1806 270 2125 286
rect 1806 222 1836 270
rect 2005 240 2124 270
rect 2005 222 2035 240
rect 2094 222 2124 240
rect 84 48 114 74
rect 171 48 201 74
rect 257 48 287 74
rect 343 48 373 74
rect 429 48 459 74
rect 515 48 545 74
rect 601 48 631 74
rect 689 48 719 74
rect 943 48 973 74
rect 1029 48 1059 74
rect 1147 48 1177 74
rect 1233 48 1263 74
rect 1353 48 1383 74
rect 1439 48 1469 74
rect 1533 48 1563 74
rect 1634 48 1664 74
rect 1720 48 1750 74
rect 1806 48 1836 74
rect 2005 48 2035 74
rect 2094 48 2124 74
<< polycont >>
rect 62 276 96 310
rect 130 276 164 310
rect 198 276 232 310
rect 465 286 499 320
rect 533 286 567 320
rect 601 286 635 320
rect 669 286 703 320
rect 917 286 951 320
rect 985 286 1019 320
rect 1053 286 1087 320
rect 1121 286 1155 320
rect 1189 286 1223 320
rect 1369 286 1403 320
rect 1437 286 1471 320
rect 1505 286 1539 320
rect 1849 286 1883 320
rect 1917 286 1951 320
rect 1985 286 2019 320
rect 2053 286 2087 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 23 406 39 440
rect 73 406 89 440
rect 23 390 89 406
rect 148 580 214 596
rect 148 546 164 580
rect 198 546 214 580
rect 148 510 214 546
rect 148 476 164 510
rect 198 476 214 510
rect 148 440 214 476
rect 248 580 314 649
rect 248 546 264 580
rect 298 546 314 580
rect 248 508 314 546
rect 248 474 264 508
rect 298 474 314 508
rect 248 458 314 474
rect 348 580 414 596
rect 348 546 364 580
rect 398 546 414 580
rect 348 497 414 546
rect 348 463 364 497
rect 398 463 414 497
rect 148 406 164 440
rect 198 424 214 440
rect 348 424 414 463
rect 448 580 781 649
rect 448 546 454 580
rect 488 546 523 580
rect 557 546 592 580
rect 626 546 662 580
rect 696 546 731 580
rect 765 546 781 580
rect 448 508 781 546
rect 448 474 454 508
rect 488 474 523 508
rect 557 474 592 508
rect 626 474 662 508
rect 696 474 731 508
rect 765 474 781 508
rect 448 458 781 474
rect 837 581 1713 615
rect 837 580 903 581
rect 837 546 853 580
rect 887 546 903 580
rect 1037 580 1103 581
rect 837 508 903 546
rect 837 474 853 508
rect 887 474 903 508
rect 837 458 903 474
rect 937 513 953 547
rect 987 513 1003 547
rect 937 479 1003 513
rect 937 445 953 479
rect 987 445 1003 479
rect 1037 546 1053 580
rect 1087 546 1103 580
rect 1257 580 1323 581
rect 1037 508 1103 546
rect 1037 474 1053 508
rect 1087 474 1103 508
rect 1037 458 1103 474
rect 1137 531 1203 547
rect 1137 497 1153 531
rect 1187 497 1203 531
rect 937 424 1003 445
rect 1137 440 1203 497
rect 1257 546 1273 580
rect 1307 546 1323 580
rect 1457 580 1523 581
rect 1257 508 1323 546
rect 1257 474 1273 508
rect 1307 474 1323 508
rect 1257 458 1323 474
rect 1357 531 1423 547
rect 1357 497 1373 531
rect 1407 497 1423 531
rect 1137 424 1153 440
rect 198 414 1153 424
rect 198 406 364 414
rect 148 390 364 406
rect 348 380 364 390
rect 398 411 1153 414
rect 398 390 953 411
rect 398 380 414 390
rect 348 364 414 380
rect 937 377 953 390
rect 987 406 1153 411
rect 1187 424 1203 440
rect 1357 440 1423 497
rect 1457 546 1473 580
rect 1507 546 1523 580
rect 1647 580 1713 581
rect 1457 508 1523 546
rect 1457 474 1473 508
rect 1507 474 1523 508
rect 1457 458 1523 474
rect 1557 531 1613 547
rect 1557 497 1573 531
rect 1607 497 1613 531
rect 1187 406 1319 424
rect 987 390 1319 406
rect 1357 406 1373 440
rect 1407 424 1423 440
rect 1557 430 1613 497
rect 1647 546 1663 580
rect 1697 546 1713 580
rect 1647 500 1713 546
rect 1647 466 1663 500
rect 1697 466 1713 500
rect 1759 580 1825 649
rect 1759 546 1775 580
rect 1809 546 1825 580
rect 1759 500 1825 546
rect 1759 466 1775 500
rect 1809 466 1825 500
rect 1859 580 1905 596
rect 1859 546 1865 580
rect 1899 546 1905 580
rect 1859 508 1905 546
rect 1859 474 1865 508
rect 1899 474 1905 508
rect 1859 430 1905 474
rect 1939 580 2005 649
rect 1939 546 1955 580
rect 1989 546 2005 580
rect 1939 500 2005 546
rect 1939 466 1955 500
rect 1989 466 2005 500
rect 2039 580 2095 596
rect 2039 546 2045 580
rect 2079 546 2095 580
rect 2039 508 2095 546
rect 2039 474 2045 508
rect 2079 474 2095 508
rect 2039 430 2095 474
rect 1557 424 2095 430
rect 1407 406 1573 424
rect 1357 390 1573 406
rect 1607 390 1865 424
rect 1899 390 2045 424
rect 2079 390 2095 424
rect 2135 580 2185 649
rect 2169 546 2185 580
rect 2135 497 2185 546
rect 2169 463 2185 497
rect 2135 414 2185 463
rect 987 377 1003 390
rect 937 364 1003 377
rect 25 310 248 356
rect 25 276 62 310
rect 96 276 130 310
rect 164 276 198 310
rect 232 276 248 310
rect 449 320 839 356
rect 1037 328 1239 356
rect 449 286 465 320
rect 499 286 533 320
rect 567 286 601 320
rect 635 286 669 320
rect 703 286 839 320
rect 897 320 1239 328
rect 897 286 917 320
rect 951 286 985 320
rect 1019 286 1053 320
rect 1087 286 1121 320
rect 1155 286 1189 320
rect 1223 286 1239 320
rect 25 260 248 276
rect 1273 252 1319 390
rect 2169 380 2185 414
rect 2135 364 2185 380
rect 1353 320 1555 356
rect 1353 286 1369 320
rect 1403 286 1437 320
rect 1471 286 1505 320
rect 1539 286 1555 320
rect 1833 320 2087 356
rect 1353 270 1555 286
rect 23 210 73 226
rect 282 220 1319 252
rect 1589 260 1795 294
rect 1833 286 1849 320
rect 1883 286 1917 320
rect 1951 286 1985 320
rect 2019 286 2053 320
rect 1833 270 2087 286
rect 1589 236 1623 260
rect 23 176 39 210
rect 23 120 73 176
rect 109 218 1319 220
rect 109 207 348 218
rect 109 204 298 207
rect 109 170 125 204
rect 159 173 298 204
rect 332 173 348 207
rect 1378 210 1623 236
rect 1745 226 1795 260
rect 1378 184 1394 210
rect 159 170 348 173
rect 109 154 348 170
rect 384 150 556 184
rect 590 150 730 184
rect 764 150 780 184
rect 814 176 1394 184
rect 1428 202 1589 210
rect 814 150 1428 176
rect 384 144 418 150
rect 23 86 39 120
rect 73 86 212 120
rect 246 110 384 120
rect 814 116 848 150
rect 984 144 1034 150
rect 246 86 418 110
rect 23 70 418 86
rect 454 82 470 116
rect 504 82 643 116
rect 677 82 848 116
rect 454 66 848 82
rect 882 82 898 116
rect 932 82 948 116
rect 882 17 948 82
rect 1018 110 1034 144
rect 1172 144 1238 150
rect 984 70 1034 110
rect 1070 100 1136 116
rect 1070 66 1086 100
rect 1120 66 1136 100
rect 1172 110 1188 144
rect 1222 110 1238 144
rect 1378 120 1428 150
rect 1172 70 1238 110
rect 1274 100 1342 116
rect 1070 17 1136 66
rect 1274 66 1291 100
rect 1325 66 1342 100
rect 1378 86 1394 120
rect 1378 70 1428 86
rect 1464 149 1530 165
rect 1464 115 1480 149
rect 1514 115 1530 149
rect 1274 17 1342 66
rect 1464 17 1530 115
rect 1589 120 1623 176
rect 1589 70 1623 86
rect 1659 210 1709 226
rect 1659 176 1675 210
rect 1659 120 1709 176
rect 1659 86 1675 120
rect 1659 17 1709 86
rect 1745 210 2083 226
rect 1745 176 1761 210
rect 1795 192 2049 210
rect 1745 120 1795 176
rect 2033 176 2049 192
rect 1745 86 1761 120
rect 1745 70 1795 86
rect 1831 142 1999 158
rect 1831 108 1847 142
rect 1881 108 1960 142
rect 1994 108 1999 142
rect 1831 17 1999 108
rect 2033 120 2083 176
rect 2033 86 2049 120
rect 2033 70 2083 86
rect 2119 210 2185 226
rect 2119 176 2135 210
rect 2169 176 2185 210
rect 2119 120 2185 176
rect 2119 86 2135 120
rect 2169 86 2185 120
rect 2119 17 2185 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o311ai_4
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 684980
string GDS_START 668068
<< end >>
