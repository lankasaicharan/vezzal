magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 207 172 845 259
rect 1 49 845 172
rect 0 0 864 49
<< scnmos >>
rect 80 62 110 146
rect 286 65 316 233
rect 372 65 402 233
rect 458 65 488 233
rect 560 65 590 233
rect 646 65 676 233
rect 732 65 762 233
<< scpmoshvt >>
rect 153 367 183 451
rect 286 367 316 619
rect 372 367 402 619
rect 474 367 504 619
rect 560 367 590 619
rect 646 367 676 619
rect 732 367 762 619
<< ndiff >>
rect 233 221 286 233
rect 233 187 241 221
rect 275 187 286 221
rect 27 124 80 146
rect 27 90 35 124
rect 69 90 80 124
rect 27 62 80 90
rect 110 121 163 146
rect 110 87 121 121
rect 155 87 163 121
rect 110 62 163 87
rect 233 111 286 187
rect 233 77 241 111
rect 275 77 286 111
rect 233 65 286 77
rect 316 225 372 233
rect 316 191 327 225
rect 361 191 372 225
rect 316 153 372 191
rect 316 119 327 153
rect 361 119 372 153
rect 316 65 372 119
rect 402 221 458 233
rect 402 187 413 221
rect 447 187 458 221
rect 402 111 458 187
rect 402 77 413 111
rect 447 77 458 111
rect 402 65 458 77
rect 488 183 560 233
rect 488 149 503 183
rect 537 149 560 183
rect 488 107 560 149
rect 488 73 503 107
rect 537 73 560 107
rect 488 65 560 73
rect 590 221 646 233
rect 590 187 601 221
rect 635 187 646 221
rect 590 111 646 187
rect 590 77 601 111
rect 635 77 646 111
rect 590 65 646 77
rect 676 183 732 233
rect 676 149 687 183
rect 721 149 732 183
rect 676 107 732 149
rect 676 73 687 107
rect 721 73 732 107
rect 676 65 732 73
rect 762 221 819 233
rect 762 187 777 221
rect 811 187 819 221
rect 762 111 819 187
rect 762 77 777 111
rect 811 77 819 111
rect 762 65 819 77
<< pdiff >>
rect 233 607 286 619
rect 233 573 241 607
rect 275 573 286 607
rect 233 502 286 573
rect 233 468 241 502
rect 275 468 286 502
rect 233 451 286 468
rect 100 426 153 451
rect 100 392 108 426
rect 142 392 153 426
rect 100 367 153 392
rect 183 413 286 451
rect 183 379 194 413
rect 228 379 286 413
rect 183 367 286 379
rect 316 599 372 619
rect 316 565 327 599
rect 361 565 372 599
rect 316 506 372 565
rect 316 472 327 506
rect 361 472 372 506
rect 316 413 372 472
rect 316 379 327 413
rect 361 379 372 413
rect 316 367 372 379
rect 402 600 474 619
rect 402 566 415 600
rect 449 566 474 600
rect 402 367 474 566
rect 504 600 560 619
rect 504 566 515 600
rect 549 566 560 600
rect 504 367 560 566
rect 590 508 646 619
rect 590 474 601 508
rect 635 474 646 508
rect 590 367 646 474
rect 676 604 732 619
rect 676 570 687 604
rect 721 570 732 604
rect 676 492 732 570
rect 676 458 687 492
rect 721 458 732 492
rect 676 367 732 458
rect 762 607 815 619
rect 762 573 773 607
rect 807 573 815 607
rect 762 506 815 573
rect 762 472 773 506
rect 807 472 815 506
rect 762 413 815 472
rect 762 379 773 413
rect 807 379 815 413
rect 762 367 815 379
<< ndiffc >>
rect 241 187 275 221
rect 35 90 69 124
rect 121 87 155 121
rect 241 77 275 111
rect 327 191 361 225
rect 327 119 361 153
rect 413 187 447 221
rect 413 77 447 111
rect 503 149 537 183
rect 503 73 537 107
rect 601 187 635 221
rect 601 77 635 111
rect 687 149 721 183
rect 687 73 721 107
rect 777 187 811 221
rect 777 77 811 111
<< pdiffc >>
rect 241 573 275 607
rect 241 468 275 502
rect 108 392 142 426
rect 194 379 228 413
rect 327 565 361 599
rect 327 472 361 506
rect 327 379 361 413
rect 415 566 449 600
rect 515 566 549 600
rect 601 474 635 508
rect 687 570 721 604
rect 687 458 721 492
rect 773 573 807 607
rect 773 472 807 506
rect 773 379 807 413
<< poly >>
rect 286 619 316 645
rect 372 619 402 645
rect 474 619 504 645
rect 560 619 590 645
rect 646 619 676 645
rect 732 619 762 645
rect 153 451 183 477
rect 153 302 183 367
rect 286 321 316 367
rect 35 286 183 302
rect 35 252 51 286
rect 85 272 183 286
rect 225 305 316 321
rect 85 252 110 272
rect 225 271 241 305
rect 275 285 316 305
rect 372 285 402 367
rect 474 335 504 367
rect 560 335 590 367
rect 646 335 676 367
rect 275 271 402 285
rect 225 255 402 271
rect 450 319 516 335
rect 450 285 466 319
rect 500 285 516 319
rect 450 269 516 285
rect 560 319 676 335
rect 560 285 576 319
rect 610 285 676 319
rect 560 269 676 285
rect 35 218 110 252
rect 286 233 316 255
rect 372 233 402 255
rect 458 233 488 269
rect 560 233 590 269
rect 646 233 676 269
rect 732 335 762 367
rect 732 319 798 335
rect 732 285 748 319
rect 782 285 798 319
rect 732 269 798 285
rect 732 233 762 269
rect 35 184 51 218
rect 85 184 110 218
rect 35 168 110 184
rect 80 146 110 168
rect 80 36 110 62
rect 286 39 316 65
rect 372 39 402 65
rect 458 39 488 65
rect 560 39 590 65
rect 646 39 676 65
rect 732 39 762 65
<< polycont >>
rect 51 252 85 286
rect 241 271 275 305
rect 466 285 500 319
rect 576 285 610 319
rect 748 285 782 319
rect 51 184 85 218
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 193 607 285 649
rect 193 573 241 607
rect 275 573 285 607
rect 193 502 285 573
rect 193 468 241 502
rect 275 468 285 502
rect 92 426 159 442
rect 92 392 108 426
rect 142 392 159 426
rect 92 351 159 392
rect 193 413 285 468
rect 193 379 194 413
rect 228 379 285 413
rect 193 363 285 379
rect 319 599 365 615
rect 319 565 327 599
rect 361 565 365 599
rect 319 524 365 565
rect 399 600 465 649
rect 399 566 415 600
rect 449 566 465 600
rect 399 558 465 566
rect 499 604 737 615
rect 499 600 687 604
rect 499 566 515 600
rect 549 570 687 600
rect 721 570 737 604
rect 549 566 737 570
rect 499 560 737 566
rect 319 508 637 524
rect 319 506 601 508
rect 319 472 327 506
rect 361 474 601 506
rect 635 474 637 508
rect 361 472 637 474
rect 319 458 637 472
rect 671 492 737 560
rect 671 458 687 492
rect 721 458 737 492
rect 773 607 823 649
rect 807 573 823 607
rect 773 506 823 573
rect 807 472 823 506
rect 319 413 369 458
rect 319 379 327 413
rect 361 379 369 413
rect 319 363 369 379
rect 119 321 159 351
rect 119 305 291 321
rect 17 286 85 302
rect 17 252 51 286
rect 17 218 85 252
rect 17 184 51 218
rect 17 168 85 184
rect 119 271 241 305
rect 275 271 291 305
rect 19 124 85 134
rect 19 90 35 124
rect 69 90 85 124
rect 19 17 85 90
rect 119 121 171 271
rect 119 87 121 121
rect 155 87 171 121
rect 119 71 171 87
rect 225 221 275 237
rect 325 229 369 363
rect 403 384 739 424
rect 403 319 516 384
rect 403 285 466 319
rect 500 285 516 319
rect 560 319 669 350
rect 560 285 576 319
rect 610 285 669 319
rect 703 329 739 384
rect 773 413 823 472
rect 807 379 823 413
rect 773 363 823 379
rect 703 319 798 329
rect 703 285 748 319
rect 782 285 798 319
rect 225 187 241 221
rect 225 111 275 187
rect 311 225 377 229
rect 311 191 327 225
rect 361 191 377 225
rect 311 153 377 191
rect 311 119 327 153
rect 361 119 377 153
rect 413 221 827 251
rect 447 217 601 221
rect 447 187 453 217
rect 225 77 241 111
rect 413 111 453 187
rect 587 187 601 217
rect 635 217 777 221
rect 635 187 637 217
rect 275 77 413 85
rect 447 77 453 111
rect 225 51 453 77
rect 487 149 503 183
rect 537 149 553 183
rect 487 107 553 149
rect 487 73 503 107
rect 537 73 553 107
rect 487 17 553 73
rect 587 111 637 187
rect 771 187 777 217
rect 811 187 827 221
rect 587 77 601 111
rect 635 77 637 111
rect 587 61 637 77
rect 671 149 687 183
rect 721 149 737 183
rect 671 107 737 149
rect 671 73 687 107
rect 721 73 737 107
rect 671 17 737 73
rect 771 111 827 187
rect 771 77 777 111
rect 811 77 827 111
rect 771 61 827 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21bai_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5202882
string GDS_START 5195074
<< end >>
