magic
tech sky130A
magscale 1 2
timestamp 1627202617
<< checkpaint >>
rect -1298 -1308 2494 1852
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1163 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 351 47 381 177
rect 435 47 465 177
rect 519 47 549 177
rect 603 47 633 177
rect 799 47 829 177
rect 883 47 913 177
rect 967 47 997 177
rect 1051 47 1081 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 351 297 381 497
rect 435 297 465 497
rect 519 297 549 497
rect 603 297 633 497
rect 799 297 829 497
rect 883 297 913 497
rect 967 297 997 497
rect 1051 297 1081 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 161 163 177
rect 109 127 119 161
rect 153 127 163 161
rect 109 47 163 127
rect 193 161 245 177
rect 193 127 203 161
rect 237 127 245 161
rect 193 93 245 127
rect 193 59 203 93
rect 237 59 245 93
rect 193 47 245 59
rect 299 93 351 177
rect 299 59 307 93
rect 341 59 351 93
rect 299 47 351 59
rect 381 161 435 177
rect 381 127 391 161
rect 425 127 435 161
rect 381 93 435 127
rect 381 59 391 93
rect 425 59 435 93
rect 381 47 435 59
rect 465 93 519 177
rect 465 59 475 93
rect 509 59 519 93
rect 465 47 519 59
rect 549 161 603 177
rect 549 127 559 161
rect 593 127 603 161
rect 549 93 603 127
rect 549 59 559 93
rect 593 59 603 93
rect 549 47 603 59
rect 633 93 689 177
rect 633 59 643 93
rect 677 59 689 93
rect 633 47 689 59
rect 743 161 799 177
rect 743 127 755 161
rect 789 127 799 161
rect 743 93 799 127
rect 743 59 755 93
rect 789 59 799 93
rect 743 47 799 59
rect 829 93 883 177
rect 829 59 839 93
rect 873 59 883 93
rect 829 47 883 59
rect 913 161 967 177
rect 913 127 923 161
rect 957 127 967 161
rect 913 93 967 127
rect 913 59 923 93
rect 957 59 967 93
rect 913 47 967 59
rect 997 93 1051 177
rect 997 59 1007 93
rect 1041 59 1051 93
rect 997 47 1051 59
rect 1081 161 1137 177
rect 1081 127 1091 161
rect 1125 127 1137 161
rect 1081 93 1137 127
rect 1081 59 1091 93
rect 1125 59 1137 93
rect 1081 47 1137 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 245 497
rect 193 451 203 485
rect 237 451 245 485
rect 193 417 245 451
rect 193 383 203 417
rect 237 383 245 417
rect 193 297 245 383
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 417 351 451
rect 299 383 307 417
rect 341 383 351 417
rect 299 297 351 383
rect 381 417 435 497
rect 381 383 391 417
rect 425 383 435 417
rect 381 349 435 383
rect 381 315 391 349
rect 425 315 435 349
rect 381 297 435 315
rect 465 477 519 497
rect 465 443 475 477
rect 509 443 519 477
rect 465 409 519 443
rect 465 375 475 409
rect 509 375 519 409
rect 465 341 519 375
rect 465 307 475 341
rect 509 307 519 341
rect 465 297 519 307
rect 549 485 603 497
rect 549 451 559 485
rect 593 451 603 485
rect 549 417 603 451
rect 549 383 559 417
rect 593 383 603 417
rect 549 297 603 383
rect 633 409 689 497
rect 633 375 643 409
rect 677 375 689 409
rect 633 341 689 375
rect 633 307 643 341
rect 677 307 689 341
rect 633 297 689 307
rect 743 407 799 497
rect 743 373 755 407
rect 789 373 799 407
rect 743 339 799 373
rect 743 305 755 339
rect 789 305 799 339
rect 743 297 799 305
rect 829 485 883 497
rect 829 451 839 485
rect 873 451 883 485
rect 829 417 883 451
rect 829 383 839 417
rect 873 383 883 417
rect 829 297 883 383
rect 913 475 967 497
rect 913 441 923 475
rect 957 441 967 475
rect 913 407 967 441
rect 913 373 923 407
rect 957 373 967 407
rect 913 339 967 373
rect 913 305 923 339
rect 957 305 967 339
rect 913 297 967 305
rect 997 485 1051 497
rect 997 451 1007 485
rect 1041 451 1051 485
rect 997 417 1051 451
rect 997 383 1007 417
rect 1041 383 1051 417
rect 997 297 1051 383
rect 1081 475 1137 497
rect 1081 441 1091 475
rect 1125 441 1137 475
rect 1081 407 1137 441
rect 1081 373 1091 407
rect 1125 373 1137 407
rect 1081 339 1137 373
rect 1081 305 1091 339
rect 1125 305 1137 339
rect 1081 297 1137 305
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 127 153 161
rect 203 127 237 161
rect 203 59 237 93
rect 307 59 341 93
rect 391 127 425 161
rect 391 59 425 93
rect 475 59 509 93
rect 559 127 593 161
rect 559 59 593 93
rect 643 59 677 93
rect 755 127 789 161
rect 755 59 789 93
rect 839 59 873 93
rect 923 127 957 161
rect 923 59 957 93
rect 1007 59 1041 93
rect 1091 127 1125 161
rect 1091 59 1125 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 307 451 341 485
rect 307 383 341 417
rect 391 383 425 417
rect 391 315 425 349
rect 475 443 509 477
rect 475 375 509 409
rect 475 307 509 341
rect 559 451 593 485
rect 559 383 593 417
rect 643 375 677 409
rect 643 307 677 341
rect 755 373 789 407
rect 755 305 789 339
rect 839 451 873 485
rect 839 383 873 417
rect 923 441 957 475
rect 923 373 957 407
rect 923 305 957 339
rect 1007 451 1041 485
rect 1007 383 1041 417
rect 1091 441 1125 475
rect 1091 373 1125 407
rect 1091 305 1125 339
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 351 497 381 523
rect 435 497 465 523
rect 519 497 549 523
rect 603 497 633 523
rect 799 497 829 523
rect 883 497 913 523
rect 967 497 997 523
rect 1051 497 1081 523
rect 79 262 109 297
rect 163 262 193 297
rect 79 261 193 262
rect 351 261 381 297
rect 435 261 465 297
rect 21 249 193 261
rect 21 215 38 249
rect 72 215 193 249
rect 21 203 193 215
rect 300 249 465 261
rect 300 215 316 249
rect 350 215 412 249
rect 446 215 465 249
rect 300 205 465 215
rect 300 203 381 205
rect 79 200 193 203
rect 79 177 109 200
rect 163 177 193 200
rect 351 177 381 203
rect 435 177 465 205
rect 519 262 549 297
rect 603 262 633 297
rect 519 249 669 262
rect 799 259 829 297
rect 883 259 913 297
rect 519 215 535 249
rect 569 215 619 249
rect 653 215 669 249
rect 519 202 669 215
rect 756 249 913 259
rect 756 215 772 249
rect 806 215 847 249
rect 881 215 913 249
rect 519 177 549 202
rect 603 177 633 202
rect 756 198 913 215
rect 799 177 829 198
rect 883 177 913 198
rect 967 259 997 297
rect 1051 259 1081 297
rect 967 249 1147 259
rect 967 215 1008 249
rect 1042 215 1097 249
rect 1131 215 1147 249
rect 967 205 1147 215
rect 967 177 997 205
rect 1051 177 1081 205
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 519 21 549 47
rect 603 21 633 47
rect 799 21 829 47
rect 883 21 913 47
rect 967 21 997 47
rect 1051 21 1081 47
<< polycont >>
rect 38 215 72 249
rect 316 215 350 249
rect 412 215 446 249
rect 535 215 569 249
rect 619 215 653 249
rect 772 215 806 249
rect 847 215 881 249
rect 1008 215 1042 249
rect 1097 215 1131 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 349 69 383
rect 17 315 35 349
rect 17 299 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 253 527
rect 237 451 253 485
rect 203 417 253 451
rect 237 383 253 417
rect 203 367 253 383
rect 291 485 509 493
rect 291 451 307 485
rect 341 477 509 485
rect 341 459 475 477
rect 291 417 341 451
rect 291 383 307 417
rect 291 367 341 383
rect 375 417 441 425
rect 375 383 391 417
rect 425 383 441 417
rect 103 315 119 349
rect 153 333 169 349
rect 375 349 441 383
rect 375 333 391 349
rect 153 315 391 333
rect 425 315 441 349
rect 103 301 441 315
rect 122 289 441 301
rect 475 409 509 443
rect 475 341 509 375
rect 543 485 889 493
rect 543 451 559 485
rect 593 459 839 485
rect 593 451 609 459
rect 543 417 609 451
rect 823 451 839 459
rect 873 451 889 485
rect 543 383 559 417
rect 593 383 609 417
rect 543 367 609 383
rect 643 409 693 425
rect 677 375 693 409
rect 643 341 693 375
rect 509 307 643 323
rect 677 307 693 341
rect 475 289 693 307
rect 739 407 789 425
rect 739 373 755 407
rect 739 339 789 373
rect 823 417 889 451
rect 823 383 839 417
rect 873 383 889 417
rect 823 367 889 383
rect 923 475 957 493
rect 923 407 957 441
rect 739 305 755 339
rect 923 339 957 373
rect 991 485 1057 527
rect 991 451 1007 485
rect 1041 451 1057 485
rect 991 417 1057 451
rect 991 383 1007 417
rect 1041 383 1057 417
rect 991 357 1057 383
rect 1091 475 1141 493
rect 1125 441 1141 475
rect 1091 407 1141 441
rect 1125 373 1141 407
rect 789 305 923 323
rect 1091 339 1141 373
rect 957 305 1091 323
rect 1125 305 1141 339
rect 739 289 1141 305
rect 21 249 88 255
rect 21 215 38 249
rect 72 215 88 249
rect 17 161 69 181
rect 122 177 169 289
rect 300 249 465 255
rect 300 215 316 249
rect 350 215 412 249
rect 446 215 465 249
rect 519 249 716 255
rect 519 215 535 249
rect 569 215 619 249
rect 653 215 716 249
rect 756 249 908 255
rect 756 215 772 249
rect 806 215 847 249
rect 881 215 908 249
rect 944 249 1179 255
rect 944 215 1008 249
rect 1042 215 1097 249
rect 1131 215 1179 249
rect 17 127 35 161
rect 103 161 169 177
rect 103 127 119 161
rect 153 127 169 161
rect 203 161 1141 181
rect 237 147 391 161
rect 237 127 253 147
rect 17 93 69 127
rect 203 93 253 127
rect 375 127 391 147
rect 425 147 559 161
rect 425 127 441 147
rect 17 59 35 93
rect 69 59 203 93
rect 237 59 253 93
rect 17 51 253 59
rect 291 93 341 109
rect 291 59 307 93
rect 291 17 341 59
rect 375 93 441 127
rect 543 127 559 147
rect 593 147 755 161
rect 593 127 609 147
rect 375 59 391 93
rect 425 59 441 93
rect 375 51 441 59
rect 475 93 509 109
rect 475 17 509 59
rect 543 93 609 127
rect 739 127 755 147
rect 789 147 923 161
rect 789 127 805 147
rect 543 59 559 93
rect 593 59 609 93
rect 543 51 609 59
rect 643 93 690 109
rect 677 59 690 93
rect 643 17 690 59
rect 739 93 805 127
rect 907 127 923 147
rect 957 147 1091 161
rect 957 127 973 147
rect 739 59 755 93
rect 789 59 805 93
rect 739 51 805 59
rect 839 93 873 109
rect 839 17 873 59
rect 907 93 973 127
rect 1075 127 1091 147
rect 1125 127 1141 161
rect 907 59 923 93
rect 957 59 973 93
rect 907 51 973 59
rect 1007 93 1041 109
rect 1007 17 1041 59
rect 1075 93 1141 127
rect 1075 59 1091 93
rect 1125 59 1141 93
rect 1075 51 1141 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 1142 221 1176 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 1050 221 1084 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 958 221 992 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 866 221 900 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 774 221 808 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 586 221 620 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 310 221 344 255 0 FreeSans 250 0 0 0 A4
port 4 nsew signal input
flabel locali s 402 221 436 255 0 FreeSans 250 0 0 0 A4
port 4 nsew signal input
flabel locali s 122 289 156 323 0 FreeSans 250 0 0 0 Y
port 10 nsew signal output
flabel locali s 122 153 156 187 0 FreeSans 250 0 0 0 Y
port 10 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 Y
port 10 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 B1
port 5 nsew signal input
flabel locali s 678 221 712 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o41ai_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 3452246
string GDS_START 3441202
string path 0.000 0.000 29.900 0.000 
<< end >>
