magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
rect 877 321 1276 331
<< pwell >>
rect 1326 241 1605 250
rect 891 229 1605 241
rect 359 203 1605 229
rect 23 49 1605 203
rect 0 0 1632 49
<< scnmos >>
rect 102 93 132 177
rect 219 93 249 177
rect 438 119 468 203
rect 524 119 554 203
rect 596 119 626 203
rect 704 119 734 203
rect 776 119 806 203
rect 970 47 1000 215
rect 1042 47 1072 215
rect 1157 131 1187 215
rect 1405 56 1435 224
rect 1494 56 1524 224
<< scpmoshvt >>
rect 102 483 132 611
rect 188 483 218 611
rect 426 481 456 609
rect 566 481 596 609
rect 638 481 668 609
rect 743 525 773 609
rect 861 525 891 609
rect 966 357 996 609
rect 1052 357 1082 609
rect 1157 357 1187 485
rect 1399 367 1429 619
rect 1485 367 1515 619
<< ndiff >>
rect 49 152 102 177
rect 49 118 57 152
rect 91 118 102 152
rect 49 93 102 118
rect 132 152 219 177
rect 132 118 159 152
rect 193 118 219 152
rect 132 93 219 118
rect 249 152 302 177
rect 249 118 260 152
rect 294 118 302 152
rect 249 93 302 118
rect 385 178 438 203
rect 385 144 393 178
rect 427 144 438 178
rect 385 119 438 144
rect 468 172 524 203
rect 468 138 479 172
rect 513 138 524 172
rect 468 119 524 138
rect 554 119 596 203
rect 626 177 704 203
rect 626 143 648 177
rect 682 143 704 177
rect 626 119 704 143
rect 734 119 776 203
rect 806 165 863 203
rect 806 131 817 165
rect 851 131 863 165
rect 806 119 863 131
rect 917 165 970 215
rect 917 131 925 165
rect 959 131 970 165
rect 917 93 970 131
rect 917 59 925 93
rect 959 59 970 93
rect 917 47 970 59
rect 1000 47 1042 215
rect 1072 131 1157 215
rect 1187 191 1240 215
rect 1187 157 1198 191
rect 1232 157 1240 191
rect 1187 131 1240 157
rect 1352 212 1405 224
rect 1352 178 1360 212
rect 1394 178 1405 212
rect 1072 97 1129 131
rect 1072 63 1083 97
rect 1117 63 1129 97
rect 1072 47 1129 63
rect 1352 102 1405 178
rect 1352 68 1360 102
rect 1394 68 1405 102
rect 1352 56 1405 68
rect 1435 196 1494 224
rect 1435 162 1449 196
rect 1483 162 1494 196
rect 1435 102 1494 162
rect 1435 68 1449 102
rect 1483 68 1494 102
rect 1435 56 1494 68
rect 1524 212 1579 224
rect 1524 178 1537 212
rect 1571 178 1579 212
rect 1524 102 1579 178
rect 1524 68 1537 102
rect 1571 68 1579 102
rect 1524 56 1579 68
<< pdiff >>
rect 49 599 102 611
rect 49 565 57 599
rect 91 565 102 599
rect 49 529 102 565
rect 49 495 57 529
rect 91 495 102 529
rect 49 483 102 495
rect 132 603 188 611
rect 132 569 143 603
rect 177 569 188 603
rect 132 535 188 569
rect 132 501 143 535
rect 177 501 188 535
rect 132 483 188 501
rect 218 597 271 611
rect 218 563 229 597
rect 263 563 271 597
rect 218 529 271 563
rect 218 495 229 529
rect 263 495 271 529
rect 218 483 271 495
rect 373 531 426 609
rect 373 497 381 531
rect 415 497 426 531
rect 373 481 426 497
rect 456 576 566 609
rect 456 542 521 576
rect 555 542 566 576
rect 456 481 566 542
rect 596 481 638 609
rect 668 531 743 609
rect 668 497 679 531
rect 713 525 743 531
rect 773 525 861 609
rect 891 578 966 609
rect 891 544 921 578
rect 955 544 966 578
rect 891 525 966 544
rect 713 497 721 525
rect 668 481 721 497
rect 913 357 966 525
rect 996 596 1052 609
rect 996 562 1007 596
rect 1041 562 1052 596
rect 996 510 1052 562
rect 996 476 1007 510
rect 1041 476 1052 510
rect 996 357 1052 476
rect 1082 567 1135 609
rect 1082 533 1093 567
rect 1127 533 1135 567
rect 1082 485 1135 533
rect 1082 357 1157 485
rect 1187 411 1240 485
rect 1187 377 1198 411
rect 1232 377 1240 411
rect 1187 357 1240 377
rect 1346 415 1399 619
rect 1346 381 1354 415
rect 1388 381 1399 415
rect 1346 367 1399 381
rect 1429 575 1485 619
rect 1429 541 1440 575
rect 1474 541 1485 575
rect 1429 367 1485 541
rect 1515 599 1568 619
rect 1515 565 1526 599
rect 1560 565 1568 599
rect 1515 503 1568 565
rect 1515 469 1526 503
rect 1560 469 1568 503
rect 1515 413 1568 469
rect 1515 379 1526 413
rect 1560 379 1568 413
rect 1515 367 1568 379
<< ndiffc >>
rect 57 118 91 152
rect 159 118 193 152
rect 260 118 294 152
rect 393 144 427 178
rect 479 138 513 172
rect 648 143 682 177
rect 817 131 851 165
rect 925 131 959 165
rect 925 59 959 93
rect 1198 157 1232 191
rect 1360 178 1394 212
rect 1083 63 1117 97
rect 1360 68 1394 102
rect 1449 162 1483 196
rect 1449 68 1483 102
rect 1537 178 1571 212
rect 1537 68 1571 102
<< pdiffc >>
rect 57 565 91 599
rect 57 495 91 529
rect 143 569 177 603
rect 143 501 177 535
rect 229 563 263 597
rect 229 495 263 529
rect 381 497 415 531
rect 521 542 555 576
rect 679 497 713 531
rect 921 544 955 578
rect 1007 562 1041 596
rect 1007 476 1041 510
rect 1093 533 1127 567
rect 1198 377 1232 411
rect 1354 381 1388 415
rect 1440 541 1474 575
rect 1526 565 1560 599
rect 1526 469 1560 503
rect 1526 379 1560 413
<< poly >>
rect 102 611 132 637
rect 188 611 218 637
rect 426 609 456 635
rect 566 609 596 635
rect 638 609 668 635
rect 743 609 773 635
rect 861 609 891 635
rect 966 609 996 635
rect 1052 609 1082 635
rect 1399 619 1429 645
rect 1485 619 1515 645
rect 102 333 132 483
rect 188 451 218 483
rect 743 493 773 525
rect 188 435 272 451
rect 188 401 204 435
rect 238 401 272 435
rect 426 424 456 481
rect 188 385 272 401
rect 102 317 177 333
rect 102 283 127 317
rect 161 283 177 317
rect 102 249 177 283
rect 102 215 127 249
rect 161 215 177 249
rect 102 199 177 215
rect 219 229 272 385
rect 399 408 468 424
rect 399 374 415 408
rect 449 374 468 408
rect 566 405 596 481
rect 399 340 468 374
rect 399 306 415 340
rect 449 306 468 340
rect 399 290 468 306
rect 219 199 370 229
rect 438 203 468 290
rect 518 389 596 405
rect 518 355 534 389
rect 568 375 596 389
rect 638 379 668 481
rect 743 477 819 493
rect 743 443 769 477
rect 803 443 819 477
rect 743 427 819 443
rect 861 385 891 525
rect 568 355 584 375
rect 518 339 584 355
rect 638 349 734 379
rect 518 271 554 339
rect 524 203 554 271
rect 596 275 662 291
rect 596 241 612 275
rect 646 241 662 275
rect 596 225 662 241
rect 596 203 626 225
rect 704 203 734 349
rect 797 369 891 385
rect 797 335 813 369
rect 847 355 891 369
rect 1157 485 1187 511
rect 847 335 863 355
rect 797 301 863 335
rect 966 303 996 357
rect 1052 308 1082 357
rect 1157 325 1187 357
rect 1156 309 1222 325
rect 797 281 813 301
rect 776 267 813 281
rect 847 267 863 301
rect 776 251 863 267
rect 905 287 996 303
rect 905 253 921 287
rect 955 267 996 287
rect 1042 292 1108 308
rect 955 253 1000 267
rect 776 203 806 251
rect 905 237 1000 253
rect 970 215 1000 237
rect 1042 258 1058 292
rect 1092 258 1108 292
rect 1156 275 1172 309
rect 1206 275 1222 309
rect 1399 287 1429 367
rect 1485 312 1515 367
rect 1477 296 1552 312
rect 1156 259 1222 275
rect 1264 271 1435 287
rect 1042 242 1108 258
rect 1042 215 1072 242
rect 1157 215 1187 259
rect 1264 237 1280 271
rect 1314 257 1435 271
rect 1314 237 1330 257
rect 102 177 132 199
rect 219 177 249 199
rect 102 67 132 93
rect 219 67 249 93
rect 340 51 370 199
rect 438 93 468 119
rect 524 93 554 119
rect 596 93 626 119
rect 704 51 734 119
rect 776 93 806 119
rect 340 21 734 51
rect 1264 203 1330 237
rect 1405 224 1435 257
rect 1477 262 1493 296
rect 1527 262 1552 296
rect 1477 246 1552 262
rect 1494 224 1524 246
rect 1264 169 1280 203
rect 1314 169 1330 203
rect 1264 153 1330 169
rect 1157 105 1187 131
rect 970 21 1000 47
rect 1042 21 1072 47
rect 1405 30 1435 56
rect 1494 30 1524 56
<< polycont >>
rect 204 401 238 435
rect 127 283 161 317
rect 127 215 161 249
rect 415 374 449 408
rect 415 306 449 340
rect 534 355 568 389
rect 769 443 803 477
rect 612 241 646 275
rect 813 335 847 369
rect 813 267 847 301
rect 921 253 955 287
rect 1058 258 1092 292
rect 1172 275 1206 309
rect 1280 237 1314 271
rect 1493 262 1527 296
rect 1280 169 1314 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 41 599 100 615
rect 41 565 57 599
rect 91 565 100 599
rect 41 529 100 565
rect 41 495 57 529
rect 91 495 100 529
rect 41 451 100 495
rect 134 603 179 649
rect 134 569 143 603
rect 177 569 179 603
rect 134 535 179 569
rect 134 501 143 535
rect 177 501 179 535
rect 134 485 179 501
rect 213 597 485 615
rect 213 563 229 597
rect 263 581 485 597
rect 263 563 309 581
rect 213 529 309 563
rect 213 495 229 529
rect 263 495 309 529
rect 213 485 309 495
rect 41 435 241 451
rect 41 401 204 435
rect 238 401 241 435
rect 41 385 241 401
rect 41 165 91 385
rect 125 317 177 351
rect 125 283 127 317
rect 161 283 177 317
rect 125 249 177 283
rect 125 215 127 249
rect 161 215 177 249
rect 125 199 177 215
rect 275 168 309 485
rect 345 531 417 547
rect 345 497 381 531
rect 415 497 417 531
rect 345 477 417 497
rect 451 492 485 581
rect 519 576 571 649
rect 519 542 521 576
rect 555 542 571 576
rect 519 526 571 542
rect 605 581 803 615
rect 605 492 639 581
rect 345 256 379 477
rect 451 458 639 492
rect 673 531 717 547
rect 673 497 679 531
rect 713 497 717 531
rect 673 477 717 497
rect 413 408 469 424
rect 413 374 415 408
rect 449 374 469 408
rect 413 340 469 374
rect 413 306 415 340
rect 449 306 469 340
rect 413 290 469 306
rect 518 389 568 405
rect 518 355 534 389
rect 518 256 568 355
rect 345 222 568 256
rect 605 291 639 458
rect 605 275 649 291
rect 605 241 612 275
rect 646 241 649 275
rect 605 225 649 241
rect 683 233 717 477
rect 751 477 803 581
rect 905 578 965 649
rect 905 544 921 578
rect 955 544 965 578
rect 905 528 965 544
rect 999 596 1043 612
rect 999 562 1007 596
rect 1041 562 1043 596
rect 999 510 1043 562
rect 1077 567 1143 649
rect 1077 533 1093 567
rect 1127 533 1143 567
rect 1424 575 1490 649
rect 1424 541 1440 575
rect 1474 541 1490 575
rect 1424 533 1490 541
rect 1524 599 1615 615
rect 1524 565 1526 599
rect 1560 565 1615 599
rect 999 494 1007 510
rect 751 443 769 477
rect 751 427 803 443
rect 837 476 1007 494
rect 1041 499 1043 510
rect 1524 503 1615 565
rect 1041 476 1490 499
rect 837 465 1490 476
rect 837 460 1162 465
rect 837 385 871 460
rect 797 369 871 385
rect 797 335 813 369
rect 847 335 871 369
rect 797 301 871 335
rect 797 267 813 301
rect 847 267 871 301
rect 905 287 955 303
rect 905 253 921 287
rect 905 233 955 253
rect 989 292 1094 424
rect 989 258 1058 292
rect 1092 258 1094 292
rect 989 242 1094 258
rect 1128 325 1162 460
rect 1198 411 1276 427
rect 1232 377 1276 411
rect 1198 361 1276 377
rect 1128 309 1206 325
rect 1128 275 1172 309
rect 1128 259 1206 275
rect 1242 287 1276 361
rect 1350 415 1411 431
rect 1350 381 1354 415
rect 1388 381 1411 415
rect 1242 271 1316 287
rect 345 217 436 222
rect 377 178 436 217
rect 683 199 955 233
rect 683 191 717 199
rect 41 152 107 165
rect 41 118 57 152
rect 91 118 107 152
rect 41 102 107 118
rect 143 152 209 165
rect 143 118 159 152
rect 193 118 209 152
rect 143 17 209 118
rect 244 152 310 168
rect 244 118 260 152
rect 294 118 310 152
rect 377 144 393 178
rect 427 144 436 178
rect 377 128 436 144
rect 470 172 529 188
rect 470 138 479 172
rect 513 138 529 172
rect 244 102 310 118
rect 470 17 529 138
rect 632 177 717 191
rect 632 143 648 177
rect 682 143 717 177
rect 1128 165 1162 259
rect 1242 237 1280 271
rect 1314 237 1316 271
rect 1242 207 1316 237
rect 632 127 717 143
rect 801 131 817 165
rect 851 131 867 165
rect 801 17 867 131
rect 909 131 925 165
rect 959 131 1162 165
rect 1196 203 1316 207
rect 1196 191 1280 203
rect 1196 157 1198 191
rect 1232 169 1280 191
rect 1314 169 1316 203
rect 1232 157 1316 169
rect 1196 141 1316 157
rect 1350 212 1411 381
rect 1445 312 1490 465
rect 1524 469 1526 503
rect 1560 469 1615 503
rect 1524 413 1615 469
rect 1524 379 1526 413
rect 1560 379 1615 413
rect 1524 348 1615 379
rect 1445 296 1529 312
rect 1445 262 1493 296
rect 1527 262 1529 296
rect 1445 246 1529 262
rect 1563 212 1615 348
rect 1350 178 1360 212
rect 1394 178 1411 212
rect 909 93 975 131
rect 1350 102 1411 178
rect 909 59 925 93
rect 959 59 975 93
rect 909 51 975 59
rect 1067 63 1083 97
rect 1117 63 1133 97
rect 1067 17 1133 63
rect 1350 68 1360 102
rect 1394 68 1411 102
rect 1350 52 1411 68
rect 1445 196 1487 212
rect 1445 162 1449 196
rect 1483 162 1487 196
rect 1445 102 1487 162
rect 1445 68 1449 102
rect 1483 68 1487 102
rect 1445 17 1487 68
rect 1521 178 1537 212
rect 1571 178 1615 212
rect 1521 102 1615 178
rect 1521 68 1537 102
rect 1571 68 1615 102
rect 1521 52 1615 68
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrbp_1
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1375 94 1409 128 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1375 168 1409 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1375 390 1409 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4305804
string GDS_START 4292276
<< end >>
