magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3122 1975
<< nwell >>
rect -38 331 1862 704
<< pwell >>
rect 353 241 936 245
rect 1 229 936 241
rect 1 157 1484 229
rect 1 49 1794 157
rect 0 0 1824 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 432 135 462 219
rect 557 51 587 219
rect 643 51 673 219
rect 751 51 781 219
rect 823 51 853 219
rect 1037 119 1067 203
rect 1109 119 1139 203
rect 1195 119 1225 203
rect 1289 119 1319 203
rect 1375 119 1405 203
rect 1599 47 1629 131
rect 1685 47 1715 131
<< scpmoshvt >>
rect 80 367 110 619
rect 167 367 197 619
rect 448 367 478 495
rect 557 367 587 619
rect 643 367 673 619
rect 760 367 790 619
rect 846 367 876 619
rect 951 503 981 587
rect 1069 503 1099 587
rect 1174 459 1204 587
rect 1246 459 1276 587
rect 1398 459 1428 587
rect 1613 483 1643 611
rect 1699 483 1729 611
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 93 80 169
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 204 166 215
rect 110 170 121 204
rect 155 170 166 204
rect 110 101 166 170
rect 110 67 121 101
rect 155 67 166 101
rect 110 47 166 67
rect 196 203 249 215
rect 196 169 207 203
rect 241 169 249 203
rect 196 93 249 169
rect 379 194 432 219
rect 379 160 387 194
rect 421 160 432 194
rect 379 135 432 160
rect 462 135 557 219
rect 196 59 207 93
rect 241 59 249 93
rect 196 47 249 59
rect 484 93 557 135
rect 484 59 496 93
rect 530 59 557 93
rect 484 51 557 59
rect 587 167 643 219
rect 587 133 598 167
rect 632 133 643 167
rect 587 95 643 133
rect 587 61 598 95
rect 632 61 643 95
rect 587 51 643 61
rect 673 167 751 219
rect 673 133 698 167
rect 732 133 751 167
rect 673 93 751 133
rect 673 59 698 93
rect 732 59 751 93
rect 673 51 751 59
rect 781 51 823 219
rect 853 187 910 219
rect 853 153 864 187
rect 898 153 910 187
rect 853 101 910 153
rect 984 178 1037 203
rect 984 144 992 178
rect 1026 144 1037 178
rect 984 119 1037 144
rect 1067 119 1109 203
rect 1139 178 1195 203
rect 1139 144 1150 178
rect 1184 144 1195 178
rect 1139 119 1195 144
rect 1225 119 1289 203
rect 1319 178 1375 203
rect 1319 144 1330 178
rect 1364 144 1375 178
rect 1319 119 1375 144
rect 1405 178 1458 203
rect 1405 144 1416 178
rect 1450 144 1458 178
rect 1405 119 1458 144
rect 853 67 864 101
rect 898 67 910 101
rect 853 51 910 67
rect 1546 106 1599 131
rect 1546 72 1554 106
rect 1588 72 1599 106
rect 1546 47 1599 72
rect 1629 106 1685 131
rect 1629 72 1640 106
rect 1674 72 1685 106
rect 1629 47 1685 72
rect 1715 106 1768 131
rect 1715 72 1726 106
rect 1760 72 1768 106
rect 1715 47 1768 72
<< pdiff >>
rect 27 607 80 619
rect 27 573 35 607
rect 69 573 80 607
rect 27 509 80 573
rect 27 475 35 509
rect 69 475 80 509
rect 27 413 80 475
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 599 167 619
rect 110 565 122 599
rect 156 565 167 599
rect 110 502 167 565
rect 110 468 122 502
rect 156 468 167 502
rect 110 409 167 468
rect 110 375 122 409
rect 156 375 167 409
rect 110 367 167 375
rect 197 607 250 619
rect 197 573 208 607
rect 242 573 250 607
rect 197 509 250 573
rect 500 575 557 619
rect 500 541 508 575
rect 542 541 557 575
rect 197 475 208 509
rect 242 475 250 509
rect 500 495 557 541
rect 197 413 250 475
rect 197 379 208 413
rect 242 379 250 413
rect 197 367 250 379
rect 391 414 448 495
rect 391 380 403 414
rect 437 380 448 414
rect 391 367 448 380
rect 478 367 557 495
rect 587 599 643 619
rect 587 565 598 599
rect 632 565 643 599
rect 587 494 643 565
rect 587 460 598 494
rect 632 460 643 494
rect 587 367 643 460
rect 673 611 760 619
rect 673 577 699 611
rect 733 577 760 611
rect 673 493 760 577
rect 673 459 699 493
rect 733 459 760 493
rect 673 367 760 459
rect 790 599 846 619
rect 790 565 801 599
rect 835 565 846 599
rect 790 506 846 565
rect 790 472 801 506
rect 835 472 846 506
rect 790 409 846 472
rect 790 375 801 409
rect 835 375 846 409
rect 790 367 846 375
rect 876 607 929 619
rect 876 573 887 607
rect 921 587 929 607
rect 921 573 951 587
rect 876 524 951 573
rect 876 490 887 524
rect 921 503 951 524
rect 981 503 1069 587
rect 1099 507 1174 587
rect 1099 503 1129 507
rect 921 490 929 503
rect 876 445 929 490
rect 876 411 887 445
rect 921 411 929 445
rect 876 367 929 411
rect 1121 473 1129 503
rect 1163 473 1174 507
rect 1121 459 1174 473
rect 1204 459 1246 587
rect 1276 579 1398 587
rect 1276 545 1289 579
rect 1323 545 1398 579
rect 1276 459 1398 545
rect 1428 512 1485 587
rect 1428 478 1443 512
rect 1477 478 1485 512
rect 1560 578 1613 611
rect 1560 544 1568 578
rect 1602 544 1613 578
rect 1560 483 1613 544
rect 1643 570 1699 611
rect 1643 536 1654 570
rect 1688 536 1699 570
rect 1643 483 1699 536
rect 1729 597 1786 611
rect 1729 563 1741 597
rect 1775 563 1786 597
rect 1729 529 1786 563
rect 1729 495 1741 529
rect 1775 495 1786 529
rect 1729 483 1786 495
rect 1428 459 1485 478
<< ndiffc >>
rect 35 169 69 203
rect 35 59 69 93
rect 121 170 155 204
rect 121 67 155 101
rect 207 169 241 203
rect 387 160 421 194
rect 207 59 241 93
rect 496 59 530 93
rect 598 133 632 167
rect 598 61 632 95
rect 698 133 732 167
rect 698 59 732 93
rect 864 153 898 187
rect 992 144 1026 178
rect 1150 144 1184 178
rect 1330 144 1364 178
rect 1416 144 1450 178
rect 864 67 898 101
rect 1554 72 1588 106
rect 1640 72 1674 106
rect 1726 72 1760 106
<< pdiffc >>
rect 35 573 69 607
rect 35 475 69 509
rect 35 379 69 413
rect 122 565 156 599
rect 122 468 156 502
rect 122 375 156 409
rect 208 573 242 607
rect 508 541 542 575
rect 208 475 242 509
rect 208 379 242 413
rect 403 380 437 414
rect 598 565 632 599
rect 598 460 632 494
rect 699 577 733 611
rect 699 459 733 493
rect 801 565 835 599
rect 801 472 835 506
rect 801 375 835 409
rect 887 573 921 607
rect 887 490 921 524
rect 887 411 921 445
rect 1129 473 1163 507
rect 1289 545 1323 579
rect 1443 478 1477 512
rect 1568 544 1602 578
rect 1654 536 1688 570
rect 1741 563 1775 597
rect 1741 495 1775 529
<< poly >>
rect 80 619 110 645
rect 167 619 197 645
rect 557 619 587 645
rect 643 619 673 645
rect 760 619 790 645
rect 846 619 876 645
rect 448 495 478 521
rect 951 587 981 613
rect 1069 587 1099 613
rect 1174 587 1204 613
rect 1246 587 1276 613
rect 1398 587 1428 613
rect 1613 611 1643 637
rect 1699 611 1729 637
rect 80 326 110 367
rect 167 326 197 367
rect 448 337 478 367
rect 557 337 587 367
rect 643 337 673 367
rect 760 343 790 367
rect 80 310 266 326
rect 80 276 216 310
rect 250 276 266 310
rect 80 260 266 276
rect 448 291 673 337
rect 448 271 555 291
rect 80 215 110 260
rect 166 215 196 260
rect 432 257 555 271
rect 589 257 623 291
rect 657 257 673 291
rect 715 319 790 343
rect 715 285 731 319
rect 765 313 790 319
rect 765 285 781 313
rect 846 307 876 367
rect 951 357 981 503
rect 1069 471 1099 503
rect 1023 455 1099 471
rect 1023 421 1039 455
rect 1073 421 1099 455
rect 1023 405 1099 421
rect 1174 369 1204 459
rect 1147 363 1204 369
rect 951 341 1027 357
rect 951 327 977 341
rect 961 307 977 327
rect 1011 321 1027 341
rect 1109 339 1204 363
rect 1246 405 1276 459
rect 1398 424 1428 459
rect 1613 451 1643 483
rect 1577 435 1643 451
rect 1367 408 1433 424
rect 1246 389 1319 405
rect 1246 355 1269 389
rect 1303 355 1319 389
rect 1246 339 1319 355
rect 1109 333 1177 339
rect 1011 307 1067 321
rect 715 269 781 285
rect 843 291 909 307
rect 961 291 1067 307
rect 843 271 859 291
rect 432 241 673 257
rect 432 219 462 241
rect 557 219 587 241
rect 643 219 673 241
rect 751 219 781 269
rect 823 257 859 271
rect 893 257 909 291
rect 823 241 909 257
rect 823 219 853 241
rect 432 109 462 135
rect 1037 203 1067 291
rect 1109 203 1139 333
rect 1181 275 1247 291
rect 1181 241 1197 275
rect 1231 241 1247 275
rect 1181 225 1247 241
rect 1195 203 1225 225
rect 1289 203 1319 339
rect 1367 374 1383 408
rect 1417 374 1433 408
rect 1367 340 1433 374
rect 1367 306 1383 340
rect 1417 306 1433 340
rect 1577 401 1593 435
rect 1627 401 1643 435
rect 1577 367 1643 401
rect 1577 333 1593 367
rect 1627 333 1643 367
rect 1577 317 1643 333
rect 1367 290 1433 306
rect 1375 203 1405 290
rect 1599 183 1629 317
rect 1699 302 1729 483
rect 1501 153 1629 183
rect 1037 93 1067 119
rect 1109 51 1139 119
rect 1195 93 1225 119
rect 1289 93 1319 119
rect 1375 93 1405 119
rect 1501 51 1531 153
rect 1599 131 1629 153
rect 1685 286 1751 302
rect 1685 252 1701 286
rect 1735 252 1751 286
rect 1685 218 1751 252
rect 1685 184 1701 218
rect 1735 184 1751 218
rect 1685 168 1751 184
rect 1685 131 1715 168
rect 80 21 110 47
rect 166 21 196 47
rect 557 25 587 51
rect 643 25 673 51
rect 751 25 781 51
rect 823 25 853 51
rect 1109 21 1531 51
rect 1599 21 1629 47
rect 1685 21 1715 47
<< polycont >>
rect 216 276 250 310
rect 555 257 589 291
rect 623 257 657 291
rect 731 285 765 319
rect 1039 421 1073 455
rect 977 307 1011 341
rect 1269 355 1303 389
rect 859 257 893 291
rect 1197 241 1231 275
rect 1383 374 1417 408
rect 1383 306 1417 340
rect 1593 401 1627 435
rect 1593 333 1627 367
rect 1701 252 1735 286
rect 1701 184 1735 218
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 19 607 77 649
rect 19 573 35 607
rect 69 573 77 607
rect 19 509 77 573
rect 19 475 35 509
rect 69 475 77 509
rect 19 413 77 475
rect 19 379 35 413
rect 69 379 77 413
rect 19 363 77 379
rect 111 599 166 615
rect 111 565 122 599
rect 156 565 166 599
rect 111 502 166 565
rect 111 468 122 502
rect 156 468 166 502
rect 111 409 166 468
rect 111 375 122 409
rect 156 375 166 409
rect 19 203 77 219
rect 19 169 35 203
rect 69 169 77 203
rect 19 93 77 169
rect 19 59 35 93
rect 69 59 77 93
rect 19 17 77 59
rect 111 204 166 375
rect 200 607 258 649
rect 200 573 208 607
rect 242 573 258 607
rect 200 509 258 573
rect 492 575 558 649
rect 492 541 508 575
rect 542 541 558 575
rect 492 532 558 541
rect 592 599 648 615
rect 592 565 598 599
rect 632 565 648 599
rect 200 475 208 509
rect 242 475 258 509
rect 592 498 648 565
rect 200 413 258 475
rect 302 494 648 498
rect 302 464 598 494
rect 487 460 598 464
rect 632 460 648 494
rect 487 452 648 460
rect 683 611 749 649
rect 683 577 699 611
rect 733 577 749 611
rect 683 493 749 577
rect 683 459 699 493
rect 733 459 749 493
rect 683 452 749 459
rect 785 599 837 615
rect 785 565 801 599
rect 835 565 837 599
rect 785 506 837 565
rect 785 472 801 506
rect 835 472 837 506
rect 200 379 208 413
rect 242 379 258 413
rect 200 363 258 379
rect 384 414 441 430
rect 384 380 403 414
rect 437 380 441 414
rect 384 326 441 380
rect 200 310 441 326
rect 200 276 216 310
rect 250 276 441 310
rect 200 260 441 276
rect 111 170 121 204
rect 155 170 166 204
rect 111 101 166 170
rect 111 67 121 101
rect 155 67 166 101
rect 111 51 166 67
rect 200 203 257 219
rect 200 169 207 203
rect 241 169 257 203
rect 200 93 257 169
rect 375 194 441 260
rect 375 160 387 194
rect 421 160 441 194
rect 375 143 441 160
rect 487 167 521 452
rect 785 418 837 472
rect 633 409 837 418
rect 871 607 937 649
rect 871 573 887 607
rect 921 573 937 607
rect 871 524 937 573
rect 871 490 887 524
rect 921 490 937 524
rect 871 445 937 490
rect 871 411 887 445
rect 921 411 937 445
rect 1023 557 1233 591
rect 1023 455 1089 557
rect 1023 421 1039 455
rect 1073 421 1089 455
rect 1023 411 1089 421
rect 1125 507 1165 523
rect 1125 473 1129 507
rect 1163 473 1165 507
rect 1125 455 1165 473
rect 1199 505 1233 557
rect 1271 579 1339 649
rect 1271 545 1289 579
rect 1323 545 1339 579
rect 1271 539 1339 545
rect 1373 578 1604 596
rect 1373 562 1568 578
rect 1373 505 1407 562
rect 1523 544 1568 562
rect 1602 544 1604 578
rect 1523 528 1604 544
rect 1638 570 1704 649
rect 1638 536 1654 570
rect 1688 536 1704 570
rect 1638 528 1704 536
rect 1738 597 1805 613
rect 1738 563 1741 597
rect 1775 563 1805 597
rect 1738 529 1805 563
rect 1199 471 1407 505
rect 1441 512 1487 528
rect 1441 478 1443 512
rect 1477 478 1487 512
rect 633 384 801 409
rect 633 307 667 384
rect 799 375 801 384
rect 835 377 837 409
rect 835 375 1027 377
rect 555 291 667 307
rect 589 257 623 291
rect 657 257 667 291
rect 701 319 765 350
rect 799 343 1027 375
rect 701 285 731 319
rect 961 341 1027 343
rect 961 307 977 341
rect 1011 307 1027 341
rect 701 269 765 285
rect 850 291 909 307
rect 961 305 1027 307
rect 555 241 667 257
rect 633 235 667 241
rect 850 257 859 291
rect 893 271 909 291
rect 1125 271 1159 455
rect 1199 291 1233 471
rect 1441 460 1487 478
rect 1353 408 1419 426
rect 893 257 1159 271
rect 850 237 1159 257
rect 633 203 816 235
rect 633 201 914 203
rect 782 187 914 201
rect 782 167 864 187
rect 487 133 598 167
rect 632 133 648 167
rect 487 131 648 133
rect 582 95 648 131
rect 200 59 207 93
rect 241 59 257 93
rect 200 17 257 59
rect 480 59 496 93
rect 530 59 546 93
rect 480 17 546 59
rect 582 61 598 95
rect 632 61 648 95
rect 582 51 648 61
rect 682 133 698 167
rect 732 133 748 167
rect 682 93 748 133
rect 682 59 698 93
rect 732 59 748 93
rect 682 17 748 59
rect 848 153 864 167
rect 898 153 914 187
rect 848 101 914 153
rect 848 67 864 101
rect 898 67 914 101
rect 848 51 914 67
rect 976 178 1042 194
rect 976 144 992 178
rect 1026 144 1042 178
rect 976 17 1042 144
rect 1125 191 1159 237
rect 1193 275 1233 291
rect 1193 241 1197 275
rect 1231 241 1233 275
rect 1193 225 1233 241
rect 1267 389 1319 405
rect 1267 355 1269 389
rect 1303 355 1319 389
rect 1267 254 1319 355
rect 1353 374 1383 408
rect 1417 374 1419 408
rect 1353 340 1419 374
rect 1353 306 1383 340
rect 1417 306 1419 340
rect 1353 290 1419 306
rect 1453 254 1487 460
rect 1267 220 1487 254
rect 1125 178 1200 191
rect 1125 144 1150 178
rect 1184 144 1200 178
rect 1125 128 1200 144
rect 1314 178 1380 186
rect 1314 144 1330 178
rect 1364 144 1380 178
rect 1314 17 1380 144
rect 1414 178 1466 220
rect 1414 144 1416 178
rect 1450 144 1466 178
rect 1414 128 1466 144
rect 1523 122 1557 528
rect 1738 495 1741 529
rect 1775 495 1805 529
rect 1738 494 1805 495
rect 1591 460 1805 494
rect 1591 435 1627 460
rect 1591 401 1593 435
rect 1591 367 1627 401
rect 1591 333 1593 367
rect 1591 317 1627 333
rect 1661 286 1735 426
rect 1661 252 1701 286
rect 1661 218 1735 252
rect 1661 184 1701 218
rect 1661 156 1735 184
rect 1769 122 1805 460
rect 1523 106 1596 122
rect 1523 72 1554 106
rect 1588 72 1596 106
rect 1523 56 1596 72
rect 1630 106 1683 122
rect 1630 72 1640 106
rect 1674 72 1683 106
rect 1630 17 1683 72
rect 1717 106 1805 122
rect 1717 72 1726 106
rect 1760 72 1805 106
rect 1717 56 1805 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrbp_2
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1375 390 1409 424 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1663 168 1697 202 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1663 390 1697 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4334612
string GDS_START 4320574
<< end >>
