magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3122 1975
<< nwell >>
rect -38 331 1862 704
<< pwell >>
rect 1 241 189 251
rect 1 49 1757 241
rect 0 0 1824 49
<< scnmos >>
rect 80 57 110 225
rect 358 47 388 215
rect 444 47 474 215
rect 530 47 560 215
rect 616 47 646 215
rect 702 47 732 215
rect 788 47 818 215
rect 874 47 904 215
rect 960 47 990 215
rect 1046 47 1076 215
rect 1132 47 1162 215
rect 1218 47 1248 215
rect 1304 47 1334 215
rect 1390 47 1420 215
rect 1476 47 1506 215
rect 1562 47 1592 215
rect 1648 47 1678 215
<< scpmoshvt >>
rect 168 367 198 619
rect 358 367 388 619
rect 444 367 474 619
rect 530 367 560 619
rect 616 367 646 619
rect 702 367 732 619
rect 788 367 818 619
rect 874 367 904 619
rect 960 367 990 619
rect 1046 367 1076 619
rect 1132 367 1162 619
rect 1218 367 1248 619
rect 1304 367 1334 619
rect 1390 367 1420 619
rect 1476 367 1506 619
rect 1562 367 1592 619
rect 1648 367 1678 619
<< ndiff >>
rect 27 192 80 225
rect 27 158 35 192
rect 69 158 80 192
rect 27 103 80 158
rect 27 69 35 103
rect 69 69 80 103
rect 27 57 80 69
rect 110 192 163 225
rect 110 158 121 192
rect 155 158 163 192
rect 110 103 163 158
rect 305 203 358 215
rect 305 169 313 203
rect 347 169 358 203
rect 110 69 121 103
rect 155 69 163 103
rect 110 57 163 69
rect 305 101 358 169
rect 305 67 313 101
rect 347 67 358 101
rect 305 47 358 67
rect 388 207 444 215
rect 388 173 399 207
rect 433 173 444 207
rect 388 93 444 173
rect 388 59 399 93
rect 433 59 444 93
rect 388 47 444 59
rect 474 203 530 215
rect 474 169 485 203
rect 519 169 530 203
rect 474 101 530 169
rect 474 67 485 101
rect 519 67 530 101
rect 474 47 530 67
rect 560 207 616 215
rect 560 173 571 207
rect 605 173 616 207
rect 560 93 616 173
rect 560 59 571 93
rect 605 59 616 93
rect 560 47 616 59
rect 646 203 702 215
rect 646 169 657 203
rect 691 169 702 203
rect 646 101 702 169
rect 646 67 657 101
rect 691 67 702 101
rect 646 47 702 67
rect 732 207 788 215
rect 732 173 743 207
rect 777 173 788 207
rect 732 93 788 173
rect 732 59 743 93
rect 777 59 788 93
rect 732 47 788 59
rect 818 203 874 215
rect 818 169 829 203
rect 863 169 874 203
rect 818 101 874 169
rect 818 67 829 101
rect 863 67 874 101
rect 818 47 874 67
rect 904 207 960 215
rect 904 173 915 207
rect 949 173 960 207
rect 904 93 960 173
rect 904 59 915 93
rect 949 59 960 93
rect 904 47 960 59
rect 990 207 1046 215
rect 990 173 1001 207
rect 1035 173 1046 207
rect 990 101 1046 173
rect 990 67 1001 101
rect 1035 67 1046 101
rect 990 47 1046 67
rect 1076 188 1132 215
rect 1076 154 1087 188
rect 1121 154 1132 188
rect 1076 47 1132 154
rect 1162 101 1218 215
rect 1162 67 1173 101
rect 1207 67 1218 101
rect 1162 47 1218 67
rect 1248 188 1304 215
rect 1248 154 1259 188
rect 1293 154 1304 188
rect 1248 47 1304 154
rect 1334 194 1390 215
rect 1334 160 1345 194
rect 1379 160 1390 194
rect 1334 94 1390 160
rect 1334 60 1345 94
rect 1379 60 1390 94
rect 1334 47 1390 60
rect 1420 169 1476 215
rect 1420 135 1431 169
rect 1465 135 1476 169
rect 1420 47 1476 135
rect 1506 194 1562 215
rect 1506 160 1517 194
rect 1551 160 1562 194
rect 1506 96 1562 160
rect 1506 62 1517 96
rect 1551 62 1562 96
rect 1506 47 1562 62
rect 1592 169 1648 215
rect 1592 135 1603 169
rect 1637 135 1648 169
rect 1592 47 1648 135
rect 1678 203 1731 215
rect 1678 169 1689 203
rect 1723 169 1731 203
rect 1678 103 1731 169
rect 1678 69 1689 103
rect 1723 69 1731 103
rect 1678 47 1731 69
<< pdiff >>
rect 115 607 168 619
rect 115 573 123 607
rect 157 573 168 607
rect 115 512 168 573
rect 115 478 123 512
rect 157 478 168 512
rect 115 413 168 478
rect 115 379 123 413
rect 157 379 168 413
rect 115 367 168 379
rect 198 599 251 619
rect 198 565 209 599
rect 243 565 251 599
rect 198 512 251 565
rect 198 478 209 512
rect 243 478 251 512
rect 198 413 251 478
rect 198 379 209 413
rect 243 379 251 413
rect 198 367 251 379
rect 305 599 358 619
rect 305 565 313 599
rect 347 565 358 599
rect 305 512 358 565
rect 305 478 313 512
rect 347 478 358 512
rect 305 413 358 478
rect 305 379 313 413
rect 347 379 358 413
rect 305 367 358 379
rect 388 607 444 619
rect 388 573 399 607
rect 433 573 444 607
rect 388 535 444 573
rect 388 501 399 535
rect 433 501 444 535
rect 388 453 444 501
rect 388 419 399 453
rect 433 419 444 453
rect 388 367 444 419
rect 474 599 530 619
rect 474 565 485 599
rect 519 565 530 599
rect 474 512 530 565
rect 474 478 485 512
rect 519 478 530 512
rect 474 413 530 478
rect 474 379 485 413
rect 519 379 530 413
rect 474 367 530 379
rect 560 607 616 619
rect 560 573 571 607
rect 605 573 616 607
rect 560 535 616 573
rect 560 501 571 535
rect 605 501 616 535
rect 560 453 616 501
rect 560 419 571 453
rect 605 419 616 453
rect 560 367 616 419
rect 646 599 702 619
rect 646 565 657 599
rect 691 565 702 599
rect 646 512 702 565
rect 646 478 657 512
rect 691 478 702 512
rect 646 413 702 478
rect 646 379 657 413
rect 691 379 702 413
rect 646 367 702 379
rect 732 607 788 619
rect 732 573 743 607
rect 777 573 788 607
rect 732 535 788 573
rect 732 501 743 535
rect 777 501 788 535
rect 732 453 788 501
rect 732 419 743 453
rect 777 419 788 453
rect 732 367 788 419
rect 818 599 874 619
rect 818 565 829 599
rect 863 565 874 599
rect 818 512 874 565
rect 818 478 829 512
rect 863 478 874 512
rect 818 413 874 478
rect 818 379 829 413
rect 863 379 874 413
rect 818 367 874 379
rect 904 607 960 619
rect 904 573 915 607
rect 949 573 960 607
rect 904 535 960 573
rect 904 501 915 535
rect 949 501 960 535
rect 904 453 960 501
rect 904 419 915 453
rect 949 419 960 453
rect 904 367 960 419
rect 990 599 1046 619
rect 990 565 1001 599
rect 1035 565 1046 599
rect 990 512 1046 565
rect 990 478 1001 512
rect 1035 478 1046 512
rect 990 413 1046 478
rect 990 379 1001 413
rect 1035 379 1046 413
rect 990 367 1046 379
rect 1076 547 1132 619
rect 1076 513 1087 547
rect 1121 513 1132 547
rect 1076 413 1132 513
rect 1076 379 1087 413
rect 1121 379 1132 413
rect 1076 367 1132 379
rect 1162 597 1218 619
rect 1162 563 1173 597
rect 1207 563 1218 597
rect 1162 529 1218 563
rect 1162 495 1173 529
rect 1207 495 1218 529
rect 1162 461 1218 495
rect 1162 427 1173 461
rect 1207 427 1218 461
rect 1162 367 1218 427
rect 1248 547 1304 619
rect 1248 513 1259 547
rect 1293 513 1304 547
rect 1248 413 1304 513
rect 1248 379 1259 413
rect 1293 379 1304 413
rect 1248 367 1304 379
rect 1334 597 1390 619
rect 1334 563 1345 597
rect 1379 563 1390 597
rect 1334 529 1390 563
rect 1334 495 1345 529
rect 1379 495 1390 529
rect 1334 461 1390 495
rect 1334 427 1345 461
rect 1379 427 1390 461
rect 1334 367 1390 427
rect 1420 547 1476 619
rect 1420 513 1431 547
rect 1465 513 1476 547
rect 1420 413 1476 513
rect 1420 379 1431 413
rect 1465 379 1476 413
rect 1420 367 1476 379
rect 1506 597 1562 619
rect 1506 563 1517 597
rect 1551 563 1562 597
rect 1506 529 1562 563
rect 1506 495 1517 529
rect 1551 495 1562 529
rect 1506 461 1562 495
rect 1506 427 1517 461
rect 1551 427 1562 461
rect 1506 367 1562 427
rect 1592 547 1648 619
rect 1592 513 1603 547
rect 1637 513 1648 547
rect 1592 413 1648 513
rect 1592 379 1603 413
rect 1637 379 1648 413
rect 1592 367 1648 379
rect 1678 599 1731 619
rect 1678 565 1689 599
rect 1723 565 1731 599
rect 1678 512 1731 565
rect 1678 478 1689 512
rect 1723 478 1731 512
rect 1678 415 1731 478
rect 1678 381 1689 415
rect 1723 381 1731 415
rect 1678 367 1731 381
<< ndiffc >>
rect 35 158 69 192
rect 35 69 69 103
rect 121 158 155 192
rect 313 169 347 203
rect 121 69 155 103
rect 313 67 347 101
rect 399 173 433 207
rect 399 59 433 93
rect 485 169 519 203
rect 485 67 519 101
rect 571 173 605 207
rect 571 59 605 93
rect 657 169 691 203
rect 657 67 691 101
rect 743 173 777 207
rect 743 59 777 93
rect 829 169 863 203
rect 829 67 863 101
rect 915 173 949 207
rect 915 59 949 93
rect 1001 173 1035 207
rect 1001 67 1035 101
rect 1087 154 1121 188
rect 1173 67 1207 101
rect 1259 154 1293 188
rect 1345 160 1379 194
rect 1345 60 1379 94
rect 1431 135 1465 169
rect 1517 160 1551 194
rect 1517 62 1551 96
rect 1603 135 1637 169
rect 1689 169 1723 203
rect 1689 69 1723 103
<< pdiffc >>
rect 123 573 157 607
rect 123 478 157 512
rect 123 379 157 413
rect 209 565 243 599
rect 209 478 243 512
rect 209 379 243 413
rect 313 565 347 599
rect 313 478 347 512
rect 313 379 347 413
rect 399 573 433 607
rect 399 501 433 535
rect 399 419 433 453
rect 485 565 519 599
rect 485 478 519 512
rect 485 379 519 413
rect 571 573 605 607
rect 571 501 605 535
rect 571 419 605 453
rect 657 565 691 599
rect 657 478 691 512
rect 657 379 691 413
rect 743 573 777 607
rect 743 501 777 535
rect 743 419 777 453
rect 829 565 863 599
rect 829 478 863 512
rect 829 379 863 413
rect 915 573 949 607
rect 915 501 949 535
rect 915 419 949 453
rect 1001 565 1035 599
rect 1001 478 1035 512
rect 1001 379 1035 413
rect 1087 513 1121 547
rect 1087 379 1121 413
rect 1173 563 1207 597
rect 1173 495 1207 529
rect 1173 427 1207 461
rect 1259 513 1293 547
rect 1259 379 1293 413
rect 1345 563 1379 597
rect 1345 495 1379 529
rect 1345 427 1379 461
rect 1431 513 1465 547
rect 1431 379 1465 413
rect 1517 563 1551 597
rect 1517 495 1551 529
rect 1517 427 1551 461
rect 1603 513 1637 547
rect 1603 379 1637 413
rect 1689 565 1723 599
rect 1689 478 1723 512
rect 1689 381 1723 415
<< poly >>
rect 168 619 198 645
rect 358 619 388 645
rect 444 619 474 645
rect 530 619 560 645
rect 616 619 646 645
rect 702 619 732 645
rect 788 619 818 645
rect 874 619 904 645
rect 960 619 990 645
rect 1046 619 1076 645
rect 1132 619 1162 645
rect 1218 619 1248 645
rect 1304 619 1334 645
rect 1390 619 1420 645
rect 1476 619 1506 645
rect 1562 619 1592 645
rect 1648 619 1678 645
rect 168 345 198 367
rect 358 345 388 367
rect 444 345 474 367
rect 530 345 560 367
rect 616 345 646 367
rect 702 345 732 367
rect 788 345 818 367
rect 874 345 904 367
rect 960 345 990 367
rect 21 311 990 345
rect 21 309 155 311
rect 21 275 37 309
rect 71 275 105 309
rect 139 275 155 309
rect 21 259 155 275
rect 1046 303 1076 367
rect 1132 303 1162 367
rect 1218 303 1248 367
rect 1304 303 1334 367
rect 1390 303 1420 367
rect 1476 303 1506 367
rect 1562 303 1592 367
rect 1648 303 1678 367
rect 1046 287 1678 303
rect 80 225 110 259
rect 197 251 990 269
rect 197 217 213 251
rect 247 237 990 251
rect 247 217 263 237
rect 197 183 263 217
rect 358 215 388 237
rect 444 215 474 237
rect 530 215 560 237
rect 616 215 646 237
rect 702 215 732 237
rect 788 215 818 237
rect 874 215 904 237
rect 960 215 990 237
rect 1046 253 1085 287
rect 1119 253 1153 287
rect 1187 253 1678 287
rect 1046 237 1678 253
rect 1046 215 1076 237
rect 1132 215 1162 237
rect 1218 215 1248 237
rect 1304 215 1334 237
rect 1390 215 1420 237
rect 1476 215 1506 237
rect 1562 215 1592 237
rect 1648 215 1678 237
rect 197 149 213 183
rect 247 149 263 183
rect 197 133 263 149
rect 80 31 110 57
rect 358 21 388 47
rect 444 21 474 47
rect 530 21 560 47
rect 616 21 646 47
rect 702 21 732 47
rect 788 21 818 47
rect 874 21 904 47
rect 960 21 990 47
rect 1046 21 1076 47
rect 1132 21 1162 47
rect 1218 21 1248 47
rect 1304 21 1334 47
rect 1390 21 1420 47
rect 1476 21 1506 47
rect 1562 21 1592 47
rect 1648 21 1678 47
<< polycont >>
rect 37 275 71 309
rect 105 275 139 309
rect 213 217 247 251
rect 1085 253 1119 287
rect 1153 253 1187 287
rect 213 149 247 183
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 119 607 161 649
rect 21 329 83 592
rect 119 573 123 607
rect 157 573 161 607
rect 119 512 161 573
rect 119 478 123 512
rect 157 478 161 512
rect 119 413 161 478
rect 119 379 123 413
rect 157 379 161 413
rect 119 363 161 379
rect 197 599 263 615
rect 197 565 209 599
rect 243 565 263 599
rect 197 512 263 565
rect 197 478 209 512
rect 243 478 263 512
rect 197 413 263 478
rect 197 379 209 413
rect 243 379 263 413
rect 21 309 155 329
rect 21 275 37 309
rect 71 275 105 309
rect 139 275 155 309
rect 21 242 155 275
rect 197 251 263 379
rect 297 599 349 615
rect 297 565 313 599
rect 347 565 349 599
rect 297 512 349 565
rect 297 478 313 512
rect 347 478 349 512
rect 297 413 349 478
rect 383 607 449 649
rect 383 573 399 607
rect 433 573 449 607
rect 383 535 449 573
rect 383 501 399 535
rect 433 501 449 535
rect 383 453 449 501
rect 383 419 399 453
rect 433 419 449 453
rect 483 599 521 615
rect 483 565 485 599
rect 519 565 521 599
rect 483 512 521 565
rect 483 478 485 512
rect 519 478 521 512
rect 297 379 313 413
rect 347 385 349 413
rect 483 413 521 478
rect 555 607 621 649
rect 555 573 571 607
rect 605 573 621 607
rect 555 535 621 573
rect 555 501 571 535
rect 605 501 621 535
rect 555 453 621 501
rect 555 419 571 453
rect 605 419 621 453
rect 655 599 693 615
rect 655 565 657 599
rect 691 565 693 599
rect 655 512 693 565
rect 655 478 657 512
rect 691 478 693 512
rect 483 385 485 413
rect 347 379 485 385
rect 519 385 521 413
rect 655 413 693 478
rect 727 607 793 649
rect 727 573 743 607
rect 777 573 793 607
rect 727 535 793 573
rect 727 501 743 535
rect 777 501 793 535
rect 727 453 793 501
rect 727 419 743 453
rect 777 419 793 453
rect 827 599 865 615
rect 827 565 829 599
rect 863 565 865 599
rect 827 512 865 565
rect 827 478 829 512
rect 863 478 865 512
rect 655 385 657 413
rect 519 379 657 385
rect 691 385 693 413
rect 827 413 865 478
rect 899 607 965 649
rect 899 573 915 607
rect 949 573 965 607
rect 899 535 965 573
rect 899 501 915 535
rect 949 501 965 535
rect 899 453 965 501
rect 899 419 915 453
rect 949 419 965 453
rect 999 599 1739 615
rect 999 565 1001 599
rect 1035 597 1689 599
rect 1035 581 1173 597
rect 1035 565 1037 581
rect 999 512 1037 565
rect 1171 563 1173 581
rect 1207 581 1345 597
rect 1207 563 1209 581
rect 999 478 1001 512
rect 1035 478 1037 512
rect 827 385 829 413
rect 691 379 829 385
rect 863 385 865 413
rect 999 413 1037 478
rect 999 385 1001 413
rect 863 379 1001 385
rect 1035 379 1037 413
rect 297 335 1037 379
rect 1071 513 1087 547
rect 1121 513 1137 547
rect 1071 413 1137 513
rect 1071 379 1087 413
rect 1121 379 1137 413
rect 1171 529 1209 563
rect 1343 563 1345 581
rect 1379 581 1517 597
rect 1379 563 1381 581
rect 1171 495 1173 529
rect 1207 495 1209 529
rect 1171 461 1209 495
rect 1171 427 1173 461
rect 1207 427 1209 461
rect 1171 411 1209 427
rect 1243 513 1259 547
rect 1293 513 1309 547
rect 1243 413 1309 513
rect 1071 375 1137 379
rect 1243 379 1259 413
rect 1293 379 1309 413
rect 1343 529 1381 563
rect 1515 563 1517 581
rect 1551 581 1689 597
rect 1551 563 1553 581
rect 1343 495 1345 529
rect 1379 495 1381 529
rect 1343 461 1381 495
rect 1343 427 1345 461
rect 1379 427 1381 461
rect 1343 411 1381 427
rect 1415 513 1431 547
rect 1465 513 1481 547
rect 1415 413 1481 513
rect 1243 375 1309 379
rect 1415 379 1431 413
rect 1465 379 1481 413
rect 1515 529 1553 563
rect 1687 565 1689 581
rect 1723 565 1739 599
rect 1515 495 1517 529
rect 1551 495 1553 529
rect 1515 461 1553 495
rect 1515 427 1517 461
rect 1551 427 1553 461
rect 1515 411 1553 427
rect 1587 513 1603 547
rect 1637 513 1653 547
rect 1587 413 1653 513
rect 1415 375 1481 379
rect 1587 379 1603 413
rect 1637 379 1653 413
rect 1587 375 1653 379
rect 1071 337 1653 375
rect 1687 512 1739 565
rect 1687 478 1689 512
rect 1723 478 1739 512
rect 1687 415 1739 478
rect 1687 381 1689 415
rect 1723 381 1739 415
rect 1687 365 1739 381
rect 1261 333 1653 337
rect 197 217 213 251
rect 247 217 263 251
rect 197 208 263 217
rect 19 192 78 208
rect 19 158 35 192
rect 69 158 78 192
rect 19 103 78 158
rect 19 69 35 103
rect 69 69 78 103
rect 19 17 78 69
rect 117 192 263 208
rect 117 158 121 192
rect 155 183 263 192
rect 155 158 213 183
rect 117 149 213 158
rect 247 149 263 183
rect 117 133 263 149
rect 297 257 1037 301
rect 297 203 356 257
rect 297 169 313 203
rect 347 169 356 203
rect 117 103 159 133
rect 117 69 121 103
rect 155 69 159 103
rect 117 53 159 69
rect 297 101 356 169
rect 297 67 313 101
rect 347 67 356 101
rect 297 51 356 67
rect 390 207 442 223
rect 390 173 399 207
rect 433 173 442 207
rect 390 93 442 173
rect 390 59 399 93
rect 433 59 442 93
rect 390 17 442 59
rect 476 203 528 257
rect 476 169 485 203
rect 519 169 528 203
rect 476 101 528 169
rect 476 67 485 101
rect 519 67 528 101
rect 476 51 528 67
rect 562 207 614 223
rect 562 173 571 207
rect 605 173 614 207
rect 562 93 614 173
rect 562 59 571 93
rect 605 59 614 93
rect 562 17 614 59
rect 648 203 700 257
rect 648 169 657 203
rect 691 169 700 203
rect 648 101 700 169
rect 648 67 657 101
rect 691 67 700 101
rect 648 51 700 67
rect 734 207 786 223
rect 734 173 743 207
rect 777 173 786 207
rect 734 93 786 173
rect 734 59 743 93
rect 777 59 786 93
rect 734 17 786 59
rect 820 203 872 257
rect 820 169 829 203
rect 863 169 872 203
rect 820 101 872 169
rect 820 67 829 101
rect 863 67 872 101
rect 820 51 872 67
rect 906 207 958 223
rect 906 173 915 207
rect 949 173 958 207
rect 906 93 958 173
rect 906 59 915 93
rect 949 59 958 93
rect 906 17 958 59
rect 992 207 1037 257
rect 1071 287 1227 303
rect 1071 253 1085 287
rect 1119 253 1153 287
rect 1187 253 1227 287
rect 1071 237 1227 253
rect 992 173 1001 207
rect 1035 173 1037 207
rect 1261 228 1645 333
rect 1261 203 1295 228
rect 992 104 1037 173
rect 1071 188 1295 203
rect 1071 154 1087 188
rect 1121 154 1259 188
rect 1293 154 1295 188
rect 1071 138 1295 154
rect 1329 160 1345 194
rect 1379 160 1395 194
rect 1329 104 1395 160
rect 1429 169 1467 228
rect 1429 135 1431 169
rect 1465 135 1467 169
rect 1429 119 1467 135
rect 1501 160 1517 194
rect 1551 160 1567 194
rect 992 101 1395 104
rect 992 67 1001 101
rect 1035 67 1173 101
rect 1207 94 1395 101
rect 1207 67 1345 94
rect 992 60 1345 67
rect 1379 85 1395 94
rect 1501 96 1567 160
rect 1601 169 1645 228
rect 1601 135 1603 169
rect 1637 135 1645 169
rect 1601 119 1645 135
rect 1679 203 1739 219
rect 1679 169 1689 203
rect 1723 169 1739 203
rect 1501 85 1517 96
rect 1379 62 1517 85
rect 1551 85 1567 96
rect 1679 103 1739 169
rect 1679 85 1689 103
rect 1551 69 1689 85
rect 1723 69 1739 103
rect 1551 62 1739 69
rect 1379 60 1739 62
rect 992 51 1739 60
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 einvn_8
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3991602
string GDS_START 3977332
<< end >>
