magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 332 1286 704
<< pwell >>
rect 4 49 1247 248
rect 0 0 1248 49
<< scpmos >>
rect 86 368 116 592
rect 186 368 216 592
rect 276 368 306 592
rect 366 368 396 592
rect 456 368 486 592
rect 546 368 576 592
rect 636 368 666 592
rect 726 368 756 592
rect 842 368 872 592
rect 942 368 972 592
rect 1032 368 1062 592
rect 1132 368 1162 592
<< nmoslvt >>
rect 87 74 117 222
rect 183 74 213 222
rect 273 74 303 222
rect 373 74 403 222
rect 459 74 489 222
rect 559 74 589 222
rect 645 74 675 222
rect 745 74 775 222
rect 845 74 875 222
rect 945 74 975 222
rect 1034 74 1064 222
rect 1134 74 1164 222
<< ndiff >>
rect 30 210 87 222
rect 30 176 42 210
rect 76 176 87 210
rect 30 120 87 176
rect 30 86 42 120
rect 76 86 87 120
rect 30 74 87 86
rect 117 136 183 222
rect 117 102 128 136
rect 162 102 183 136
rect 117 74 183 102
rect 213 210 273 222
rect 213 176 228 210
rect 262 176 273 210
rect 213 120 273 176
rect 213 86 228 120
rect 262 86 273 120
rect 213 74 273 86
rect 303 131 373 222
rect 303 97 328 131
rect 362 97 373 131
rect 303 74 373 97
rect 403 210 459 222
rect 403 176 414 210
rect 448 176 459 210
rect 403 120 459 176
rect 403 86 414 120
rect 448 86 459 120
rect 403 74 459 86
rect 489 126 559 222
rect 489 92 500 126
rect 534 92 559 126
rect 489 74 559 92
rect 589 210 645 222
rect 589 176 600 210
rect 634 176 645 210
rect 589 120 645 176
rect 589 86 600 120
rect 634 86 645 120
rect 589 74 645 86
rect 675 142 745 222
rect 675 108 700 142
rect 734 108 745 142
rect 675 74 745 108
rect 775 210 845 222
rect 775 176 800 210
rect 834 176 845 210
rect 775 120 845 176
rect 775 86 800 120
rect 834 86 845 120
rect 775 74 845 86
rect 875 126 945 222
rect 875 92 900 126
rect 934 92 945 126
rect 875 74 945 92
rect 975 210 1034 222
rect 975 176 987 210
rect 1021 176 1034 210
rect 975 120 1034 176
rect 975 86 987 120
rect 1021 86 1034 120
rect 975 74 1034 86
rect 1064 126 1134 222
rect 1064 92 1075 126
rect 1109 92 1134 126
rect 1064 74 1134 92
rect 1164 210 1221 222
rect 1164 176 1175 210
rect 1209 176 1221 210
rect 1164 120 1221 176
rect 1164 86 1175 120
rect 1209 86 1221 120
rect 1164 74 1221 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 440 86 476
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 566 186 592
rect 116 532 139 566
rect 173 532 186 566
rect 116 368 186 532
rect 216 414 276 592
rect 216 380 229 414
rect 263 380 276 414
rect 216 368 276 380
rect 306 566 366 592
rect 306 532 319 566
rect 353 532 366 566
rect 306 368 366 532
rect 396 414 456 592
rect 396 380 409 414
rect 443 380 456 414
rect 396 368 456 380
rect 486 566 546 592
rect 486 532 499 566
rect 533 532 546 566
rect 486 368 546 532
rect 576 414 636 592
rect 576 380 589 414
rect 623 380 636 414
rect 576 368 636 380
rect 666 566 726 592
rect 666 532 679 566
rect 713 532 726 566
rect 666 368 726 532
rect 756 414 842 592
rect 756 380 782 414
rect 816 380 842 414
rect 756 368 842 380
rect 872 566 942 592
rect 872 532 885 566
rect 919 532 942 566
rect 872 368 942 532
rect 972 580 1032 592
rect 972 546 985 580
rect 1019 546 1032 580
rect 972 478 1032 546
rect 972 444 985 478
rect 1019 444 1032 478
rect 972 368 1032 444
rect 1062 546 1132 592
rect 1062 512 1085 546
rect 1119 512 1132 546
rect 1062 368 1132 512
rect 1162 580 1221 592
rect 1162 546 1175 580
rect 1209 546 1221 580
rect 1162 497 1221 546
rect 1162 463 1175 497
rect 1209 463 1221 497
rect 1162 414 1221 463
rect 1162 380 1175 414
rect 1209 380 1221 414
rect 1162 368 1221 380
<< ndiffc >>
rect 42 176 76 210
rect 42 86 76 120
rect 128 102 162 136
rect 228 176 262 210
rect 228 86 262 120
rect 328 97 362 131
rect 414 176 448 210
rect 414 86 448 120
rect 500 92 534 126
rect 600 176 634 210
rect 600 86 634 120
rect 700 108 734 142
rect 800 176 834 210
rect 800 86 834 120
rect 900 92 934 126
rect 987 176 1021 210
rect 987 86 1021 120
rect 1075 92 1109 126
rect 1175 176 1209 210
rect 1175 86 1209 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 139 532 173 566
rect 229 380 263 414
rect 319 532 353 566
rect 409 380 443 414
rect 499 532 533 566
rect 589 380 623 414
rect 679 532 713 566
rect 782 380 816 414
rect 885 532 919 566
rect 985 546 1019 580
rect 985 444 1019 478
rect 1085 512 1119 546
rect 1175 546 1209 580
rect 1175 463 1209 497
rect 1175 380 1209 414
<< poly >>
rect 86 592 116 618
rect 186 592 216 618
rect 276 592 306 618
rect 366 592 396 618
rect 456 592 486 618
rect 546 592 576 618
rect 636 592 666 618
rect 726 592 756 618
rect 842 592 872 618
rect 942 592 972 618
rect 1032 592 1062 618
rect 1132 592 1162 618
rect 86 353 116 368
rect 186 353 216 368
rect 276 353 306 368
rect 366 353 396 368
rect 456 353 486 368
rect 546 353 576 368
rect 636 353 666 368
rect 726 353 756 368
rect 842 353 872 368
rect 942 353 972 368
rect 1032 353 1062 368
rect 1132 353 1162 368
rect 83 336 119 353
rect 44 320 119 336
rect 44 286 60 320
rect 94 286 119 320
rect 44 270 119 286
rect 183 326 219 353
rect 273 326 309 353
rect 363 326 399 353
rect 453 326 489 353
rect 543 326 579 353
rect 633 326 669 353
rect 723 326 759 353
rect 839 326 875 353
rect 942 330 975 353
rect 1029 330 1065 353
rect 1129 330 1165 353
rect 183 310 875 326
rect 183 276 349 310
rect 383 276 417 310
rect 451 276 485 310
rect 519 276 553 310
rect 587 276 621 310
rect 655 276 689 310
rect 723 276 757 310
rect 791 276 825 310
rect 859 276 875 310
rect 87 222 117 270
rect 183 260 875 276
rect 183 222 213 260
rect 273 222 303 260
rect 373 222 403 260
rect 459 222 489 260
rect 559 222 589 260
rect 645 222 675 260
rect 745 222 775 260
rect 845 222 875 260
rect 945 314 1165 330
rect 945 280 1010 314
rect 1044 280 1078 314
rect 1112 294 1165 314
rect 1112 280 1164 294
rect 945 264 1164 280
rect 945 222 975 264
rect 1034 222 1064 264
rect 1134 222 1164 264
rect 87 48 117 74
rect 183 48 213 74
rect 273 48 303 74
rect 373 48 403 74
rect 459 48 489 74
rect 559 48 589 74
rect 645 48 675 74
rect 745 48 775 74
rect 845 48 875 74
rect 945 48 975 74
rect 1034 48 1064 74
rect 1134 48 1164 74
<< polycont >>
rect 60 286 94 320
rect 349 276 383 310
rect 417 276 451 310
rect 485 276 519 310
rect 553 276 587 310
rect 621 276 655 310
rect 689 276 723 310
rect 757 276 791 310
rect 825 276 859 310
rect 1010 280 1044 314
rect 1078 280 1112 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 123 566 189 649
rect 123 532 139 566
rect 173 532 189 566
rect 123 516 189 532
rect 303 566 369 649
rect 303 532 319 566
rect 353 532 369 566
rect 303 516 369 532
rect 483 566 549 649
rect 483 532 499 566
rect 533 532 549 566
rect 483 516 549 532
rect 663 566 729 649
rect 663 532 679 566
rect 713 532 729 566
rect 663 516 729 532
rect 869 566 935 649
rect 869 532 885 566
rect 919 532 935 566
rect 869 516 935 532
rect 969 580 1035 596
rect 969 546 985 580
rect 1019 546 1035 580
rect 23 476 39 510
rect 73 482 89 510
rect 73 476 913 482
rect 23 448 913 476
rect 23 440 89 448
rect 23 406 39 440
rect 73 406 89 440
rect 23 390 89 406
rect 25 320 110 356
rect 25 286 60 320
rect 94 286 110 320
rect 25 270 110 286
rect 144 236 178 448
rect 26 210 178 236
rect 26 176 42 210
rect 76 202 178 210
rect 212 380 229 414
rect 263 380 409 414
rect 443 380 589 414
rect 623 380 782 414
rect 816 380 845 414
rect 212 360 845 380
rect 879 394 913 448
rect 969 478 1035 546
rect 1069 546 1135 649
rect 1069 512 1085 546
rect 1119 512 1135 546
rect 1069 496 1135 512
rect 1169 580 1225 596
rect 1169 546 1175 580
rect 1209 546 1225 580
rect 1169 497 1225 546
rect 969 444 985 478
rect 1019 462 1035 478
rect 1169 463 1175 497
rect 1209 463 1225 497
rect 1169 462 1225 463
rect 1019 444 1225 462
rect 969 428 1225 444
rect 1159 414 1225 428
rect 879 360 1121 394
rect 212 226 278 360
rect 333 310 964 326
rect 333 276 349 310
rect 383 276 417 310
rect 451 276 485 310
rect 519 276 553 310
rect 587 276 621 310
rect 655 276 689 310
rect 723 276 757 310
rect 791 276 825 310
rect 859 276 964 310
rect 333 260 964 276
rect 998 314 1121 360
rect 998 280 1010 314
rect 1044 280 1078 314
rect 1112 280 1121 314
rect 998 264 1121 280
rect 1159 380 1175 414
rect 1209 380 1225 414
rect 930 226 964 260
rect 1159 226 1225 380
rect 212 210 850 226
rect 26 120 76 176
rect 212 176 228 210
rect 262 176 414 210
rect 448 176 600 210
rect 634 192 800 210
rect 634 176 650 192
rect 26 86 42 120
rect 26 70 76 86
rect 112 136 178 168
rect 112 102 128 136
rect 162 102 178 136
rect 112 17 178 102
rect 212 120 278 176
rect 212 86 228 120
rect 262 86 278 120
rect 212 70 278 86
rect 312 131 378 142
rect 312 97 328 131
rect 362 97 378 131
rect 312 17 378 97
rect 412 120 450 176
rect 412 86 414 120
rect 448 86 450 120
rect 412 70 450 86
rect 484 126 550 142
rect 484 92 500 126
rect 534 92 550 126
rect 484 17 550 92
rect 584 120 650 176
rect 784 176 800 192
rect 834 176 850 210
rect 930 210 1225 226
rect 930 176 987 210
rect 1021 176 1175 210
rect 1209 176 1225 210
rect 584 86 600 120
rect 634 86 650 120
rect 584 70 650 86
rect 684 142 750 158
rect 684 108 700 142
rect 734 108 750 142
rect 684 17 750 108
rect 784 120 850 176
rect 784 86 800 120
rect 834 86 850 120
rect 784 70 850 86
rect 884 126 950 142
rect 884 92 900 126
rect 934 92 950 126
rect 884 17 950 92
rect 984 120 1025 176
rect 984 86 987 120
rect 1021 86 1025 120
rect 984 70 1025 86
rect 1059 126 1125 142
rect 1059 92 1075 126
rect 1109 92 1125 126
rect 1059 17 1125 92
rect 1159 120 1225 176
rect 1159 86 1175 120
rect 1209 86 1225 120
rect 1159 70 1225 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
rlabel comment s 0 0 0 0 4 bufinv_8
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 609050
string GDS_START 599878
<< end >>
