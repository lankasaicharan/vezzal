magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 34 49 926 241
rect 0 0 960 49
<< scnmos >>
rect 113 47 143 215
rect 215 47 245 215
rect 301 47 331 215
rect 387 47 417 215
rect 473 47 503 215
rect 559 47 589 215
rect 645 47 675 215
rect 731 47 761 215
rect 817 47 847 215
<< scpmoshvt >>
rect 113 367 143 619
rect 215 367 245 619
rect 301 367 331 619
rect 387 367 417 619
rect 473 367 503 619
rect 559 367 589 619
rect 645 367 675 619
rect 731 367 761 619
rect 817 367 847 619
<< ndiff >>
rect 60 203 113 215
rect 60 169 68 203
rect 102 169 113 203
rect 60 101 113 169
rect 60 67 68 101
rect 102 67 113 101
rect 60 47 113 67
rect 143 167 215 215
rect 143 133 154 167
rect 188 133 215 167
rect 143 93 215 133
rect 143 59 154 93
rect 188 59 215 93
rect 143 47 215 59
rect 245 179 301 215
rect 245 145 256 179
rect 290 145 301 179
rect 245 101 301 145
rect 245 67 256 101
rect 290 67 301 101
rect 245 47 301 67
rect 331 99 387 215
rect 331 65 342 99
rect 376 65 387 99
rect 331 47 387 65
rect 417 179 473 215
rect 417 145 428 179
rect 462 145 473 179
rect 417 101 473 145
rect 417 67 428 101
rect 462 67 473 101
rect 417 47 473 67
rect 503 99 559 215
rect 503 65 514 99
rect 548 65 559 99
rect 503 47 559 65
rect 589 175 645 215
rect 589 141 600 175
rect 634 141 645 175
rect 589 101 645 141
rect 589 67 600 101
rect 634 67 645 101
rect 589 47 645 67
rect 675 99 731 215
rect 675 65 686 99
rect 720 65 731 99
rect 675 47 731 65
rect 761 203 817 215
rect 761 169 772 203
rect 806 169 817 203
rect 761 101 817 169
rect 761 67 772 101
rect 806 67 817 101
rect 761 47 817 67
rect 847 161 900 215
rect 847 127 858 161
rect 892 127 900 161
rect 847 93 900 127
rect 847 59 858 93
rect 892 59 900 93
rect 847 47 900 59
<< pdiff >>
rect 60 599 113 619
rect 60 565 68 599
rect 102 565 113 599
rect 60 518 113 565
rect 60 484 68 518
rect 102 484 113 518
rect 60 436 113 484
rect 60 402 68 436
rect 102 402 113 436
rect 60 367 113 402
rect 143 607 215 619
rect 143 573 166 607
rect 200 573 215 607
rect 143 493 215 573
rect 143 459 166 493
rect 200 459 215 493
rect 143 367 215 459
rect 245 607 301 619
rect 245 573 256 607
rect 290 573 301 607
rect 245 367 301 573
rect 331 447 387 619
rect 331 413 342 447
rect 376 413 387 447
rect 331 367 387 413
rect 417 607 473 619
rect 417 573 428 607
rect 462 573 473 607
rect 417 367 473 573
rect 503 527 559 619
rect 503 493 514 527
rect 548 493 559 527
rect 503 367 559 493
rect 589 597 645 619
rect 589 563 600 597
rect 634 563 645 597
rect 589 525 645 563
rect 589 491 600 525
rect 634 491 645 525
rect 589 367 645 491
rect 675 527 731 619
rect 675 493 686 527
rect 720 493 731 527
rect 675 459 731 493
rect 675 425 686 459
rect 720 425 731 459
rect 675 367 731 425
rect 761 597 817 619
rect 761 563 772 597
rect 806 563 817 597
rect 761 525 817 563
rect 761 491 772 525
rect 806 491 817 525
rect 761 367 817 491
rect 847 607 900 619
rect 847 573 858 607
rect 892 573 900 607
rect 847 512 900 573
rect 847 478 858 512
rect 892 478 900 512
rect 847 367 900 478
<< ndiffc >>
rect 68 169 102 203
rect 68 67 102 101
rect 154 133 188 167
rect 154 59 188 93
rect 256 145 290 179
rect 256 67 290 101
rect 342 65 376 99
rect 428 145 462 179
rect 428 67 462 101
rect 514 65 548 99
rect 600 141 634 175
rect 600 67 634 101
rect 686 65 720 99
rect 772 169 806 203
rect 772 67 806 101
rect 858 127 892 161
rect 858 59 892 93
<< pdiffc >>
rect 68 565 102 599
rect 68 484 102 518
rect 68 402 102 436
rect 166 573 200 607
rect 166 459 200 493
rect 256 573 290 607
rect 342 413 376 447
rect 428 573 462 607
rect 514 493 548 527
rect 600 563 634 597
rect 600 491 634 525
rect 686 493 720 527
rect 686 425 720 459
rect 772 563 806 597
rect 772 491 806 525
rect 858 573 892 607
rect 858 478 892 512
<< poly >>
rect 113 619 143 645
rect 215 619 245 645
rect 301 619 331 645
rect 387 619 417 645
rect 473 619 503 645
rect 559 619 589 645
rect 645 619 675 645
rect 731 619 761 645
rect 817 619 847 645
rect 113 325 143 367
rect 215 335 245 367
rect 21 309 143 325
rect 21 275 37 309
rect 71 275 143 309
rect 21 259 143 275
rect 193 319 259 335
rect 193 285 209 319
rect 243 285 259 319
rect 193 269 259 285
rect 301 303 331 367
rect 387 303 417 367
rect 301 287 417 303
rect 113 215 143 259
rect 215 215 245 269
rect 301 253 329 287
rect 363 253 417 287
rect 301 237 417 253
rect 301 215 331 237
rect 387 215 417 237
rect 473 335 503 367
rect 559 335 589 367
rect 473 319 589 335
rect 473 285 489 319
rect 523 285 589 319
rect 473 269 589 285
rect 473 215 503 269
rect 559 215 589 269
rect 645 303 675 367
rect 731 303 761 367
rect 817 335 847 367
rect 645 287 761 303
rect 645 253 677 287
rect 711 253 761 287
rect 809 319 875 335
rect 809 285 825 319
rect 859 285 875 319
rect 809 269 875 285
rect 645 237 761 253
rect 645 215 675 237
rect 731 215 761 237
rect 817 215 847 269
rect 113 21 143 47
rect 215 21 245 47
rect 301 21 331 47
rect 387 21 417 47
rect 473 21 503 47
rect 559 21 589 47
rect 645 21 675 47
rect 731 21 761 47
rect 817 21 847 47
<< polycont >>
rect 37 275 71 309
rect 209 285 243 319
rect 329 253 363 287
rect 489 285 523 319
rect 677 253 711 287
rect 825 285 859 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 52 599 106 615
rect 52 565 68 599
rect 102 565 106 599
rect 52 518 106 565
rect 52 484 68 518
rect 102 484 106 518
rect 52 436 106 484
rect 150 607 206 649
rect 150 573 166 607
rect 200 573 206 607
rect 150 531 206 573
rect 240 607 808 613
rect 240 573 256 607
rect 290 573 428 607
rect 462 597 808 607
rect 462 573 600 597
rect 240 565 600 573
rect 598 563 600 565
rect 634 577 772 597
rect 634 563 638 577
rect 150 527 564 531
rect 150 493 514 527
rect 548 493 564 527
rect 150 459 166 493
rect 200 485 564 493
rect 598 525 638 563
rect 768 563 772 577
rect 806 563 808 597
rect 598 491 600 525
rect 634 491 638 525
rect 200 459 216 485
rect 598 475 638 491
rect 682 527 724 543
rect 682 493 686 527
rect 720 493 724 527
rect 150 454 216 459
rect 682 459 724 493
rect 768 525 808 563
rect 768 491 772 525
rect 806 491 808 525
rect 768 475 808 491
rect 842 607 908 649
rect 842 573 858 607
rect 892 573 908 607
rect 842 512 908 573
rect 842 478 858 512
rect 892 478 908 512
rect 842 475 908 478
rect 52 402 68 436
rect 102 420 106 436
rect 326 447 392 451
rect 102 402 157 420
rect 326 413 342 447
rect 376 441 392 447
rect 682 441 686 459
rect 376 425 686 441
rect 720 441 724 459
rect 720 425 940 441
rect 376 413 940 425
rect 326 407 940 413
rect 52 386 157 402
rect 21 309 87 352
rect 21 275 37 309
rect 71 275 87 309
rect 21 269 87 275
rect 123 251 157 386
rect 193 339 861 373
rect 193 319 259 339
rect 193 285 209 319
rect 243 285 259 319
rect 413 319 641 339
rect 313 287 379 303
rect 313 253 329 287
rect 363 253 379 287
rect 413 285 489 319
rect 523 285 641 319
rect 809 319 861 339
rect 675 287 727 303
rect 313 251 379 253
rect 675 253 677 287
rect 711 253 727 287
rect 809 285 825 319
rect 859 285 861 319
rect 809 269 861 285
rect 675 251 727 253
rect 123 235 727 251
rect 895 235 940 407
rect 52 217 727 235
rect 52 203 157 217
rect 52 169 68 203
rect 102 201 157 203
rect 768 203 940 235
rect 102 169 104 201
rect 768 183 772 203
rect 52 101 104 169
rect 240 179 772 183
rect 52 67 68 101
rect 102 67 104 101
rect 52 51 104 67
rect 138 133 154 167
rect 188 133 204 167
rect 138 93 204 133
rect 138 59 154 93
rect 188 59 204 93
rect 138 17 204 59
rect 240 145 256 179
rect 290 149 428 179
rect 290 145 306 149
rect 240 101 306 145
rect 412 145 428 149
rect 462 175 772 179
rect 462 149 600 175
rect 462 145 478 149
rect 240 67 256 101
rect 290 67 306 101
rect 240 51 306 67
rect 340 99 378 115
rect 340 65 342 99
rect 376 65 378 99
rect 340 17 378 65
rect 412 101 478 145
rect 584 141 600 149
rect 634 169 772 175
rect 806 201 940 203
rect 634 149 806 169
rect 634 141 650 149
rect 412 67 428 101
rect 462 67 478 101
rect 412 51 478 67
rect 512 99 550 115
rect 512 65 514 99
rect 548 65 550 99
rect 512 17 550 65
rect 584 101 650 141
rect 584 67 600 101
rect 634 67 650 101
rect 584 51 650 67
rect 684 99 736 115
rect 684 65 686 99
rect 720 65 736 99
rect 684 17 736 65
rect 770 101 806 149
rect 770 67 772 101
rect 770 51 806 67
rect 842 161 908 167
rect 842 127 858 161
rect 892 127 908 161
rect 842 93 908 127
rect 842 59 858 93
rect 892 59 908 93
rect 842 17 908 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor2b_4
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5259928
string GDS_START 5251846
<< end >>
