magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 1 259 839 263
rect 1 49 1631 259
rect 0 0 1632 49
<< scnmos >>
rect 80 69 110 237
rect 166 69 196 237
rect 252 69 282 237
rect 338 69 368 237
rect 424 69 454 237
rect 510 69 540 237
rect 612 69 642 237
rect 714 69 744 237
rect 920 65 950 233
rect 1006 65 1036 233
rect 1092 65 1122 233
rect 1178 65 1208 233
rect 1264 65 1294 233
rect 1350 65 1380 233
rect 1436 65 1466 233
rect 1522 65 1552 233
<< scpmoshvt >>
rect 94 367 124 619
rect 180 367 210 619
rect 266 367 296 619
rect 352 367 382 619
rect 438 367 468 619
rect 524 367 554 619
rect 610 367 640 619
rect 804 367 834 619
rect 890 367 920 619
rect 976 367 1006 619
rect 1062 367 1092 619
rect 1148 367 1178 619
rect 1250 367 1280 619
rect 1336 367 1366 619
rect 1422 367 1452 619
rect 1508 367 1538 619
<< ndiff >>
rect 27 225 80 237
rect 27 191 35 225
rect 69 191 80 225
rect 27 115 80 191
rect 27 81 35 115
rect 69 81 80 115
rect 27 69 80 81
rect 110 183 166 237
rect 110 149 121 183
rect 155 149 166 183
rect 110 111 166 149
rect 110 77 121 111
rect 155 77 166 111
rect 110 69 166 77
rect 196 225 252 237
rect 196 191 207 225
rect 241 191 252 225
rect 196 115 252 191
rect 196 81 207 115
rect 241 81 252 115
rect 196 69 252 81
rect 282 183 338 237
rect 282 149 293 183
rect 327 149 338 183
rect 282 111 338 149
rect 282 77 293 111
rect 327 77 338 111
rect 282 69 338 77
rect 368 225 424 237
rect 368 191 379 225
rect 413 191 424 225
rect 368 115 424 191
rect 368 81 379 115
rect 413 81 424 115
rect 368 69 424 81
rect 454 183 510 237
rect 454 149 465 183
rect 499 149 510 183
rect 454 111 510 149
rect 454 77 465 111
rect 499 77 510 111
rect 454 69 510 77
rect 540 229 612 237
rect 540 195 567 229
rect 601 195 612 229
rect 540 155 612 195
rect 540 121 567 155
rect 601 121 612 155
rect 540 69 612 121
rect 642 183 714 237
rect 642 149 669 183
rect 703 149 714 183
rect 642 111 714 149
rect 642 77 669 111
rect 703 77 714 111
rect 642 69 714 77
rect 744 225 813 237
rect 744 191 771 225
rect 805 191 813 225
rect 744 155 813 191
rect 744 121 771 155
rect 805 121 813 155
rect 744 69 813 121
rect 867 218 920 233
rect 867 184 875 218
rect 909 184 920 218
rect 867 65 920 184
rect 950 118 1006 233
rect 950 84 961 118
rect 995 84 1006 118
rect 950 65 1006 84
rect 1036 225 1092 233
rect 1036 191 1047 225
rect 1081 191 1092 225
rect 1036 153 1092 191
rect 1036 119 1047 153
rect 1081 119 1092 153
rect 1036 65 1092 119
rect 1122 160 1178 233
rect 1122 126 1133 160
rect 1167 126 1178 160
rect 1122 65 1178 126
rect 1208 221 1264 233
rect 1208 187 1219 221
rect 1253 187 1264 221
rect 1208 107 1264 187
rect 1208 73 1219 107
rect 1253 73 1264 107
rect 1208 65 1264 73
rect 1294 181 1350 233
rect 1294 147 1305 181
rect 1339 147 1350 181
rect 1294 107 1350 147
rect 1294 73 1305 107
rect 1339 73 1350 107
rect 1294 65 1350 73
rect 1380 221 1436 233
rect 1380 187 1391 221
rect 1425 187 1436 221
rect 1380 107 1436 187
rect 1380 73 1391 107
rect 1425 73 1436 107
rect 1380 65 1436 73
rect 1466 181 1522 233
rect 1466 147 1477 181
rect 1511 147 1522 181
rect 1466 107 1522 147
rect 1466 73 1477 107
rect 1511 73 1522 107
rect 1466 65 1522 73
rect 1552 221 1605 233
rect 1552 187 1563 221
rect 1597 187 1605 221
rect 1552 111 1605 187
rect 1552 77 1563 111
rect 1597 77 1605 111
rect 1552 65 1605 77
<< pdiff >>
rect 41 599 94 619
rect 41 565 49 599
rect 83 565 94 599
rect 41 518 94 565
rect 41 484 49 518
rect 83 484 94 518
rect 41 436 94 484
rect 41 402 49 436
rect 83 402 94 436
rect 41 367 94 402
rect 124 607 180 619
rect 124 573 135 607
rect 169 573 180 607
rect 124 496 180 573
rect 124 462 135 496
rect 169 462 180 496
rect 124 367 180 462
rect 210 599 266 619
rect 210 565 221 599
rect 255 565 266 599
rect 210 523 266 565
rect 210 489 221 523
rect 255 489 266 523
rect 210 436 266 489
rect 210 402 221 436
rect 255 402 266 436
rect 210 367 266 402
rect 296 607 352 619
rect 296 573 307 607
rect 341 573 352 607
rect 296 496 352 573
rect 296 462 307 496
rect 341 462 352 496
rect 296 367 352 462
rect 382 599 438 619
rect 382 565 393 599
rect 427 565 438 599
rect 382 523 438 565
rect 382 489 393 523
rect 427 489 438 523
rect 382 436 438 489
rect 382 402 393 436
rect 427 402 438 436
rect 382 367 438 402
rect 468 607 524 619
rect 468 573 479 607
rect 513 573 524 607
rect 468 496 524 573
rect 468 462 479 496
rect 513 462 524 496
rect 468 367 524 462
rect 554 599 610 619
rect 554 565 565 599
rect 599 565 610 599
rect 554 528 610 565
rect 554 494 565 528
rect 599 494 610 528
rect 554 436 610 494
rect 554 402 565 436
rect 599 402 610 436
rect 554 367 610 402
rect 640 607 804 619
rect 640 573 651 607
rect 685 573 759 607
rect 793 573 804 607
rect 640 488 804 573
rect 640 454 651 488
rect 685 454 719 488
rect 753 454 804 488
rect 640 367 804 454
rect 834 599 890 619
rect 834 565 845 599
rect 879 565 890 599
rect 834 508 890 565
rect 834 474 845 508
rect 879 474 890 508
rect 834 367 890 474
rect 920 567 976 619
rect 920 533 931 567
rect 965 533 976 567
rect 920 367 976 533
rect 1006 599 1062 619
rect 1006 565 1017 599
rect 1051 565 1062 599
rect 1006 508 1062 565
rect 1006 474 1017 508
rect 1051 474 1062 508
rect 1006 367 1062 474
rect 1092 567 1148 619
rect 1092 533 1103 567
rect 1137 533 1148 567
rect 1092 367 1148 533
rect 1178 599 1250 619
rect 1178 565 1189 599
rect 1223 565 1250 599
rect 1178 508 1250 565
rect 1178 474 1189 508
rect 1223 474 1250 508
rect 1178 367 1250 474
rect 1280 541 1336 619
rect 1280 507 1291 541
rect 1325 507 1336 541
rect 1280 440 1336 507
rect 1280 406 1291 440
rect 1325 406 1336 440
rect 1280 367 1336 406
rect 1366 599 1422 619
rect 1366 565 1377 599
rect 1411 565 1422 599
rect 1366 508 1422 565
rect 1366 474 1377 508
rect 1411 474 1422 508
rect 1366 367 1422 474
rect 1452 542 1508 619
rect 1452 508 1463 542
rect 1497 508 1508 542
rect 1452 440 1508 508
rect 1452 406 1463 440
rect 1497 406 1508 440
rect 1452 367 1508 406
rect 1538 599 1591 619
rect 1538 565 1549 599
rect 1583 565 1591 599
rect 1538 518 1591 565
rect 1538 484 1549 518
rect 1583 484 1591 518
rect 1538 440 1591 484
rect 1538 406 1549 440
rect 1583 406 1591 440
rect 1538 367 1591 406
<< ndiffc >>
rect 35 191 69 225
rect 35 81 69 115
rect 121 149 155 183
rect 121 77 155 111
rect 207 191 241 225
rect 207 81 241 115
rect 293 149 327 183
rect 293 77 327 111
rect 379 191 413 225
rect 379 81 413 115
rect 465 149 499 183
rect 465 77 499 111
rect 567 195 601 229
rect 567 121 601 155
rect 669 149 703 183
rect 669 77 703 111
rect 771 191 805 225
rect 771 121 805 155
rect 875 184 909 218
rect 961 84 995 118
rect 1047 191 1081 225
rect 1047 119 1081 153
rect 1133 126 1167 160
rect 1219 187 1253 221
rect 1219 73 1253 107
rect 1305 147 1339 181
rect 1305 73 1339 107
rect 1391 187 1425 221
rect 1391 73 1425 107
rect 1477 147 1511 181
rect 1477 73 1511 107
rect 1563 187 1597 221
rect 1563 77 1597 111
<< pdiffc >>
rect 49 565 83 599
rect 49 484 83 518
rect 49 402 83 436
rect 135 573 169 607
rect 135 462 169 496
rect 221 565 255 599
rect 221 489 255 523
rect 221 402 255 436
rect 307 573 341 607
rect 307 462 341 496
rect 393 565 427 599
rect 393 489 427 523
rect 393 402 427 436
rect 479 573 513 607
rect 479 462 513 496
rect 565 565 599 599
rect 565 494 599 528
rect 565 402 599 436
rect 651 573 685 607
rect 759 573 793 607
rect 651 454 685 488
rect 719 454 753 488
rect 845 565 879 599
rect 845 474 879 508
rect 931 533 965 567
rect 1017 565 1051 599
rect 1017 474 1051 508
rect 1103 533 1137 567
rect 1189 565 1223 599
rect 1189 474 1223 508
rect 1291 507 1325 541
rect 1291 406 1325 440
rect 1377 565 1411 599
rect 1377 474 1411 508
rect 1463 508 1497 542
rect 1463 406 1497 440
rect 1549 565 1583 599
rect 1549 484 1583 518
rect 1549 406 1583 440
<< poly >>
rect 94 619 124 645
rect 180 619 210 645
rect 266 619 296 645
rect 352 619 382 645
rect 438 619 468 645
rect 524 619 554 645
rect 610 619 640 645
rect 804 619 834 645
rect 890 619 920 645
rect 976 619 1006 645
rect 1062 619 1092 645
rect 1148 619 1178 645
rect 1250 619 1280 645
rect 1336 619 1366 645
rect 1422 619 1452 645
rect 1508 619 1538 645
rect 94 335 124 367
rect 180 335 210 367
rect 266 335 296 367
rect 352 335 382 367
rect 44 319 382 335
rect 44 285 60 319
rect 94 285 128 319
rect 162 285 196 319
rect 230 285 264 319
rect 298 285 332 319
rect 366 285 382 319
rect 438 335 468 367
rect 524 335 554 367
rect 610 335 640 367
rect 804 335 834 367
rect 438 319 834 335
rect 438 299 602 319
rect 44 269 382 285
rect 424 285 602 299
rect 636 285 670 319
rect 704 285 738 319
rect 772 285 834 319
rect 890 335 920 367
rect 976 335 1006 367
rect 1062 335 1092 367
rect 1148 335 1178 367
rect 1250 337 1280 367
rect 1336 337 1366 367
rect 1422 337 1452 367
rect 1508 337 1538 367
rect 890 319 1208 335
rect 890 305 1007 319
rect 424 269 834 285
rect 920 285 1007 305
rect 1041 285 1075 319
rect 1109 285 1143 319
rect 1177 285 1208 319
rect 1250 319 1552 337
rect 1250 307 1366 319
rect 80 237 110 269
rect 166 237 196 269
rect 252 237 282 269
rect 338 237 368 269
rect 424 237 454 269
rect 510 237 540 269
rect 612 237 642 269
rect 714 237 744 269
rect 920 259 1208 285
rect 920 233 950 259
rect 1006 233 1036 259
rect 1092 233 1122 259
rect 1178 233 1208 259
rect 1264 285 1366 307
rect 1400 285 1434 319
rect 1468 285 1502 319
rect 1536 285 1552 319
rect 1264 269 1552 285
rect 1264 233 1294 269
rect 1350 233 1380 269
rect 1436 233 1466 269
rect 1522 233 1552 269
rect 80 43 110 69
rect 166 43 196 69
rect 252 43 282 69
rect 338 43 368 69
rect 424 43 454 69
rect 510 43 540 69
rect 612 43 642 69
rect 714 43 744 69
rect 920 39 950 65
rect 1006 39 1036 65
rect 1092 39 1122 65
rect 1178 39 1208 65
rect 1264 39 1294 65
rect 1350 39 1380 65
rect 1436 39 1466 65
rect 1522 39 1552 65
<< polycont >>
rect 60 285 94 319
rect 128 285 162 319
rect 196 285 230 319
rect 264 285 298 319
rect 332 285 366 319
rect 602 285 636 319
rect 670 285 704 319
rect 738 285 772 319
rect 1007 285 1041 319
rect 1075 285 1109 319
rect 1143 285 1177 319
rect 1366 285 1400 319
rect 1434 285 1468 319
rect 1502 285 1536 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 33 599 85 615
rect 33 565 49 599
rect 83 565 85 599
rect 33 518 85 565
rect 33 484 49 518
rect 83 484 85 518
rect 33 436 85 484
rect 119 607 185 649
rect 119 573 135 607
rect 169 573 185 607
rect 119 496 185 573
rect 119 462 135 496
rect 169 462 185 496
rect 119 454 185 462
rect 219 599 257 615
rect 219 565 221 599
rect 255 565 257 599
rect 219 523 257 565
rect 219 489 221 523
rect 255 489 257 523
rect 33 402 49 436
rect 83 420 85 436
rect 219 436 257 489
rect 291 607 357 649
rect 291 573 307 607
rect 341 573 357 607
rect 291 496 357 573
rect 291 462 307 496
rect 341 462 357 496
rect 291 454 357 462
rect 391 599 429 615
rect 391 565 393 599
rect 427 565 429 599
rect 391 523 429 565
rect 391 489 393 523
rect 427 489 429 523
rect 219 420 221 436
rect 83 402 221 420
rect 255 420 257 436
rect 391 436 429 489
rect 463 607 529 649
rect 463 573 479 607
rect 513 573 529 607
rect 463 496 529 573
rect 463 462 479 496
rect 513 462 529 496
rect 463 454 529 462
rect 563 599 601 615
rect 563 565 565 599
rect 599 565 601 599
rect 563 528 601 565
rect 563 494 565 528
rect 599 494 601 528
rect 391 420 393 436
rect 255 402 393 420
rect 427 420 429 436
rect 563 436 601 494
rect 635 607 803 649
rect 635 573 651 607
rect 685 573 759 607
rect 793 573 803 607
rect 635 528 803 573
rect 837 599 881 615
rect 837 565 845 599
rect 879 565 881 599
rect 635 488 769 528
rect 837 508 881 565
rect 915 567 981 649
rect 915 533 931 567
rect 965 533 981 567
rect 915 526 981 533
rect 1015 599 1053 615
rect 1015 565 1017 599
rect 1051 565 1053 599
rect 837 494 845 508
rect 635 454 651 488
rect 685 454 719 488
rect 753 454 769 488
rect 803 474 845 494
rect 879 492 881 508
rect 1015 508 1053 565
rect 1087 567 1153 649
rect 1087 533 1103 567
rect 1137 533 1153 567
rect 1087 526 1153 533
rect 1187 599 1599 615
rect 1187 565 1189 599
rect 1223 581 1377 599
rect 1223 565 1241 581
rect 1015 492 1017 508
rect 879 474 1017 492
rect 1051 492 1053 508
rect 1187 508 1241 565
rect 1375 565 1377 581
rect 1411 581 1549 599
rect 1411 565 1413 581
rect 1187 492 1189 508
rect 1051 474 1189 492
rect 1223 474 1241 508
rect 803 458 1241 474
rect 1275 541 1341 547
rect 1275 507 1291 541
rect 1325 507 1341 541
rect 563 420 565 436
rect 427 402 565 420
rect 599 420 601 436
rect 803 420 837 458
rect 1275 440 1341 507
rect 1375 508 1413 565
rect 1583 565 1599 599
rect 1375 474 1377 508
rect 1411 474 1413 508
rect 1375 458 1413 474
rect 1447 542 1513 547
rect 1447 508 1463 542
rect 1497 508 1513 542
rect 1275 424 1291 440
rect 599 402 837 420
rect 33 386 837 402
rect 871 406 1291 424
rect 1325 424 1341 440
rect 1447 440 1513 508
rect 1447 424 1463 440
rect 1325 406 1463 424
rect 1497 406 1513 440
rect 871 390 1513 406
rect 1549 518 1599 565
rect 1583 484 1599 518
rect 1549 440 1599 484
rect 1583 406 1599 440
rect 1549 390 1599 406
rect 31 319 545 352
rect 31 285 60 319
rect 94 285 128 319
rect 162 285 196 319
rect 230 285 264 319
rect 298 285 332 319
rect 366 285 545 319
rect 586 319 833 352
rect 586 285 602 319
rect 636 285 670 319
rect 704 285 738 319
rect 772 285 833 319
rect 871 251 941 390
rect 975 319 1313 356
rect 975 285 1007 319
rect 1041 285 1075 319
rect 1109 285 1143 319
rect 1177 285 1313 319
rect 1350 319 1612 356
rect 1350 285 1366 319
rect 1400 285 1434 319
rect 1468 285 1502 319
rect 1536 285 1612 319
rect 19 229 821 251
rect 19 225 567 229
rect 19 191 35 225
rect 69 217 207 225
rect 19 115 69 191
rect 205 191 207 217
rect 241 217 379 225
rect 241 191 243 217
rect 19 81 35 115
rect 19 65 69 81
rect 105 149 121 183
rect 155 149 171 183
rect 105 111 171 149
rect 105 77 121 111
rect 155 77 171 111
rect 105 17 171 77
rect 205 115 243 191
rect 377 191 379 217
rect 413 217 567 225
rect 413 191 415 217
rect 205 81 207 115
rect 241 81 243 115
rect 205 65 243 81
rect 277 149 293 183
rect 327 149 343 183
rect 277 111 343 149
rect 277 77 293 111
rect 327 77 343 111
rect 277 17 343 77
rect 377 115 415 191
rect 551 195 567 217
rect 601 225 821 229
rect 601 217 771 225
rect 601 195 617 217
rect 377 81 379 115
rect 413 81 415 115
rect 377 65 415 81
rect 449 149 465 183
rect 499 149 515 183
rect 449 111 515 149
rect 551 155 617 195
rect 755 191 771 217
rect 805 191 821 225
rect 551 121 567 155
rect 601 121 617 155
rect 551 119 617 121
rect 653 149 669 183
rect 703 149 719 183
rect 449 77 465 111
rect 499 85 515 111
rect 653 111 719 149
rect 755 155 821 191
rect 871 225 1613 251
rect 871 218 1047 225
rect 871 184 875 218
rect 909 191 1047 218
rect 1081 221 1613 225
rect 1081 210 1219 221
rect 1081 191 1097 210
rect 909 184 1097 191
rect 871 168 1097 184
rect 1215 187 1219 210
rect 1253 215 1391 221
rect 1253 187 1255 215
rect 755 121 771 155
rect 805 121 821 155
rect 1031 153 1097 168
rect 755 119 821 121
rect 653 85 669 111
rect 499 77 669 85
rect 703 85 719 111
rect 945 118 997 134
rect 1031 119 1047 153
rect 1081 119 1097 153
rect 1131 160 1171 176
rect 1131 126 1133 160
rect 1167 126 1171 160
rect 945 85 961 118
rect 703 84 961 85
rect 995 85 997 118
rect 1131 85 1171 126
rect 995 84 1171 85
rect 703 77 1171 84
rect 449 51 1171 77
rect 1215 107 1255 187
rect 1389 187 1391 215
rect 1425 215 1563 221
rect 1425 187 1427 215
rect 1215 73 1219 107
rect 1253 73 1255 107
rect 1215 57 1255 73
rect 1289 147 1305 181
rect 1339 147 1355 181
rect 1289 107 1355 147
rect 1289 73 1305 107
rect 1339 73 1355 107
rect 1289 17 1355 73
rect 1389 107 1427 187
rect 1597 187 1613 221
rect 1389 73 1391 107
rect 1425 73 1427 107
rect 1389 57 1427 73
rect 1461 147 1477 181
rect 1511 147 1527 181
rect 1461 107 1527 147
rect 1461 73 1477 107
rect 1511 73 1527 107
rect 1461 17 1527 73
rect 1563 111 1613 187
rect 1597 77 1613 111
rect 1563 61 1613 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a31oi_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3418222
string GDS_START 3403704
<< end >>
