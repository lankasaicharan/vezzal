magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 1 172 189 250
rect 566 172 937 256
rect 1 49 937 172
rect 0 0 960 49
<< scnmos >>
rect 80 56 110 224
rect 277 62 307 146
rect 363 62 393 146
rect 449 62 479 146
rect 645 146 675 230
rect 723 146 753 230
rect 828 62 858 230
<< scpmoshvt >>
rect 108 367 138 619
rect 285 428 315 512
rect 371 428 401 512
rect 477 428 507 512
rect 645 428 675 512
rect 731 428 761 512
rect 844 367 874 619
<< ndiff >>
rect 27 212 80 224
rect 27 178 35 212
rect 69 178 80 212
rect 27 102 80 178
rect 27 68 35 102
rect 69 68 80 102
rect 27 56 80 68
rect 110 196 163 224
rect 110 162 121 196
rect 155 162 163 196
rect 110 102 163 162
rect 592 201 645 230
rect 110 68 121 102
rect 155 68 163 102
rect 110 56 163 68
rect 224 121 277 146
rect 224 87 232 121
rect 266 87 277 121
rect 224 62 277 87
rect 307 121 363 146
rect 307 87 318 121
rect 352 87 363 121
rect 307 62 363 87
rect 393 121 449 146
rect 393 87 404 121
rect 438 87 449 121
rect 393 62 449 87
rect 479 121 532 146
rect 479 87 490 121
rect 524 87 532 121
rect 479 62 532 87
rect 592 167 600 201
rect 634 167 645 201
rect 592 146 645 167
rect 675 146 723 230
rect 753 202 828 230
rect 753 168 774 202
rect 808 168 828 202
rect 753 146 828 168
rect 775 108 828 146
rect 775 74 783 108
rect 817 74 828 108
rect 775 62 828 74
rect 858 202 911 230
rect 858 168 869 202
rect 903 168 911 202
rect 858 108 911 168
rect 858 74 869 108
rect 903 74 911 108
rect 858 62 911 74
<< pdiff >>
rect 55 599 108 619
rect 55 565 63 599
rect 97 565 108 599
rect 55 503 108 565
rect 55 469 63 503
rect 97 469 108 503
rect 55 413 108 469
rect 55 379 63 413
rect 97 379 108 413
rect 55 367 108 379
rect 138 607 191 619
rect 138 573 149 607
rect 183 573 191 607
rect 138 512 191 573
rect 791 607 844 619
rect 791 573 799 607
rect 833 573 844 607
rect 791 512 844 573
rect 138 478 149 512
rect 183 478 285 512
rect 138 428 285 478
rect 315 485 371 512
rect 315 451 326 485
rect 360 451 371 485
rect 315 428 371 451
rect 401 428 477 512
rect 507 504 645 512
rect 507 470 528 504
rect 562 470 600 504
rect 634 470 645 504
rect 507 428 645 470
rect 675 485 731 512
rect 675 451 686 485
rect 720 451 731 485
rect 675 428 731 451
rect 761 503 844 512
rect 761 469 772 503
rect 806 469 844 503
rect 761 428 844 469
rect 138 413 191 428
rect 138 379 149 413
rect 183 379 191 413
rect 138 367 191 379
rect 791 413 844 428
rect 791 379 799 413
rect 833 379 844 413
rect 791 367 844 379
rect 874 599 927 619
rect 874 565 885 599
rect 919 565 927 599
rect 874 502 927 565
rect 874 468 885 502
rect 919 468 927 502
rect 874 413 927 468
rect 874 379 885 413
rect 919 379 927 413
rect 874 367 927 379
<< ndiffc >>
rect 35 178 69 212
rect 35 68 69 102
rect 121 162 155 196
rect 121 68 155 102
rect 232 87 266 121
rect 318 87 352 121
rect 404 87 438 121
rect 490 87 524 121
rect 600 167 634 201
rect 774 168 808 202
rect 783 74 817 108
rect 869 168 903 202
rect 869 74 903 108
<< pdiffc >>
rect 63 565 97 599
rect 63 469 97 503
rect 63 379 97 413
rect 149 573 183 607
rect 799 573 833 607
rect 149 478 183 512
rect 326 451 360 485
rect 528 470 562 504
rect 600 470 634 504
rect 686 451 720 485
rect 772 469 806 503
rect 149 379 183 413
rect 799 379 833 413
rect 885 565 919 599
rect 885 468 919 502
rect 885 379 919 413
<< poly >>
rect 108 619 138 645
rect 844 619 874 645
rect 285 512 315 538
rect 371 512 401 538
rect 477 512 507 538
rect 645 512 675 538
rect 731 512 761 538
rect 285 386 315 428
rect 223 370 315 386
rect 371 380 401 428
rect 108 312 138 367
rect 223 336 239 370
rect 273 356 315 370
rect 273 336 307 356
rect 223 320 307 336
rect 80 296 159 312
rect 80 262 109 296
rect 143 262 159 296
rect 80 246 159 262
rect 80 224 110 246
rect 277 146 307 320
rect 363 354 429 380
rect 363 320 379 354
rect 413 320 429 354
rect 363 286 429 320
rect 363 252 379 286
rect 413 252 429 286
rect 363 236 429 252
rect 477 366 507 428
rect 477 350 543 366
rect 477 316 493 350
rect 527 316 543 350
rect 645 318 675 428
rect 731 396 761 428
rect 477 300 543 316
rect 591 302 675 318
rect 363 146 393 236
rect 477 198 507 300
rect 591 268 607 302
rect 641 268 675 302
rect 591 252 675 268
rect 645 230 675 252
rect 723 366 761 396
rect 723 230 753 366
rect 844 318 874 367
rect 795 302 874 318
rect 795 268 811 302
rect 845 268 874 302
rect 795 252 874 268
rect 828 230 858 252
rect 449 168 577 198
rect 449 146 479 168
rect 547 72 577 168
rect 645 120 675 146
rect 723 72 753 146
rect 80 30 110 56
rect 277 36 307 62
rect 363 36 393 62
rect 449 36 479 62
rect 547 42 753 72
rect 828 36 858 62
<< polycont >>
rect 239 336 273 370
rect 109 262 143 296
rect 379 320 413 354
rect 379 252 413 286
rect 493 316 527 350
rect 607 268 641 302
rect 811 268 845 302
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 19 599 101 615
rect 19 565 63 599
rect 97 565 101 599
rect 19 503 101 565
rect 19 469 63 503
rect 97 469 101 503
rect 19 413 101 469
rect 19 379 63 413
rect 97 379 101 413
rect 19 348 101 379
rect 145 607 205 649
rect 145 573 149 607
rect 183 573 205 607
rect 145 512 205 573
rect 145 478 149 512
rect 183 478 205 512
rect 145 413 205 478
rect 145 379 149 413
rect 183 379 205 413
rect 145 363 205 379
rect 239 535 494 577
rect 239 370 273 535
rect 19 212 73 348
rect 239 320 273 336
rect 309 485 376 501
rect 309 451 326 485
rect 360 451 376 485
rect 309 435 376 451
rect 107 296 159 312
rect 107 262 109 296
rect 143 280 159 296
rect 309 280 343 435
rect 460 420 494 535
rect 528 504 650 649
rect 562 470 600 504
rect 634 470 650 504
rect 770 607 845 649
rect 770 573 799 607
rect 833 573 845 607
rect 770 503 845 573
rect 528 454 650 470
rect 684 485 736 501
rect 684 451 686 485
rect 720 451 736 485
rect 684 420 736 451
rect 460 386 736 420
rect 143 262 343 280
rect 107 246 343 262
rect 377 354 429 370
rect 377 320 379 354
rect 413 320 429 354
rect 377 286 429 320
rect 463 350 558 352
rect 463 316 493 350
rect 527 316 558 350
rect 463 314 558 316
rect 377 252 379 286
rect 413 280 429 286
rect 592 302 654 352
rect 592 280 607 302
rect 413 268 607 280
rect 641 268 654 302
rect 413 252 654 268
rect 377 246 654 252
rect 688 318 736 386
rect 770 469 772 503
rect 806 469 845 503
rect 770 413 845 469
rect 770 379 799 413
rect 833 379 845 413
rect 770 363 845 379
rect 879 599 943 615
rect 879 565 885 599
rect 919 565 943 599
rect 879 502 943 565
rect 879 468 885 502
rect 919 468 943 502
rect 879 413 943 468
rect 879 379 885 413
rect 919 379 943 413
rect 688 302 845 318
rect 688 268 811 302
rect 688 252 845 268
rect 19 178 35 212
rect 69 178 73 212
rect 19 102 73 178
rect 19 68 35 102
rect 69 68 73 102
rect 19 52 73 68
rect 107 196 171 212
rect 107 162 121 196
rect 155 162 171 196
rect 107 102 171 162
rect 107 68 121 102
rect 155 68 171 102
rect 216 121 274 246
rect 377 236 429 246
rect 688 212 724 252
rect 879 218 943 379
rect 216 87 232 121
rect 266 87 274 121
rect 216 71 274 87
rect 308 168 540 202
rect 308 121 354 168
rect 308 87 318 121
rect 352 87 354 121
rect 308 71 354 87
rect 388 121 454 134
rect 388 87 404 121
rect 438 87 454 121
rect 107 17 171 68
rect 388 17 454 87
rect 488 121 540 168
rect 584 201 724 212
rect 584 167 600 201
rect 634 167 724 201
rect 584 151 724 167
rect 758 202 831 218
rect 758 168 774 202
rect 808 168 831 202
rect 488 87 490 121
rect 524 87 540 121
rect 488 71 540 87
rect 758 108 831 168
rect 758 74 783 108
rect 817 74 831 108
rect 758 17 831 74
rect 865 202 943 218
rect 865 168 869 202
rect 903 168 943 202
rect 865 108 943 168
rect 865 74 869 108
rect 903 74 943 108
rect 865 58 943 74
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ha_1
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 895 94 929 128 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 895 464 929 498 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 895 538 929 572 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6678532
string GDS_START 6669326
<< end >>
