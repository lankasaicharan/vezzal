magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4370 1975
<< nwell >>
rect -38 331 3110 704
<< pwell >>
rect 1735 229 1999 273
rect 2761 260 3071 272
rect 1050 228 1999 229
rect 2269 228 3071 260
rect 1050 183 3071 228
rect 831 157 3071 183
rect 57 49 3071 157
rect 0 0 3072 49
<< scnmos >>
rect 136 47 166 131
rect 222 47 252 131
rect 294 47 324 131
rect 448 47 478 131
rect 533 47 563 131
rect 619 47 649 131
rect 910 73 940 157
rect 1129 119 1159 203
rect 1215 119 1245 203
rect 1287 119 1317 203
rect 1545 119 1575 203
rect 1617 119 1647 203
rect 1818 119 1848 247
rect 1890 119 1920 247
rect 1995 118 2025 202
rect 2067 118 2097 202
rect 2139 118 2169 202
rect 2348 150 2378 234
rect 2552 150 2582 234
rect 2844 78 2874 246
rect 2962 78 2992 246
<< scpmoshvt >>
rect 87 481 117 609
rect 173 481 203 609
rect 245 481 275 609
rect 353 481 383 609
rect 425 481 455 609
rect 610 481 640 609
rect 871 441 901 569
rect 1116 463 1146 547
rect 1202 463 1232 547
rect 1274 463 1304 547
rect 1405 463 1435 547
rect 1491 463 1521 547
rect 1788 379 1818 547
rect 1890 404 1920 572
rect 1995 488 2025 572
rect 2067 488 2097 572
rect 2240 488 2270 572
rect 2464 484 2494 568
rect 2618 440 2648 568
rect 2844 367 2874 619
rect 2930 367 2960 619
<< ndiff >>
rect 1076 167 1129 203
rect 83 106 136 131
rect 83 72 91 106
rect 125 72 136 106
rect 83 47 136 72
rect 166 106 222 131
rect 166 72 177 106
rect 211 72 222 106
rect 166 47 222 72
rect 252 47 294 131
rect 324 106 448 131
rect 324 72 335 106
rect 369 72 403 106
rect 437 72 448 106
rect 324 47 448 72
rect 478 47 533 131
rect 563 92 619 131
rect 563 58 574 92
rect 608 58 619 92
rect 563 47 619 58
rect 649 116 702 131
rect 649 82 660 116
rect 694 82 702 116
rect 649 47 702 82
rect 857 130 910 157
rect 857 96 865 130
rect 899 96 910 130
rect 857 73 910 96
rect 940 130 993 157
rect 940 96 951 130
rect 985 96 993 130
rect 1076 133 1084 167
rect 1118 133 1129 167
rect 1076 119 1129 133
rect 1159 178 1215 203
rect 1159 144 1170 178
rect 1204 144 1215 178
rect 1159 119 1215 144
rect 1245 119 1287 203
rect 1317 165 1370 203
rect 1317 131 1328 165
rect 1362 131 1370 165
rect 1317 119 1370 131
rect 1761 203 1818 247
rect 940 73 993 96
rect 1492 165 1545 203
rect 1492 131 1500 165
rect 1534 131 1545 165
rect 1492 119 1545 131
rect 1575 119 1617 203
rect 1647 166 1818 203
rect 1647 132 1773 166
rect 1807 132 1818 166
rect 1647 119 1818 132
rect 1848 119 1890 247
rect 1920 202 1973 247
rect 2295 209 2348 234
rect 1920 178 1995 202
rect 1920 144 1931 178
rect 1965 144 1995 178
rect 1920 119 1995 144
rect 1945 118 1995 119
rect 2025 118 2067 202
rect 2097 118 2139 202
rect 2169 176 2222 202
rect 2169 142 2180 176
rect 2214 142 2222 176
rect 2295 175 2303 209
rect 2337 175 2348 209
rect 2295 150 2348 175
rect 2378 200 2552 234
rect 2378 166 2389 200
rect 2423 166 2457 200
rect 2491 166 2552 200
rect 2378 150 2552 166
rect 2582 208 2635 234
rect 2787 238 2844 246
rect 2582 174 2593 208
rect 2627 174 2635 208
rect 2787 204 2799 238
rect 2833 204 2844 238
rect 2582 150 2635 174
rect 2169 118 2222 142
rect 2787 78 2844 204
rect 2874 98 2962 246
rect 2874 78 2901 98
rect 2889 64 2901 78
rect 2935 78 2962 98
rect 2992 234 3045 246
rect 2992 200 3003 234
rect 3037 200 3045 234
rect 2992 126 3045 200
rect 2992 92 3003 126
rect 3037 92 3045 126
rect 2992 78 3045 92
rect 2935 64 2947 78
rect 2889 56 2947 64
<< pdiff >>
rect 799 627 849 639
rect 34 597 87 609
rect 34 563 42 597
rect 76 563 87 597
rect 34 527 87 563
rect 34 493 42 527
rect 76 493 87 527
rect 34 481 87 493
rect 117 601 173 609
rect 117 567 128 601
rect 162 567 173 601
rect 117 527 173 567
rect 117 493 128 527
rect 162 493 173 527
rect 117 481 173 493
rect 203 481 245 609
rect 275 601 353 609
rect 275 567 308 601
rect 342 567 353 601
rect 275 533 353 567
rect 275 499 308 533
rect 342 499 353 533
rect 275 481 353 499
rect 383 481 425 609
rect 455 601 610 609
rect 455 567 497 601
rect 531 567 610 601
rect 455 481 610 567
rect 640 529 693 609
rect 640 495 651 529
rect 685 495 693 529
rect 640 481 693 495
rect 799 593 807 627
rect 841 593 849 627
rect 799 569 849 593
rect 799 441 871 569
rect 901 487 954 569
rect 1536 562 1773 572
rect 1536 547 1548 562
rect 901 453 912 487
rect 946 453 954 487
rect 1063 522 1116 547
rect 1063 488 1071 522
rect 1105 488 1116 522
rect 1063 463 1116 488
rect 1146 522 1202 547
rect 1146 488 1157 522
rect 1191 488 1202 522
rect 1146 463 1202 488
rect 1232 463 1274 547
rect 1304 522 1405 547
rect 1304 488 1317 522
rect 1351 488 1405 522
rect 1304 463 1405 488
rect 1435 522 1491 547
rect 1435 488 1446 522
rect 1480 488 1491 522
rect 1435 463 1491 488
rect 1521 528 1548 547
rect 1582 528 1638 562
rect 1672 528 1727 562
rect 1761 547 1773 562
rect 2791 599 2844 619
rect 1840 547 1890 572
rect 1761 528 1788 547
rect 1521 463 1788 528
rect 901 441 954 453
rect 1738 379 1788 463
rect 1818 404 1890 547
rect 1920 560 1995 572
rect 1920 526 1941 560
rect 1975 526 1995 560
rect 1920 488 1995 526
rect 2025 488 2067 572
rect 2097 562 2240 572
rect 2097 528 2108 562
rect 2142 528 2195 562
rect 2229 528 2240 562
rect 2097 488 2240 528
rect 2270 548 2323 572
rect 2270 514 2281 548
rect 2315 514 2323 548
rect 2270 488 2323 514
rect 2411 543 2464 568
rect 2411 509 2419 543
rect 2453 509 2464 543
rect 1920 474 1973 488
rect 1920 440 1931 474
rect 1965 440 1973 474
rect 1920 404 1973 440
rect 1818 379 1868 404
rect 2411 484 2464 509
rect 2494 556 2618 568
rect 2494 522 2573 556
rect 2607 522 2618 556
rect 2494 486 2618 522
rect 2494 484 2573 486
rect 2565 452 2573 484
rect 2607 452 2618 486
rect 2565 440 2618 452
rect 2648 556 2701 568
rect 2648 522 2659 556
rect 2693 522 2701 556
rect 2648 486 2701 522
rect 2648 452 2659 486
rect 2693 452 2701 486
rect 2648 440 2701 452
rect 2791 565 2799 599
rect 2833 565 2844 599
rect 2791 506 2844 565
rect 2791 472 2799 506
rect 2833 472 2844 506
rect 2791 413 2844 472
rect 2791 379 2799 413
rect 2833 379 2844 413
rect 2791 367 2844 379
rect 2874 611 2930 619
rect 2874 577 2885 611
rect 2919 577 2930 611
rect 2874 511 2930 577
rect 2874 477 2885 511
rect 2919 477 2930 511
rect 2874 418 2930 477
rect 2874 384 2885 418
rect 2919 384 2930 418
rect 2874 367 2930 384
rect 2960 599 3013 619
rect 2960 565 2971 599
rect 3005 565 3013 599
rect 2960 506 3013 565
rect 2960 472 2971 506
rect 3005 472 3013 506
rect 2960 418 3013 472
rect 2960 384 2971 418
rect 3005 384 3013 418
rect 2960 367 3013 384
<< ndiffc >>
rect 91 72 125 106
rect 177 72 211 106
rect 335 72 369 106
rect 403 72 437 106
rect 574 58 608 92
rect 660 82 694 116
rect 865 96 899 130
rect 951 96 985 130
rect 1084 133 1118 167
rect 1170 144 1204 178
rect 1328 131 1362 165
rect 1500 131 1534 165
rect 1773 132 1807 166
rect 1931 144 1965 178
rect 2180 142 2214 176
rect 2303 175 2337 209
rect 2389 166 2423 200
rect 2457 166 2491 200
rect 2593 174 2627 208
rect 2799 204 2833 238
rect 2901 64 2935 98
rect 3003 200 3037 234
rect 3003 92 3037 126
<< pdiffc >>
rect 42 563 76 597
rect 42 493 76 527
rect 128 567 162 601
rect 128 493 162 527
rect 308 567 342 601
rect 308 499 342 533
rect 497 567 531 601
rect 651 495 685 529
rect 807 593 841 627
rect 912 453 946 487
rect 1071 488 1105 522
rect 1157 488 1191 522
rect 1317 488 1351 522
rect 1446 488 1480 522
rect 1548 528 1582 562
rect 1638 528 1672 562
rect 1727 528 1761 562
rect 1941 526 1975 560
rect 2108 528 2142 562
rect 2195 528 2229 562
rect 2281 514 2315 548
rect 2419 509 2453 543
rect 1931 440 1965 474
rect 2573 522 2607 556
rect 2573 452 2607 486
rect 2659 522 2693 556
rect 2659 452 2693 486
rect 2799 565 2833 599
rect 2799 472 2833 506
rect 2799 379 2833 413
rect 2885 577 2919 611
rect 2885 477 2919 511
rect 2885 384 2919 418
rect 2971 565 3005 599
rect 2971 472 3005 506
rect 2971 384 3005 418
<< poly >>
rect 87 609 117 635
rect 173 609 203 635
rect 245 609 275 635
rect 353 609 383 635
rect 425 609 455 635
rect 610 609 640 635
rect 871 615 1920 645
rect 2844 619 2874 645
rect 2930 619 2960 645
rect 871 569 901 615
rect 87 449 117 481
rect 173 449 203 481
rect 43 433 203 449
rect 43 399 127 433
rect 161 399 203 433
rect 43 383 203 399
rect 245 405 275 481
rect 245 389 311 405
rect 43 183 73 383
rect 245 355 261 389
rect 295 355 311 389
rect 245 339 311 355
rect 353 291 383 481
rect 425 441 455 481
rect 425 425 563 441
rect 425 411 511 425
rect 495 391 511 411
rect 545 391 563 425
rect 495 375 563 391
rect 121 275 383 291
rect 121 241 137 275
rect 171 261 383 275
rect 425 317 491 333
rect 425 283 441 317
rect 475 283 491 317
rect 171 241 252 261
rect 121 225 252 241
rect 43 153 166 183
rect 136 131 166 153
rect 222 131 252 225
rect 425 249 491 283
rect 294 203 383 219
rect 294 169 333 203
rect 367 169 383 203
rect 425 215 441 249
rect 475 215 491 249
rect 425 199 491 215
rect 294 153 383 169
rect 294 131 324 153
rect 448 131 478 199
rect 533 131 563 375
rect 610 332 640 481
rect 1116 547 1146 573
rect 1202 547 1232 615
rect 1274 547 1304 573
rect 1405 547 1435 573
rect 1491 547 1521 573
rect 1788 547 1818 573
rect 1890 572 1920 615
rect 1995 572 2025 598
rect 2067 572 2097 598
rect 2240 572 2270 598
rect 610 302 649 332
rect 871 313 901 441
rect 1116 409 1146 463
rect 1202 437 1232 463
rect 619 286 721 302
rect 619 252 671 286
rect 705 252 721 286
rect 619 218 721 252
rect 619 184 671 218
rect 705 184 721 218
rect 619 168 721 184
rect 775 297 901 313
rect 775 263 791 297
rect 825 283 901 297
rect 969 393 1146 409
rect 1274 431 1304 463
rect 1274 415 1357 431
rect 1274 401 1307 415
rect 969 359 985 393
rect 1019 359 1146 393
rect 969 341 1146 359
rect 1287 381 1307 401
rect 1341 381 1357 415
rect 1287 365 1357 381
rect 969 325 1245 341
rect 969 291 985 325
rect 1019 291 1195 325
rect 1229 291 1245 325
rect 825 263 841 283
rect 969 275 1245 291
rect 775 229 841 263
rect 775 195 791 229
rect 825 209 841 229
rect 825 195 940 209
rect 1129 203 1159 229
rect 1215 203 1245 275
rect 1287 203 1317 365
rect 1405 255 1435 463
rect 1491 424 1521 463
rect 1477 408 1647 424
rect 1477 374 1493 408
rect 1527 374 1647 408
rect 2464 568 2494 594
rect 2618 568 2648 594
rect 1477 358 1647 374
rect 1398 225 1575 255
rect 1398 223 1464 225
rect 775 179 940 195
rect 619 131 649 168
rect 910 157 940 179
rect 1398 189 1414 223
rect 1448 189 1464 223
rect 1545 203 1575 225
rect 1617 203 1647 358
rect 1788 336 1818 379
rect 1890 378 1920 404
rect 1995 336 2025 488
rect 1689 320 1818 336
rect 1689 286 1705 320
rect 1739 300 1818 320
rect 1890 320 2025 336
rect 1739 286 1848 300
rect 1689 270 1848 286
rect 1818 247 1848 270
rect 1890 286 1908 320
rect 1942 306 2025 320
rect 2067 366 2097 488
rect 2240 440 2270 488
rect 2464 452 2494 484
rect 2240 424 2306 440
rect 2240 390 2256 424
rect 2290 390 2306 424
rect 2240 374 2306 390
rect 2464 436 2533 452
rect 2464 402 2483 436
rect 2517 425 2533 436
rect 2618 425 2648 440
rect 2517 402 2648 425
rect 2464 395 2648 402
rect 2067 350 2198 366
rect 2067 316 2148 350
rect 2182 316 2198 350
rect 1942 286 1998 306
rect 1890 270 1998 286
rect 2067 300 2198 316
rect 1890 247 1920 270
rect 1398 155 1464 189
rect 1398 121 1414 155
rect 1448 121 1464 155
rect 910 51 940 73
rect 1129 51 1159 119
rect 1215 93 1245 119
rect 1287 93 1317 119
rect 1398 105 1464 121
rect 1995 202 2025 228
rect 2067 202 2097 300
rect 2246 258 2276 374
rect 2464 368 2533 395
rect 2464 348 2483 368
rect 2139 228 2276 258
rect 2348 334 2483 348
rect 2517 348 2533 368
rect 2679 350 2745 366
rect 2517 334 2582 348
rect 2348 318 2582 334
rect 2348 234 2378 318
rect 2552 234 2582 318
rect 2679 316 2695 350
rect 2729 316 2745 350
rect 2679 298 2745 316
rect 2844 298 2874 367
rect 2930 334 2960 367
rect 2679 282 2874 298
rect 2679 248 2695 282
rect 2729 268 2874 282
rect 2917 318 2992 334
rect 2917 284 2933 318
rect 2967 284 2992 318
rect 2917 268 2992 284
rect 2729 248 2745 268
rect 2139 202 2169 228
rect 1545 93 1575 119
rect 1617 93 1647 119
rect 1818 93 1848 119
rect 1890 93 1920 119
rect 2679 232 2745 248
rect 2844 246 2874 268
rect 2962 246 2992 268
rect 2681 168 2747 184
rect 2348 124 2378 150
rect 2552 135 2582 150
rect 2681 135 2697 168
rect 2552 134 2697 135
rect 2731 134 2747 168
rect 1995 51 2025 118
rect 2067 92 2097 118
rect 2139 92 2169 118
rect 2552 105 2747 134
rect 2681 100 2747 105
rect 136 21 166 47
rect 222 21 252 47
rect 294 21 324 47
rect 448 21 478 47
rect 533 21 563 47
rect 619 21 649 47
rect 910 21 2025 51
rect 2681 66 2697 100
rect 2731 66 2747 100
rect 2681 50 2747 66
rect 2844 52 2874 78
rect 2962 52 2992 78
<< polycont >>
rect 127 399 161 433
rect 261 355 295 389
rect 511 391 545 425
rect 137 241 171 275
rect 441 283 475 317
rect 333 169 367 203
rect 441 215 475 249
rect 671 252 705 286
rect 671 184 705 218
rect 791 263 825 297
rect 985 359 1019 393
rect 1307 381 1341 415
rect 985 291 1019 325
rect 1195 291 1229 325
rect 791 195 825 229
rect 1493 374 1527 408
rect 1414 189 1448 223
rect 1705 286 1739 320
rect 1908 286 1942 320
rect 2256 390 2290 424
rect 2483 402 2517 436
rect 2148 316 2182 350
rect 1414 121 1448 155
rect 2483 334 2517 368
rect 2695 316 2729 350
rect 2695 248 2729 282
rect 2933 284 2967 318
rect 2697 134 2731 168
rect 2697 66 2731 100
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 26 597 78 613
rect 26 563 42 597
rect 76 563 78 597
rect 26 527 78 563
rect 26 493 42 527
rect 76 493 78 527
rect 112 601 178 649
rect 112 567 128 601
rect 162 567 178 601
rect 112 527 178 567
rect 112 493 128 527
rect 162 493 178 527
rect 292 601 358 605
rect 292 567 308 601
rect 342 567 358 601
rect 292 533 358 567
rect 481 601 547 649
rect 791 627 857 649
rect 481 567 497 601
rect 531 567 547 601
rect 481 563 547 567
rect 581 579 755 613
rect 791 593 807 627
rect 841 593 857 627
rect 791 591 857 593
rect 292 499 308 533
rect 342 529 358 533
rect 581 529 615 579
rect 721 557 755 579
rect 342 499 615 529
rect 292 495 615 499
rect 26 291 78 493
rect 112 433 475 459
rect 112 399 127 433
rect 161 425 475 433
rect 161 399 187 425
rect 112 383 187 399
rect 221 355 261 389
rect 295 355 311 389
rect 26 275 187 291
rect 26 241 137 275
rect 171 241 187 275
rect 26 225 187 241
rect 26 122 76 225
rect 221 203 383 355
rect 221 169 333 203
rect 367 169 383 203
rect 425 317 475 425
rect 425 283 441 317
rect 425 249 475 283
rect 425 215 441 249
rect 509 425 547 441
rect 509 391 511 425
rect 545 391 547 425
rect 509 216 547 391
rect 425 199 475 215
rect 221 153 383 169
rect 581 165 615 495
rect 649 529 687 545
rect 649 495 651 529
rect 685 495 687 529
rect 721 523 1115 557
rect 649 487 687 495
rect 1055 522 1115 523
rect 1055 488 1071 522
rect 1105 488 1115 522
rect 649 446 825 487
rect 655 286 751 377
rect 655 252 671 286
rect 705 252 751 286
rect 655 218 751 252
rect 655 184 671 218
rect 705 184 751 218
rect 655 166 751 184
rect 785 297 825 446
rect 785 263 791 297
rect 896 453 912 487
rect 946 453 1021 487
rect 896 393 1021 453
rect 896 359 985 393
rect 1019 359 1021 393
rect 896 325 1021 359
rect 896 291 985 325
rect 1019 291 1021 325
rect 896 275 1021 291
rect 1055 472 1115 488
rect 1149 522 1207 538
rect 1149 488 1157 522
rect 1191 488 1207 522
rect 785 229 825 263
rect 785 195 791 229
rect 474 131 615 165
rect 785 132 825 195
rect 26 106 127 122
rect 474 119 508 131
rect 26 72 91 106
rect 125 72 127 106
rect 26 56 127 72
rect 161 106 227 119
rect 161 72 177 106
rect 211 72 227 106
rect 161 17 227 72
rect 319 106 508 119
rect 319 72 335 106
rect 369 72 403 106
rect 437 72 508 106
rect 658 116 825 132
rect 319 56 508 72
rect 558 92 624 97
rect 558 58 574 92
rect 608 58 624 92
rect 658 82 660 116
rect 694 82 825 116
rect 658 66 825 82
rect 859 130 907 146
rect 859 96 865 130
rect 899 96 907 130
rect 558 17 624 58
rect 859 17 907 96
rect 941 130 1001 275
rect 1055 207 1091 472
rect 1149 411 1207 488
rect 1301 522 1367 649
rect 1530 562 1777 649
rect 1301 488 1317 522
rect 1351 488 1367 522
rect 1301 472 1367 488
rect 1401 522 1496 538
rect 1530 528 1548 562
rect 1582 528 1638 562
rect 1672 528 1727 562
rect 1761 528 1777 562
rect 1929 560 2030 576
rect 1401 488 1446 522
rect 1480 494 1496 522
rect 1929 526 1941 560
rect 1975 526 2030 560
rect 2092 562 2245 649
rect 2092 528 2108 562
rect 2142 528 2195 562
rect 2229 528 2245 562
rect 2279 581 2537 615
rect 2279 548 2331 581
rect 1929 494 2030 526
rect 2279 514 2281 548
rect 2315 514 2331 548
rect 2279 494 2331 514
rect 1480 488 1895 494
rect 1401 460 1895 488
rect 1401 438 1435 460
rect 1125 377 1207 411
rect 1291 415 1435 438
rect 1291 381 1307 415
rect 1341 381 1435 415
rect 1469 424 1529 426
rect 1469 390 1471 424
rect 1505 408 1529 424
rect 1125 241 1159 377
rect 1469 374 1493 390
rect 1527 374 1529 408
rect 1861 390 1895 460
rect 1929 474 2331 494
rect 1929 440 1931 474
rect 1965 460 2331 474
rect 2395 543 2469 547
rect 2395 509 2419 543
rect 2453 509 2469 543
rect 2395 493 2469 509
rect 1965 440 2096 460
rect 1929 424 2096 440
rect 1469 358 1529 374
rect 1563 356 1825 390
rect 1861 356 2026 390
rect 1193 325 1245 341
rect 1193 291 1195 325
rect 1229 309 1245 325
rect 1563 309 1597 356
rect 1791 322 1825 356
rect 1229 291 1597 309
rect 1193 275 1597 291
rect 1633 320 1755 322
rect 1633 286 1705 320
rect 1739 286 1755 320
rect 1633 284 1755 286
rect 1791 320 1958 322
rect 1791 286 1908 320
rect 1942 286 1958 320
rect 1791 284 1958 286
rect 1633 241 1667 284
rect 1992 250 2026 356
rect 1125 223 1667 241
rect 1125 207 1414 223
rect 941 96 951 130
rect 985 96 1001 130
rect 1051 173 1091 207
rect 1168 205 1414 207
rect 1168 178 1220 205
rect 1051 167 1134 173
rect 1051 133 1084 167
rect 1118 133 1134 167
rect 1051 117 1134 133
rect 1168 144 1170 178
rect 1204 144 1220 178
rect 1412 189 1414 205
rect 1448 205 1667 223
rect 1703 216 2026 250
rect 1448 189 1450 205
rect 1168 128 1220 144
rect 1312 165 1378 171
rect 1312 131 1328 165
rect 1362 131 1378 165
rect 941 80 1001 96
rect 1312 17 1378 131
rect 1412 155 1450 189
rect 1703 171 1737 216
rect 2062 182 2096 424
rect 2130 424 2306 426
rect 2130 390 2143 424
rect 2177 390 2256 424
rect 2290 390 2306 424
rect 2130 384 2306 390
rect 2395 350 2430 493
rect 2503 452 2537 581
rect 2132 316 2148 350
rect 2182 316 2430 350
rect 2464 436 2537 452
rect 2571 556 2623 649
rect 2783 599 2850 615
rect 2571 522 2573 556
rect 2607 522 2623 556
rect 2571 486 2623 522
rect 2571 452 2573 486
rect 2607 452 2623 486
rect 2571 436 2623 452
rect 2657 556 2709 572
rect 2657 522 2659 556
rect 2693 522 2709 556
rect 2657 486 2709 522
rect 2657 452 2659 486
rect 2693 452 2709 486
rect 2464 402 2483 436
rect 2517 402 2537 436
rect 2464 368 2559 402
rect 2464 334 2483 368
rect 2517 334 2559 368
rect 2464 318 2559 334
rect 2132 299 2430 316
rect 2275 209 2346 299
rect 1412 121 1414 155
rect 1448 121 1450 155
rect 1484 165 1737 171
rect 1484 131 1500 165
rect 1534 131 1737 165
rect 1484 127 1737 131
rect 1771 166 1811 182
rect 1771 132 1773 166
rect 1807 132 1811 166
rect 1412 105 1450 121
rect 1771 17 1811 132
rect 1915 178 2096 182
rect 1915 144 1931 178
rect 1965 144 2096 178
rect 1915 128 2096 144
rect 2164 176 2230 192
rect 2164 142 2180 176
rect 2214 142 2230 176
rect 2275 175 2303 209
rect 2337 175 2346 209
rect 2275 159 2346 175
rect 2380 200 2491 216
rect 2380 166 2389 200
rect 2423 166 2457 200
rect 2164 17 2230 142
rect 2380 17 2491 166
rect 2525 124 2559 318
rect 2657 366 2709 452
rect 2783 565 2799 599
rect 2833 565 2850 599
rect 2783 506 2850 565
rect 2783 472 2799 506
rect 2833 472 2850 506
rect 2783 413 2850 472
rect 2783 379 2799 413
rect 2833 379 2850 413
rect 2657 350 2733 366
rect 2657 316 2695 350
rect 2729 316 2733 350
rect 2657 282 2733 316
rect 2657 266 2695 282
rect 2593 248 2695 266
rect 2729 248 2733 282
rect 2593 232 2733 248
rect 2783 238 2850 379
rect 2885 611 2923 649
rect 2919 577 2923 611
rect 2885 511 2923 577
rect 2919 477 2923 511
rect 2885 418 2923 477
rect 2919 384 2923 418
rect 2885 368 2923 384
rect 2967 599 3055 615
rect 2967 565 2971 599
rect 3005 565 3055 599
rect 2967 506 3055 565
rect 2967 472 2971 506
rect 3005 472 3055 506
rect 2967 418 3055 472
rect 2967 384 2971 418
rect 3005 384 3055 418
rect 2967 368 3055 384
rect 2593 208 2647 232
rect 2627 174 2647 208
rect 2783 204 2799 238
rect 2833 204 2850 238
rect 2933 318 2967 334
rect 2593 158 2647 174
rect 2933 170 2967 284
rect 2681 168 2967 170
rect 2681 134 2697 168
rect 2731 136 2967 168
rect 3001 234 3055 368
rect 3001 200 3003 234
rect 3037 200 3055 234
rect 2731 134 2747 136
rect 2681 124 2747 134
rect 2525 100 2747 124
rect 3001 126 3055 200
rect 2525 90 2697 100
rect 2681 66 2697 90
rect 2731 66 2747 100
rect 2885 98 2951 102
rect 2885 64 2901 98
rect 2935 64 2951 98
rect 3001 92 3003 126
rect 3037 92 3055 126
rect 3001 76 3055 92
rect 2885 17 2951 64
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 1471 408 1505 424
rect 1471 390 1493 408
rect 1493 390 1505 408
rect 2143 390 2177 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 683 3072 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 0 617 3072 649
rect 1459 424 1517 430
rect 1459 390 1471 424
rect 1505 421 1517 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1505 393 2143 421
rect 1505 390 1517 393
rect 1459 384 1517 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 3072 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
rect 0 -49 3072 -17
<< labels >>
flabel pwell s 0 0 3072 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 3072 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfsbp_1
flabel comment s 1080 312 1080 312 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 2143 390 2177 424 0 FreeSans 200 0 0 0 SET_B
port 5 nsew signal input
flabel metal1 s 0 617 3072 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 3072 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2815 242 2849 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2815 316 2849 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2815 390 2849 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2815 464 2849 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2815 538 2849 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3007 94 3041 128 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3007 168 3041 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3007 242 3041 276 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3007 316 3041 350 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3007 390 3041 424 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3007 464 3041 498 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3007 538 3041 572 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3072 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5572168
string GDS_START 5550242
<< end >>
