magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 1 49 1337 243
rect 0 0 1344 49
<< scnmos >>
rect 80 49 110 217
rect 271 49 301 217
rect 357 49 387 217
rect 443 49 473 217
rect 529 49 559 217
rect 626 49 656 217
rect 712 49 742 217
rect 798 49 828 217
rect 884 49 914 217
rect 970 49 1000 217
rect 1056 49 1086 217
rect 1142 49 1172 217
rect 1228 49 1258 217
<< scpmoshvt >>
rect 91 367 121 619
rect 271 367 301 619
rect 357 367 387 619
rect 443 367 473 619
rect 529 367 559 619
rect 623 367 653 619
rect 709 367 739 619
rect 795 367 825 619
rect 881 367 911 619
rect 967 367 997 619
rect 1053 367 1083 619
rect 1139 367 1169 619
rect 1225 367 1255 619
<< ndiff >>
rect 27 205 80 217
rect 27 171 35 205
rect 69 171 80 205
rect 27 101 80 171
rect 27 67 35 101
rect 69 67 80 101
rect 27 49 80 67
rect 110 181 163 217
rect 110 147 121 181
rect 155 147 163 181
rect 110 95 163 147
rect 110 61 121 95
rect 155 61 163 95
rect 110 49 163 61
rect 218 187 271 217
rect 218 153 226 187
rect 260 153 271 187
rect 218 95 271 153
rect 218 61 226 95
rect 260 61 271 95
rect 218 49 271 61
rect 301 205 357 217
rect 301 171 312 205
rect 346 171 357 205
rect 301 49 357 171
rect 387 103 443 217
rect 387 69 398 103
rect 432 69 443 103
rect 387 49 443 69
rect 473 205 529 217
rect 473 171 484 205
rect 518 171 529 205
rect 473 49 529 171
rect 559 205 626 217
rect 559 171 581 205
rect 615 171 626 205
rect 559 101 626 171
rect 559 67 581 101
rect 615 67 626 101
rect 559 49 626 67
rect 656 177 712 217
rect 656 143 667 177
rect 701 143 712 177
rect 656 91 712 143
rect 656 57 667 91
rect 701 57 712 91
rect 656 49 712 57
rect 742 205 798 217
rect 742 171 753 205
rect 787 171 798 205
rect 742 101 798 171
rect 742 67 753 101
rect 787 67 798 101
rect 742 49 798 67
rect 828 177 884 217
rect 828 143 839 177
rect 873 143 884 177
rect 828 95 884 143
rect 828 61 839 95
rect 873 61 884 95
rect 828 49 884 61
rect 914 205 970 217
rect 914 171 925 205
rect 959 171 970 205
rect 914 101 970 171
rect 914 67 925 101
rect 959 67 970 101
rect 914 49 970 67
rect 1000 169 1056 217
rect 1000 135 1011 169
rect 1045 135 1056 169
rect 1000 95 1056 135
rect 1000 61 1011 95
rect 1045 61 1056 95
rect 1000 49 1056 61
rect 1086 205 1142 217
rect 1086 171 1097 205
rect 1131 171 1142 205
rect 1086 101 1142 171
rect 1086 67 1097 101
rect 1131 67 1142 101
rect 1086 49 1142 67
rect 1172 173 1228 217
rect 1172 139 1183 173
rect 1217 139 1228 173
rect 1172 95 1228 139
rect 1172 61 1183 95
rect 1217 61 1228 95
rect 1172 49 1228 61
rect 1258 205 1311 217
rect 1258 171 1269 205
rect 1303 171 1311 205
rect 1258 101 1311 171
rect 1258 67 1269 101
rect 1303 67 1311 101
rect 1258 49 1311 67
<< pdiff >>
rect 38 599 91 619
rect 38 565 46 599
rect 80 565 91 599
rect 38 517 91 565
rect 38 483 46 517
rect 80 483 91 517
rect 38 436 91 483
rect 38 402 46 436
rect 80 402 91 436
rect 38 367 91 402
rect 121 611 271 619
rect 121 577 132 611
rect 166 607 271 611
rect 166 577 226 607
rect 121 573 226 577
rect 260 573 271 607
rect 121 509 271 573
rect 121 504 226 509
rect 121 470 132 504
rect 166 475 226 504
rect 260 475 271 509
rect 166 470 271 475
rect 121 415 271 470
rect 121 381 226 415
rect 260 381 271 415
rect 121 367 271 381
rect 301 599 357 619
rect 301 565 312 599
rect 346 565 357 599
rect 301 505 357 565
rect 301 471 312 505
rect 346 471 357 505
rect 301 413 357 471
rect 301 379 312 413
rect 346 379 357 413
rect 301 367 357 379
rect 387 607 443 619
rect 387 573 398 607
rect 432 573 443 607
rect 387 533 443 573
rect 387 499 398 533
rect 432 499 443 533
rect 387 455 443 499
rect 387 421 398 455
rect 432 421 443 455
rect 387 367 443 421
rect 473 599 529 619
rect 473 565 484 599
rect 518 565 529 599
rect 473 505 529 565
rect 473 471 484 505
rect 518 471 529 505
rect 473 413 529 471
rect 473 379 484 413
rect 518 379 529 413
rect 473 367 529 379
rect 559 590 623 619
rect 559 556 574 590
rect 608 556 623 590
rect 559 367 623 556
rect 653 596 709 619
rect 653 562 664 596
rect 698 562 709 596
rect 653 367 709 562
rect 739 506 795 619
rect 739 472 750 506
rect 784 472 795 506
rect 739 367 795 472
rect 825 596 881 619
rect 825 562 836 596
rect 870 562 881 596
rect 825 367 881 562
rect 911 506 967 619
rect 911 472 922 506
rect 956 472 967 506
rect 911 367 967 472
rect 997 599 1053 619
rect 997 565 1008 599
rect 1042 565 1053 599
rect 997 491 1053 565
rect 997 457 1008 491
rect 1042 457 1053 491
rect 997 367 1053 457
rect 1083 570 1139 619
rect 1083 536 1094 570
rect 1128 536 1139 570
rect 1083 367 1139 536
rect 1169 599 1225 619
rect 1169 565 1180 599
rect 1214 565 1225 599
rect 1169 513 1225 565
rect 1169 479 1180 513
rect 1214 479 1225 513
rect 1169 436 1225 479
rect 1169 402 1180 436
rect 1214 402 1225 436
rect 1169 367 1225 402
rect 1255 607 1308 619
rect 1255 573 1266 607
rect 1300 573 1308 607
rect 1255 511 1308 573
rect 1255 477 1266 511
rect 1300 477 1308 511
rect 1255 420 1308 477
rect 1255 386 1266 420
rect 1300 386 1308 420
rect 1255 367 1308 386
<< ndiffc >>
rect 35 171 69 205
rect 35 67 69 101
rect 121 147 155 181
rect 121 61 155 95
rect 226 153 260 187
rect 226 61 260 95
rect 312 171 346 205
rect 398 69 432 103
rect 484 171 518 205
rect 581 171 615 205
rect 581 67 615 101
rect 667 143 701 177
rect 667 57 701 91
rect 753 171 787 205
rect 753 67 787 101
rect 839 143 873 177
rect 839 61 873 95
rect 925 171 959 205
rect 925 67 959 101
rect 1011 135 1045 169
rect 1011 61 1045 95
rect 1097 171 1131 205
rect 1097 67 1131 101
rect 1183 139 1217 173
rect 1183 61 1217 95
rect 1269 171 1303 205
rect 1269 67 1303 101
<< pdiffc >>
rect 46 565 80 599
rect 46 483 80 517
rect 46 402 80 436
rect 132 577 166 611
rect 226 573 260 607
rect 132 470 166 504
rect 226 475 260 509
rect 226 381 260 415
rect 312 565 346 599
rect 312 471 346 505
rect 312 379 346 413
rect 398 573 432 607
rect 398 499 432 533
rect 398 421 432 455
rect 484 565 518 599
rect 484 471 518 505
rect 484 379 518 413
rect 574 556 608 590
rect 664 562 698 596
rect 750 472 784 506
rect 836 562 870 596
rect 922 472 956 506
rect 1008 565 1042 599
rect 1008 457 1042 491
rect 1094 536 1128 570
rect 1180 565 1214 599
rect 1180 479 1214 513
rect 1180 402 1214 436
rect 1266 573 1300 607
rect 1266 477 1300 511
rect 1266 386 1300 420
<< poly >>
rect 91 619 121 645
rect 271 619 301 645
rect 357 619 387 645
rect 443 619 473 645
rect 529 619 559 645
rect 623 619 653 645
rect 709 619 739 645
rect 795 619 825 645
rect 881 619 911 645
rect 967 619 997 645
rect 1053 619 1083 645
rect 1139 619 1169 645
rect 1225 619 1255 645
rect 91 335 121 367
rect 271 345 301 367
rect 357 345 387 367
rect 443 345 473 367
rect 529 345 559 367
rect 44 319 121 335
rect 44 285 60 319
rect 94 299 121 319
rect 163 315 559 345
rect 623 335 653 367
rect 709 335 739 367
rect 795 335 825 367
rect 881 335 911 367
rect 967 335 997 367
rect 94 285 110 299
rect 44 269 110 285
rect 80 217 110 269
rect 163 281 179 315
rect 213 281 247 315
rect 281 281 315 315
rect 349 281 383 315
rect 417 281 559 315
rect 163 265 559 281
rect 601 319 667 335
rect 601 285 617 319
rect 651 285 667 319
rect 709 319 997 335
rect 709 305 728 319
rect 601 269 667 285
rect 712 285 728 305
rect 762 285 796 319
rect 830 285 864 319
rect 898 285 932 319
rect 966 299 997 319
rect 1053 325 1083 367
rect 1139 325 1169 367
rect 1225 325 1255 367
rect 1053 309 1323 325
rect 966 285 1000 299
rect 712 269 1000 285
rect 271 217 301 265
rect 357 217 387 265
rect 443 217 473 265
rect 529 217 559 265
rect 626 217 656 269
rect 712 217 742 269
rect 798 217 828 269
rect 884 217 914 269
rect 970 217 1000 269
rect 1053 275 1069 309
rect 1103 275 1137 309
rect 1171 275 1205 309
rect 1239 275 1273 309
rect 1307 275 1323 309
rect 1053 259 1323 275
rect 1056 217 1086 259
rect 1142 217 1172 259
rect 1228 217 1258 259
rect 80 23 110 49
rect 271 23 301 49
rect 357 23 387 49
rect 443 23 473 49
rect 529 23 559 49
rect 626 23 656 49
rect 712 23 742 49
rect 798 23 828 49
rect 884 23 914 49
rect 970 23 1000 49
rect 1056 23 1086 49
rect 1142 23 1172 49
rect 1228 23 1258 49
<< polycont >>
rect 60 285 94 319
rect 179 281 213 315
rect 247 281 281 315
rect 315 281 349 315
rect 383 281 417 315
rect 617 285 651 319
rect 728 285 762 319
rect 796 285 830 319
rect 864 285 898 319
rect 932 285 966 319
rect 1069 275 1103 309
rect 1137 275 1171 309
rect 1205 275 1239 309
rect 1273 275 1307 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 30 599 89 615
rect 30 565 46 599
rect 80 565 89 599
rect 30 517 89 565
rect 30 483 46 517
rect 80 483 89 517
rect 30 436 89 483
rect 123 611 268 649
rect 123 577 132 611
rect 166 607 268 611
rect 166 577 226 607
rect 123 573 226 577
rect 260 573 268 607
rect 123 509 268 573
rect 123 504 226 509
rect 123 470 132 504
rect 166 475 226 504
rect 260 475 268 509
rect 166 470 268 475
rect 123 454 268 470
rect 30 402 46 436
rect 80 420 89 436
rect 80 402 186 420
rect 30 386 186 402
rect 31 319 110 352
rect 31 285 60 319
rect 94 285 110 319
rect 31 283 110 285
rect 152 331 186 386
rect 220 415 268 454
rect 220 381 226 415
rect 260 381 268 415
rect 220 365 268 381
rect 302 599 348 615
rect 302 565 312 599
rect 346 565 348 599
rect 302 505 348 565
rect 302 471 312 505
rect 346 471 348 505
rect 302 413 348 471
rect 382 607 448 649
rect 382 573 398 607
rect 432 573 448 607
rect 382 533 448 573
rect 382 499 398 533
rect 432 499 448 533
rect 382 455 448 499
rect 382 421 398 455
rect 432 421 448 455
rect 482 599 520 615
rect 482 565 484 599
rect 518 565 520 599
rect 482 506 520 565
rect 554 590 614 649
rect 554 556 574 590
rect 608 556 614 590
rect 648 599 1044 615
rect 648 596 1008 599
rect 648 562 664 596
rect 698 562 836 596
rect 870 565 1008 596
rect 1042 565 1044 599
rect 870 562 1044 565
rect 648 558 1044 562
rect 554 540 614 556
rect 648 506 958 522
rect 482 505 750 506
rect 482 471 484 505
rect 518 472 750 505
rect 784 472 922 506
rect 956 472 958 506
rect 518 471 958 472
rect 482 456 958 471
rect 992 492 1044 558
rect 1078 570 1144 649
rect 1078 536 1094 570
rect 1128 536 1144 570
rect 1078 526 1144 536
rect 1178 599 1216 615
rect 1178 565 1180 599
rect 1214 565 1216 599
rect 1178 513 1216 565
rect 1178 492 1180 513
rect 992 491 1180 492
rect 992 457 1008 491
rect 1042 479 1180 491
rect 1214 479 1216 513
rect 1042 457 1216 479
rect 302 379 312 413
rect 346 385 348 413
rect 482 413 545 456
rect 992 454 1216 457
rect 1176 436 1216 454
rect 482 385 484 413
rect 346 379 484 385
rect 518 379 545 413
rect 302 351 545 379
rect 152 317 268 331
rect 152 315 433 317
rect 152 281 179 315
rect 213 281 247 315
rect 281 281 315 315
rect 349 281 383 315
rect 417 281 433 315
rect 152 271 433 281
rect 152 265 276 271
rect 152 249 186 265
rect 19 215 186 249
rect 467 237 545 351
rect 601 386 1087 420
rect 1176 402 1180 436
rect 1214 402 1216 436
rect 1176 386 1216 402
rect 1250 607 1316 649
rect 1250 573 1266 607
rect 1300 573 1316 607
rect 1250 511 1316 573
rect 1250 477 1266 511
rect 1300 477 1316 511
rect 1250 420 1316 477
rect 1250 386 1266 420
rect 1300 386 1316 420
rect 601 319 667 386
rect 1053 352 1087 386
rect 601 285 617 319
rect 651 285 667 319
rect 703 319 982 350
rect 703 285 728 319
rect 762 285 796 319
rect 830 285 864 319
rect 898 285 932 319
rect 966 285 982 319
rect 1053 309 1323 352
rect 1053 275 1069 309
rect 1103 275 1137 309
rect 1171 275 1205 309
rect 1239 275 1273 309
rect 1307 275 1323 309
rect 19 205 71 215
rect 19 171 35 205
rect 69 171 71 205
rect 310 205 545 237
rect 210 187 276 189
rect 19 101 71 171
rect 19 67 35 101
rect 69 67 71 101
rect 19 51 71 67
rect 105 147 121 181
rect 155 147 171 181
rect 105 95 171 147
rect 105 61 121 95
rect 155 61 171 95
rect 105 17 171 61
rect 210 153 226 187
rect 260 153 276 187
rect 310 171 312 205
rect 346 171 484 205
rect 518 171 545 205
rect 310 155 545 171
rect 579 241 959 245
rect 579 211 1319 241
rect 579 205 617 211
rect 579 171 581 205
rect 615 171 617 205
rect 751 205 789 211
rect 210 119 276 153
rect 579 119 617 171
rect 210 103 617 119
rect 210 95 398 103
rect 210 61 226 95
rect 260 69 398 95
rect 432 101 617 103
rect 432 69 581 101
rect 260 67 581 69
rect 615 67 617 101
rect 260 61 617 67
rect 210 51 617 61
rect 651 143 667 177
rect 701 143 717 177
rect 651 91 717 143
rect 651 57 667 91
rect 701 57 717 91
rect 651 17 717 57
rect 751 171 753 205
rect 787 171 789 205
rect 923 207 1319 211
rect 923 205 1133 207
rect 751 101 789 171
rect 751 67 753 101
rect 787 67 789 101
rect 751 51 789 67
rect 823 143 839 177
rect 873 143 889 177
rect 823 95 889 143
rect 823 61 839 95
rect 873 61 889 95
rect 823 17 889 61
rect 923 171 925 205
rect 959 203 1097 205
rect 959 171 961 203
rect 923 101 961 171
rect 1095 171 1097 203
rect 1131 171 1133 205
rect 1267 205 1319 207
rect 923 67 925 101
rect 959 67 961 101
rect 923 51 961 67
rect 995 135 1011 169
rect 1045 135 1061 169
rect 995 95 1061 135
rect 995 61 1011 95
rect 1045 61 1061 95
rect 995 17 1061 61
rect 1095 101 1133 171
rect 1095 67 1097 101
rect 1131 67 1133 101
rect 1095 51 1133 67
rect 1167 139 1183 173
rect 1217 139 1233 173
rect 1167 95 1233 139
rect 1167 61 1183 95
rect 1217 61 1233 95
rect 1167 17 1233 61
rect 1267 171 1269 205
rect 1303 171 1319 205
rect 1267 101 1319 171
rect 1267 67 1269 101
rect 1303 67 1319 101
rect 1267 51 1319 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21bai_4
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5174282
string GDS_START 5162718
<< end >>
