magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 6 49 1088 241
rect 0 0 1152 49
<< scnmos >>
rect 85 47 115 215
rect 171 47 201 215
rect 257 47 287 215
rect 365 47 395 215
rect 460 47 490 215
rect 568 47 598 215
rect 654 47 684 215
rect 794 47 824 215
rect 893 47 923 215
rect 979 47 1009 215
<< scpmoshvt >>
rect 85 367 115 619
rect 171 367 201 619
rect 257 367 287 619
rect 343 367 373 619
rect 437 367 467 619
rect 523 367 553 619
rect 713 367 743 619
rect 799 367 829 619
rect 885 367 915 619
rect 979 367 1009 619
<< ndiff >>
rect 32 192 85 215
rect 32 158 40 192
rect 74 158 85 192
rect 32 103 85 158
rect 32 69 40 103
rect 74 69 85 103
rect 32 47 85 69
rect 115 132 171 215
rect 115 98 126 132
rect 160 98 171 132
rect 115 47 171 98
rect 201 192 257 215
rect 201 158 212 192
rect 246 158 257 192
rect 201 103 257 158
rect 201 69 212 103
rect 246 69 257 103
rect 201 47 257 69
rect 287 132 365 215
rect 287 98 309 132
rect 343 98 365 132
rect 287 47 365 98
rect 395 203 460 215
rect 395 169 412 203
rect 446 169 460 203
rect 395 101 460 169
rect 395 67 412 101
rect 446 67 460 101
rect 395 47 460 67
rect 490 183 568 215
rect 490 149 509 183
rect 543 149 568 183
rect 490 93 568 149
rect 490 59 509 93
rect 543 59 568 93
rect 490 47 568 59
rect 598 203 654 215
rect 598 169 609 203
rect 643 169 654 203
rect 598 92 654 169
rect 598 58 609 92
rect 643 58 654 92
rect 598 47 654 58
rect 684 203 794 215
rect 684 169 722 203
rect 756 169 794 203
rect 684 92 794 169
rect 684 58 722 92
rect 756 58 794 92
rect 684 47 794 58
rect 824 132 893 215
rect 824 98 841 132
rect 875 98 893 132
rect 824 47 893 98
rect 923 192 979 215
rect 923 158 934 192
rect 968 158 979 192
rect 923 101 979 158
rect 923 67 934 101
rect 968 67 979 101
rect 923 47 979 67
rect 1009 203 1062 215
rect 1009 169 1020 203
rect 1054 169 1062 203
rect 1009 101 1062 169
rect 1009 67 1020 101
rect 1054 67 1062 101
rect 1009 47 1062 67
<< pdiff >>
rect 32 599 85 619
rect 32 565 40 599
rect 74 565 85 599
rect 32 523 85 565
rect 32 489 40 523
rect 74 489 85 523
rect 32 441 85 489
rect 32 407 40 441
rect 74 407 85 441
rect 32 367 85 407
rect 115 523 171 619
rect 115 489 126 523
rect 160 489 171 523
rect 115 441 171 489
rect 115 407 126 441
rect 160 407 171 441
rect 115 367 171 407
rect 201 455 257 619
rect 201 421 212 455
rect 246 421 257 455
rect 201 367 257 421
rect 287 509 343 619
rect 287 475 298 509
rect 332 475 343 509
rect 287 367 343 475
rect 373 599 437 619
rect 373 565 384 599
rect 418 565 437 599
rect 373 509 437 565
rect 373 475 384 509
rect 418 475 437 509
rect 373 367 437 475
rect 467 513 523 619
rect 467 479 478 513
rect 512 479 523 513
rect 467 367 523 479
rect 553 603 606 619
rect 553 569 564 603
rect 598 569 606 603
rect 553 367 606 569
rect 660 599 713 619
rect 660 565 668 599
rect 702 565 713 599
rect 660 493 713 565
rect 660 459 668 493
rect 702 459 713 493
rect 660 367 713 459
rect 743 569 799 619
rect 743 535 754 569
rect 788 535 799 569
rect 743 367 799 535
rect 829 599 885 619
rect 829 565 840 599
rect 874 565 885 599
rect 829 493 885 565
rect 829 459 840 493
rect 874 459 885 493
rect 829 367 885 459
rect 915 569 979 619
rect 915 535 930 569
rect 964 535 979 569
rect 915 367 979 535
rect 1009 599 1062 619
rect 1009 565 1020 599
rect 1054 565 1062 599
rect 1009 493 1062 565
rect 1009 459 1020 493
rect 1054 459 1062 493
rect 1009 367 1062 459
<< ndiffc >>
rect 40 158 74 192
rect 40 69 74 103
rect 126 98 160 132
rect 212 158 246 192
rect 212 69 246 103
rect 309 98 343 132
rect 412 169 446 203
rect 412 67 446 101
rect 509 149 543 183
rect 509 59 543 93
rect 609 169 643 203
rect 609 58 643 92
rect 722 169 756 203
rect 722 58 756 92
rect 841 98 875 132
rect 934 158 968 192
rect 934 67 968 101
rect 1020 169 1054 203
rect 1020 67 1054 101
<< pdiffc >>
rect 40 565 74 599
rect 40 489 74 523
rect 40 407 74 441
rect 126 489 160 523
rect 126 407 160 441
rect 212 421 246 455
rect 298 475 332 509
rect 384 565 418 599
rect 384 475 418 509
rect 478 479 512 513
rect 564 569 598 603
rect 668 565 702 599
rect 668 459 702 493
rect 754 535 788 569
rect 840 565 874 599
rect 840 459 874 493
rect 930 535 964 569
rect 1020 565 1054 599
rect 1020 459 1054 493
<< poly >>
rect 85 619 115 645
rect 171 619 201 645
rect 257 619 287 645
rect 343 619 373 645
rect 437 619 467 645
rect 523 619 553 645
rect 713 619 743 645
rect 799 619 829 645
rect 885 619 915 645
rect 979 619 1009 645
rect 85 325 115 367
rect 25 309 115 325
rect 25 275 41 309
rect 75 275 115 309
rect 25 259 115 275
rect 85 215 115 259
rect 171 303 201 367
rect 257 303 287 367
rect 343 325 373 367
rect 437 335 467 367
rect 523 335 553 367
rect 713 335 743 367
rect 171 287 287 303
rect 171 253 187 287
rect 221 253 287 287
rect 329 309 395 325
rect 329 275 345 309
rect 379 275 395 309
rect 329 259 395 275
rect 437 319 598 335
rect 437 285 453 319
rect 487 285 521 319
rect 555 285 598 319
rect 437 269 598 285
rect 171 237 287 253
rect 171 215 201 237
rect 257 215 287 237
rect 365 215 395 259
rect 460 215 490 269
rect 568 215 598 269
rect 654 319 743 335
rect 654 285 693 319
rect 727 285 743 319
rect 654 269 743 285
rect 654 215 684 269
rect 799 267 829 367
rect 885 303 915 367
rect 979 335 1009 367
rect 979 319 1045 335
rect 871 287 937 303
rect 871 267 887 287
rect 794 253 887 267
rect 921 253 937 287
rect 794 237 937 253
rect 979 285 995 319
rect 1029 285 1045 319
rect 979 269 1045 285
rect 794 215 824 237
rect 893 215 923 237
rect 979 215 1009 269
rect 85 21 115 47
rect 171 21 201 47
rect 257 21 287 47
rect 365 21 395 47
rect 460 21 490 47
rect 568 21 598 47
rect 654 21 684 47
rect 794 21 824 47
rect 893 21 923 47
rect 979 21 1009 47
<< polycont >>
rect 41 275 75 309
rect 187 253 221 287
rect 345 275 379 309
rect 453 285 487 319
rect 521 285 555 319
rect 693 285 727 319
rect 887 253 921 287
rect 995 285 1029 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 24 603 614 615
rect 24 599 564 603
rect 24 565 40 599
rect 74 573 384 599
rect 74 565 80 573
rect 24 523 80 565
rect 374 565 384 573
rect 418 569 564 599
rect 598 569 614 603
rect 418 565 614 569
rect 374 563 614 565
rect 652 599 704 615
rect 652 565 668 599
rect 702 565 704 599
rect 24 489 40 523
rect 74 489 80 523
rect 24 441 80 489
rect 24 407 40 441
rect 74 407 80 441
rect 24 391 80 407
rect 114 523 340 539
rect 114 489 126 523
rect 160 509 340 523
rect 160 505 298 509
rect 160 489 166 505
rect 114 441 166 489
rect 290 475 298 505
rect 332 475 340 509
rect 114 407 126 441
rect 160 407 166 441
rect 114 391 166 407
rect 200 455 253 471
rect 290 459 340 475
rect 374 509 433 563
rect 652 529 704 565
rect 374 475 384 509
rect 418 475 433 509
rect 374 459 433 475
rect 467 513 704 529
rect 738 569 804 649
rect 738 535 754 569
rect 788 535 804 569
rect 738 527 804 535
rect 838 599 880 615
rect 838 565 840 599
rect 874 565 880 599
rect 467 479 478 513
rect 512 493 704 513
rect 838 493 880 565
rect 914 569 980 649
rect 914 535 930 569
rect 964 535 980 569
rect 914 527 980 535
rect 1014 599 1070 615
rect 1014 565 1020 599
rect 1054 565 1070 599
rect 1014 493 1070 565
rect 512 479 668 493
rect 467 459 668 479
rect 702 459 840 493
rect 874 459 1020 493
rect 1054 459 1070 493
rect 200 421 212 455
rect 246 425 253 455
rect 246 421 1132 425
rect 200 391 1132 421
rect 200 389 659 391
rect 25 321 379 355
rect 25 309 91 321
rect 25 275 41 309
rect 75 275 91 309
rect 305 309 379 321
rect 25 259 91 275
rect 125 253 187 287
rect 221 253 271 287
rect 305 275 345 309
rect 413 319 571 355
rect 413 285 453 319
rect 487 285 521 319
rect 555 285 571 319
rect 305 259 379 275
rect 125 242 271 253
rect 605 251 659 389
rect 693 323 1031 357
rect 693 319 837 323
rect 727 285 837 319
rect 979 319 1031 323
rect 693 269 837 285
rect 413 217 659 251
rect 871 253 887 287
rect 921 253 945 287
rect 979 285 995 319
rect 1029 285 1031 319
rect 979 269 1031 285
rect 871 242 945 253
rect 1065 219 1132 391
rect 413 208 459 217
rect 24 203 459 208
rect 24 192 412 203
rect 24 158 40 192
rect 74 174 212 192
rect 74 158 76 174
rect 24 103 76 158
rect 210 158 212 174
rect 246 174 412 192
rect 246 158 259 174
rect 24 69 40 103
rect 74 69 76 103
rect 24 51 76 69
rect 110 132 176 140
rect 110 98 126 132
rect 160 98 176 132
rect 110 17 176 98
rect 210 103 259 158
rect 393 169 412 174
rect 446 169 459 203
rect 593 203 659 217
rect 210 69 212 103
rect 246 69 259 103
rect 210 53 259 69
rect 293 132 359 140
rect 293 98 309 132
rect 343 98 359 132
rect 293 17 359 98
rect 393 101 459 169
rect 393 67 412 101
rect 446 67 459 101
rect 393 51 459 67
rect 493 149 509 183
rect 543 149 559 183
rect 493 93 559 149
rect 493 59 509 93
rect 543 59 559 93
rect 493 17 559 59
rect 593 169 609 203
rect 643 169 659 203
rect 593 92 659 169
rect 593 58 609 92
rect 643 58 659 92
rect 593 51 659 58
rect 706 203 970 208
rect 706 169 722 203
rect 756 192 970 203
rect 756 174 934 192
rect 756 169 772 174
rect 706 92 772 169
rect 925 158 934 174
rect 968 158 970 192
rect 706 58 722 92
rect 756 58 772 92
rect 706 51 772 58
rect 825 132 891 140
rect 825 98 841 132
rect 875 98 891 132
rect 825 17 891 98
rect 925 101 970 158
rect 925 67 934 101
rect 968 67 970 101
rect 925 51 970 67
rect 1004 203 1132 219
rect 1004 169 1020 203
rect 1054 169 1132 203
rect 1004 101 1132 169
rect 1004 67 1020 101
rect 1054 67 1132 101
rect 1004 51 1132 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2111oi_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4793088
string GDS_START 4783382
<< end >>
