magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
rect 518 325 1328 331
<< pwell >>
rect 166 49 2096 241
rect 0 0 2112 49
<< scnmos >>
rect 245 47 275 215
rect 331 47 361 215
rect 417 47 447 215
rect 503 47 533 215
rect 605 47 635 215
rect 707 47 737 215
rect 793 47 823 215
rect 897 47 927 215
rect 997 47 1027 215
rect 1099 47 1129 215
rect 1185 47 1215 215
rect 1271 47 1301 215
rect 1357 47 1387 215
rect 1443 47 1473 215
rect 1529 47 1559 215
rect 1642 47 1672 215
rect 1729 47 1759 215
rect 1815 47 1845 215
rect 1901 47 1931 215
rect 1987 47 2017 215
<< scpmoshvt >>
rect 159 367 189 619
rect 245 367 275 619
rect 331 367 361 619
rect 417 367 447 619
rect 607 361 637 613
rect 693 361 723 613
rect 779 361 809 613
rect 865 361 895 613
rect 951 361 981 613
rect 1037 361 1067 613
rect 1123 361 1153 613
rect 1209 361 1239 613
rect 1399 367 1429 619
rect 1485 367 1515 619
rect 1571 367 1601 619
rect 1657 367 1687 619
rect 1743 367 1773 619
rect 1829 367 1859 619
rect 1915 367 1945 619
rect 2001 367 2031 619
<< ndiff >>
rect 192 203 245 215
rect 192 169 200 203
rect 234 169 245 203
rect 192 105 245 169
rect 192 71 200 105
rect 234 71 245 105
rect 192 47 245 71
rect 275 169 331 215
rect 275 135 286 169
rect 320 135 331 169
rect 275 47 331 135
rect 361 167 417 215
rect 361 133 372 167
rect 406 133 417 167
rect 361 93 417 133
rect 361 59 372 93
rect 406 59 417 93
rect 361 47 417 59
rect 447 169 503 215
rect 447 135 458 169
rect 492 135 503 169
rect 447 47 503 135
rect 533 167 605 215
rect 533 133 544 167
rect 578 133 605 167
rect 533 93 605 133
rect 533 59 544 93
rect 578 59 605 93
rect 533 47 605 59
rect 635 93 707 215
rect 635 59 646 93
rect 680 59 707 93
rect 635 47 707 59
rect 737 167 793 215
rect 737 133 748 167
rect 782 133 793 167
rect 737 93 793 133
rect 737 59 748 93
rect 782 59 793 93
rect 737 47 793 59
rect 823 93 897 215
rect 823 59 850 93
rect 884 59 897 93
rect 823 47 897 59
rect 927 167 997 215
rect 927 133 952 167
rect 986 133 997 167
rect 927 93 997 133
rect 927 59 952 93
rect 986 59 997 93
rect 927 47 997 59
rect 1027 161 1099 215
rect 1027 127 1053 161
rect 1087 127 1099 161
rect 1027 93 1099 127
rect 1027 59 1053 93
rect 1087 59 1099 93
rect 1027 47 1099 59
rect 1129 203 1185 215
rect 1129 169 1140 203
rect 1174 169 1185 203
rect 1129 101 1185 169
rect 1129 67 1140 101
rect 1174 67 1185 101
rect 1129 47 1185 67
rect 1215 167 1271 215
rect 1215 133 1226 167
rect 1260 133 1271 167
rect 1215 93 1271 133
rect 1215 59 1226 93
rect 1260 59 1271 93
rect 1215 47 1271 59
rect 1301 203 1357 215
rect 1301 169 1312 203
rect 1346 169 1357 203
rect 1301 101 1357 169
rect 1301 67 1312 101
rect 1346 67 1357 101
rect 1301 47 1357 67
rect 1387 167 1443 215
rect 1387 133 1398 167
rect 1432 133 1443 167
rect 1387 93 1443 133
rect 1387 59 1398 93
rect 1432 59 1443 93
rect 1387 47 1443 59
rect 1473 203 1529 215
rect 1473 169 1484 203
rect 1518 169 1529 203
rect 1473 101 1529 169
rect 1473 67 1484 101
rect 1518 67 1529 101
rect 1473 47 1529 67
rect 1559 167 1642 215
rect 1559 133 1584 167
rect 1618 133 1642 167
rect 1559 93 1642 133
rect 1559 59 1584 93
rect 1618 59 1642 93
rect 1559 47 1642 59
rect 1672 203 1729 215
rect 1672 169 1683 203
rect 1717 169 1729 203
rect 1672 101 1729 169
rect 1672 67 1683 101
rect 1717 67 1729 101
rect 1672 47 1729 67
rect 1759 124 1815 215
rect 1759 90 1770 124
rect 1804 90 1815 124
rect 1759 47 1815 90
rect 1845 192 1901 215
rect 1845 158 1856 192
rect 1890 158 1901 192
rect 1845 101 1901 158
rect 1845 67 1856 101
rect 1890 67 1901 101
rect 1845 47 1901 67
rect 1931 124 1987 215
rect 1931 90 1942 124
rect 1976 90 1987 124
rect 1931 47 1987 90
rect 2017 192 2070 215
rect 2017 158 2028 192
rect 2062 158 2070 192
rect 2017 101 2070 158
rect 2017 67 2028 101
rect 2062 67 2070 101
rect 2017 47 2070 67
<< pdiff >>
rect 106 607 159 619
rect 106 573 114 607
rect 148 573 159 607
rect 106 510 159 573
rect 106 476 114 510
rect 148 476 159 510
rect 106 420 159 476
rect 106 386 114 420
rect 148 386 159 420
rect 106 367 159 386
rect 189 599 245 619
rect 189 565 200 599
rect 234 565 245 599
rect 189 523 245 565
rect 189 489 200 523
rect 234 489 245 523
rect 189 436 245 489
rect 189 402 200 436
rect 234 402 245 436
rect 189 367 245 402
rect 275 607 331 619
rect 275 573 286 607
rect 320 573 331 607
rect 275 496 331 573
rect 275 462 286 496
rect 320 462 331 496
rect 275 367 331 462
rect 361 599 417 619
rect 361 565 372 599
rect 406 565 417 599
rect 361 517 417 565
rect 361 483 372 517
rect 406 483 417 517
rect 361 420 417 483
rect 361 386 372 420
rect 406 386 417 420
rect 361 367 417 386
rect 447 607 500 619
rect 447 573 458 607
rect 492 573 500 607
rect 447 496 500 573
rect 447 462 458 496
rect 492 462 500 496
rect 447 367 500 462
rect 554 599 607 613
rect 554 565 562 599
rect 596 565 607 599
rect 554 504 607 565
rect 554 470 562 504
rect 596 470 607 504
rect 554 361 607 470
rect 637 539 693 613
rect 637 505 648 539
rect 682 505 693 539
rect 637 426 693 505
rect 637 392 648 426
rect 682 392 693 426
rect 637 361 693 392
rect 723 599 779 613
rect 723 565 734 599
rect 768 565 779 599
rect 723 504 779 565
rect 723 470 734 504
rect 768 470 779 504
rect 723 361 779 470
rect 809 545 865 613
rect 809 511 820 545
rect 854 511 865 545
rect 809 471 865 511
rect 809 437 820 471
rect 854 437 865 471
rect 809 403 865 437
rect 809 369 820 403
rect 854 369 865 403
rect 809 361 865 369
rect 895 599 951 613
rect 895 565 906 599
rect 940 565 951 599
rect 895 529 951 565
rect 895 495 906 529
rect 940 495 951 529
rect 895 459 951 495
rect 895 425 906 459
rect 940 425 951 459
rect 895 361 951 425
rect 981 605 1037 613
rect 981 571 992 605
rect 1026 571 1037 605
rect 981 513 1037 571
rect 981 479 992 513
rect 1026 479 1037 513
rect 981 361 1037 479
rect 1067 521 1123 613
rect 1067 487 1078 521
rect 1112 487 1123 521
rect 1067 434 1123 487
rect 1067 400 1078 434
rect 1112 400 1123 434
rect 1067 361 1123 400
rect 1153 605 1209 613
rect 1153 571 1164 605
rect 1198 571 1209 605
rect 1153 513 1209 571
rect 1153 479 1164 513
rect 1198 479 1209 513
rect 1153 361 1209 479
rect 1239 521 1292 613
rect 1239 487 1250 521
rect 1284 487 1292 521
rect 1239 418 1292 487
rect 1239 384 1250 418
rect 1284 384 1292 418
rect 1239 361 1292 384
rect 1346 521 1399 619
rect 1346 487 1354 521
rect 1388 487 1399 521
rect 1346 418 1399 487
rect 1346 384 1354 418
rect 1388 384 1399 418
rect 1346 367 1399 384
rect 1429 597 1485 619
rect 1429 563 1440 597
rect 1474 563 1485 597
rect 1429 488 1485 563
rect 1429 454 1440 488
rect 1474 454 1485 488
rect 1429 367 1485 454
rect 1515 482 1571 619
rect 1515 448 1526 482
rect 1560 448 1571 482
rect 1515 413 1571 448
rect 1515 379 1526 413
rect 1560 379 1571 413
rect 1515 367 1571 379
rect 1601 599 1657 619
rect 1601 565 1612 599
rect 1646 565 1657 599
rect 1601 529 1657 565
rect 1601 495 1612 529
rect 1646 495 1657 529
rect 1601 459 1657 495
rect 1601 425 1612 459
rect 1646 425 1657 459
rect 1601 367 1657 425
rect 1687 599 1743 619
rect 1687 565 1698 599
rect 1732 565 1743 599
rect 1687 511 1743 565
rect 1687 477 1698 511
rect 1732 477 1743 511
rect 1687 413 1743 477
rect 1687 379 1698 413
rect 1732 379 1743 413
rect 1687 367 1743 379
rect 1773 607 1829 619
rect 1773 573 1784 607
rect 1818 573 1829 607
rect 1773 526 1829 573
rect 1773 492 1784 526
rect 1818 492 1829 526
rect 1773 443 1829 492
rect 1773 409 1784 443
rect 1818 409 1829 443
rect 1773 367 1829 409
rect 1859 599 1915 619
rect 1859 565 1870 599
rect 1904 565 1915 599
rect 1859 511 1915 565
rect 1859 477 1870 511
rect 1904 477 1915 511
rect 1859 413 1915 477
rect 1859 379 1870 413
rect 1904 379 1915 413
rect 1859 367 1915 379
rect 1945 607 2001 619
rect 1945 573 1956 607
rect 1990 573 2001 607
rect 1945 526 2001 573
rect 1945 492 1956 526
rect 1990 492 2001 526
rect 1945 443 2001 492
rect 1945 409 1956 443
rect 1990 409 2001 443
rect 1945 367 2001 409
rect 2031 599 2084 619
rect 2031 565 2042 599
rect 2076 565 2084 599
rect 2031 511 2084 565
rect 2031 477 2042 511
rect 2076 477 2084 511
rect 2031 413 2084 477
rect 2031 379 2042 413
rect 2076 379 2084 413
rect 2031 367 2084 379
<< ndiffc >>
rect 200 169 234 203
rect 200 71 234 105
rect 286 135 320 169
rect 372 133 406 167
rect 372 59 406 93
rect 458 135 492 169
rect 544 133 578 167
rect 544 59 578 93
rect 646 59 680 93
rect 748 133 782 167
rect 748 59 782 93
rect 850 59 884 93
rect 952 133 986 167
rect 952 59 986 93
rect 1053 127 1087 161
rect 1053 59 1087 93
rect 1140 169 1174 203
rect 1140 67 1174 101
rect 1226 133 1260 167
rect 1226 59 1260 93
rect 1312 169 1346 203
rect 1312 67 1346 101
rect 1398 133 1432 167
rect 1398 59 1432 93
rect 1484 169 1518 203
rect 1484 67 1518 101
rect 1584 133 1618 167
rect 1584 59 1618 93
rect 1683 169 1717 203
rect 1683 67 1717 101
rect 1770 90 1804 124
rect 1856 158 1890 192
rect 1856 67 1890 101
rect 1942 90 1976 124
rect 2028 158 2062 192
rect 2028 67 2062 101
<< pdiffc >>
rect 114 573 148 607
rect 114 476 148 510
rect 114 386 148 420
rect 200 565 234 599
rect 200 489 234 523
rect 200 402 234 436
rect 286 573 320 607
rect 286 462 320 496
rect 372 565 406 599
rect 372 483 406 517
rect 372 386 406 420
rect 458 573 492 607
rect 458 462 492 496
rect 562 565 596 599
rect 562 470 596 504
rect 648 505 682 539
rect 648 392 682 426
rect 734 565 768 599
rect 734 470 768 504
rect 820 511 854 545
rect 820 437 854 471
rect 820 369 854 403
rect 906 565 940 599
rect 906 495 940 529
rect 906 425 940 459
rect 992 571 1026 605
rect 992 479 1026 513
rect 1078 487 1112 521
rect 1078 400 1112 434
rect 1164 571 1198 605
rect 1164 479 1198 513
rect 1250 487 1284 521
rect 1250 384 1284 418
rect 1354 487 1388 521
rect 1354 384 1388 418
rect 1440 563 1474 597
rect 1440 454 1474 488
rect 1526 448 1560 482
rect 1526 379 1560 413
rect 1612 565 1646 599
rect 1612 495 1646 529
rect 1612 425 1646 459
rect 1698 565 1732 599
rect 1698 477 1732 511
rect 1698 379 1732 413
rect 1784 573 1818 607
rect 1784 492 1818 526
rect 1784 409 1818 443
rect 1870 565 1904 599
rect 1870 477 1904 511
rect 1870 379 1904 413
rect 1956 573 1990 607
rect 1956 492 1990 526
rect 1956 409 1990 443
rect 2042 565 2076 599
rect 2042 477 2076 511
rect 2042 379 2076 413
<< poly >>
rect 159 619 189 645
rect 245 619 275 645
rect 331 619 361 645
rect 417 619 447 645
rect 607 613 637 639
rect 693 613 723 639
rect 779 613 809 639
rect 865 613 895 639
rect 951 613 981 639
rect 1037 613 1067 639
rect 1123 613 1153 639
rect 1209 613 1239 639
rect 1399 619 1429 645
rect 1485 619 1515 645
rect 1571 619 1601 645
rect 1657 619 1687 645
rect 1743 619 1773 645
rect 1829 619 1859 645
rect 1915 619 1945 645
rect 2001 619 2031 645
rect 159 325 189 367
rect 245 325 275 367
rect 331 325 361 367
rect 417 325 447 367
rect 21 309 563 325
rect 607 321 637 361
rect 693 321 723 361
rect 779 321 809 361
rect 865 321 895 361
rect 21 275 37 309
rect 71 275 105 309
rect 139 275 173 309
rect 207 275 241 309
rect 275 275 309 309
rect 343 275 377 309
rect 411 275 445 309
rect 479 275 513 309
rect 547 275 563 309
rect 21 259 563 275
rect 605 305 895 321
rect 951 339 981 361
rect 1037 339 1067 361
rect 1123 339 1153 361
rect 1209 339 1239 361
rect 951 313 1307 339
rect 1399 321 1429 367
rect 1485 321 1515 367
rect 1571 321 1601 367
rect 1657 321 1687 367
rect 951 309 985 313
rect 605 271 623 305
rect 657 271 712 305
rect 746 271 801 305
rect 835 271 895 305
rect 605 267 895 271
rect 969 279 985 309
rect 1019 279 1053 313
rect 1087 279 1121 313
rect 1155 279 1189 313
rect 1223 279 1257 313
rect 1291 279 1307 313
rect 245 215 275 259
rect 331 215 361 259
rect 417 215 447 259
rect 503 215 533 259
rect 605 237 927 267
rect 969 263 1307 279
rect 1349 305 1687 321
rect 1349 271 1365 305
rect 1399 271 1433 305
rect 1467 271 1501 305
rect 1535 271 1569 305
rect 1603 271 1637 305
rect 1671 271 1687 305
rect 1743 303 1773 367
rect 1829 303 1859 367
rect 1915 303 1945 367
rect 2001 303 2031 367
rect 605 215 635 237
rect 707 215 737 237
rect 793 215 823 237
rect 897 215 927 237
rect 997 215 1027 263
rect 1099 215 1129 263
rect 1185 215 1215 263
rect 1271 215 1301 263
rect 1349 255 1687 271
rect 1729 287 2091 303
rect 1357 215 1387 255
rect 1443 215 1473 255
rect 1529 215 1559 255
rect 1642 215 1672 255
rect 1729 253 1769 287
rect 1803 253 1837 287
rect 1871 253 1905 287
rect 1939 253 1973 287
rect 2007 253 2041 287
rect 2075 253 2091 287
rect 1729 237 2091 253
rect 1729 215 1759 237
rect 1815 215 1845 237
rect 1901 215 1931 237
rect 1987 215 2017 237
rect 245 21 275 47
rect 331 21 361 47
rect 417 21 447 47
rect 503 21 533 47
rect 605 21 635 47
rect 707 21 737 47
rect 793 21 823 47
rect 897 21 927 47
rect 997 21 1027 47
rect 1099 21 1129 47
rect 1185 21 1215 47
rect 1271 21 1301 47
rect 1357 21 1387 47
rect 1443 21 1473 47
rect 1529 21 1559 47
rect 1642 21 1672 47
rect 1729 21 1759 47
rect 1815 21 1845 47
rect 1901 21 1931 47
rect 1987 21 2017 47
<< polycont >>
rect 37 275 71 309
rect 105 275 139 309
rect 173 275 207 309
rect 241 275 275 309
rect 309 275 343 309
rect 377 275 411 309
rect 445 275 479 309
rect 513 275 547 309
rect 623 271 657 305
rect 712 271 746 305
rect 801 271 835 305
rect 985 279 1019 313
rect 1053 279 1087 313
rect 1121 279 1155 313
rect 1189 279 1223 313
rect 1257 279 1291 313
rect 1365 271 1399 305
rect 1433 271 1467 305
rect 1501 271 1535 305
rect 1569 271 1603 305
rect 1637 271 1671 305
rect 1769 253 1803 287
rect 1837 253 1871 287
rect 1905 253 1939 287
rect 1973 253 2007 287
rect 2041 253 2075 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 98 607 164 649
rect 98 573 114 607
rect 148 573 164 607
rect 98 510 164 573
rect 98 476 114 510
rect 148 476 164 510
rect 98 420 164 476
rect 98 386 114 420
rect 148 386 164 420
rect 198 599 236 615
rect 198 565 200 599
rect 234 565 236 599
rect 198 523 236 565
rect 198 489 200 523
rect 234 489 236 523
rect 198 436 236 489
rect 270 607 336 649
rect 270 573 286 607
rect 320 573 336 607
rect 270 496 336 573
rect 270 462 286 496
rect 320 462 336 496
rect 270 454 336 462
rect 372 599 408 615
rect 406 565 408 599
rect 372 517 408 565
rect 406 483 408 517
rect 198 402 200 436
rect 234 420 236 436
rect 372 420 408 483
rect 442 607 508 649
rect 442 573 458 607
rect 492 573 508 607
rect 442 496 508 573
rect 442 462 458 496
rect 492 462 508 496
rect 442 454 508 462
rect 546 599 942 615
rect 546 565 562 599
rect 596 579 734 599
rect 596 565 598 579
rect 546 504 598 565
rect 732 565 734 579
rect 768 579 906 599
rect 768 565 770 579
rect 546 470 562 504
rect 596 470 598 504
rect 546 454 598 470
rect 632 539 698 545
rect 632 505 648 539
rect 682 505 698 539
rect 632 426 698 505
rect 732 504 770 565
rect 904 565 906 579
rect 940 565 942 599
rect 732 470 734 504
rect 768 470 770 504
rect 732 454 770 470
rect 804 511 820 545
rect 854 511 870 545
rect 804 471 870 511
rect 632 420 648 426
rect 234 402 372 420
rect 198 386 372 402
rect 406 392 648 420
rect 682 420 698 426
rect 804 437 820 471
rect 854 437 870 471
rect 804 420 870 437
rect 682 403 870 420
rect 904 529 942 565
rect 904 495 906 529
rect 940 495 942 529
rect 904 459 942 495
rect 976 605 1662 615
rect 976 571 992 605
rect 1026 571 1164 605
rect 1198 599 1662 605
rect 1198 597 1612 599
rect 1198 571 1440 597
rect 976 513 1042 571
rect 976 479 992 513
rect 1026 479 1042 513
rect 1076 521 1114 537
rect 1076 487 1078 521
rect 1112 487 1114 521
rect 904 425 906 459
rect 940 445 942 459
rect 1076 445 1114 487
rect 1148 513 1214 571
rect 1424 563 1440 571
rect 1474 565 1612 597
rect 1646 565 1662 599
rect 1474 563 1662 565
rect 1424 547 1662 563
rect 1148 479 1164 513
rect 1198 479 1214 513
rect 1248 521 1300 537
rect 1248 487 1250 521
rect 1284 487 1300 521
rect 1248 445 1300 487
rect 940 434 1300 445
rect 940 425 1078 434
rect 904 409 1078 425
rect 682 392 820 403
rect 406 386 820 392
rect 804 369 820 386
rect 854 375 870 403
rect 969 400 1078 409
rect 1112 418 1300 434
rect 1112 400 1250 418
rect 969 384 1250 400
rect 1284 384 1300 418
rect 1338 521 1390 537
rect 1338 487 1354 521
rect 1388 487 1390 521
rect 1338 420 1390 487
rect 1424 488 1490 547
rect 1610 529 1662 547
rect 1424 454 1440 488
rect 1474 454 1490 488
rect 1524 482 1576 498
rect 1524 448 1526 482
rect 1560 448 1576 482
rect 1524 420 1576 448
rect 1338 418 1576 420
rect 1338 384 1354 418
rect 1388 413 1576 418
rect 1388 384 1526 413
rect 1524 379 1526 384
rect 1560 379 1576 413
rect 1610 495 1612 529
rect 1646 495 1662 529
rect 1610 459 1662 495
rect 1610 425 1612 459
rect 1646 425 1662 459
rect 1610 409 1662 425
rect 1696 599 1734 615
rect 1696 565 1698 599
rect 1732 565 1734 599
rect 1696 511 1734 565
rect 1696 477 1698 511
rect 1732 477 1734 511
rect 1696 413 1734 477
rect 1524 375 1576 379
rect 1696 379 1698 413
rect 1732 379 1734 413
rect 1768 607 1834 649
rect 1768 573 1784 607
rect 1818 573 1834 607
rect 1768 526 1834 573
rect 1768 492 1784 526
rect 1818 492 1834 526
rect 1768 443 1834 492
rect 1768 409 1784 443
rect 1818 409 1834 443
rect 1868 599 1906 615
rect 1868 565 1870 599
rect 1904 565 1906 599
rect 1868 511 1906 565
rect 1868 477 1870 511
rect 1904 477 1906 511
rect 1868 413 1906 477
rect 1696 375 1734 379
rect 1868 379 1870 413
rect 1904 379 1906 413
rect 1940 607 2006 649
rect 1940 573 1956 607
rect 1990 573 2006 607
rect 1940 526 2006 573
rect 1940 492 1956 526
rect 1990 492 2006 526
rect 1940 443 2006 492
rect 1940 409 1956 443
rect 1990 409 2006 443
rect 2040 599 2092 615
rect 2040 565 2042 599
rect 2076 565 2092 599
rect 2040 511 2092 565
rect 2040 477 2042 511
rect 2076 477 2092 511
rect 2040 413 2092 477
rect 1868 375 1906 379
rect 2040 379 2042 413
rect 2076 379 2092 413
rect 2040 375 2092 379
rect 854 369 935 375
rect 17 309 563 352
rect 17 275 37 309
rect 71 275 105 309
rect 139 275 173 309
rect 207 275 241 309
rect 275 275 309 309
rect 343 275 377 309
rect 411 275 445 309
rect 479 275 513 309
rect 547 275 563 309
rect 597 305 737 352
rect 804 341 935 369
rect 597 271 623 305
rect 657 271 712 305
rect 746 271 801 305
rect 835 271 851 305
rect 885 237 935 341
rect 969 313 1315 350
rect 969 279 985 313
rect 1019 279 1053 313
rect 1087 279 1121 313
rect 1155 279 1189 313
rect 1223 279 1257 313
rect 1291 279 1315 313
rect 969 269 1315 279
rect 1349 305 1467 350
rect 1524 339 2092 375
rect 1349 271 1365 305
rect 1399 271 1433 305
rect 1467 271 1501 305
rect 1535 271 1569 305
rect 1603 271 1637 305
rect 1671 271 1687 305
rect 1349 269 1687 271
rect 1753 287 2095 305
rect 1753 253 1769 287
rect 1803 253 1837 287
rect 1871 253 1905 287
rect 1939 253 1973 287
rect 2007 253 2041 287
rect 2075 253 2095 287
rect 1753 242 2095 253
rect 184 203 243 219
rect 184 169 200 203
rect 234 169 243 203
rect 184 105 243 169
rect 277 203 935 237
rect 969 208 1717 235
rect 969 203 2078 208
rect 277 169 322 203
rect 456 169 494 203
rect 969 201 1140 203
rect 969 169 1003 201
rect 277 135 286 169
rect 320 135 322 169
rect 277 119 322 135
rect 356 167 422 169
rect 356 133 372 167
rect 406 133 422 167
rect 184 71 200 105
rect 234 85 243 105
rect 356 93 422 133
rect 456 135 458 169
rect 492 135 494 169
rect 456 119 494 135
rect 528 167 1003 169
rect 1138 169 1140 201
rect 1174 201 1312 203
rect 1174 169 1176 201
rect 528 133 544 167
rect 578 135 748 167
rect 578 133 594 135
rect 356 85 372 93
rect 234 71 372 85
rect 184 59 372 71
rect 406 85 422 93
rect 528 93 594 133
rect 732 133 748 135
rect 782 135 952 167
rect 782 133 798 135
rect 528 85 544 93
rect 406 59 544 85
rect 578 59 594 93
rect 184 51 594 59
rect 630 93 696 101
rect 630 59 646 93
rect 680 59 696 93
rect 630 17 696 59
rect 732 93 798 133
rect 936 133 952 135
rect 986 133 1003 167
rect 732 59 748 93
rect 782 59 798 93
rect 732 51 798 59
rect 834 93 900 101
rect 834 59 850 93
rect 884 59 900 93
rect 834 17 900 59
rect 936 93 1003 133
rect 936 59 952 93
rect 986 59 1003 93
rect 936 51 1003 59
rect 1037 161 1103 167
rect 1037 127 1053 161
rect 1087 127 1103 161
rect 1037 93 1103 127
rect 1037 59 1053 93
rect 1087 59 1103 93
rect 1037 17 1103 59
rect 1138 101 1176 169
rect 1310 169 1312 201
rect 1346 201 1484 203
rect 1346 169 1348 201
rect 1138 67 1140 101
rect 1174 67 1176 101
rect 1138 51 1176 67
rect 1210 133 1226 167
rect 1260 133 1276 167
rect 1210 93 1276 133
rect 1210 59 1226 93
rect 1260 59 1276 93
rect 1210 17 1276 59
rect 1310 101 1348 169
rect 1482 169 1484 201
rect 1518 201 1683 203
rect 1518 169 1534 201
rect 1310 67 1312 101
rect 1346 67 1348 101
rect 1310 51 1348 67
rect 1382 133 1398 167
rect 1432 133 1448 167
rect 1382 93 1448 133
rect 1382 59 1398 93
rect 1432 59 1448 93
rect 1382 17 1448 59
rect 1482 101 1534 169
rect 1668 169 1683 201
rect 1717 192 2078 203
rect 1717 174 1856 192
rect 1717 169 1725 174
rect 1482 67 1484 101
rect 1518 67 1534 101
rect 1482 51 1534 67
rect 1568 133 1584 167
rect 1618 133 1634 167
rect 1568 93 1634 133
rect 1568 59 1584 93
rect 1618 59 1634 93
rect 1568 17 1634 59
rect 1668 101 1725 169
rect 1848 158 1856 174
rect 1890 174 2028 192
rect 1890 158 1898 174
rect 1668 67 1683 101
rect 1717 67 1725 101
rect 1668 51 1725 67
rect 1759 124 1814 140
rect 1759 90 1770 124
rect 1804 90 1814 124
rect 1759 17 1814 90
rect 1848 101 1898 158
rect 2022 158 2028 174
rect 2062 158 2078 192
rect 1848 67 1856 101
rect 1890 67 1898 101
rect 1848 51 1898 67
rect 1932 124 1988 140
rect 1932 90 1942 124
rect 1976 90 1988 124
rect 1932 17 1988 90
rect 2022 101 2078 158
rect 2022 67 2028 101
rect 2062 67 2078 101
rect 2022 51 2078 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o41ai_4
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6574754
string GDS_START 6556806
<< end >>
