magic
tech sky130A
magscale 1 2
timestamp 1627201166
<< checkpaint >>
rect -1260 -1349 1554 1995
<< nwell >>
rect 0 0 294 672
<< pmos >>
rect 89 36 119 636
rect 175 36 205 636
<< pdiff >>
rect 36 605 89 636
rect 36 571 44 605
rect 78 571 89 605
rect 36 533 89 571
rect 36 499 44 533
rect 78 499 89 533
rect 36 461 89 499
rect 36 427 44 461
rect 78 427 89 461
rect 36 389 89 427
rect 36 355 44 389
rect 78 355 89 389
rect 36 317 89 355
rect 36 283 44 317
rect 78 283 89 317
rect 36 245 89 283
rect 36 211 44 245
rect 78 211 89 245
rect 36 173 89 211
rect 36 139 44 173
rect 78 139 89 173
rect 36 101 89 139
rect 36 67 44 101
rect 78 67 89 101
rect 36 36 89 67
rect 119 605 175 636
rect 119 571 130 605
rect 164 571 175 605
rect 119 533 175 571
rect 119 499 130 533
rect 164 499 175 533
rect 119 461 175 499
rect 119 427 130 461
rect 164 427 175 461
rect 119 389 175 427
rect 119 355 130 389
rect 164 355 175 389
rect 119 317 175 355
rect 119 283 130 317
rect 164 283 175 317
rect 119 245 175 283
rect 119 211 130 245
rect 164 211 175 245
rect 119 173 175 211
rect 119 139 130 173
rect 164 139 175 173
rect 119 101 175 139
rect 119 67 130 101
rect 164 67 175 101
rect 119 36 175 67
rect 205 605 258 636
rect 205 571 216 605
rect 250 571 258 605
rect 205 533 258 571
rect 205 499 216 533
rect 250 499 258 533
rect 205 461 258 499
rect 205 427 216 461
rect 250 427 258 461
rect 205 389 258 427
rect 205 355 216 389
rect 250 355 258 389
rect 205 317 258 355
rect 205 283 216 317
rect 250 283 258 317
rect 205 245 258 283
rect 205 211 216 245
rect 250 211 258 245
rect 205 173 258 211
rect 205 139 216 173
rect 250 139 258 173
rect 205 101 258 139
rect 205 67 216 101
rect 250 67 258 101
rect 205 36 258 67
<< pdiffc >>
rect 44 571 78 605
rect 44 499 78 533
rect 44 427 78 461
rect 44 355 78 389
rect 44 283 78 317
rect 44 211 78 245
rect 44 139 78 173
rect 44 67 78 101
rect 130 571 164 605
rect 130 499 164 533
rect 130 427 164 461
rect 130 355 164 389
rect 130 283 164 317
rect 130 211 164 245
rect 130 139 164 173
rect 130 67 164 101
rect 216 571 250 605
rect 216 499 250 533
rect 216 427 250 461
rect 216 355 250 389
rect 216 283 250 317
rect 216 211 250 245
rect 216 139 250 173
rect 216 67 250 101
<< poly >>
rect 80 719 214 735
rect 80 685 96 719
rect 130 685 164 719
rect 198 685 214 719
rect 80 667 214 685
rect 89 662 205 667
rect 89 636 119 662
rect 175 636 205 662
rect 89 10 119 36
rect 175 10 205 36
<< polycont >>
rect 96 685 130 719
rect 164 685 198 719
<< locali >>
rect 80 719 214 735
rect 80 685 94 719
rect 130 685 164 719
rect 200 685 214 719
rect 80 667 214 685
rect 44 605 78 621
rect 44 533 78 571
rect 44 461 78 499
rect 44 389 78 427
rect 44 317 78 355
rect 44 245 78 283
rect 44 173 78 211
rect 44 101 78 139
rect 44 47 78 67
rect 130 605 164 621
rect 130 533 164 571
rect 130 461 164 499
rect 130 389 164 427
rect 130 317 164 355
rect 130 245 164 283
rect 130 173 164 211
rect 130 101 164 139
rect 130 51 164 67
rect 216 605 250 621
rect 216 533 250 571
rect 216 461 250 499
rect 216 389 250 427
rect 216 317 250 355
rect 216 245 250 283
rect 216 173 250 211
rect 216 101 250 139
rect 216 51 250 67
<< viali >>
rect 94 685 96 719
rect 96 685 128 719
rect 166 685 198 719
rect 198 685 200 719
rect 44 571 78 605
rect 44 499 78 533
rect 44 427 78 461
rect 44 355 78 389
rect 44 283 78 317
rect 44 211 78 245
rect 44 139 78 173
rect 44 67 78 101
rect 130 571 164 605
rect 130 499 164 533
rect 130 427 164 461
rect 130 355 164 389
rect 130 283 164 317
rect 130 211 164 245
rect 130 139 164 173
rect 130 67 164 101
rect 216 571 250 605
rect 216 499 250 533
rect 216 427 250 461
rect 216 355 250 389
rect 216 283 250 317
rect 216 211 250 245
rect 216 139 250 173
rect 216 67 250 101
<< metal1 >>
rect 82 719 212 731
rect 82 685 94 719
rect 128 685 166 719
rect 200 685 212 719
rect 82 673 212 685
rect 38 605 84 621
rect 38 571 44 605
rect 78 571 84 605
rect 38 533 84 571
rect 38 499 44 533
rect 78 499 84 533
rect 38 461 84 499
rect 38 427 44 461
rect 78 427 84 461
rect 38 389 84 427
rect 38 355 44 389
rect 78 355 84 389
rect 38 317 84 355
rect 38 283 44 317
rect 78 283 84 317
rect 38 245 84 283
rect 38 211 44 245
rect 78 211 84 245
rect 38 173 84 211
rect 38 139 44 173
rect 78 139 84 173
rect 38 101 84 139
rect 38 67 44 101
rect 78 67 84 101
rect 38 -29 84 67
rect 121 610 173 621
rect 121 546 173 558
rect 121 461 173 494
rect 121 427 130 461
rect 164 427 173 461
rect 121 389 173 427
rect 121 355 130 389
rect 164 355 173 389
rect 121 317 173 355
rect 121 283 130 317
rect 164 283 173 317
rect 121 245 173 283
rect 121 211 130 245
rect 164 211 173 245
rect 121 173 173 211
rect 121 139 130 173
rect 164 139 173 173
rect 121 101 173 139
rect 121 67 130 101
rect 164 67 173 101
rect 121 51 173 67
rect 210 605 256 621
rect 210 571 216 605
rect 250 571 256 605
rect 210 533 256 571
rect 210 499 216 533
rect 250 499 256 533
rect 210 461 256 499
rect 210 427 216 461
rect 250 427 256 461
rect 210 389 256 427
rect 210 355 216 389
rect 250 355 256 389
rect 210 317 256 355
rect 210 283 216 317
rect 250 283 256 317
rect 210 245 256 283
rect 210 211 216 245
rect 250 211 256 245
rect 210 173 256 211
rect 210 139 216 173
rect 250 139 256 173
rect 210 101 256 139
rect 210 67 216 101
rect 250 67 256 101
rect 210 -29 256 67
rect 38 -89 256 -29
<< via1 >>
rect 121 605 173 610
rect 121 571 130 605
rect 130 571 164 605
rect 164 571 173 605
rect 121 558 173 571
rect 121 533 173 546
rect 121 499 130 533
rect 130 499 164 533
rect 164 499 173 533
rect 121 494 173 499
<< metal2 >>
rect 121 610 173 616
rect 121 546 173 558
rect 121 488 173 494
<< labels >>
flabel metal2 s 121 488 173 616 0 FreeSans 400 0 0 0 DRAIN
port 2 nsew
flabel metal1 s 38 -89 256 -29 0 FreeSans 400 0 0 0 SOURCE
port 4 nsew
flabel metal1 s 82 673 212 731 0 FreeSans 400 0 0 0 GATE
port 3 nsew
flabel nwell s 75 663 79 670 0 FreeSans 400 0 0 0 BULK
port 1 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9176582
string GDS_START 9170258
string path 0.950 -1.475 6.400 -1.475 
<< end >>
