magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 4 241 391 263
rect 4 49 767 241
rect 0 0 768 49
<< scnmos >>
rect 83 69 113 237
rect 169 69 199 237
rect 274 153 304 237
rect 478 47 508 215
rect 564 47 594 215
rect 658 47 688 215
<< scpmoshvt >>
rect 83 367 113 619
rect 169 367 199 619
rect 278 367 308 451
rect 478 367 508 619
rect 564 367 594 619
rect 658 367 688 619
<< ndiff >>
rect 30 225 83 237
rect 30 191 38 225
rect 72 191 83 225
rect 30 115 83 191
rect 30 81 38 115
rect 72 81 83 115
rect 30 69 83 81
rect 113 212 169 237
rect 113 178 124 212
rect 158 178 169 212
rect 113 115 169 178
rect 113 81 124 115
rect 158 81 169 115
rect 113 69 169 81
rect 199 192 274 237
rect 199 158 210 192
rect 244 158 274 192
rect 199 153 274 158
rect 304 202 365 237
rect 304 168 315 202
rect 349 168 365 202
rect 304 153 365 168
rect 199 115 252 153
rect 199 81 210 115
rect 244 81 252 115
rect 199 69 252 81
rect 425 125 478 215
rect 425 91 433 125
rect 467 91 478 125
rect 425 47 478 91
rect 508 190 564 215
rect 508 156 519 190
rect 553 156 564 190
rect 508 101 564 156
rect 508 67 519 101
rect 553 67 564 101
rect 508 47 564 67
rect 594 47 658 215
rect 688 203 741 215
rect 688 169 699 203
rect 733 169 741 203
rect 688 93 741 169
rect 688 59 699 93
rect 733 59 741 93
rect 688 47 741 59
<< pdiff >>
rect 30 574 83 619
rect 30 540 38 574
rect 72 540 83 574
rect 30 367 83 540
rect 113 413 169 619
rect 113 379 124 413
rect 158 379 169 413
rect 113 367 169 379
rect 199 574 252 619
rect 199 540 210 574
rect 244 540 252 574
rect 199 451 252 540
rect 425 599 478 619
rect 425 565 433 599
rect 467 565 478 599
rect 425 506 478 565
rect 425 472 433 506
rect 467 472 478 506
rect 199 367 278 451
rect 308 415 369 451
rect 308 381 327 415
rect 361 381 369 415
rect 308 367 369 381
rect 425 413 478 472
rect 425 379 433 413
rect 467 379 478 413
rect 425 367 478 379
rect 508 599 564 619
rect 508 565 519 599
rect 553 565 564 599
rect 508 506 564 565
rect 508 472 519 506
rect 553 472 564 506
rect 508 413 564 472
rect 508 379 519 413
rect 553 379 564 413
rect 508 367 564 379
rect 594 607 658 619
rect 594 573 609 607
rect 643 573 658 607
rect 594 519 658 573
rect 594 485 609 519
rect 643 485 658 519
rect 594 439 658 485
rect 594 405 609 439
rect 643 405 658 439
rect 594 367 658 405
rect 688 599 741 619
rect 688 565 699 599
rect 733 565 741 599
rect 688 509 741 565
rect 688 475 699 509
rect 733 475 741 509
rect 688 413 741 475
rect 688 379 699 413
rect 733 379 741 413
rect 688 367 741 379
<< ndiffc >>
rect 38 191 72 225
rect 38 81 72 115
rect 124 178 158 212
rect 124 81 158 115
rect 210 158 244 192
rect 315 168 349 202
rect 210 81 244 115
rect 433 91 467 125
rect 519 156 553 190
rect 519 67 553 101
rect 699 169 733 203
rect 699 59 733 93
<< pdiffc >>
rect 38 540 72 574
rect 124 379 158 413
rect 210 540 244 574
rect 433 565 467 599
rect 433 472 467 506
rect 327 381 361 415
rect 433 379 467 413
rect 519 565 553 599
rect 519 472 553 506
rect 519 379 553 413
rect 609 573 643 607
rect 609 485 643 519
rect 609 405 643 439
rect 699 565 733 599
rect 699 475 733 509
rect 699 379 733 413
<< poly >>
rect 83 619 113 645
rect 169 619 199 645
rect 478 619 508 645
rect 564 619 594 645
rect 658 619 688 645
rect 278 451 308 477
rect 83 325 113 367
rect 22 309 113 325
rect 22 275 38 309
rect 72 289 113 309
rect 169 289 199 367
rect 278 325 308 367
rect 72 275 199 289
rect 22 259 199 275
rect 241 309 308 325
rect 241 275 257 309
rect 291 275 308 309
rect 241 259 308 275
rect 350 309 416 325
rect 350 275 366 309
rect 400 289 416 309
rect 478 289 508 367
rect 564 303 594 367
rect 658 303 688 367
rect 400 275 508 289
rect 350 259 508 275
rect 83 237 113 259
rect 169 237 199 259
rect 274 237 304 259
rect 478 215 508 259
rect 550 287 616 303
rect 550 253 566 287
rect 600 253 616 287
rect 550 237 616 253
rect 658 287 727 303
rect 658 253 677 287
rect 711 253 727 287
rect 658 237 727 253
rect 564 215 594 237
rect 658 215 688 237
rect 274 127 304 153
rect 83 43 113 69
rect 169 43 199 69
rect 478 21 508 47
rect 564 21 594 47
rect 658 21 688 47
<< polycont >>
rect 38 275 72 309
rect 257 275 291 309
rect 366 275 400 309
rect 566 253 600 287
rect 677 253 711 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 22 574 88 649
rect 22 540 38 574
rect 72 540 88 574
rect 22 533 88 540
rect 194 574 260 649
rect 194 540 210 574
rect 244 540 260 574
rect 194 533 260 540
rect 417 599 472 615
rect 417 565 433 599
rect 467 565 472 599
rect 417 506 472 565
rect 417 499 433 506
rect 22 472 433 499
rect 467 472 472 506
rect 22 465 472 472
rect 22 309 88 465
rect 22 275 38 309
rect 72 275 88 309
rect 122 413 165 431
rect 122 379 124 413
rect 158 379 165 413
rect 22 225 88 241
rect 22 191 38 225
rect 72 191 88 225
rect 22 115 88 191
rect 22 81 38 115
rect 72 81 88 115
rect 22 17 88 81
rect 122 212 165 379
rect 212 309 291 424
rect 212 275 257 309
rect 212 242 291 275
rect 325 415 377 431
rect 325 381 327 415
rect 361 381 377 415
rect 325 325 377 381
rect 417 413 472 465
rect 417 379 433 413
rect 467 379 472 413
rect 417 363 472 379
rect 325 309 403 325
rect 325 275 366 309
rect 400 275 403 309
rect 122 178 124 212
rect 158 178 165 212
rect 325 211 403 275
rect 325 208 383 211
rect 122 115 165 178
rect 122 81 124 115
rect 158 81 165 115
rect 122 65 165 81
rect 199 192 260 208
rect 199 158 210 192
rect 244 158 260 192
rect 299 202 383 208
rect 299 168 315 202
rect 349 168 383 202
rect 437 206 472 363
rect 506 599 559 615
rect 506 565 519 599
rect 553 565 559 599
rect 506 506 559 565
rect 506 472 519 506
rect 553 472 559 506
rect 506 413 559 472
rect 506 379 519 413
rect 553 379 559 413
rect 593 607 659 649
rect 593 573 609 607
rect 643 573 659 607
rect 593 519 659 573
rect 593 485 609 519
rect 643 485 659 519
rect 593 439 659 485
rect 593 405 609 439
rect 643 405 659 439
rect 693 599 749 615
rect 693 565 699 599
rect 733 565 749 599
rect 693 509 749 565
rect 693 475 699 509
rect 733 475 749 509
rect 693 413 749 475
rect 506 371 559 379
rect 693 379 699 413
rect 733 379 749 413
rect 693 371 749 379
rect 506 337 749 371
rect 506 287 641 303
rect 506 253 566 287
rect 600 253 641 287
rect 506 240 641 253
rect 677 287 737 303
rect 711 253 737 287
rect 677 237 737 253
rect 437 190 569 206
rect 437 172 519 190
rect 299 159 383 168
rect 199 115 260 158
rect 517 156 519 172
rect 553 156 569 190
rect 199 81 210 115
rect 244 81 260 115
rect 199 17 260 81
rect 417 125 483 138
rect 417 91 433 125
rect 467 91 483 125
rect 417 17 483 91
rect 517 101 569 156
rect 517 67 519 101
rect 553 67 569 101
rect 517 51 569 67
rect 683 169 699 203
rect 733 169 749 203
rect 683 93 749 169
rect 683 59 699 93
rect 733 59 749 93
rect 683 17 749 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21bo_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3744544
string GDS_START 3736946
<< end >>
