magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 332 1094 704
<< pwell >>
rect 288 49 1055 248
rect 0 0 1056 49
<< scnmos >>
rect 371 74 401 222
rect 473 74 503 222
rect 571 74 601 222
rect 671 74 701 222
rect 758 74 788 222
rect 856 74 886 222
rect 942 74 972 222
<< scpmoshvt >>
rect 86 388 116 588
rect 176 388 206 588
rect 272 388 302 588
rect 362 388 392 588
rect 463 388 493 588
rect 563 388 593 588
rect 670 368 700 592
rect 760 368 790 592
rect 850 368 880 592
rect 940 368 970 592
<< ndiff >>
rect 314 188 371 222
rect 314 154 326 188
rect 360 154 371 188
rect 314 120 371 154
rect 314 86 326 120
rect 360 86 371 120
rect 314 74 371 86
rect 401 120 473 222
rect 401 86 426 120
rect 460 86 473 120
rect 401 74 473 86
rect 503 188 571 222
rect 503 154 526 188
rect 560 154 571 188
rect 503 120 571 154
rect 503 86 526 120
rect 560 86 571 120
rect 503 74 571 86
rect 601 120 671 222
rect 601 86 626 120
rect 660 86 671 120
rect 601 74 671 86
rect 701 210 758 222
rect 701 176 713 210
rect 747 176 758 210
rect 701 120 758 176
rect 701 86 713 120
rect 747 86 758 120
rect 701 74 758 86
rect 788 131 856 222
rect 788 97 799 131
rect 833 97 856 131
rect 788 74 856 97
rect 886 210 942 222
rect 886 176 897 210
rect 931 176 942 210
rect 886 120 942 176
rect 886 86 897 120
rect 931 86 942 120
rect 886 74 942 86
rect 972 139 1029 222
rect 972 105 983 139
rect 1017 105 1029 139
rect 972 74 1029 105
<< pdiff >>
rect 611 588 670 592
rect 27 576 86 588
rect 27 542 39 576
rect 73 542 86 576
rect 27 505 86 542
rect 27 471 39 505
rect 73 471 86 505
rect 27 434 86 471
rect 27 400 39 434
rect 73 400 86 434
rect 27 388 86 400
rect 116 576 176 588
rect 116 542 129 576
rect 163 542 176 576
rect 116 508 176 542
rect 116 474 129 508
rect 163 474 176 508
rect 116 440 176 474
rect 116 406 129 440
rect 163 406 176 440
rect 116 388 176 406
rect 206 576 272 588
rect 206 542 222 576
rect 256 542 272 576
rect 206 388 272 542
rect 302 437 362 588
rect 302 403 315 437
rect 349 403 362 437
rect 302 388 362 403
rect 392 576 463 588
rect 392 542 410 576
rect 444 542 463 576
rect 392 388 463 542
rect 493 576 563 588
rect 493 542 516 576
rect 550 542 563 576
rect 493 508 563 542
rect 493 474 516 508
rect 550 474 563 508
rect 493 388 563 474
rect 593 580 670 588
rect 593 546 623 580
rect 657 546 670 580
rect 593 508 670 546
rect 593 474 623 508
rect 657 474 670 508
rect 593 388 670 474
rect 617 368 670 388
rect 700 580 760 592
rect 700 546 713 580
rect 747 546 760 580
rect 700 497 760 546
rect 700 463 713 497
rect 747 463 760 497
rect 700 414 760 463
rect 700 380 713 414
rect 747 380 760 414
rect 700 368 760 380
rect 790 580 850 592
rect 790 546 803 580
rect 837 546 850 580
rect 790 478 850 546
rect 790 444 803 478
rect 837 444 850 478
rect 790 368 850 444
rect 880 580 940 592
rect 880 546 893 580
rect 927 546 940 580
rect 880 497 940 546
rect 880 463 893 497
rect 927 463 940 497
rect 880 414 940 463
rect 880 380 893 414
rect 927 380 940 414
rect 880 368 940 380
rect 970 580 1029 592
rect 970 546 983 580
rect 1017 546 1029 580
rect 970 478 1029 546
rect 970 444 983 478
rect 1017 444 1029 478
rect 970 368 1029 444
<< ndiffc >>
rect 326 154 360 188
rect 326 86 360 120
rect 426 86 460 120
rect 526 154 560 188
rect 526 86 560 120
rect 626 86 660 120
rect 713 176 747 210
rect 713 86 747 120
rect 799 97 833 131
rect 897 176 931 210
rect 897 86 931 120
rect 983 105 1017 139
<< pdiffc >>
rect 39 542 73 576
rect 39 471 73 505
rect 39 400 73 434
rect 129 542 163 576
rect 129 474 163 508
rect 129 406 163 440
rect 222 542 256 576
rect 315 403 349 437
rect 410 542 444 576
rect 516 542 550 576
rect 516 474 550 508
rect 623 546 657 580
rect 623 474 657 508
rect 713 546 747 580
rect 713 463 747 497
rect 713 380 747 414
rect 803 546 837 580
rect 803 444 837 478
rect 893 546 927 580
rect 893 463 927 497
rect 893 380 927 414
rect 983 546 1017 580
rect 983 444 1017 478
<< poly >>
rect 86 588 116 614
rect 176 588 206 614
rect 272 588 302 614
rect 362 588 392 614
rect 463 588 493 614
rect 563 588 593 614
rect 670 592 700 618
rect 760 592 790 618
rect 850 592 880 618
rect 940 592 970 618
rect 86 373 116 388
rect 176 373 206 388
rect 272 373 302 388
rect 362 373 392 388
rect 463 373 493 388
rect 563 373 593 388
rect 83 326 119 373
rect 173 356 209 373
rect 21 310 119 326
rect 21 276 37 310
rect 71 276 119 310
rect 161 340 227 356
rect 161 306 177 340
rect 211 306 227 340
rect 161 290 227 306
rect 269 301 305 373
rect 359 301 395 373
rect 460 356 496 373
rect 21 242 119 276
rect 269 267 395 301
rect 443 340 509 356
rect 443 306 459 340
rect 493 306 509 340
rect 560 310 596 373
rect 670 353 700 368
rect 760 353 790 368
rect 850 353 880 368
rect 940 353 970 368
rect 667 326 703 353
rect 757 326 793 353
rect 847 326 883 353
rect 937 326 973 353
rect 667 310 973 326
rect 443 290 509 306
rect 551 294 617 310
rect 269 248 401 267
rect 21 208 37 242
rect 71 208 119 242
rect 21 174 119 208
rect 21 140 37 174
rect 71 140 119 174
rect 21 106 119 140
rect 21 72 37 106
rect 71 72 119 106
rect 21 56 119 72
rect 210 237 401 248
rect 210 172 299 237
rect 371 222 401 237
rect 473 222 503 290
rect 551 260 567 294
rect 601 260 617 294
rect 667 276 683 310
rect 717 276 751 310
rect 785 276 819 310
rect 853 276 887 310
rect 921 276 973 310
rect 667 260 973 276
rect 551 244 617 260
rect 571 222 601 244
rect 671 222 701 260
rect 758 222 788 260
rect 856 222 886 260
rect 942 222 972 260
rect 210 138 226 172
rect 260 138 299 172
rect 210 104 299 138
rect 210 70 226 104
rect 260 70 299 104
rect 210 54 299 70
rect 371 48 401 74
rect 473 48 503 74
rect 571 48 601 74
rect 671 48 701 74
rect 758 48 788 74
rect 856 48 886 74
rect 942 48 972 74
<< polycont >>
rect 37 276 71 310
rect 177 306 211 340
rect 459 306 493 340
rect 37 208 71 242
rect 37 140 71 174
rect 37 72 71 106
rect 567 260 601 294
rect 683 276 717 310
rect 751 276 785 310
rect 819 276 853 310
rect 887 276 921 310
rect 226 138 260 172
rect 226 70 260 104
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 576 73 649
rect 23 542 39 576
rect 23 505 73 542
rect 23 471 39 505
rect 23 434 73 471
rect 23 400 39 434
rect 23 384 73 400
rect 113 576 163 592
rect 113 542 129 576
rect 203 576 466 592
rect 203 542 222 576
rect 256 542 410 576
rect 444 542 466 576
rect 500 576 566 592
rect 500 542 516 576
rect 550 542 566 576
rect 113 508 163 542
rect 500 508 566 542
rect 113 474 129 508
rect 163 474 516 508
rect 550 474 566 508
rect 113 440 163 474
rect 500 458 566 474
rect 607 580 673 649
rect 607 546 623 580
rect 657 546 673 580
rect 607 508 673 546
rect 607 474 623 508
rect 657 474 673 508
rect 607 458 673 474
rect 713 580 747 596
rect 713 497 747 546
rect 113 406 129 440
rect 113 390 163 406
rect 299 437 365 440
rect 299 403 315 437
rect 349 424 365 437
rect 349 403 679 424
rect 299 390 679 403
rect 121 340 509 356
rect 21 310 87 326
rect 21 276 37 310
rect 71 276 87 310
rect 121 306 177 340
rect 211 306 459 340
rect 493 306 509 340
rect 645 326 679 390
rect 713 414 747 463
rect 787 580 837 649
rect 787 546 803 580
rect 787 478 837 546
rect 787 444 803 478
rect 787 428 837 444
rect 877 580 943 596
rect 877 546 893 580
rect 927 546 943 580
rect 877 497 943 546
rect 877 463 893 497
rect 927 463 943 497
rect 877 414 943 463
rect 983 580 1033 649
rect 1017 546 1033 580
rect 983 478 1033 546
rect 1017 444 1033 478
rect 983 428 1033 444
rect 877 394 893 414
rect 747 380 893 394
rect 927 394 943 414
rect 927 380 1031 394
rect 713 360 1031 380
rect 645 310 937 326
rect 121 290 509 306
rect 551 294 611 310
rect 21 256 87 276
rect 551 260 567 294
rect 601 260 611 294
rect 551 256 611 260
rect 21 242 611 256
rect 21 208 37 242
rect 71 222 611 242
rect 645 276 683 310
rect 717 276 751 310
rect 785 276 819 310
rect 853 276 887 310
rect 921 276 937 310
rect 645 260 937 276
rect 71 208 87 222
rect 21 174 87 208
rect 645 188 679 260
rect 985 226 1031 360
rect 21 140 37 174
rect 71 140 87 174
rect 21 106 87 140
rect 21 72 37 106
rect 71 72 87 106
rect 21 56 87 72
rect 210 172 276 188
rect 210 138 226 172
rect 260 138 276 172
rect 210 104 276 138
rect 210 70 226 104
rect 260 70 276 104
rect 310 154 326 188
rect 360 154 526 188
rect 560 154 679 188
rect 713 210 1031 226
rect 747 192 897 210
rect 310 120 376 154
rect 510 120 576 154
rect 713 120 747 176
rect 881 176 897 192
rect 931 192 1031 210
rect 310 86 326 120
rect 360 86 376 120
rect 310 70 376 86
rect 410 86 426 120
rect 460 86 476 120
rect 210 54 276 70
rect 410 17 476 86
rect 510 86 526 120
rect 560 86 576 120
rect 510 70 576 86
rect 610 86 626 120
rect 660 86 676 120
rect 610 17 676 86
rect 713 70 747 86
rect 783 131 833 158
rect 783 97 799 131
rect 783 17 833 97
rect 881 120 931 176
rect 881 86 897 120
rect 881 70 931 86
rect 967 139 1033 158
rect 967 105 983 139
rect 1017 105 1033 139
rect 967 17 1033 105
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or3_4
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 1665080
string GDS_START 1655644
<< end >>
