magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 4 49 664 241
rect 0 0 672 49
<< scnmos >>
rect 151 47 181 215
rect 239 47 269 215
rect 331 47 361 215
rect 441 47 471 215
rect 555 47 585 215
<< scpmoshvt >>
rect 151 367 181 619
rect 259 367 289 619
rect 369 367 399 619
rect 483 367 513 619
rect 555 367 585 619
<< ndiff >>
rect 30 203 151 215
rect 30 169 38 203
rect 72 169 151 203
rect 30 118 151 169
rect 30 101 106 118
rect 30 67 38 101
rect 72 84 106 101
rect 140 84 151 118
rect 72 67 151 84
rect 30 47 151 67
rect 181 47 239 215
rect 269 47 331 215
rect 361 203 441 215
rect 361 169 384 203
rect 418 169 441 203
rect 361 101 441 169
rect 361 67 384 101
rect 418 67 441 101
rect 361 47 441 67
rect 471 157 555 215
rect 471 123 496 157
rect 530 123 555 157
rect 471 89 555 123
rect 471 55 496 89
rect 530 55 555 89
rect 471 47 555 55
rect 585 203 638 215
rect 585 169 596 203
rect 630 169 638 203
rect 585 101 638 169
rect 585 67 596 101
rect 630 67 638 101
rect 585 47 638 67
<< pdiff >>
rect 98 607 151 619
rect 98 573 106 607
rect 140 573 151 607
rect 98 533 151 573
rect 98 499 106 533
rect 140 499 151 533
rect 98 453 151 499
rect 98 419 106 453
rect 140 419 151 453
rect 98 367 151 419
rect 181 599 259 619
rect 181 565 203 599
rect 237 565 259 599
rect 181 506 259 565
rect 181 472 203 506
rect 237 472 259 506
rect 181 413 259 472
rect 181 379 203 413
rect 237 379 259 413
rect 181 367 259 379
rect 289 607 369 619
rect 289 573 312 607
rect 346 573 369 607
rect 289 504 369 573
rect 289 470 312 504
rect 346 470 369 504
rect 289 367 369 470
rect 399 607 483 619
rect 399 573 423 607
rect 457 573 483 607
rect 399 514 483 573
rect 399 480 423 514
rect 457 480 483 514
rect 399 420 483 480
rect 399 386 423 420
rect 457 386 483 420
rect 399 367 483 386
rect 513 367 555 619
rect 585 607 638 619
rect 585 573 596 607
rect 630 573 638 607
rect 585 514 638 573
rect 585 480 596 514
rect 630 480 638 514
rect 585 419 638 480
rect 585 385 596 419
rect 630 385 638 419
rect 585 367 638 385
<< ndiffc >>
rect 38 169 72 203
rect 38 67 72 101
rect 106 84 140 118
rect 384 169 418 203
rect 384 67 418 101
rect 496 123 530 157
rect 496 55 530 89
rect 596 169 630 203
rect 596 67 630 101
<< pdiffc >>
rect 106 573 140 607
rect 106 499 140 533
rect 106 419 140 453
rect 203 565 237 599
rect 203 472 237 506
rect 203 379 237 413
rect 312 573 346 607
rect 312 470 346 504
rect 423 573 457 607
rect 423 480 457 514
rect 423 386 457 420
rect 596 573 630 607
rect 596 480 630 514
rect 596 385 630 419
<< poly >>
rect 151 619 181 645
rect 259 619 289 645
rect 369 619 399 645
rect 483 619 513 645
rect 555 619 585 645
rect 151 303 181 367
rect 259 303 289 367
rect 369 335 399 367
rect 483 335 513 367
rect 111 287 181 303
rect 111 253 127 287
rect 161 253 181 287
rect 111 237 181 253
rect 223 287 289 303
rect 223 253 239 287
rect 273 253 289 287
rect 223 237 289 253
rect 331 319 399 335
rect 331 285 347 319
rect 381 285 399 319
rect 331 269 399 285
rect 441 319 513 335
rect 441 285 463 319
rect 497 285 513 319
rect 441 269 513 285
rect 555 325 585 367
rect 555 309 647 325
rect 555 275 597 309
rect 631 275 647 309
rect 151 215 181 237
rect 239 215 269 237
rect 331 215 361 269
rect 441 215 471 269
rect 555 259 647 275
rect 555 215 585 259
rect 151 21 181 47
rect 239 21 269 47
rect 331 21 361 47
rect 441 21 471 47
rect 555 21 585 47
<< polycont >>
rect 127 253 161 287
rect 239 253 273 287
rect 347 285 381 319
rect 463 285 497 319
rect 597 275 631 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 86 607 156 649
rect 86 573 106 607
rect 140 573 156 607
rect 86 533 156 573
rect 86 499 106 533
rect 140 499 156 533
rect 86 453 156 499
rect 86 419 106 453
rect 140 419 156 453
rect 190 599 257 615
rect 190 565 203 599
rect 237 565 257 599
rect 190 506 257 565
rect 190 472 203 506
rect 237 472 257 506
rect 190 420 257 472
rect 296 607 362 649
rect 296 573 312 607
rect 346 573 362 607
rect 296 504 362 573
rect 296 470 312 504
rect 346 470 362 504
rect 296 454 362 470
rect 407 607 473 615
rect 407 573 423 607
rect 457 573 473 607
rect 407 514 473 573
rect 407 480 423 514
rect 457 480 473 514
rect 407 420 473 480
rect 190 413 423 420
rect 190 385 203 413
rect 22 379 203 385
rect 237 386 423 413
rect 457 386 473 420
rect 580 607 646 649
rect 580 573 596 607
rect 630 573 646 607
rect 580 514 646 573
rect 580 480 596 514
rect 630 480 646 514
rect 580 419 646 480
rect 237 379 273 386
rect 580 385 596 419
rect 630 385 646 419
rect 22 337 273 379
rect 22 203 88 337
rect 307 319 381 352
rect 22 169 38 203
rect 72 169 88 203
rect 22 134 88 169
rect 122 287 177 303
rect 122 253 127 287
rect 161 253 177 287
rect 122 168 177 253
rect 211 287 273 303
rect 211 253 239 287
rect 307 285 347 319
rect 307 269 381 285
rect 415 319 547 352
rect 415 285 463 319
rect 497 285 547 319
rect 415 269 547 285
rect 581 309 647 351
rect 581 275 597 309
rect 631 275 647 309
rect 581 269 647 275
rect 22 118 156 134
rect 22 101 106 118
rect 22 67 38 101
rect 72 84 106 101
rect 140 84 156 118
rect 72 67 156 84
rect 211 76 273 253
rect 368 203 646 235
rect 368 169 384 203
rect 418 201 596 203
rect 418 169 434 201
rect 368 101 434 169
rect 580 169 596 201
rect 630 169 646 203
rect 22 51 156 67
rect 368 67 384 101
rect 418 67 434 101
rect 368 51 434 67
rect 480 157 546 161
rect 480 123 496 157
rect 530 123 546 157
rect 480 89 546 123
rect 480 55 496 89
rect 530 55 546 89
rect 480 17 546 55
rect 580 101 646 169
rect 580 67 596 101
rect 630 67 646 101
rect 580 51 646 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2111ai_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4765800
string GDS_START 4758896
<< end >>
