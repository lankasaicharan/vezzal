magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
<< pwell >>
rect 1625 241 1871 289
rect 1625 235 2111 241
rect 221 231 738 233
rect 33 219 738 231
rect 1135 219 2111 235
rect 33 49 2111 219
rect 0 0 2112 49
<< scnmos >>
rect 112 121 142 205
rect 184 121 214 205
rect 320 123 350 207
rect 408 123 438 207
rect 510 123 540 207
rect 609 123 639 207
rect 847 109 877 193
rect 989 65 1019 193
rect 1107 65 1137 193
rect 1245 125 1275 209
rect 1317 125 1347 209
rect 1435 125 1465 209
rect 1507 125 1537 209
rect 1704 179 1734 263
rect 1897 47 1927 131
rect 2002 47 2032 215
<< scpmoshvt >>
rect 80 463 110 547
rect 212 463 242 547
rect 306 463 336 547
rect 417 463 447 547
rect 525 463 555 547
rect 643 463 673 547
rect 847 392 877 520
rect 983 447 1013 615
rect 1069 447 1099 615
rect 1199 531 1229 615
rect 1307 531 1337 615
rect 1427 531 1457 615
rect 1559 485 1589 569
rect 1676 485 1706 613
rect 1885 367 1915 495
rect 2002 367 2032 619
<< ndiff >>
rect 247 205 320 207
rect 59 180 112 205
rect 59 146 67 180
rect 101 146 112 180
rect 59 121 112 146
rect 142 121 184 205
rect 214 180 320 205
rect 214 146 246 180
rect 280 146 320 180
rect 214 123 320 146
rect 350 185 408 207
rect 350 151 361 185
rect 395 151 408 185
rect 350 123 408 151
rect 438 123 510 207
rect 540 123 609 207
rect 639 123 712 207
rect 214 121 267 123
rect 654 108 712 123
rect 654 74 666 108
rect 700 74 712 108
rect 654 66 712 74
rect 1161 193 1245 209
rect 787 160 847 193
rect 787 126 799 160
rect 833 126 847 160
rect 787 109 847 126
rect 877 109 989 193
rect 898 81 989 109
rect 898 47 910 81
rect 944 65 989 81
rect 1019 169 1107 193
rect 1019 135 1062 169
rect 1096 135 1107 169
rect 1019 65 1107 135
rect 1137 171 1245 193
rect 1137 137 1200 171
rect 1234 137 1245 171
rect 1137 125 1245 137
rect 1275 125 1317 209
rect 1347 140 1435 209
rect 1347 125 1374 140
rect 1137 65 1187 125
rect 1362 106 1374 125
rect 1408 125 1435 140
rect 1465 125 1507 209
rect 1537 182 1590 209
rect 1537 148 1548 182
rect 1582 148 1590 182
rect 1537 125 1590 148
rect 1408 106 1420 125
rect 1362 98 1420 106
rect 1651 238 1704 263
rect 1651 204 1659 238
rect 1693 204 1704 238
rect 1651 179 1704 204
rect 1734 248 1845 263
rect 1734 214 1803 248
rect 1837 214 1845 248
rect 1734 198 1845 214
rect 1734 179 1784 198
rect 1949 202 2002 215
rect 1949 168 1957 202
rect 1991 168 2002 202
rect 1949 131 2002 168
rect 944 47 958 65
rect 898 39 958 47
rect 1844 106 1897 131
rect 1844 72 1852 106
rect 1886 72 1897 106
rect 1844 47 1897 72
rect 1927 93 2002 131
rect 1927 59 1950 93
rect 1984 59 2002 93
rect 1927 47 2002 59
rect 2032 203 2085 215
rect 2032 169 2043 203
rect 2077 169 2085 203
rect 2032 101 2085 169
rect 2032 67 2043 101
rect 2077 67 2085 101
rect 2032 47 2085 67
<< pdiff >>
rect 909 629 968 639
rect 125 562 197 578
rect 125 547 144 562
rect 27 522 80 547
rect 27 488 35 522
rect 69 488 80 522
rect 27 463 80 488
rect 110 528 144 547
rect 178 547 197 562
rect 570 558 628 574
rect 570 547 582 558
rect 178 528 212 547
rect 110 463 212 528
rect 242 531 306 547
rect 242 497 253 531
rect 287 497 306 531
rect 242 463 306 497
rect 336 520 417 547
rect 336 486 363 520
rect 397 486 417 520
rect 336 463 417 486
rect 447 463 525 547
rect 555 524 582 547
rect 616 547 628 558
rect 616 524 643 547
rect 555 463 643 524
rect 673 520 726 547
rect 909 595 921 629
rect 955 615 968 629
rect 955 595 983 615
rect 909 520 983 595
rect 673 486 684 520
rect 718 486 726 520
rect 673 463 726 486
rect 782 420 847 520
rect 782 386 790 420
rect 824 392 847 420
rect 877 447 983 520
rect 1013 489 1069 615
rect 1013 455 1024 489
rect 1058 455 1069 489
rect 1013 447 1069 455
rect 1099 531 1199 615
rect 1229 531 1307 615
rect 1337 607 1427 615
rect 1337 573 1348 607
rect 1382 573 1427 607
rect 1337 531 1427 573
rect 1457 569 1537 615
rect 1623 601 1676 613
rect 1623 569 1631 601
rect 1457 531 1559 569
rect 1099 501 1152 531
rect 1099 467 1110 501
rect 1144 467 1152 501
rect 1099 447 1152 467
rect 877 392 968 447
rect 824 386 832 392
rect 782 367 832 386
rect 1479 527 1559 531
rect 1479 493 1493 527
rect 1527 493 1559 527
rect 1479 485 1559 493
rect 1589 567 1631 569
rect 1665 567 1676 601
rect 1589 485 1676 567
rect 1706 599 1759 613
rect 1706 565 1717 599
rect 1751 565 1759 599
rect 1706 531 1759 565
rect 1706 497 1717 531
rect 1751 497 1759 531
rect 1949 607 2002 619
rect 1949 573 1957 607
rect 1991 573 2002 607
rect 1706 485 1759 497
rect 1949 509 2002 573
rect 1949 495 1957 509
rect 1832 483 1885 495
rect 1832 449 1840 483
rect 1874 449 1885 483
rect 1832 413 1885 449
rect 1832 379 1840 413
rect 1874 379 1885 413
rect 1832 367 1885 379
rect 1915 475 1957 495
rect 1991 475 2002 509
rect 1915 413 2002 475
rect 1915 379 1937 413
rect 1971 379 2002 413
rect 1915 367 2002 379
rect 2032 599 2085 619
rect 2032 565 2043 599
rect 2077 565 2085 599
rect 2032 502 2085 565
rect 2032 468 2043 502
rect 2077 468 2085 502
rect 2032 419 2085 468
rect 2032 385 2043 419
rect 2077 385 2085 419
rect 2032 367 2085 385
<< ndiffc >>
rect 67 146 101 180
rect 246 146 280 180
rect 361 151 395 185
rect 666 74 700 108
rect 799 126 833 160
rect 910 47 944 81
rect 1062 135 1096 169
rect 1200 137 1234 171
rect 1374 106 1408 140
rect 1548 148 1582 182
rect 1659 204 1693 238
rect 1803 214 1837 248
rect 1957 168 1991 202
rect 1852 72 1886 106
rect 1950 59 1984 93
rect 2043 169 2077 203
rect 2043 67 2077 101
<< pdiffc >>
rect 35 488 69 522
rect 144 528 178 562
rect 253 497 287 531
rect 363 486 397 520
rect 582 524 616 558
rect 921 595 955 629
rect 684 486 718 520
rect 790 386 824 420
rect 1024 455 1058 489
rect 1348 573 1382 607
rect 1110 467 1144 501
rect 1493 493 1527 527
rect 1631 567 1665 601
rect 1717 565 1751 599
rect 1717 497 1751 531
rect 1957 573 1991 607
rect 1840 449 1874 483
rect 1840 379 1874 413
rect 1957 475 1991 509
rect 1937 379 1971 413
rect 2043 565 2077 599
rect 2043 468 2077 502
rect 2043 385 2077 419
<< poly >>
rect 80 615 673 645
rect 80 547 110 615
rect 212 547 242 573
rect 306 547 336 573
rect 417 547 447 573
rect 525 547 555 573
rect 643 547 673 615
rect 805 602 877 618
rect 805 568 821 602
rect 855 568 877 602
rect 805 552 877 568
rect 847 520 877 552
rect 983 615 1013 641
rect 1069 615 1099 641
rect 1199 615 1229 641
rect 1307 615 1337 641
rect 1427 615 1457 641
rect 80 434 110 463
rect 70 415 136 434
rect 70 381 86 415
rect 120 381 136 415
rect 70 347 136 381
rect 70 313 86 347
rect 120 330 136 347
rect 120 313 142 330
rect 70 297 142 313
rect 112 205 142 297
rect 212 293 242 463
rect 306 307 336 463
rect 417 415 447 463
rect 417 399 483 415
rect 417 365 433 399
rect 467 365 483 399
rect 417 349 483 365
rect 184 277 250 293
rect 306 277 424 307
rect 525 295 555 463
rect 643 448 673 463
rect 609 363 673 448
rect 1676 613 1706 639
rect 2002 619 2032 645
rect 1559 569 1589 595
rect 1199 499 1229 531
rect 1169 483 1250 499
rect 1169 449 1200 483
rect 1234 449 1250 483
rect 609 347 675 363
rect 609 313 625 347
rect 659 313 675 347
rect 609 297 675 313
rect 184 243 200 277
rect 234 243 250 277
rect 184 227 250 243
rect 394 252 424 277
rect 501 279 567 295
rect 184 205 214 227
rect 320 207 350 235
rect 394 222 438 252
rect 501 245 517 279
rect 551 245 567 279
rect 501 229 567 245
rect 408 207 438 222
rect 510 207 540 229
rect 609 207 639 297
rect 847 238 877 392
rect 983 321 1013 447
rect 1069 362 1099 447
rect 1169 433 1250 449
rect 919 305 1013 321
rect 919 271 935 305
rect 969 304 1013 305
rect 1061 346 1127 362
rect 1061 312 1077 346
rect 1111 312 1127 346
rect 969 271 1019 304
rect 1061 296 1127 312
rect 919 255 1019 271
rect 727 208 877 238
rect 112 44 142 121
rect 184 44 214 121
rect 320 101 350 123
rect 294 85 360 101
rect 294 51 310 85
rect 344 51 360 85
rect 294 35 360 51
rect 408 51 438 123
rect 510 97 540 123
rect 609 97 639 123
rect 727 51 772 208
rect 847 193 877 208
rect 989 193 1019 255
rect 1169 254 1199 433
rect 1307 410 1337 531
rect 1427 450 1457 531
rect 1885 495 1915 521
rect 1409 434 1475 450
rect 1287 394 1353 410
rect 1287 360 1303 394
rect 1337 360 1353 394
rect 1287 326 1353 360
rect 1287 292 1303 326
rect 1337 292 1353 326
rect 1409 400 1425 434
rect 1459 400 1475 434
rect 1409 366 1475 400
rect 1409 332 1425 366
rect 1459 332 1475 366
rect 1409 316 1475 332
rect 1287 276 1353 292
rect 1107 224 1199 254
rect 1107 193 1137 224
rect 1245 209 1275 235
rect 1317 209 1347 276
rect 1435 209 1465 316
rect 1559 261 1589 485
rect 1676 443 1706 485
rect 1631 427 1734 443
rect 1631 393 1647 427
rect 1681 393 1734 427
rect 1631 359 1734 393
rect 1631 325 1647 359
rect 1681 325 1734 359
rect 1631 309 1734 325
rect 1704 263 1734 309
rect 1507 231 1636 261
rect 1507 209 1537 231
rect 847 83 877 109
rect 408 21 772 51
rect 1245 103 1275 125
rect 1209 87 1275 103
rect 1317 99 1347 125
rect 1435 99 1465 125
rect 1507 99 1537 125
rect 1606 103 1636 231
rect 1885 183 1915 367
rect 2002 335 2032 367
rect 1957 319 2032 335
rect 1957 285 1973 319
rect 2007 285 2032 319
rect 1957 269 2032 285
rect 2002 215 2032 269
rect 1704 153 1734 179
rect 1799 153 1927 183
rect 1799 103 1829 153
rect 1897 131 1927 153
rect 989 39 1019 65
rect 1107 39 1137 65
rect 1209 53 1225 87
rect 1259 53 1275 87
rect 1209 37 1275 53
rect 1606 87 1829 103
rect 1606 53 1622 87
rect 1656 73 1829 87
rect 1656 53 1672 73
rect 1606 37 1672 53
rect 1897 21 1927 47
rect 2002 21 2032 47
<< polycont >>
rect 821 568 855 602
rect 86 381 120 415
rect 86 313 120 347
rect 433 365 467 399
rect 1200 449 1234 483
rect 625 313 659 347
rect 200 243 234 277
rect 517 245 551 279
rect 935 271 969 305
rect 1077 312 1111 346
rect 310 51 344 85
rect 1303 360 1337 394
rect 1303 292 1337 326
rect 1425 400 1459 434
rect 1425 332 1459 366
rect 1647 393 1681 427
rect 1647 325 1681 359
rect 1973 285 2007 319
rect 1225 53 1259 87
rect 1622 53 1656 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 128 562 194 649
rect 20 522 94 547
rect 128 528 144 562
rect 178 528 194 562
rect 566 558 632 649
rect 905 629 971 649
rect 128 526 194 528
rect 232 531 313 547
rect 20 488 35 522
rect 69 492 94 522
rect 232 497 253 531
rect 287 497 313 531
rect 232 492 313 497
rect 69 488 313 492
rect 20 458 313 488
rect 19 415 136 424
rect 19 381 86 415
rect 120 381 136 415
rect 19 350 136 381
rect 19 316 31 350
rect 65 347 136 350
rect 65 316 86 347
rect 19 313 86 316
rect 120 313 136 347
rect 232 364 313 458
rect 347 520 408 547
rect 566 524 582 558
rect 616 524 632 558
rect 805 602 871 613
rect 805 568 821 602
rect 855 568 871 602
rect 905 595 921 629
rect 955 595 971 629
rect 905 593 971 595
rect 1344 607 1384 649
rect 805 559 871 568
rect 1040 559 1249 587
rect 805 553 1249 559
rect 1344 573 1348 607
rect 1382 573 1384 607
rect 1344 557 1384 573
rect 1418 579 1595 613
rect 566 522 632 524
rect 347 486 363 520
rect 397 488 408 520
rect 666 520 729 547
rect 805 525 1074 553
rect 666 488 684 520
rect 397 486 684 488
rect 718 488 729 520
rect 1184 520 1249 553
rect 1418 520 1452 579
rect 1108 501 1144 517
rect 1005 489 1074 491
rect 718 486 969 488
rect 347 454 969 486
rect 347 417 397 454
rect 232 313 327 364
rect 19 277 259 279
rect 19 243 200 277
rect 234 243 259 277
rect 19 230 259 243
rect 293 196 327 313
rect 51 180 117 196
rect 51 146 67 180
rect 101 146 117 180
rect 51 17 117 146
rect 230 180 327 196
rect 230 146 246 180
rect 280 146 327 180
rect 230 130 327 146
rect 361 185 397 417
rect 395 151 397 185
rect 361 135 397 151
rect 431 399 790 420
rect 431 365 433 399
rect 467 386 790 399
rect 824 386 855 420
rect 467 384 855 386
rect 431 176 467 365
rect 545 347 675 350
rect 545 316 625 347
rect 511 313 625 316
rect 659 313 675 347
rect 935 305 969 454
rect 501 245 517 279
rect 551 245 567 279
rect 935 255 969 271
rect 1005 455 1024 489
rect 1058 455 1074 489
rect 1005 449 1074 455
rect 1108 467 1110 501
rect 501 244 567 245
rect 501 221 901 244
rect 1005 241 1041 449
rect 1108 431 1144 467
rect 1184 486 1452 520
rect 1493 527 1527 545
rect 1184 483 1250 486
rect 1184 449 1200 483
rect 1234 449 1250 483
rect 1409 434 1459 450
rect 1108 423 1154 431
rect 1108 420 1160 423
rect 1108 415 1166 420
rect 1108 396 1234 415
rect 1122 395 1234 396
rect 1125 393 1234 395
rect 1128 392 1234 393
rect 1131 390 1234 392
rect 1136 387 1234 390
rect 1140 381 1234 387
rect 1077 347 1111 362
rect 1077 346 1166 347
rect 1111 312 1166 346
rect 1077 296 1166 312
rect 1005 221 1096 241
rect 501 210 1096 221
rect 867 187 1096 210
rect 431 160 833 176
rect 431 142 799 160
rect 431 96 467 142
rect 783 126 799 142
rect 1062 169 1096 187
rect 833 126 1028 153
rect 783 117 1028 126
rect 1062 119 1096 135
rect 783 110 849 117
rect 294 85 467 96
rect 294 51 310 85
rect 344 51 467 85
rect 650 74 666 108
rect 700 74 716 108
rect 994 85 1028 117
rect 1132 87 1166 296
rect 1200 212 1234 381
rect 1303 394 1337 410
rect 1409 400 1425 434
rect 1409 367 1459 400
rect 1303 326 1337 360
rect 1371 366 1459 367
rect 1371 350 1425 366
rect 1371 316 1375 350
rect 1409 332 1425 350
rect 1409 316 1459 332
rect 1303 280 1337 292
rect 1493 280 1527 493
rect 1561 515 1595 579
rect 1629 601 1667 649
rect 1629 567 1631 601
rect 1665 567 1667 601
rect 1629 549 1667 567
rect 1701 599 1769 615
rect 1701 565 1717 599
rect 1751 565 1769 599
rect 1701 531 1769 565
rect 1701 515 1717 531
rect 1561 497 1717 515
rect 1751 497 1769 531
rect 1921 607 1995 649
rect 1921 573 1957 607
rect 1991 573 1995 607
rect 1921 509 1995 573
rect 1561 481 1769 497
rect 1561 427 1701 443
rect 1561 393 1647 427
rect 1681 393 1701 427
rect 1561 359 1701 393
rect 1561 325 1647 359
rect 1681 325 1701 359
rect 1561 314 1701 325
rect 1735 280 1769 481
rect 1824 483 1887 499
rect 1824 449 1840 483
rect 1874 449 1887 483
rect 1824 413 1887 449
rect 1824 379 1840 413
rect 1874 379 1887 413
rect 1824 335 1887 379
rect 1921 475 1957 509
rect 1991 475 1995 509
rect 1921 413 1995 475
rect 1921 379 1937 413
rect 1971 379 1995 413
rect 1921 369 1995 379
rect 2029 599 2095 615
rect 2029 565 2043 599
rect 2077 565 2095 599
rect 2029 502 2095 565
rect 2029 468 2043 502
rect 2077 468 2095 502
rect 2029 419 2095 468
rect 2029 385 2043 419
rect 2077 385 2095 419
rect 2029 369 2095 385
rect 1824 319 2007 335
rect 1824 301 1973 319
rect 1303 246 1598 280
rect 1200 176 1498 212
rect 1200 171 1245 176
rect 1234 137 1245 171
rect 1200 121 1245 137
rect 1358 140 1424 142
rect 1358 106 1374 140
rect 1408 106 1424 140
rect 1132 85 1225 87
rect 650 17 716 74
rect 894 81 960 83
rect 894 47 910 81
rect 944 47 960 81
rect 994 53 1225 85
rect 1259 53 1275 87
rect 994 51 1275 53
rect 894 17 960 47
rect 1358 17 1424 106
rect 1462 98 1498 176
rect 1532 182 1598 246
rect 1643 246 1769 280
rect 1877 285 1973 301
rect 1877 269 2007 285
rect 1803 248 1843 264
rect 1643 238 1695 246
rect 1643 204 1659 238
rect 1693 204 1695 238
rect 1837 214 1843 248
rect 1803 212 1843 214
rect 1643 188 1695 204
rect 1532 148 1548 182
rect 1582 148 1598 182
rect 1532 132 1598 148
rect 1752 178 1843 212
rect 1462 87 1672 98
rect 1462 53 1622 87
rect 1656 53 1672 87
rect 1752 17 1786 178
rect 1877 122 1911 269
rect 2041 218 2095 369
rect 1836 106 1911 122
rect 1836 72 1852 106
rect 1886 72 1911 106
rect 1836 56 1911 72
rect 1945 202 1997 218
rect 1945 168 1957 202
rect 1991 168 1997 202
rect 1945 93 1997 168
rect 1945 59 1950 93
rect 1984 59 1997 93
rect 1945 17 1997 59
rect 2031 203 2095 218
rect 2031 169 2043 203
rect 2077 169 2095 203
rect 2031 101 2095 169
rect 2031 67 2043 101
rect 2077 67 2095 101
rect 2031 51 2095 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 316 65 350
rect 511 316 545 350
rect 1375 316 1409 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 19 350 77 356
rect 19 316 31 350
rect 65 347 77 350
rect 499 350 557 356
rect 499 347 511 350
rect 65 319 511 347
rect 65 316 77 319
rect 19 310 77 316
rect 499 316 511 319
rect 545 347 557 350
rect 1363 350 1421 356
rect 1363 347 1375 350
rect 545 319 1375 347
rect 545 316 557 319
rect 499 310 557 316
rect 1363 316 1375 319
rect 1409 316 1421 350
rect 1363 310 1421 316
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfrtn_1
flabel metal1 s 31 316 65 350 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 1663 390 1697 424 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 2047 94 2081 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 168 2081 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 464 2081 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 538 2081 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry R90
string GDS_END 6425384
string GDS_START 6408722
<< end >>
