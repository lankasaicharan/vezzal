magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 260 248 726 290
rect 147 49 726 248
rect 0 0 768 49
<< scpmos >>
rect 81 368 117 592
rect 331 392 367 592
rect 427 392 463 592
rect 517 392 553 592
rect 595 392 631 592
<< nmoslvt >>
rect 226 74 256 222
rect 336 136 366 264
rect 431 136 461 264
rect 517 136 547 264
rect 617 136 647 264
<< ndiff >>
rect 286 222 336 264
rect 173 210 226 222
rect 173 176 181 210
rect 215 176 226 210
rect 173 120 226 176
rect 173 86 181 120
rect 215 86 226 120
rect 173 74 226 86
rect 256 184 336 222
rect 256 150 291 184
rect 325 150 336 184
rect 256 136 336 150
rect 366 136 431 264
rect 461 221 517 264
rect 461 187 472 221
rect 506 187 517 221
rect 461 136 517 187
rect 547 182 617 264
rect 547 148 572 182
rect 606 148 617 182
rect 547 136 617 148
rect 647 251 700 264
rect 647 217 658 251
rect 692 217 700 251
rect 647 136 700 217
rect 256 116 313 136
rect 256 82 267 116
rect 301 82 313 116
rect 256 74 313 82
<< pdiff >>
rect 29 580 81 592
rect 29 546 37 580
rect 71 546 81 580
rect 29 497 81 546
rect 29 463 37 497
rect 71 463 81 497
rect 29 414 81 463
rect 29 380 37 414
rect 71 380 81 414
rect 29 368 81 380
rect 117 580 169 592
rect 117 546 127 580
rect 161 546 169 580
rect 117 497 169 546
rect 117 463 127 497
rect 161 463 169 497
rect 117 414 169 463
rect 117 380 127 414
rect 161 380 169 414
rect 279 580 331 592
rect 279 546 287 580
rect 321 546 331 580
rect 279 510 331 546
rect 279 476 287 510
rect 321 476 331 510
rect 279 440 331 476
rect 279 406 287 440
rect 321 406 331 440
rect 279 392 331 406
rect 367 580 427 592
rect 367 546 380 580
rect 414 546 427 580
rect 367 508 427 546
rect 367 474 380 508
rect 414 474 427 508
rect 367 392 427 474
rect 463 580 517 592
rect 463 546 473 580
rect 507 546 517 580
rect 463 510 517 546
rect 463 476 473 510
rect 507 476 517 510
rect 463 440 517 476
rect 463 406 473 440
rect 507 406 517 440
rect 463 392 517 406
rect 553 392 595 592
rect 631 580 683 592
rect 631 546 641 580
rect 675 546 683 580
rect 631 509 683 546
rect 631 475 641 509
rect 675 475 683 509
rect 631 438 683 475
rect 631 404 641 438
rect 675 404 683 438
rect 631 392 683 404
rect 117 368 169 380
<< ndiffc >>
rect 181 176 215 210
rect 181 86 215 120
rect 291 150 325 184
rect 472 187 506 221
rect 572 148 606 182
rect 658 217 692 251
rect 267 82 301 116
<< pdiffc >>
rect 37 546 71 580
rect 37 463 71 497
rect 37 380 71 414
rect 127 546 161 580
rect 127 463 161 497
rect 127 380 161 414
rect 287 546 321 580
rect 287 476 321 510
rect 287 406 321 440
rect 380 546 414 580
rect 380 474 414 508
rect 473 546 507 580
rect 473 476 507 510
rect 473 406 507 440
rect 641 546 675 580
rect 641 475 675 509
rect 641 404 675 438
<< poly >>
rect 81 592 117 618
rect 331 592 367 618
rect 427 592 463 618
rect 517 592 553 618
rect 595 592 631 618
rect 81 330 117 368
rect 331 356 367 392
rect 427 356 463 392
rect 301 340 367 356
rect 81 314 256 330
rect 81 280 101 314
rect 135 280 206 314
rect 240 280 256 314
rect 301 306 317 340
rect 351 306 367 340
rect 301 290 367 306
rect 409 340 475 356
rect 409 306 425 340
rect 459 306 475 340
rect 409 290 475 306
rect 81 264 256 280
rect 336 264 366 290
rect 431 264 461 290
rect 517 279 553 392
rect 595 309 631 392
rect 595 279 647 309
rect 517 264 547 279
rect 617 264 647 279
rect 226 222 256 264
rect 336 110 366 136
rect 431 110 461 136
rect 517 114 547 136
rect 617 114 647 136
rect 509 98 575 114
rect 226 48 256 74
rect 509 64 525 98
rect 559 64 575 98
rect 509 48 575 64
rect 617 98 743 114
rect 617 64 693 98
rect 727 64 743 98
rect 617 48 743 64
<< polycont >>
rect 101 280 135 314
rect 206 280 240 314
rect 317 306 351 340
rect 425 306 459 340
rect 525 64 559 98
rect 693 64 727 98
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 580 87 596
rect 17 546 37 580
rect 71 546 87 580
rect 17 497 87 546
rect 17 463 37 497
rect 71 463 87 497
rect 17 414 87 463
rect 17 380 37 414
rect 71 380 87 414
rect 17 364 87 380
rect 127 580 177 649
rect 161 546 177 580
rect 127 497 177 546
rect 161 463 177 497
rect 127 414 177 463
rect 161 380 177 414
rect 271 580 337 596
rect 271 546 287 580
rect 321 546 337 580
rect 271 510 337 546
rect 271 476 287 510
rect 321 476 337 510
rect 271 440 337 476
rect 377 580 417 649
rect 377 546 380 580
rect 414 546 417 580
rect 377 508 417 546
rect 377 474 380 508
rect 414 474 417 508
rect 377 458 417 474
rect 457 580 523 596
rect 457 546 473 580
rect 507 546 523 580
rect 457 510 523 546
rect 457 476 473 510
rect 507 476 523 510
rect 271 406 287 440
rect 321 424 337 440
rect 457 440 523 476
rect 457 424 473 440
rect 321 406 473 424
rect 507 406 523 440
rect 271 390 523 406
rect 625 580 708 596
rect 625 546 641 580
rect 675 546 708 580
rect 625 509 708 546
rect 625 475 641 509
rect 675 475 708 509
rect 625 438 708 475
rect 625 404 641 438
rect 675 404 708 438
rect 127 364 177 380
rect 17 226 51 364
rect 317 340 367 356
rect 85 314 283 330
rect 85 280 101 314
rect 135 280 206 314
rect 240 280 283 314
rect 351 306 367 340
rect 317 290 367 306
rect 409 340 551 356
rect 409 306 425 340
rect 459 306 551 340
rect 409 290 551 306
rect 249 256 283 280
rect 625 256 708 404
rect 249 251 708 256
rect 17 210 215 226
rect 249 222 658 251
rect 17 176 181 210
rect 456 221 658 222
rect 17 120 215 176
rect 17 87 181 120
rect 165 86 181 87
rect 165 69 215 86
rect 251 184 341 188
rect 251 150 291 184
rect 325 150 341 184
rect 456 187 472 221
rect 506 217 658 221
rect 692 217 708 251
rect 506 216 708 217
rect 506 187 522 216
rect 456 168 522 187
rect 251 116 341 150
rect 556 148 572 182
rect 606 148 643 182
rect 251 82 267 116
rect 301 82 341 116
rect 251 17 341 82
rect 409 114 455 134
rect 409 98 575 114
rect 409 64 525 98
rect 559 64 575 98
rect 409 51 575 64
rect 609 17 643 148
rect 677 98 743 134
rect 677 64 693 98
rect 727 64 743 98
rect 677 51 743 64
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a211o_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 1001478
string GDS_START 994456
<< end >>
