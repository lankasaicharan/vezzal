magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 332 1958 704
<< pwell >>
rect 1 228 527 272
rect 1465 228 1919 248
rect 1 184 820 228
rect 1009 184 1919 228
rect 1 49 1919 184
rect 0 0 1920 49
<< scpmos >>
rect 89 394 125 562
rect 199 394 235 562
rect 404 392 440 560
rect 528 392 564 592
rect 606 392 642 592
rect 714 504 750 588
rect 888 504 924 588
rect 1068 420 1104 588
rect 1158 420 1194 588
rect 1258 420 1294 588
rect 1362 420 1398 588
rect 1479 368 1515 592
rect 1569 368 1605 592
rect 1669 368 1705 592
rect 1779 368 1815 592
<< nmoslvt >>
rect 84 136 114 246
rect 202 98 232 246
rect 421 98 451 246
rect 636 74 666 202
rect 714 74 744 202
rect 809 74 839 158
rect 894 74 924 158
rect 1092 74 1122 202
rect 1178 74 1208 202
rect 1264 74 1294 202
rect 1350 74 1380 202
rect 1548 74 1578 222
rect 1634 74 1664 222
rect 1720 74 1750 222
rect 1806 74 1836 222
<< ndiff >>
rect 27 208 84 246
rect 27 174 39 208
rect 73 174 84 208
rect 27 136 84 174
rect 114 136 202 246
rect 129 98 202 136
rect 232 234 310 246
rect 232 200 253 234
rect 287 200 310 234
rect 232 98 310 200
rect 364 234 421 246
rect 364 200 376 234
rect 410 200 421 234
rect 364 98 421 200
rect 451 202 501 246
rect 451 98 636 202
rect 129 82 187 98
rect 129 48 141 82
rect 175 48 187 82
rect 466 82 636 98
rect 129 36 187 48
rect 466 48 478 82
rect 512 48 575 82
rect 609 74 636 82
rect 666 74 714 202
rect 744 158 794 202
rect 1035 188 1092 202
rect 744 130 809 158
rect 744 96 764 130
rect 798 96 809 130
rect 744 74 809 96
rect 839 74 894 158
rect 924 120 981 158
rect 924 86 935 120
rect 969 86 981 120
rect 924 74 981 86
rect 1035 154 1047 188
rect 1081 154 1092 188
rect 1035 116 1092 154
rect 1035 82 1047 116
rect 1081 82 1092 116
rect 1035 74 1092 82
rect 1122 179 1178 202
rect 1122 145 1133 179
rect 1167 145 1178 179
rect 1122 74 1178 145
rect 1208 190 1264 202
rect 1208 156 1219 190
rect 1253 156 1264 190
rect 1208 116 1264 156
rect 1208 82 1219 116
rect 1253 82 1264 116
rect 1208 74 1264 82
rect 1294 120 1350 202
rect 1294 86 1305 120
rect 1339 86 1350 120
rect 1294 74 1350 86
rect 1380 189 1437 202
rect 1380 155 1391 189
rect 1425 155 1437 189
rect 1380 121 1437 155
rect 1380 87 1391 121
rect 1425 87 1437 121
rect 1380 74 1437 87
rect 1491 190 1548 222
rect 1491 156 1503 190
rect 1537 156 1548 190
rect 1491 122 1548 156
rect 1491 88 1503 122
rect 1537 88 1548 122
rect 1491 74 1548 88
rect 1578 210 1634 222
rect 1578 176 1589 210
rect 1623 176 1634 210
rect 1578 122 1634 176
rect 1578 88 1589 122
rect 1623 88 1634 122
rect 1578 74 1634 88
rect 1664 142 1720 222
rect 1664 108 1675 142
rect 1709 108 1720 142
rect 1664 74 1720 108
rect 1750 210 1806 222
rect 1750 176 1761 210
rect 1795 176 1806 210
rect 1750 122 1806 176
rect 1750 88 1761 122
rect 1795 88 1806 122
rect 1750 74 1806 88
rect 1836 123 1893 222
rect 1836 89 1847 123
rect 1881 89 1893 123
rect 1836 74 1893 89
rect 609 48 621 74
rect 466 36 621 48
<< pdiff >>
rect 455 622 513 634
rect 455 588 467 622
rect 501 592 513 622
rect 501 588 528 592
rect 33 550 89 562
rect 33 516 45 550
rect 79 516 89 550
rect 33 440 89 516
rect 33 406 45 440
rect 79 406 89 440
rect 33 394 89 406
rect 125 550 199 562
rect 125 516 145 550
rect 179 516 199 550
rect 125 440 199 516
rect 125 406 145 440
rect 179 406 199 440
rect 125 394 199 406
rect 235 550 291 562
rect 455 560 528 588
rect 235 516 245 550
rect 279 516 291 550
rect 235 440 291 516
rect 235 406 245 440
rect 279 406 291 440
rect 235 394 291 406
rect 348 454 404 560
rect 348 420 360 454
rect 394 420 404 454
rect 348 392 404 420
rect 440 392 528 560
rect 564 392 606 592
rect 642 588 692 592
rect 1413 588 1479 592
rect 642 504 714 588
rect 750 504 888 588
rect 924 576 1068 588
rect 924 542 934 576
rect 968 542 1014 576
rect 1048 542 1068 576
rect 924 504 1068 542
rect 642 486 699 504
rect 642 452 652 486
rect 686 452 699 486
rect 642 392 699 452
rect 1018 420 1068 504
rect 1104 576 1158 588
rect 1104 542 1114 576
rect 1148 542 1158 576
rect 1104 466 1158 542
rect 1104 432 1114 466
rect 1148 432 1158 466
rect 1104 420 1158 432
rect 1194 576 1258 588
rect 1194 542 1214 576
rect 1248 542 1258 576
rect 1194 466 1258 542
rect 1194 432 1214 466
rect 1248 432 1258 466
rect 1194 420 1258 432
rect 1294 576 1362 588
rect 1294 542 1314 576
rect 1348 542 1362 576
rect 1294 466 1362 542
rect 1294 432 1314 466
rect 1348 432 1362 466
rect 1294 420 1362 432
rect 1398 576 1479 588
rect 1398 542 1425 576
rect 1459 542 1479 576
rect 1398 466 1479 542
rect 1398 432 1425 466
rect 1459 432 1479 466
rect 1398 420 1479 432
rect 1429 368 1479 420
rect 1515 580 1569 592
rect 1515 546 1525 580
rect 1559 546 1569 580
rect 1515 511 1569 546
rect 1515 477 1525 511
rect 1559 477 1569 511
rect 1515 442 1569 477
rect 1515 408 1525 442
rect 1559 408 1569 442
rect 1515 368 1569 408
rect 1605 580 1669 592
rect 1605 546 1625 580
rect 1659 546 1669 580
rect 1605 510 1669 546
rect 1605 476 1625 510
rect 1659 476 1669 510
rect 1605 368 1669 476
rect 1705 580 1779 592
rect 1705 546 1725 580
rect 1759 546 1779 580
rect 1705 497 1779 546
rect 1705 463 1725 497
rect 1759 463 1779 497
rect 1705 414 1779 463
rect 1705 380 1725 414
rect 1759 380 1779 414
rect 1705 368 1779 380
rect 1815 580 1871 592
rect 1815 546 1825 580
rect 1859 546 1871 580
rect 1815 478 1871 546
rect 1815 444 1825 478
rect 1859 444 1871 478
rect 1815 368 1871 444
<< ndiffc >>
rect 39 174 73 208
rect 253 200 287 234
rect 376 200 410 234
rect 141 48 175 82
rect 478 48 512 82
rect 575 48 609 82
rect 764 96 798 130
rect 935 86 969 120
rect 1047 154 1081 188
rect 1047 82 1081 116
rect 1133 145 1167 179
rect 1219 156 1253 190
rect 1219 82 1253 116
rect 1305 86 1339 120
rect 1391 155 1425 189
rect 1391 87 1425 121
rect 1503 156 1537 190
rect 1503 88 1537 122
rect 1589 176 1623 210
rect 1589 88 1623 122
rect 1675 108 1709 142
rect 1761 176 1795 210
rect 1761 88 1795 122
rect 1847 89 1881 123
<< pdiffc >>
rect 467 588 501 622
rect 45 516 79 550
rect 45 406 79 440
rect 145 516 179 550
rect 145 406 179 440
rect 245 516 279 550
rect 245 406 279 440
rect 360 420 394 454
rect 934 542 968 576
rect 1014 542 1048 576
rect 652 452 686 486
rect 1114 542 1148 576
rect 1114 432 1148 466
rect 1214 542 1248 576
rect 1214 432 1248 466
rect 1314 542 1348 576
rect 1314 432 1348 466
rect 1425 542 1459 576
rect 1425 432 1459 466
rect 1525 546 1559 580
rect 1525 477 1559 511
rect 1525 408 1559 442
rect 1625 546 1659 580
rect 1625 476 1659 510
rect 1725 546 1759 580
rect 1725 463 1759 497
rect 1725 380 1759 414
rect 1825 546 1859 580
rect 1825 444 1859 478
<< poly >>
rect 528 592 564 618
rect 606 592 642 618
rect 89 562 125 588
rect 199 562 235 588
rect 404 560 440 586
rect 89 356 125 394
rect 199 356 235 394
rect 714 588 750 614
rect 888 588 924 614
rect 1068 588 1104 614
rect 1158 588 1194 614
rect 1258 588 1294 614
rect 1362 588 1398 614
rect 1479 592 1515 618
rect 1569 592 1605 618
rect 1669 592 1705 618
rect 1779 592 1815 618
rect 714 472 750 504
rect 888 472 924 504
rect 714 456 840 472
rect 714 422 790 456
rect 824 422 840 456
rect 714 406 840 422
rect 888 456 954 472
rect 888 422 904 456
rect 938 422 954 456
rect 888 406 954 422
rect 84 340 151 356
rect 84 306 101 340
rect 135 306 151 340
rect 84 290 151 306
rect 193 340 259 356
rect 404 350 440 392
rect 193 306 209 340
rect 243 306 259 340
rect 193 290 259 306
rect 307 334 440 350
rect 528 334 564 392
rect 307 300 323 334
rect 357 314 440 334
rect 498 318 564 334
rect 357 300 451 314
rect 84 246 114 290
rect 202 246 232 290
rect 307 284 451 300
rect 421 246 451 284
rect 498 284 514 318
rect 548 284 564 318
rect 606 355 642 392
rect 606 339 672 355
rect 606 305 622 339
rect 656 305 672 339
rect 606 289 672 305
rect 498 268 564 284
rect 534 247 564 268
rect 84 110 114 136
rect 534 217 666 247
rect 636 202 666 217
rect 714 202 744 406
rect 894 347 930 406
rect 1068 358 1104 420
rect 1158 358 1194 420
rect 786 288 852 304
rect 786 254 802 288
rect 836 254 852 288
rect 786 238 852 254
rect 202 72 232 98
rect 421 72 451 98
rect 809 158 839 238
rect 894 158 924 347
rect 978 342 1194 358
rect 978 308 994 342
rect 1028 308 1194 342
rect 978 274 1194 308
rect 1258 318 1294 420
rect 1362 318 1398 420
rect 1258 290 1398 318
rect 1479 326 1515 368
rect 1569 326 1605 368
rect 1669 326 1705 368
rect 1779 326 1815 368
rect 1479 310 1815 326
rect 1479 296 1629 310
rect 978 240 994 274
rect 1028 254 1194 274
rect 1264 274 1398 290
rect 1028 240 1208 254
rect 978 224 1208 240
rect 1092 202 1122 224
rect 1178 202 1208 224
rect 1264 240 1280 274
rect 1314 240 1348 274
rect 1382 240 1398 274
rect 1264 224 1398 240
rect 1548 276 1629 296
rect 1663 276 1697 310
rect 1731 276 1765 310
rect 1799 290 1815 310
rect 1799 276 1836 290
rect 1548 260 1836 276
rect 1264 202 1294 224
rect 1350 202 1380 224
rect 1548 222 1578 260
rect 1634 222 1664 260
rect 1720 222 1750 260
rect 1806 222 1836 260
rect 636 48 666 74
rect 714 48 744 74
rect 809 48 839 74
rect 894 48 924 74
rect 1092 48 1122 74
rect 1178 48 1208 74
rect 1264 48 1294 74
rect 1350 48 1380 74
rect 1548 48 1578 74
rect 1634 48 1664 74
rect 1720 48 1750 74
rect 1806 48 1836 74
<< polycont >>
rect 790 422 824 456
rect 904 422 938 456
rect 101 306 135 340
rect 209 306 243 340
rect 323 300 357 334
rect 514 284 548 318
rect 622 305 656 339
rect 802 254 836 288
rect 994 308 1028 342
rect 994 240 1028 274
rect 1280 240 1314 274
rect 1348 240 1382 274
rect 1629 276 1663 310
rect 1697 276 1731 310
rect 1765 276 1799 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 17 550 95 566
rect 17 516 45 550
rect 79 516 95 550
rect 17 440 95 516
rect 17 406 45 440
rect 79 406 95 440
rect 17 390 95 406
rect 129 550 195 649
rect 451 622 517 649
rect 451 588 467 622
rect 501 588 517 622
rect 918 576 1064 649
rect 129 516 145 550
rect 179 516 195 550
rect 129 440 195 516
rect 129 406 145 440
rect 179 406 195 440
rect 129 390 195 406
rect 229 554 326 566
rect 229 550 840 554
rect 229 516 245 550
rect 279 520 840 550
rect 918 542 934 576
rect 968 542 1014 576
rect 1048 542 1064 576
rect 918 526 1064 542
rect 1098 576 1164 592
rect 1098 542 1114 576
rect 1148 542 1164 576
rect 279 516 326 520
rect 229 440 326 516
rect 229 406 245 440
rect 279 406 326 440
rect 229 390 326 406
rect 17 250 51 390
rect 85 340 161 356
rect 85 306 101 340
rect 135 306 161 340
rect 85 290 161 306
rect 195 340 258 356
rect 195 306 209 340
rect 243 306 258 340
rect 195 290 258 306
rect 292 350 326 390
rect 360 454 441 486
rect 394 420 441 454
rect 636 452 652 486
rect 686 452 740 486
rect 360 418 441 420
rect 360 384 672 418
rect 292 334 373 350
rect 292 300 323 334
rect 357 300 373 334
rect 292 284 373 300
rect 292 250 326 284
rect 407 250 441 384
rect 606 339 672 384
rect 17 208 89 250
rect 17 174 39 208
rect 73 174 89 208
rect 227 234 326 250
rect 227 200 253 234
rect 287 200 326 234
rect 360 234 441 250
rect 360 200 376 234
rect 410 200 441 234
rect 498 318 564 334
rect 498 284 514 318
rect 548 284 564 318
rect 17 166 89 174
rect 498 166 564 284
rect 606 305 622 339
rect 656 305 672 339
rect 706 372 740 452
rect 774 456 840 520
rect 1098 472 1164 542
rect 774 422 790 456
rect 824 422 840 456
rect 774 406 840 422
rect 888 466 1164 472
rect 888 456 1114 466
rect 888 422 904 456
rect 938 432 1114 456
rect 1148 432 1164 466
rect 938 422 1164 432
rect 888 406 1164 422
rect 1198 576 1264 649
rect 1198 542 1214 576
rect 1248 542 1264 576
rect 1198 466 1264 542
rect 1198 432 1214 466
rect 1248 432 1264 466
rect 1198 416 1264 432
rect 1298 576 1364 592
rect 1298 542 1314 576
rect 1348 542 1364 576
rect 1298 466 1364 542
rect 1298 432 1314 466
rect 1348 432 1364 466
rect 706 342 1044 372
rect 706 338 994 342
rect 606 304 672 305
rect 963 308 994 338
rect 1028 308 1044 342
rect 1098 358 1164 406
rect 1298 358 1364 432
rect 1409 576 1475 649
rect 1409 542 1425 576
rect 1459 542 1475 576
rect 1409 466 1475 542
rect 1409 432 1425 466
rect 1459 432 1475 466
rect 1409 416 1475 432
rect 1509 580 1575 596
rect 1509 546 1525 580
rect 1559 546 1575 580
rect 1509 511 1575 546
rect 1509 477 1525 511
rect 1559 477 1575 511
rect 1509 442 1575 477
rect 1609 580 1675 649
rect 1609 546 1625 580
rect 1659 546 1675 580
rect 1609 510 1675 546
rect 1609 476 1625 510
rect 1659 476 1675 510
rect 1609 460 1675 476
rect 1709 580 1775 596
rect 1709 546 1725 580
rect 1759 546 1775 580
rect 1709 497 1775 546
rect 1709 463 1725 497
rect 1759 463 1775 497
rect 1509 408 1525 442
rect 1559 426 1575 442
rect 1709 426 1775 463
rect 1809 580 1875 649
rect 1809 546 1825 580
rect 1859 546 1875 580
rect 1809 478 1875 546
rect 1809 444 1825 478
rect 1859 444 1875 478
rect 1809 428 1875 444
rect 1559 414 1775 426
rect 1559 408 1725 414
rect 1509 392 1725 408
rect 1709 380 1725 392
rect 1759 394 1775 414
rect 1759 380 1895 394
rect 1709 360 1895 380
rect 1098 326 1579 358
rect 1098 324 1815 326
rect 606 288 852 304
rect 606 254 802 288
rect 836 254 852 288
rect 606 238 852 254
rect 963 274 1044 308
rect 963 240 994 274
rect 1028 240 1044 274
rect 963 224 1044 240
rect 963 204 997 224
rect 17 132 564 166
rect 748 170 997 204
rect 1031 188 1097 190
rect 748 130 814 170
rect 1031 154 1047 188
rect 1081 154 1097 188
rect 125 82 191 98
rect 125 48 141 82
rect 175 48 191 82
rect 125 17 191 48
rect 462 82 625 98
rect 462 48 478 82
rect 512 48 575 82
rect 609 48 625 82
rect 748 96 764 130
rect 798 96 814 130
rect 748 80 814 96
rect 919 120 985 136
rect 919 86 935 120
rect 969 86 985 120
rect 462 17 625 48
rect 919 17 985 86
rect 1031 116 1097 154
rect 1133 179 1167 324
rect 1545 310 1815 324
rect 1264 274 1511 290
rect 1264 240 1280 274
rect 1314 240 1348 274
rect 1382 240 1511 274
rect 1545 276 1629 310
rect 1663 276 1697 310
rect 1731 276 1765 310
rect 1799 276 1815 310
rect 1545 260 1815 276
rect 1264 224 1511 240
rect 1849 226 1895 360
rect 1587 210 1895 226
rect 1133 119 1167 145
rect 1203 156 1219 190
rect 1253 189 1441 190
rect 1253 156 1391 189
rect 1203 155 1391 156
rect 1425 155 1441 189
rect 1203 154 1441 155
rect 1031 82 1047 116
rect 1081 85 1097 116
rect 1203 116 1253 154
rect 1389 121 1441 154
rect 1203 85 1219 116
rect 1081 82 1219 85
rect 1031 51 1253 82
rect 1289 86 1305 120
rect 1339 86 1355 120
rect 1289 17 1355 86
rect 1389 87 1391 121
rect 1425 87 1441 121
rect 1389 71 1441 87
rect 1487 156 1503 190
rect 1537 156 1553 190
rect 1487 122 1553 156
rect 1487 88 1503 122
rect 1537 88 1553 122
rect 1487 17 1553 88
rect 1587 176 1589 210
rect 1623 192 1761 210
rect 1623 176 1625 192
rect 1587 122 1625 176
rect 1759 176 1761 192
rect 1795 176 1895 210
rect 1759 160 1895 176
rect 1587 88 1589 122
rect 1623 88 1625 122
rect 1587 72 1625 88
rect 1659 142 1725 158
rect 1659 108 1675 142
rect 1709 108 1725 142
rect 1659 17 1725 108
rect 1759 122 1797 160
rect 1759 88 1761 122
rect 1795 88 1797 122
rect 1759 72 1797 88
rect 1831 123 1897 126
rect 1831 89 1847 123
rect 1881 89 1897 123
rect 1831 17 1897 89
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrtn_4
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1855 168 1889 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 1641100
string GDS_START 1627336
<< end >>
