magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 26 49 817 242
rect 0 0 864 49
<< scnmos >>
rect 105 48 135 216
rect 236 132 266 216
rect 330 132 360 216
rect 416 132 446 216
rect 488 132 518 216
rect 704 132 734 216
<< scpmoshvt >>
rect 105 367 135 619
rect 258 434 288 518
rect 330 434 360 518
rect 488 434 518 518
rect 596 434 626 518
rect 704 434 734 518
<< ndiff >>
rect 52 204 105 216
rect 52 170 60 204
rect 94 170 105 204
rect 52 101 105 170
rect 52 67 60 101
rect 94 67 105 101
rect 52 48 105 67
rect 135 164 236 216
rect 135 130 146 164
rect 180 132 236 164
rect 266 132 330 216
rect 360 191 416 216
rect 360 157 371 191
rect 405 157 416 191
rect 360 132 416 157
rect 446 132 488 216
rect 518 191 704 216
rect 518 157 581 191
rect 615 157 659 191
rect 693 157 704 191
rect 518 132 704 157
rect 734 191 791 216
rect 734 157 749 191
rect 783 157 791 191
rect 734 132 791 157
rect 180 130 188 132
rect 135 94 188 130
rect 135 60 146 94
rect 180 60 188 94
rect 135 48 188 60
<< pdiff >>
rect 52 599 105 619
rect 52 565 60 599
rect 94 565 105 599
rect 52 506 105 565
rect 52 472 60 506
rect 94 472 105 506
rect 52 413 105 472
rect 52 379 60 413
rect 94 379 105 413
rect 52 367 105 379
rect 135 607 188 619
rect 135 573 146 607
rect 180 573 188 607
rect 135 518 188 573
rect 135 505 258 518
rect 135 471 170 505
rect 204 471 258 505
rect 135 434 258 471
rect 288 434 330 518
rect 360 492 488 518
rect 360 458 420 492
rect 454 458 488 492
rect 360 434 488 458
rect 518 434 596 518
rect 626 510 704 518
rect 626 476 653 510
rect 687 476 704 510
rect 626 434 704 476
rect 734 498 787 518
rect 734 464 745 498
rect 779 464 787 498
rect 734 434 787 464
rect 135 413 188 434
rect 135 379 146 413
rect 180 379 188 413
rect 135 367 188 379
<< ndiffc >>
rect 60 170 94 204
rect 60 67 94 101
rect 146 130 180 164
rect 371 157 405 191
rect 581 157 615 191
rect 659 157 693 191
rect 749 157 783 191
rect 146 60 180 94
<< pdiffc >>
rect 60 565 94 599
rect 60 472 94 506
rect 60 379 94 413
rect 146 573 180 607
rect 170 471 204 505
rect 420 458 454 492
rect 653 476 687 510
rect 745 464 779 498
rect 146 379 180 413
<< poly >>
rect 105 619 135 645
rect 258 518 288 544
rect 330 518 360 544
rect 488 518 518 544
rect 596 518 626 544
rect 704 518 734 544
rect 258 402 288 434
rect 222 386 288 402
rect 105 304 135 367
rect 222 352 238 386
rect 272 352 288 386
rect 222 318 288 352
rect 105 288 180 304
rect 105 254 130 288
rect 164 254 180 288
rect 222 284 238 318
rect 272 284 288 318
rect 330 382 360 434
rect 488 402 518 434
rect 488 386 554 402
rect 330 366 446 382
rect 330 332 346 366
rect 380 332 446 366
rect 488 352 504 386
rect 538 352 554 386
rect 488 336 554 352
rect 330 316 446 332
rect 222 268 288 284
rect 105 238 180 254
rect 105 216 135 238
rect 236 216 266 268
rect 330 216 360 242
rect 416 216 446 316
rect 596 310 626 434
rect 704 402 734 434
rect 704 386 770 402
rect 704 352 720 386
rect 754 352 770 386
rect 704 336 770 352
rect 596 294 662 310
rect 596 274 612 294
rect 488 260 612 274
rect 646 260 662 294
rect 488 244 662 260
rect 488 216 518 244
rect 704 216 734 336
rect 236 106 266 132
rect 330 110 360 132
rect 308 94 374 110
rect 416 106 446 132
rect 488 106 518 132
rect 704 106 734 132
rect 308 60 324 94
rect 358 60 374 94
rect 105 22 135 48
rect 308 44 374 60
<< polycont >>
rect 238 352 272 386
rect 130 254 164 288
rect 238 284 272 318
rect 346 332 380 366
rect 504 352 538 386
rect 720 352 754 386
rect 612 260 646 294
rect 324 60 358 94
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 17 599 94 615
rect 17 565 60 599
rect 17 506 94 565
rect 17 472 60 506
rect 17 413 94 472
rect 17 379 60 413
rect 17 204 94 379
rect 142 607 204 649
rect 142 573 146 607
rect 180 573 204 607
rect 142 505 204 573
rect 142 471 170 505
rect 142 413 204 471
rect 142 379 146 413
rect 180 379 204 413
rect 142 363 204 379
rect 238 577 615 611
rect 238 386 272 577
rect 238 318 272 352
rect 17 170 60 204
rect 128 288 180 304
rect 128 254 130 288
rect 164 254 180 288
rect 306 366 380 516
rect 306 332 346 366
rect 306 298 380 332
rect 414 492 458 508
rect 414 458 420 492
rect 454 458 458 492
rect 238 268 272 284
rect 128 232 180 254
rect 414 232 458 458
rect 128 198 458 232
rect 492 386 547 523
rect 492 352 504 386
rect 538 352 547 386
rect 17 101 94 170
rect 355 191 421 198
rect 17 67 60 101
rect 17 51 94 67
rect 130 130 146 164
rect 180 130 196 164
rect 355 157 371 191
rect 405 157 421 191
rect 355 141 421 157
rect 130 94 196 130
rect 492 107 547 352
rect 581 426 615 577
rect 649 510 695 649
rect 649 476 653 510
rect 687 476 695 510
rect 649 460 695 476
rect 729 498 840 514
rect 729 464 745 498
rect 779 464 840 498
rect 729 460 840 464
rect 581 386 770 426
rect 581 352 720 386
rect 754 352 770 386
rect 581 344 770 352
rect 806 310 840 460
rect 596 294 840 310
rect 596 260 612 294
rect 646 276 840 294
rect 646 260 812 276
rect 596 244 812 260
rect 130 60 146 94
rect 180 60 196 94
rect 130 17 196 60
rect 308 94 547 107
rect 308 60 324 94
rect 358 60 547 94
rect 308 51 547 60
rect 581 191 699 207
rect 615 157 659 191
rect 693 157 699 191
rect 581 17 699 157
rect 733 191 812 244
rect 733 157 749 191
rect 783 157 812 191
rect 733 141 812 157
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1708760
string GDS_START 1700622
<< end >>
