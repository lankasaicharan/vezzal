magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 6 266 195 275
rect 6 248 311 266
rect 6 190 817 248
rect 6 49 853 190
rect 0 0 864 49
<< scpmos >>
rect 86 398 116 566
rect 196 398 226 566
rect 398 368 428 592
rect 516 368 546 592
rect 616 368 646 592
rect 726 368 756 592
<< nmoslvt >>
rect 89 139 119 249
rect 205 130 235 240
rect 405 74 435 222
rect 483 74 513 222
rect 597 74 627 222
rect 711 74 741 222
<< ndiff >>
rect 32 227 89 249
rect 32 193 44 227
rect 78 193 89 227
rect 32 172 89 193
rect 39 139 89 172
rect 119 240 169 249
rect 119 176 205 240
rect 119 142 146 176
rect 180 142 205 176
rect 119 139 205 142
rect 134 130 205 139
rect 235 188 285 240
rect 235 176 294 188
rect 235 142 247 176
rect 281 142 294 176
rect 235 130 294 142
rect 355 136 405 222
rect 348 122 405 136
rect 348 88 360 122
rect 394 88 405 122
rect 348 74 405 88
rect 435 74 483 222
rect 513 74 597 222
rect 627 74 711 222
rect 741 164 791 222
rect 741 136 827 164
rect 741 102 781 136
rect 815 102 827 136
rect 741 74 827 102
<< pdiff >>
rect 339 580 398 592
rect 27 554 86 566
rect 27 520 39 554
rect 73 520 86 554
rect 27 444 86 520
rect 27 410 39 444
rect 73 410 86 444
rect 27 398 86 410
rect 116 554 196 566
rect 116 520 139 554
rect 173 520 196 554
rect 116 444 196 520
rect 116 410 139 444
rect 173 410 196 444
rect 116 398 196 410
rect 226 554 285 566
rect 226 520 239 554
rect 273 520 285 554
rect 226 444 285 520
rect 226 410 239 444
rect 273 410 285 444
rect 226 398 285 410
rect 339 546 351 580
rect 385 546 398 580
rect 339 512 398 546
rect 339 478 351 512
rect 385 478 398 512
rect 339 368 398 478
rect 428 580 516 592
rect 428 546 460 580
rect 494 546 516 580
rect 428 368 516 546
rect 546 580 616 592
rect 546 546 569 580
rect 603 546 616 580
rect 546 497 616 546
rect 546 463 569 497
rect 603 463 616 497
rect 546 414 616 463
rect 546 380 569 414
rect 603 380 616 414
rect 546 368 616 380
rect 646 580 726 592
rect 646 546 669 580
rect 703 546 726 580
rect 646 508 726 546
rect 646 474 669 508
rect 703 474 726 508
rect 646 368 726 474
rect 756 580 815 592
rect 756 546 769 580
rect 803 546 815 580
rect 756 510 815 546
rect 756 476 769 510
rect 803 476 815 510
rect 756 440 815 476
rect 756 406 769 440
rect 803 406 815 440
rect 756 368 815 406
<< ndiffc >>
rect 44 193 78 227
rect 146 142 180 176
rect 247 142 281 176
rect 360 88 394 122
rect 781 102 815 136
<< pdiffc >>
rect 39 520 73 554
rect 39 410 73 444
rect 139 520 173 554
rect 139 410 173 444
rect 239 520 273 554
rect 239 410 273 444
rect 351 546 385 580
rect 351 478 385 512
rect 460 546 494 580
rect 569 546 603 580
rect 569 463 603 497
rect 569 380 603 414
rect 669 546 703 580
rect 669 474 703 508
rect 769 546 803 580
rect 769 476 803 510
rect 769 406 803 440
<< poly >>
rect 398 592 428 618
rect 516 592 546 618
rect 616 592 646 618
rect 726 592 756 618
rect 86 566 116 592
rect 196 566 226 592
rect 86 383 116 398
rect 196 383 226 398
rect 83 275 119 383
rect 193 360 229 383
rect 169 344 235 360
rect 398 353 428 368
rect 516 353 546 368
rect 616 353 646 368
rect 726 353 756 368
rect 169 310 185 344
rect 219 310 235 344
rect 395 310 431 353
rect 513 310 549 353
rect 613 310 649 353
rect 723 336 759 353
rect 711 320 777 336
rect 169 294 235 310
rect 89 249 119 275
rect 205 240 235 294
rect 337 294 435 310
rect 337 260 353 294
rect 387 260 435 294
rect 337 244 435 260
rect 89 117 119 139
rect 405 222 435 244
rect 483 294 549 310
rect 483 260 499 294
rect 533 260 549 294
rect 483 244 549 260
rect 597 294 663 310
rect 597 260 613 294
rect 647 260 663 294
rect 597 244 663 260
rect 711 286 727 320
rect 761 286 777 320
rect 711 270 777 286
rect 483 222 513 244
rect 597 222 627 244
rect 711 222 741 270
rect 30 101 119 117
rect 205 104 235 130
rect 30 67 46 101
rect 80 67 119 101
rect 30 51 119 67
rect 405 48 435 74
rect 483 48 513 74
rect 597 48 627 74
rect 711 48 741 74
<< polycont >>
rect 185 310 219 344
rect 353 260 387 294
rect 499 260 533 294
rect 613 260 647 294
rect 727 286 761 320
rect 46 67 80 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 554 89 570
rect 23 520 39 554
rect 73 520 89 554
rect 23 444 89 520
rect 23 410 39 444
rect 73 410 89 444
rect 23 394 89 410
rect 123 554 189 649
rect 335 580 401 596
rect 123 520 139 554
rect 173 520 189 554
rect 123 444 189 520
rect 123 410 139 444
rect 173 410 189 444
rect 123 394 189 410
rect 223 554 289 570
rect 223 520 239 554
rect 273 520 289 554
rect 223 444 289 520
rect 335 546 351 580
rect 385 546 401 580
rect 335 512 401 546
rect 435 580 519 649
rect 435 546 460 580
rect 494 546 519 580
rect 435 530 519 546
rect 553 580 619 596
rect 553 546 569 580
rect 603 546 619 580
rect 335 478 351 512
rect 385 496 401 512
rect 553 497 619 546
rect 553 496 569 497
rect 385 478 569 496
rect 335 463 569 478
rect 603 463 619 497
rect 335 462 619 463
rect 223 410 239 444
rect 273 428 289 444
rect 273 410 471 428
rect 223 394 471 410
rect 23 260 57 394
rect 121 344 263 360
rect 121 310 185 344
rect 219 310 263 344
rect 437 310 471 394
rect 505 424 619 462
rect 653 580 719 649
rect 653 546 669 580
rect 703 546 719 580
rect 653 508 719 546
rect 653 474 669 508
rect 703 474 719 508
rect 653 458 719 474
rect 753 580 845 596
rect 753 546 769 580
rect 803 546 845 580
rect 753 510 845 546
rect 753 476 769 510
rect 803 476 845 510
rect 753 440 845 476
rect 753 424 769 440
rect 505 414 769 424
rect 505 380 569 414
rect 603 406 769 414
rect 803 406 845 440
rect 603 390 845 406
rect 603 380 619 390
rect 505 364 619 380
rect 697 320 777 356
rect 121 294 263 310
rect 337 294 403 310
rect 337 260 353 294
rect 387 260 403 294
rect 23 227 403 260
rect 23 193 44 227
rect 78 226 403 227
rect 437 294 549 310
rect 437 260 499 294
rect 533 260 549 294
rect 437 244 549 260
rect 597 294 663 310
rect 597 260 613 294
rect 647 260 663 294
rect 697 286 727 320
rect 761 286 777 320
rect 697 270 777 286
rect 78 193 94 226
rect 23 168 94 193
rect 437 192 471 244
rect 130 176 196 192
rect 130 142 146 176
rect 180 142 196 176
rect 25 101 96 134
rect 25 67 46 101
rect 80 67 96 101
rect 25 51 96 67
rect 130 17 196 142
rect 230 176 471 192
rect 230 142 247 176
rect 281 158 471 176
rect 597 162 663 260
rect 811 236 845 390
rect 697 202 845 236
rect 281 142 298 158
rect 230 126 298 142
rect 697 124 731 202
rect 344 122 731 124
rect 344 88 360 122
rect 394 88 731 122
rect 344 70 731 88
rect 765 136 831 168
rect 765 102 781 136
rect 815 102 831 136
rect 765 17 831 102
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 nand4bb_1
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 3751750
string GDS_START 3744222
<< end >>
