magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 331 1958 704
<< pwell >>
rect 783 229 971 273
rect 1731 268 1919 273
rect 1430 229 1919 268
rect 214 192 1919 229
rect 1 49 1919 192
rect 0 0 1920 49
<< scnmos >>
rect 80 82 110 166
rect 293 119 323 203
rect 453 119 483 203
rect 539 119 569 203
rect 625 119 655 203
rect 697 119 727 203
rect 862 119 892 247
rect 967 119 997 203
rect 1075 119 1105 203
rect 1149 119 1179 203
rect 1287 75 1317 203
rect 1509 158 1539 242
rect 1618 74 1648 242
rect 1810 79 1840 247
<< scpmoshvt >>
rect 80 468 110 596
rect 270 463 300 591
rect 410 463 440 547
rect 496 463 526 547
rect 620 499 650 583
rect 722 463 752 547
rect 862 379 892 547
rect 1002 379 1032 547
rect 1107 379 1137 463
rect 1179 379 1209 463
rect 1287 379 1317 547
rect 1513 367 1543 495
rect 1618 367 1648 619
rect 1810 367 1840 619
<< ndiff >>
rect 809 203 862 247
rect 240 178 293 203
rect 27 130 80 166
rect 27 96 35 130
rect 69 96 80 130
rect 27 82 80 96
rect 110 140 167 166
rect 110 106 125 140
rect 159 106 167 140
rect 240 144 248 178
rect 282 144 293 178
rect 240 119 293 144
rect 323 179 453 203
rect 323 145 367 179
rect 401 145 453 179
rect 323 119 453 145
rect 483 177 539 203
rect 483 143 494 177
rect 528 143 539 177
rect 483 119 539 143
rect 569 177 625 203
rect 569 143 580 177
rect 614 143 625 177
rect 569 119 625 143
rect 655 119 697 203
rect 727 174 862 203
rect 727 140 738 174
rect 772 140 817 174
rect 851 140 862 174
rect 727 119 862 140
rect 892 235 945 247
rect 892 201 903 235
rect 937 203 945 235
rect 1456 204 1509 242
rect 937 201 967 203
rect 892 167 967 201
rect 892 133 903 167
rect 937 133 967 167
rect 892 119 967 133
rect 997 178 1075 203
rect 997 144 1018 178
rect 1052 144 1075 178
rect 997 119 1075 144
rect 1105 119 1149 203
rect 1179 189 1287 203
rect 1179 155 1226 189
rect 1260 155 1287 189
rect 1179 121 1287 155
rect 1179 119 1226 121
rect 110 82 167 106
rect 1218 87 1226 119
rect 1260 87 1287 121
rect 1218 75 1287 87
rect 1317 189 1370 203
rect 1317 155 1328 189
rect 1362 155 1370 189
rect 1456 170 1464 204
rect 1498 170 1509 204
rect 1456 158 1509 170
rect 1539 230 1618 242
rect 1539 196 1565 230
rect 1599 196 1618 230
rect 1539 158 1618 196
rect 1317 121 1370 155
rect 1317 87 1328 121
rect 1362 87 1370 121
rect 1317 75 1370 87
rect 1561 116 1618 158
rect 1561 82 1573 116
rect 1607 82 1618 116
rect 1561 74 1618 82
rect 1648 230 1701 242
rect 1648 196 1659 230
rect 1693 196 1701 230
rect 1648 121 1701 196
rect 1648 87 1659 121
rect 1693 87 1701 121
rect 1648 74 1701 87
rect 1757 235 1810 247
rect 1757 201 1765 235
rect 1799 201 1810 235
rect 1757 125 1810 201
rect 1757 91 1765 125
rect 1799 91 1810 125
rect 1757 79 1810 91
rect 1840 235 1893 247
rect 1840 201 1851 235
rect 1885 201 1893 235
rect 1840 125 1893 201
rect 1840 91 1851 125
rect 1885 91 1893 125
rect 1840 79 1893 91
<< pdiff >>
rect 27 584 80 596
rect 27 550 35 584
rect 69 550 80 584
rect 27 514 80 550
rect 27 480 35 514
rect 69 480 80 514
rect 27 468 80 480
rect 110 582 163 596
rect 110 548 121 582
rect 155 548 163 582
rect 110 514 163 548
rect 110 480 121 514
rect 155 480 163 514
rect 110 468 163 480
rect 217 577 270 591
rect 217 543 225 577
rect 259 543 270 577
rect 217 509 270 543
rect 217 475 225 509
rect 259 475 270 509
rect 217 463 270 475
rect 300 581 357 591
rect 797 587 847 599
rect 300 547 311 581
rect 345 547 357 581
rect 548 547 620 583
rect 300 463 410 547
rect 440 523 496 547
rect 440 489 451 523
rect 485 489 496 523
rect 440 463 496 489
rect 526 523 620 547
rect 526 489 556 523
rect 590 499 620 523
rect 650 547 700 583
rect 797 553 805 587
rect 839 553 847 587
rect 797 547 847 553
rect 1565 585 1618 619
rect 1565 551 1573 585
rect 1607 551 1618 585
rect 650 499 722 547
rect 590 489 598 499
rect 526 463 598 489
rect 672 463 722 499
rect 752 463 862 547
rect 797 379 862 463
rect 892 431 1002 547
rect 892 397 903 431
rect 937 397 1002 431
rect 892 379 1002 397
rect 1032 534 1085 547
rect 1032 500 1043 534
rect 1077 500 1085 534
rect 1032 463 1085 500
rect 1234 535 1287 547
rect 1234 501 1242 535
rect 1276 501 1287 535
rect 1234 463 1287 501
rect 1032 425 1107 463
rect 1032 391 1043 425
rect 1077 391 1107 425
rect 1032 379 1107 391
rect 1137 379 1179 463
rect 1209 430 1287 463
rect 1209 396 1232 430
rect 1266 396 1287 430
rect 1209 379 1287 396
rect 1317 535 1370 547
rect 1317 501 1328 535
rect 1362 501 1370 535
rect 1317 425 1370 501
rect 1565 495 1618 551
rect 1317 391 1328 425
rect 1362 391 1370 425
rect 1317 379 1370 391
rect 1460 425 1513 495
rect 1460 391 1468 425
rect 1502 391 1513 425
rect 1460 367 1513 391
rect 1543 367 1618 495
rect 1648 425 1701 619
rect 1648 391 1659 425
rect 1693 391 1701 425
rect 1648 367 1701 391
rect 1757 607 1810 619
rect 1757 573 1765 607
rect 1799 573 1810 607
rect 1757 367 1810 573
rect 1840 599 1893 619
rect 1840 565 1851 599
rect 1885 565 1893 599
rect 1840 504 1893 565
rect 1840 470 1851 504
rect 1885 470 1893 504
rect 1840 413 1893 470
rect 1840 379 1851 413
rect 1885 379 1893 413
rect 1840 367 1893 379
<< ndiffc >>
rect 35 96 69 130
rect 125 106 159 140
rect 248 144 282 178
rect 367 145 401 179
rect 494 143 528 177
rect 580 143 614 177
rect 738 140 772 174
rect 817 140 851 174
rect 903 201 937 235
rect 903 133 937 167
rect 1018 144 1052 178
rect 1226 155 1260 189
rect 1226 87 1260 121
rect 1328 155 1362 189
rect 1464 170 1498 204
rect 1565 196 1599 230
rect 1328 87 1362 121
rect 1573 82 1607 116
rect 1659 196 1693 230
rect 1659 87 1693 121
rect 1765 201 1799 235
rect 1765 91 1799 125
rect 1851 201 1885 235
rect 1851 91 1885 125
<< pdiffc >>
rect 35 550 69 584
rect 35 480 69 514
rect 121 548 155 582
rect 121 480 155 514
rect 225 543 259 577
rect 225 475 259 509
rect 311 547 345 581
rect 451 489 485 523
rect 556 489 590 523
rect 805 553 839 587
rect 1573 551 1607 585
rect 903 397 937 431
rect 1043 500 1077 534
rect 1242 501 1276 535
rect 1043 391 1077 425
rect 1232 396 1266 430
rect 1328 501 1362 535
rect 1328 391 1362 425
rect 1468 391 1502 425
rect 1659 391 1693 425
rect 1765 573 1799 607
rect 1851 565 1885 599
rect 1851 470 1885 504
rect 1851 379 1885 413
<< poly >>
rect 80 596 110 622
rect 270 615 1032 645
rect 1618 619 1648 645
rect 1810 619 1840 645
rect 270 591 300 615
rect 80 322 110 468
rect 620 583 650 615
rect 410 547 440 573
rect 496 547 526 573
rect 722 547 752 573
rect 862 547 892 573
rect 1002 547 1032 615
rect 1287 547 1317 573
rect 620 473 650 499
rect 35 306 110 322
rect 35 272 51 306
rect 85 272 110 306
rect 35 238 110 272
rect 158 361 224 377
rect 158 327 174 361
rect 208 327 224 361
rect 158 293 224 327
rect 158 259 174 293
rect 208 273 224 293
rect 270 273 300 463
rect 410 376 440 463
rect 365 360 440 376
rect 496 431 526 463
rect 722 431 752 463
rect 496 415 655 431
rect 496 381 605 415
rect 639 381 655 415
rect 496 365 655 381
rect 699 415 765 431
rect 699 381 715 415
rect 749 381 765 415
rect 699 365 765 381
rect 1107 463 1137 489
rect 1179 463 1209 489
rect 1513 495 1543 521
rect 365 326 381 360
rect 415 326 440 360
rect 365 292 440 326
rect 208 259 323 273
rect 158 243 323 259
rect 35 204 51 238
rect 85 204 110 238
rect 35 188 110 204
rect 293 203 323 243
rect 365 258 381 292
rect 415 272 440 292
rect 415 258 483 272
rect 365 242 483 258
rect 453 203 483 242
rect 539 203 569 229
rect 625 203 655 365
rect 735 291 765 365
rect 862 347 892 379
rect 1002 353 1032 379
rect 826 331 892 347
rect 1107 333 1137 379
rect 826 297 842 331
rect 876 297 892 331
rect 1077 311 1137 333
rect 697 275 775 291
rect 826 281 892 297
rect 697 241 725 275
rect 759 241 775 275
rect 862 247 892 281
rect 967 303 1137 311
rect 1179 347 1209 379
rect 1179 331 1245 347
rect 967 295 1107 303
rect 967 261 983 295
rect 1017 281 1107 295
rect 1179 297 1195 331
rect 1229 297 1245 331
rect 1179 281 1245 297
rect 1287 291 1317 379
rect 1513 330 1543 367
rect 1401 314 1543 330
rect 1017 261 1033 281
rect 697 225 775 241
rect 697 203 727 225
rect 80 166 110 188
rect 967 245 1033 261
rect 1179 255 1215 281
rect 967 203 997 245
rect 1075 203 1105 229
rect 1149 225 1215 255
rect 1287 275 1353 291
rect 1287 241 1303 275
rect 1337 241 1353 275
rect 1401 280 1417 314
rect 1451 300 1543 314
rect 1451 280 1539 300
rect 1401 264 1539 280
rect 1509 242 1539 264
rect 1618 242 1648 367
rect 1810 335 1840 367
rect 1744 319 1840 335
rect 1744 285 1760 319
rect 1794 285 1840 319
rect 1744 269 1840 285
rect 1810 247 1840 269
rect 1287 225 1353 241
rect 1149 203 1179 225
rect 1287 203 1317 225
rect 80 56 110 82
rect 293 51 323 119
rect 453 93 483 119
rect 539 51 569 119
rect 625 93 655 119
rect 697 93 727 119
rect 862 93 892 119
rect 967 93 997 119
rect 1075 51 1105 119
rect 1149 93 1179 119
rect 1509 132 1539 158
rect 1401 103 1467 119
rect 293 21 1105 51
rect 1287 49 1317 75
rect 1401 69 1417 103
rect 1451 69 1467 103
rect 1401 52 1467 69
rect 1618 52 1648 74
rect 1810 53 1840 79
rect 1401 22 1648 52
<< polycont >>
rect 51 272 85 306
rect 174 327 208 361
rect 174 259 208 293
rect 605 381 639 415
rect 715 381 749 415
rect 381 326 415 360
rect 51 204 85 238
rect 381 258 415 292
rect 842 297 876 331
rect 725 241 759 275
rect 983 261 1017 295
rect 1195 297 1229 331
rect 1303 241 1337 275
rect 1417 280 1451 314
rect 1760 285 1794 319
rect 1417 69 1451 103
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 19 584 78 649
rect 19 550 35 584
rect 69 550 78 584
rect 19 514 78 550
rect 19 480 35 514
rect 69 480 78 514
rect 19 464 78 480
rect 112 582 159 598
rect 112 548 121 582
rect 155 548 159 582
rect 112 514 159 548
rect 112 480 121 514
rect 155 480 159 514
rect 112 464 159 480
rect 17 306 85 430
rect 17 272 51 306
rect 17 238 85 272
rect 17 204 51 238
rect 17 168 85 204
rect 119 377 159 464
rect 209 577 265 593
rect 209 543 225 577
rect 259 543 265 577
rect 209 509 265 543
rect 299 581 347 649
rect 299 547 311 581
rect 345 547 347 581
rect 299 531 347 547
rect 381 573 660 615
rect 209 475 225 509
rect 259 497 265 509
rect 381 497 415 573
rect 259 475 415 497
rect 209 463 415 475
rect 449 523 487 539
rect 449 489 451 523
rect 485 489 487 523
rect 209 459 284 463
rect 119 361 208 377
rect 119 327 174 361
rect 119 293 208 327
rect 119 259 174 293
rect 119 243 208 259
rect 119 140 175 243
rect 19 130 85 134
rect 19 96 35 130
rect 69 96 85 130
rect 19 17 85 96
rect 119 106 125 140
rect 159 106 175 140
rect 242 178 284 459
rect 318 360 415 429
rect 318 326 381 360
rect 318 292 415 326
rect 318 258 381 292
rect 318 242 415 258
rect 242 144 248 178
rect 282 144 284 178
rect 242 128 284 144
rect 351 179 415 195
rect 351 145 367 179
rect 401 145 415 179
rect 119 90 175 106
rect 351 17 415 145
rect 449 193 487 489
rect 521 523 592 539
rect 521 489 556 523
rect 590 489 592 523
rect 521 473 592 489
rect 626 517 660 573
rect 789 587 855 649
rect 789 553 805 587
rect 839 553 855 587
rect 1041 534 1093 550
rect 626 483 1007 517
rect 521 345 555 473
rect 626 431 660 483
rect 589 415 660 431
rect 589 381 605 415
rect 639 381 660 415
rect 589 379 660 381
rect 699 431 939 447
rect 699 415 903 431
rect 699 381 715 415
rect 749 397 903 415
rect 937 397 939 431
rect 749 381 939 397
rect 699 379 939 381
rect 521 331 892 345
rect 521 311 842 331
rect 449 177 539 193
rect 449 143 494 177
rect 528 143 539 177
rect 449 127 539 143
rect 573 177 632 311
rect 826 297 842 311
rect 876 297 892 331
rect 826 285 892 297
rect 973 311 1007 483
rect 1041 500 1043 534
rect 1077 500 1093 534
rect 1041 425 1093 500
rect 1041 391 1043 425
rect 1077 391 1093 425
rect 1216 535 1282 649
rect 1557 585 1623 649
rect 1557 551 1573 585
rect 1607 551 1623 585
rect 1761 607 1803 649
rect 1761 573 1765 607
rect 1799 573 1803 607
rect 1761 557 1803 573
rect 1847 599 1901 615
rect 1847 565 1851 599
rect 1885 565 1901 599
rect 1216 501 1242 535
rect 1276 501 1282 535
rect 1216 430 1282 501
rect 1216 396 1232 430
rect 1266 396 1282 430
rect 1216 395 1282 396
rect 1316 535 1375 551
rect 1557 543 1623 551
rect 1316 501 1328 535
rect 1362 509 1375 535
rect 1362 501 1810 509
rect 1316 475 1810 501
rect 1316 425 1407 475
rect 1041 375 1093 391
rect 973 295 1019 311
rect 709 275 775 277
rect 709 241 725 275
rect 759 251 775 275
rect 973 261 983 295
rect 1017 261 1019 295
rect 759 241 939 251
rect 973 245 1019 261
rect 1053 259 1093 375
rect 1316 391 1328 425
rect 1362 391 1407 425
rect 1316 361 1407 391
rect 1452 425 1521 441
rect 1452 391 1468 425
rect 1502 391 1521 425
rect 1452 375 1521 391
rect 1179 331 1407 361
rect 1179 297 1195 331
rect 1229 330 1407 331
rect 1229 327 1453 330
rect 1229 297 1245 327
rect 1373 314 1453 327
rect 1287 275 1337 291
rect 1287 259 1303 275
rect 709 235 939 241
rect 709 217 903 235
rect 901 201 903 217
rect 937 201 939 235
rect 573 143 580 177
rect 614 143 632 177
rect 573 127 632 143
rect 722 174 867 183
rect 722 140 738 174
rect 772 140 817 174
rect 851 140 867 174
rect 722 17 867 140
rect 901 167 939 201
rect 1053 241 1303 259
rect 1053 225 1337 241
rect 1373 280 1417 314
rect 1451 280 1453 314
rect 1373 264 1453 280
rect 1053 199 1087 225
rect 901 133 903 167
rect 937 133 939 167
rect 901 117 939 133
rect 1002 178 1087 199
rect 1373 191 1407 264
rect 1487 208 1521 375
rect 1651 425 1709 441
rect 1651 391 1659 425
rect 1693 391 1709 425
rect 1002 144 1018 178
rect 1052 144 1087 178
rect 1002 128 1087 144
rect 1210 189 1276 191
rect 1210 155 1226 189
rect 1260 155 1276 189
rect 1210 121 1276 155
rect 1210 87 1226 121
rect 1260 87 1276 121
rect 1210 17 1276 87
rect 1310 189 1407 191
rect 1310 155 1328 189
rect 1362 155 1407 189
rect 1443 204 1521 208
rect 1443 170 1464 204
rect 1498 170 1521 204
rect 1443 166 1521 170
rect 1555 230 1617 246
rect 1555 196 1565 230
rect 1599 196 1617 230
rect 1310 121 1378 155
rect 1310 87 1328 121
rect 1362 87 1378 121
rect 1443 119 1477 166
rect 1310 71 1378 87
rect 1412 103 1477 119
rect 1412 69 1417 103
rect 1451 69 1477 103
rect 1412 53 1477 69
rect 1555 116 1617 196
rect 1555 82 1573 116
rect 1607 82 1617 116
rect 1555 17 1617 82
rect 1651 230 1709 391
rect 1744 319 1810 475
rect 1744 285 1760 319
rect 1794 285 1810 319
rect 1847 504 1901 565
rect 1847 470 1851 504
rect 1885 470 1901 504
rect 1847 413 1901 470
rect 1847 379 1851 413
rect 1885 379 1901 413
rect 1651 196 1659 230
rect 1693 196 1709 230
rect 1651 121 1709 196
rect 1651 87 1659 121
rect 1693 87 1709 121
rect 1651 71 1709 87
rect 1749 235 1803 251
rect 1749 201 1765 235
rect 1799 201 1803 235
rect 1749 125 1803 201
rect 1749 91 1765 125
rect 1799 91 1803 125
rect 1749 17 1803 91
rect 1847 235 1901 379
rect 1847 201 1851 235
rect 1885 201 1901 235
rect 1847 125 1901 201
rect 1847 91 1851 125
rect 1885 91 1901 125
rect 1847 75 1901 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfxbp_1
flabel comment s 746 335 746 335 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 1663 168 1697 202 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1663 390 1697 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1855 94 1889 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1855 168 1889 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1855 390 1889 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1855 464 1889 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1855 538 1889 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2378898
string GDS_START 2363712
<< end >>
