magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 245 381 248
rect 1 49 765 245
rect 0 0 768 49
<< scnmos >>
rect 84 54 114 222
rect 251 138 281 222
rect 464 51 494 219
rect 550 51 580 219
rect 656 51 686 219
<< scpmoshvt >>
rect 124 367 154 619
rect 251 367 281 451
rect 464 367 494 619
rect 554 367 584 619
rect 656 367 686 619
<< ndiff >>
rect 27 212 84 222
rect 27 178 39 212
rect 73 178 84 212
rect 27 101 84 178
rect 27 67 39 101
rect 73 67 84 101
rect 27 54 84 67
rect 114 138 251 222
rect 281 210 355 222
rect 281 176 313 210
rect 347 176 355 210
rect 281 138 355 176
rect 411 207 464 219
rect 411 173 419 207
rect 453 173 464 207
rect 114 131 175 138
rect 114 97 128 131
rect 162 97 175 131
rect 114 54 175 97
rect 411 103 464 173
rect 411 69 419 103
rect 453 69 464 103
rect 411 51 464 69
rect 494 207 550 219
rect 494 173 505 207
rect 539 173 550 207
rect 494 103 550 173
rect 494 69 505 103
rect 539 69 550 103
rect 494 51 550 69
rect 580 173 656 219
rect 580 139 597 173
rect 631 139 656 173
rect 580 97 656 139
rect 580 63 597 97
rect 631 63 656 97
rect 580 51 656 63
rect 686 207 739 219
rect 686 173 697 207
rect 731 173 739 207
rect 686 97 739 173
rect 686 63 697 97
rect 731 63 739 97
rect 686 51 739 63
<< pdiff >>
rect 71 599 124 619
rect 71 565 79 599
rect 113 565 124 599
rect 71 508 124 565
rect 71 474 79 508
rect 113 474 124 508
rect 71 413 124 474
rect 71 379 79 413
rect 113 379 124 413
rect 71 367 124 379
rect 154 607 207 619
rect 154 573 165 607
rect 199 573 207 607
rect 154 517 207 573
rect 154 483 165 517
rect 199 483 207 517
rect 154 451 207 483
rect 411 607 464 619
rect 411 573 419 607
rect 453 573 464 607
rect 411 493 464 573
rect 411 459 419 493
rect 453 459 464 493
rect 154 419 251 451
rect 154 385 186 419
rect 220 385 251 419
rect 154 367 251 385
rect 281 426 347 451
rect 281 392 301 426
rect 335 392 347 426
rect 281 367 347 392
rect 411 367 464 459
rect 494 599 554 619
rect 494 565 509 599
rect 543 565 554 599
rect 494 504 554 565
rect 494 470 509 504
rect 543 470 554 504
rect 494 419 554 470
rect 494 385 509 419
rect 543 385 554 419
rect 494 367 554 385
rect 584 367 656 619
rect 686 607 739 619
rect 686 573 697 607
rect 731 573 739 607
rect 686 512 739 573
rect 686 478 697 512
rect 731 478 739 512
rect 686 418 739 478
rect 686 384 697 418
rect 731 384 739 418
rect 686 367 739 384
<< ndiffc >>
rect 39 178 73 212
rect 39 67 73 101
rect 313 176 347 210
rect 419 173 453 207
rect 128 97 162 131
rect 419 69 453 103
rect 505 173 539 207
rect 505 69 539 103
rect 597 139 631 173
rect 597 63 631 97
rect 697 173 731 207
rect 697 63 731 97
<< pdiffc >>
rect 79 565 113 599
rect 79 474 113 508
rect 79 379 113 413
rect 165 573 199 607
rect 165 483 199 517
rect 419 573 453 607
rect 419 459 453 493
rect 186 385 220 419
rect 301 392 335 426
rect 509 565 543 599
rect 509 470 543 504
rect 509 385 543 419
rect 697 573 731 607
rect 697 478 731 512
rect 697 384 731 418
<< poly >>
rect 124 619 154 645
rect 464 619 494 645
rect 554 619 584 645
rect 656 619 686 645
rect 251 451 281 477
rect 124 310 154 367
rect 251 310 281 367
rect 464 310 494 367
rect 554 335 584 367
rect 84 294 163 310
rect 84 260 113 294
rect 147 260 163 294
rect 84 244 163 260
rect 211 294 281 310
rect 211 260 227 294
rect 261 260 281 294
rect 211 244 281 260
rect 329 294 494 310
rect 329 260 345 294
rect 379 260 494 294
rect 542 319 608 335
rect 542 285 558 319
rect 592 285 608 319
rect 542 269 608 285
rect 656 325 686 367
rect 656 309 743 325
rect 656 275 693 309
rect 727 275 743 309
rect 329 244 494 260
rect 84 222 114 244
rect 251 222 281 244
rect 464 219 494 244
rect 550 219 580 269
rect 656 259 743 275
rect 656 219 686 259
rect 251 112 281 138
rect 84 28 114 54
rect 464 25 494 51
rect 550 25 580 51
rect 656 25 686 51
<< polycont >>
rect 113 260 147 294
rect 227 260 261 294
rect 345 260 379 294
rect 558 285 592 319
rect 693 275 727 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 599 115 615
rect 17 565 79 599
rect 113 565 115 599
rect 17 508 115 565
rect 17 474 79 508
rect 113 474 115 508
rect 17 413 115 474
rect 17 379 79 413
rect 113 379 115 413
rect 149 607 251 649
rect 149 573 165 607
rect 199 573 251 607
rect 149 517 251 573
rect 149 483 165 517
rect 199 483 251 517
rect 149 419 251 483
rect 403 607 469 649
rect 403 573 419 607
rect 453 573 469 607
rect 403 493 469 573
rect 403 459 419 493
rect 453 459 469 493
rect 403 454 469 459
rect 505 599 559 615
rect 505 565 509 599
rect 543 565 559 599
rect 505 504 559 565
rect 505 470 509 504
rect 543 470 559 504
rect 149 385 186 419
rect 220 385 251 419
rect 285 426 351 442
rect 285 392 301 426
rect 335 392 351 426
rect 505 420 559 470
rect 285 385 351 392
rect 17 363 115 379
rect 17 212 77 363
rect 113 294 187 310
rect 147 260 187 294
rect 113 244 187 260
rect 17 178 39 212
rect 73 178 77 212
rect 17 101 77 178
rect 153 208 187 244
rect 221 294 261 350
rect 221 260 227 294
rect 221 242 261 260
rect 295 310 351 385
rect 415 419 559 420
rect 415 385 509 419
rect 543 385 559 419
rect 681 607 747 649
rect 681 573 697 607
rect 731 573 747 607
rect 681 512 747 573
rect 681 478 697 512
rect 731 478 747 512
rect 681 418 747 478
rect 295 294 381 310
rect 295 260 345 294
rect 379 260 381 294
rect 295 210 381 260
rect 153 174 261 208
rect 17 67 39 101
rect 73 67 77 101
rect 17 51 77 67
rect 111 131 183 140
rect 111 97 128 131
rect 162 97 183 131
rect 111 17 183 97
rect 227 85 261 174
rect 295 176 313 210
rect 347 176 381 210
rect 295 172 381 176
rect 415 207 462 385
rect 681 384 697 418
rect 731 384 747 418
rect 496 319 643 350
rect 496 285 558 319
rect 592 285 643 319
rect 677 309 751 350
rect 677 275 693 309
rect 727 275 751 309
rect 415 173 419 207
rect 453 173 462 207
rect 415 103 462 173
rect 415 85 419 103
rect 227 69 419 85
rect 453 69 462 103
rect 227 51 462 69
rect 496 207 747 241
rect 496 173 505 207
rect 539 173 543 207
rect 681 173 697 207
rect 731 173 747 207
rect 496 103 543 173
rect 496 69 505 103
rect 539 69 543 103
rect 496 51 543 69
rect 581 139 597 173
rect 631 139 647 173
rect 581 97 647 139
rect 581 63 597 97
rect 631 63 647 97
rect 581 17 647 63
rect 681 97 747 173
rect 681 63 697 97
rect 731 63 747 97
rect 681 51 747 63
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21ba_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6526466
string GDS_START 6518840
<< end >>
