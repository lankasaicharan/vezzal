magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 79 49 1129 243
rect 0 0 1152 49
<< scnmos >>
rect 158 49 188 217
rect 244 49 274 217
rect 330 49 360 217
rect 416 49 446 217
rect 582 49 612 217
rect 668 49 698 217
rect 762 49 792 217
rect 848 49 878 217
rect 934 49 964 217
rect 1020 49 1050 217
<< scpmoshvt >>
rect 134 367 164 619
rect 220 367 250 619
rect 306 367 336 619
rect 392 367 422 619
rect 582 367 612 619
rect 668 367 698 619
rect 754 367 784 619
rect 848 367 878 619
rect 934 367 964 619
rect 1020 367 1050 619
<< ndiff >>
rect 105 181 158 217
rect 105 147 113 181
rect 147 147 158 181
rect 105 95 158 147
rect 105 61 113 95
rect 147 61 158 95
rect 105 49 158 61
rect 188 205 244 217
rect 188 171 199 205
rect 233 171 244 205
rect 188 101 244 171
rect 188 67 199 101
rect 233 67 244 101
rect 188 49 244 67
rect 274 181 330 217
rect 274 147 285 181
rect 319 147 330 181
rect 274 95 330 147
rect 274 61 285 95
rect 319 61 330 95
rect 274 49 330 61
rect 360 205 416 217
rect 360 171 371 205
rect 405 171 416 205
rect 360 101 416 171
rect 360 67 371 101
rect 405 67 416 101
rect 360 49 416 67
rect 446 124 582 217
rect 446 90 457 124
rect 491 90 537 124
rect 571 90 582 124
rect 446 49 582 90
rect 612 190 668 217
rect 612 156 623 190
rect 657 156 668 190
rect 612 101 668 156
rect 612 67 623 101
rect 657 67 668 101
rect 612 49 668 67
rect 698 122 762 217
rect 698 88 713 122
rect 747 88 762 122
rect 698 49 762 88
rect 792 122 848 217
rect 792 88 803 122
rect 837 88 848 122
rect 792 49 848 88
rect 878 171 934 217
rect 878 137 889 171
rect 923 137 934 171
rect 878 49 934 137
rect 964 205 1020 217
rect 964 171 975 205
rect 1009 171 1020 205
rect 964 101 1020 171
rect 964 67 975 101
rect 1009 67 1020 101
rect 964 49 1020 67
rect 1050 205 1103 217
rect 1050 171 1061 205
rect 1095 171 1103 205
rect 1050 95 1103 171
rect 1050 61 1061 95
rect 1095 61 1103 95
rect 1050 49 1103 61
<< pdiff >>
rect 81 607 134 619
rect 81 573 89 607
rect 123 573 134 607
rect 81 537 134 573
rect 81 503 89 537
rect 123 503 134 537
rect 81 465 134 503
rect 81 431 89 465
rect 123 431 134 465
rect 81 367 134 431
rect 164 599 220 619
rect 164 565 175 599
rect 209 565 220 599
rect 164 507 220 565
rect 164 473 175 507
rect 209 473 220 507
rect 164 413 220 473
rect 164 379 175 413
rect 209 379 220 413
rect 164 367 220 379
rect 250 607 306 619
rect 250 573 261 607
rect 295 573 306 607
rect 250 537 306 573
rect 250 503 261 537
rect 295 503 306 537
rect 250 465 306 503
rect 250 431 261 465
rect 295 431 306 465
rect 250 367 306 431
rect 336 599 392 619
rect 336 565 347 599
rect 381 565 392 599
rect 336 507 392 565
rect 336 473 347 507
rect 381 473 392 507
rect 336 413 392 473
rect 336 379 347 413
rect 381 379 392 413
rect 336 367 392 379
rect 422 607 475 619
rect 422 573 433 607
rect 467 573 475 607
rect 422 509 475 573
rect 422 475 433 509
rect 467 475 475 509
rect 422 413 475 475
rect 422 379 433 413
rect 467 379 475 413
rect 422 367 475 379
rect 529 607 582 619
rect 529 573 537 607
rect 571 573 582 607
rect 529 524 582 573
rect 529 490 537 524
rect 571 490 582 524
rect 529 436 582 490
rect 529 402 537 436
rect 571 402 582 436
rect 529 367 582 402
rect 612 547 668 619
rect 612 513 623 547
rect 657 513 668 547
rect 612 479 668 513
rect 612 445 623 479
rect 657 445 668 479
rect 612 411 668 445
rect 612 377 623 411
rect 657 377 668 411
rect 612 367 668 377
rect 698 599 754 619
rect 698 565 709 599
rect 743 565 754 599
rect 698 507 754 565
rect 698 473 709 507
rect 743 473 754 507
rect 698 413 754 473
rect 698 379 709 413
rect 743 379 754 413
rect 698 367 754 379
rect 784 578 848 619
rect 784 544 799 578
rect 833 544 848 578
rect 784 367 848 544
rect 878 599 934 619
rect 878 565 889 599
rect 923 565 934 599
rect 878 510 934 565
rect 878 476 889 510
rect 923 476 934 510
rect 878 367 934 476
rect 964 578 1020 619
rect 964 544 975 578
rect 1009 544 1020 578
rect 964 367 1020 544
rect 1050 599 1103 619
rect 1050 565 1061 599
rect 1095 565 1103 599
rect 1050 507 1103 565
rect 1050 473 1061 507
rect 1095 473 1103 507
rect 1050 413 1103 473
rect 1050 379 1061 413
rect 1095 379 1103 413
rect 1050 367 1103 379
<< ndiffc >>
rect 113 147 147 181
rect 113 61 147 95
rect 199 171 233 205
rect 199 67 233 101
rect 285 147 319 181
rect 285 61 319 95
rect 371 171 405 205
rect 371 67 405 101
rect 457 90 491 124
rect 537 90 571 124
rect 623 156 657 190
rect 623 67 657 101
rect 713 88 747 122
rect 803 88 837 122
rect 889 137 923 171
rect 975 171 1009 205
rect 975 67 1009 101
rect 1061 171 1095 205
rect 1061 61 1095 95
<< pdiffc >>
rect 89 573 123 607
rect 89 503 123 537
rect 89 431 123 465
rect 175 565 209 599
rect 175 473 209 507
rect 175 379 209 413
rect 261 573 295 607
rect 261 503 295 537
rect 261 431 295 465
rect 347 565 381 599
rect 347 473 381 507
rect 347 379 381 413
rect 433 573 467 607
rect 433 475 467 509
rect 433 379 467 413
rect 537 573 571 607
rect 537 490 571 524
rect 537 402 571 436
rect 623 513 657 547
rect 623 445 657 479
rect 623 377 657 411
rect 709 565 743 599
rect 709 473 743 507
rect 709 379 743 413
rect 799 544 833 578
rect 889 565 923 599
rect 889 476 923 510
rect 975 544 1009 578
rect 1061 565 1095 599
rect 1061 473 1095 507
rect 1061 379 1095 413
<< poly >>
rect 134 619 164 645
rect 220 619 250 645
rect 306 619 336 645
rect 392 619 422 645
rect 582 619 612 645
rect 668 619 698 645
rect 754 619 784 645
rect 848 619 878 645
rect 934 619 964 645
rect 1020 619 1050 645
rect 134 335 164 367
rect 220 335 250 367
rect 306 335 336 367
rect 392 335 422 367
rect 134 319 467 335
rect 134 285 213 319
rect 247 285 281 319
rect 315 285 349 319
rect 383 285 417 319
rect 451 285 467 319
rect 582 308 612 367
rect 134 269 467 285
rect 537 292 612 308
rect 158 217 188 269
rect 244 217 274 269
rect 330 217 360 269
rect 416 217 446 269
rect 537 258 553 292
rect 587 272 612 292
rect 668 272 698 367
rect 754 325 784 367
rect 587 258 698 272
rect 740 309 806 325
rect 740 275 756 309
rect 790 275 806 309
rect 740 259 806 275
rect 848 305 878 367
rect 934 305 964 367
rect 848 289 964 305
rect 537 242 698 258
rect 582 217 612 242
rect 668 217 698 242
rect 762 217 792 259
rect 848 255 869 289
rect 903 255 964 289
rect 848 239 964 255
rect 848 217 878 239
rect 934 217 964 239
rect 1020 335 1050 367
rect 1020 319 1086 335
rect 1020 285 1036 319
rect 1070 285 1086 319
rect 1020 269 1086 285
rect 1020 217 1050 269
rect 158 23 188 49
rect 244 23 274 49
rect 330 23 360 49
rect 416 23 446 49
rect 582 23 612 49
rect 668 23 698 49
rect 762 23 792 49
rect 848 23 878 49
rect 934 23 964 49
rect 1020 23 1050 49
<< polycont >>
rect 213 285 247 319
rect 281 285 315 319
rect 349 285 383 319
rect 417 285 451 319
rect 553 258 587 292
rect 756 275 790 309
rect 869 255 903 289
rect 1036 285 1070 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 73 607 139 649
rect 73 573 89 607
rect 123 573 139 607
rect 73 537 139 573
rect 73 503 89 537
rect 123 503 139 537
rect 73 465 139 503
rect 73 431 89 465
rect 123 431 139 465
rect 173 599 211 615
rect 173 565 175 599
rect 209 565 211 599
rect 173 507 211 565
rect 173 473 175 507
rect 209 473 211 507
rect 173 413 211 473
rect 245 607 311 649
rect 245 573 261 607
rect 295 573 311 607
rect 245 537 311 573
rect 245 503 261 537
rect 295 503 311 537
rect 245 465 311 503
rect 245 431 261 465
rect 295 431 311 465
rect 345 599 383 615
rect 345 565 347 599
rect 381 565 383 599
rect 345 507 383 565
rect 345 473 347 507
rect 381 473 383 507
rect 173 397 175 413
rect 31 379 175 397
rect 209 397 211 413
rect 345 413 383 473
rect 345 397 347 413
rect 209 379 347 397
rect 381 379 383 413
rect 31 356 383 379
rect 417 607 477 649
rect 417 573 433 607
rect 467 573 477 607
rect 417 509 477 573
rect 417 475 433 509
rect 467 475 477 509
rect 417 413 477 475
rect 417 379 433 413
rect 467 379 477 413
rect 521 607 747 615
rect 521 573 537 607
rect 571 599 747 607
rect 571 581 709 599
rect 571 573 573 581
rect 521 524 573 573
rect 707 565 709 581
rect 743 565 747 599
rect 521 490 537 524
rect 571 490 573 524
rect 521 436 573 490
rect 521 402 537 436
rect 571 402 573 436
rect 521 386 573 402
rect 607 513 623 547
rect 657 513 673 547
rect 607 479 673 513
rect 607 445 623 479
rect 657 445 673 479
rect 607 411 673 445
rect 607 382 623 411
rect 417 363 477 379
rect 621 377 623 382
rect 657 377 673 411
rect 31 249 161 356
rect 197 319 475 322
rect 197 285 213 319
rect 247 285 281 319
rect 315 285 349 319
rect 383 285 417 319
rect 451 285 475 319
rect 197 283 475 285
rect 31 215 407 249
rect 197 205 235 215
rect 97 147 113 181
rect 147 147 163 181
rect 97 95 163 147
rect 97 61 113 95
rect 147 61 163 95
rect 97 17 163 61
rect 197 171 199 205
rect 233 171 235 205
rect 369 205 407 215
rect 197 101 235 171
rect 197 67 199 101
rect 233 67 235 101
rect 197 51 235 67
rect 269 147 285 181
rect 319 147 335 181
rect 269 95 335 147
rect 269 61 285 95
rect 319 61 335 95
rect 269 17 335 61
rect 369 171 371 205
rect 405 171 407 205
rect 441 208 475 283
rect 511 292 587 352
rect 511 258 553 292
rect 511 242 587 258
rect 621 208 673 377
rect 707 507 747 565
rect 783 578 849 649
rect 783 544 799 578
rect 833 544 849 578
rect 783 528 849 544
rect 883 599 925 615
rect 883 565 889 599
rect 923 565 925 599
rect 707 473 709 507
rect 743 494 747 507
rect 883 510 925 565
rect 959 578 1025 649
rect 959 544 975 578
rect 1009 544 1025 578
rect 959 528 1025 544
rect 1059 599 1099 615
rect 1059 565 1061 599
rect 1095 565 1099 599
rect 883 494 889 510
rect 743 476 889 494
rect 923 494 925 510
rect 1059 507 1099 565
rect 1059 494 1061 507
rect 923 476 1061 494
rect 743 473 1061 476
rect 1095 473 1099 507
rect 707 460 1099 473
rect 707 413 749 460
rect 707 379 709 413
rect 743 379 749 413
rect 707 363 749 379
rect 783 390 1025 424
rect 783 325 817 390
rect 740 309 817 325
rect 740 275 756 309
rect 790 275 817 309
rect 740 259 817 275
rect 853 289 929 350
rect 853 255 869 289
rect 903 255 929 289
rect 991 329 1025 390
rect 1059 413 1099 460
rect 1059 379 1061 413
rect 1095 379 1099 413
rect 1059 363 1099 379
rect 991 319 1086 329
rect 991 285 1036 319
rect 1070 285 1086 319
rect 991 269 1086 285
rect 853 242 929 255
rect 441 206 673 208
rect 441 190 925 206
rect 441 174 623 190
rect 369 101 407 171
rect 613 156 623 174
rect 657 172 925 190
rect 657 156 661 172
rect 369 67 371 101
rect 405 67 407 101
rect 369 51 407 67
rect 448 124 579 140
rect 448 90 457 124
rect 491 90 537 124
rect 571 90 579 124
rect 448 17 579 90
rect 613 101 661 156
rect 881 171 925 172
rect 613 67 623 101
rect 657 67 661 101
rect 613 51 661 67
rect 695 122 763 138
rect 695 88 713 122
rect 747 88 763 122
rect 695 17 763 88
rect 797 122 847 138
rect 797 88 803 122
rect 837 88 847 122
rect 881 137 889 171
rect 923 137 925 171
rect 881 121 925 137
rect 959 205 1018 221
rect 959 171 975 205
rect 1009 171 1018 205
rect 797 87 847 88
rect 959 101 1018 171
rect 959 87 975 101
rect 797 67 975 87
rect 1009 67 1018 101
rect 797 51 1018 67
rect 1052 205 1111 221
rect 1052 171 1061 205
rect 1095 171 1111 205
rect 1052 95 1111 171
rect 1052 61 1061 95
rect 1095 61 1111 95
rect 1052 17 1111 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21o_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2561416
string GDS_START 2551374
<< end >>
