magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 817 259 1615 261
rect 1 49 1615 259
rect 0 0 1632 49
<< scnmos >>
rect 80 65 110 233
rect 166 65 196 233
rect 252 65 282 233
rect 338 65 368 233
rect 424 65 454 233
rect 510 65 540 233
rect 596 65 626 233
rect 682 65 712 233
rect 900 67 930 235
rect 986 67 1016 235
rect 1072 67 1102 235
rect 1158 67 1188 235
rect 1244 67 1274 235
rect 1330 67 1360 235
rect 1416 67 1446 235
rect 1502 67 1532 235
<< scpmoshvt >>
rect 90 367 120 619
rect 176 367 206 619
rect 262 367 292 619
rect 348 367 378 619
rect 466 367 496 619
rect 552 367 582 619
rect 638 367 668 619
rect 724 367 754 619
rect 810 367 840 619
rect 896 367 926 619
rect 982 367 1012 619
rect 1068 367 1098 619
rect 1244 367 1274 619
rect 1330 367 1360 619
rect 1416 367 1446 619
rect 1502 367 1532 619
<< ndiff >>
rect 27 221 80 233
rect 27 187 35 221
rect 69 187 80 221
rect 27 111 80 187
rect 27 77 35 111
rect 69 77 80 111
rect 27 65 80 77
rect 110 183 166 233
rect 110 149 121 183
rect 155 149 166 183
rect 110 107 166 149
rect 110 73 121 107
rect 155 73 166 107
rect 110 65 166 73
rect 196 221 252 233
rect 196 187 207 221
rect 241 187 252 221
rect 196 111 252 187
rect 196 77 207 111
rect 241 77 252 111
rect 196 65 252 77
rect 282 183 338 233
rect 282 149 293 183
rect 327 149 338 183
rect 282 107 338 149
rect 282 73 293 107
rect 327 73 338 107
rect 282 65 338 73
rect 368 221 424 233
rect 368 187 379 221
rect 413 187 424 221
rect 368 107 424 187
rect 368 73 379 107
rect 413 73 424 107
rect 368 65 424 73
rect 454 225 510 233
rect 454 191 465 225
rect 499 191 510 225
rect 454 155 510 191
rect 454 121 465 155
rect 499 121 510 155
rect 454 65 510 121
rect 540 157 596 233
rect 540 123 551 157
rect 585 123 596 157
rect 540 65 596 123
rect 626 225 682 233
rect 626 191 637 225
rect 671 191 682 225
rect 626 155 682 191
rect 626 121 637 155
rect 671 121 682 155
rect 626 65 682 121
rect 712 107 785 233
rect 712 73 739 107
rect 773 73 785 107
rect 712 65 785 73
rect 843 109 900 235
rect 843 75 855 109
rect 889 75 900 109
rect 843 67 900 75
rect 930 183 986 235
rect 930 149 941 183
rect 975 149 986 183
rect 930 67 986 149
rect 1016 109 1072 235
rect 1016 75 1027 109
rect 1061 75 1072 109
rect 1016 67 1072 75
rect 1102 183 1158 235
rect 1102 149 1113 183
rect 1147 149 1158 183
rect 1102 67 1158 149
rect 1188 167 1244 235
rect 1188 133 1199 167
rect 1233 133 1244 167
rect 1188 67 1244 133
rect 1274 227 1330 235
rect 1274 193 1285 227
rect 1319 193 1330 227
rect 1274 159 1330 193
rect 1274 125 1285 159
rect 1319 125 1330 159
rect 1274 67 1330 125
rect 1360 167 1416 235
rect 1360 133 1371 167
rect 1405 133 1416 167
rect 1360 67 1416 133
rect 1446 227 1502 235
rect 1446 193 1457 227
rect 1491 193 1502 227
rect 1446 159 1502 193
rect 1446 125 1457 159
rect 1491 125 1502 159
rect 1446 67 1502 125
rect 1532 223 1589 235
rect 1532 189 1543 223
rect 1577 189 1589 223
rect 1532 113 1589 189
rect 1532 79 1543 113
rect 1577 79 1589 113
rect 1532 67 1589 79
<< pdiff >>
rect 37 607 90 619
rect 37 573 45 607
rect 79 573 90 607
rect 37 516 90 573
rect 37 482 45 516
rect 79 482 90 516
rect 37 434 90 482
rect 37 400 45 434
rect 79 400 90 434
rect 37 367 90 400
rect 120 599 176 619
rect 120 565 131 599
rect 165 565 176 599
rect 120 516 176 565
rect 120 482 131 516
rect 165 482 176 516
rect 120 434 176 482
rect 120 400 131 434
rect 165 400 176 434
rect 120 367 176 400
rect 206 607 262 619
rect 206 573 217 607
rect 251 573 262 607
rect 206 495 262 573
rect 206 461 217 495
rect 251 461 262 495
rect 206 367 262 461
rect 292 599 348 619
rect 292 565 303 599
rect 337 565 348 599
rect 292 516 348 565
rect 292 482 303 516
rect 337 482 348 516
rect 292 434 348 482
rect 292 400 303 434
rect 337 400 348 434
rect 292 367 348 400
rect 378 607 466 619
rect 378 573 405 607
rect 439 573 466 607
rect 378 489 466 573
rect 378 455 405 489
rect 439 455 466 489
rect 378 367 466 455
rect 496 599 552 619
rect 496 565 507 599
rect 541 565 552 599
rect 496 516 552 565
rect 496 482 507 516
rect 541 482 552 516
rect 496 434 552 482
rect 496 400 507 434
rect 541 400 552 434
rect 496 367 552 400
rect 582 607 638 619
rect 582 573 593 607
rect 627 573 638 607
rect 582 489 638 573
rect 582 455 593 489
rect 627 455 638 489
rect 582 367 638 455
rect 668 599 724 619
rect 668 565 679 599
rect 713 565 724 599
rect 668 516 724 565
rect 668 482 679 516
rect 713 482 724 516
rect 668 434 724 482
rect 668 400 679 434
rect 713 400 724 434
rect 668 367 724 400
rect 754 607 810 619
rect 754 573 765 607
rect 799 573 810 607
rect 754 489 810 573
rect 754 455 765 489
rect 799 455 810 489
rect 754 367 810 455
rect 840 599 896 619
rect 840 565 851 599
rect 885 565 896 599
rect 840 516 896 565
rect 840 482 851 516
rect 885 482 896 516
rect 840 434 896 482
rect 840 400 851 434
rect 885 400 896 434
rect 840 367 896 400
rect 926 607 982 619
rect 926 573 937 607
rect 971 573 982 607
rect 926 489 982 573
rect 926 455 937 489
rect 971 455 982 489
rect 926 367 982 455
rect 1012 599 1068 619
rect 1012 565 1023 599
rect 1057 565 1068 599
rect 1012 516 1068 565
rect 1012 482 1023 516
rect 1057 482 1068 516
rect 1012 434 1068 482
rect 1012 400 1023 434
rect 1057 400 1068 434
rect 1012 367 1068 400
rect 1098 607 1244 619
rect 1098 573 1109 607
rect 1143 573 1199 607
rect 1233 573 1244 607
rect 1098 489 1244 573
rect 1098 455 1109 489
rect 1143 455 1199 489
rect 1233 455 1244 489
rect 1098 367 1244 455
rect 1274 599 1330 619
rect 1274 565 1285 599
rect 1319 565 1330 599
rect 1274 516 1330 565
rect 1274 482 1285 516
rect 1319 482 1330 516
rect 1274 434 1330 482
rect 1274 400 1285 434
rect 1319 400 1330 434
rect 1274 367 1330 400
rect 1360 607 1416 619
rect 1360 573 1371 607
rect 1405 573 1416 607
rect 1360 489 1416 573
rect 1360 455 1371 489
rect 1405 455 1416 489
rect 1360 367 1416 455
rect 1446 599 1502 619
rect 1446 565 1457 599
rect 1491 565 1502 599
rect 1446 516 1502 565
rect 1446 482 1457 516
rect 1491 482 1502 516
rect 1446 434 1502 482
rect 1446 400 1457 434
rect 1491 400 1502 434
rect 1446 367 1502 400
rect 1532 607 1585 619
rect 1532 573 1543 607
rect 1577 573 1585 607
rect 1532 514 1585 573
rect 1532 480 1543 514
rect 1577 480 1585 514
rect 1532 419 1585 480
rect 1532 385 1543 419
rect 1577 385 1585 419
rect 1532 367 1585 385
<< ndiffc >>
rect 35 187 69 221
rect 35 77 69 111
rect 121 149 155 183
rect 121 73 155 107
rect 207 187 241 221
rect 207 77 241 111
rect 293 149 327 183
rect 293 73 327 107
rect 379 187 413 221
rect 379 73 413 107
rect 465 191 499 225
rect 465 121 499 155
rect 551 123 585 157
rect 637 191 671 225
rect 637 121 671 155
rect 739 73 773 107
rect 855 75 889 109
rect 941 149 975 183
rect 1027 75 1061 109
rect 1113 149 1147 183
rect 1199 133 1233 167
rect 1285 193 1319 227
rect 1285 125 1319 159
rect 1371 133 1405 167
rect 1457 193 1491 227
rect 1457 125 1491 159
rect 1543 189 1577 223
rect 1543 79 1577 113
<< pdiffc >>
rect 45 573 79 607
rect 45 482 79 516
rect 45 400 79 434
rect 131 565 165 599
rect 131 482 165 516
rect 131 400 165 434
rect 217 573 251 607
rect 217 461 251 495
rect 303 565 337 599
rect 303 482 337 516
rect 303 400 337 434
rect 405 573 439 607
rect 405 455 439 489
rect 507 565 541 599
rect 507 482 541 516
rect 507 400 541 434
rect 593 573 627 607
rect 593 455 627 489
rect 679 565 713 599
rect 679 482 713 516
rect 679 400 713 434
rect 765 573 799 607
rect 765 455 799 489
rect 851 565 885 599
rect 851 482 885 516
rect 851 400 885 434
rect 937 573 971 607
rect 937 455 971 489
rect 1023 565 1057 599
rect 1023 482 1057 516
rect 1023 400 1057 434
rect 1109 573 1143 607
rect 1199 573 1233 607
rect 1109 455 1143 489
rect 1199 455 1233 489
rect 1285 565 1319 599
rect 1285 482 1319 516
rect 1285 400 1319 434
rect 1371 573 1405 607
rect 1371 455 1405 489
rect 1457 565 1491 599
rect 1457 482 1491 516
rect 1457 400 1491 434
rect 1543 573 1577 607
rect 1543 480 1577 514
rect 1543 385 1577 419
<< poly >>
rect 90 619 120 645
rect 176 619 206 645
rect 262 619 292 645
rect 348 619 378 645
rect 466 619 496 645
rect 552 619 582 645
rect 638 619 668 645
rect 724 619 754 645
rect 810 619 840 645
rect 896 619 926 645
rect 982 619 1012 645
rect 1068 619 1098 645
rect 1244 619 1274 645
rect 1330 619 1360 645
rect 1416 619 1446 645
rect 1502 619 1532 645
rect 90 335 120 367
rect 176 335 206 367
rect 262 335 292 367
rect 348 335 378 367
rect 466 335 496 367
rect 552 335 582 367
rect 638 335 668 367
rect 724 335 754 367
rect 810 335 840 367
rect 896 335 926 367
rect 982 335 1012 367
rect 1068 335 1098 367
rect 1244 345 1274 367
rect 1330 345 1360 367
rect 1416 345 1446 367
rect 1502 345 1532 367
rect 1244 335 1532 345
rect 80 319 378 335
rect 80 285 96 319
rect 130 285 164 319
rect 198 285 232 319
rect 266 285 300 319
rect 334 305 378 319
rect 420 319 754 335
rect 334 285 368 305
rect 80 269 368 285
rect 420 285 436 319
rect 470 285 504 319
rect 538 285 572 319
rect 606 285 640 319
rect 674 305 754 319
rect 796 319 1202 335
rect 674 285 712 305
rect 420 269 712 285
rect 796 285 812 319
rect 846 285 880 319
rect 914 285 948 319
rect 982 285 1016 319
rect 1050 285 1084 319
rect 1118 285 1152 319
rect 1186 285 1202 319
rect 796 269 1202 285
rect 1244 319 1582 335
rect 1244 285 1260 319
rect 1294 285 1328 319
rect 1362 285 1396 319
rect 1430 285 1464 319
rect 1498 285 1532 319
rect 1566 285 1582 319
rect 1244 269 1582 285
rect 80 233 110 269
rect 166 233 196 269
rect 252 233 282 269
rect 338 233 368 269
rect 424 233 454 269
rect 510 233 540 269
rect 596 233 626 269
rect 682 233 712 269
rect 900 235 930 269
rect 986 235 1016 269
rect 1072 235 1102 269
rect 1158 235 1188 269
rect 1244 235 1274 269
rect 1330 235 1360 269
rect 1416 235 1446 269
rect 1502 235 1532 269
rect 80 39 110 65
rect 166 39 196 65
rect 252 39 282 65
rect 338 39 368 65
rect 424 39 454 65
rect 510 39 540 65
rect 596 39 626 65
rect 682 39 712 65
rect 900 41 930 67
rect 986 41 1016 67
rect 1072 41 1102 67
rect 1158 41 1188 67
rect 1244 41 1274 67
rect 1330 41 1360 67
rect 1416 41 1446 67
rect 1502 41 1532 67
<< polycont >>
rect 96 285 130 319
rect 164 285 198 319
rect 232 285 266 319
rect 300 285 334 319
rect 436 285 470 319
rect 504 285 538 319
rect 572 285 606 319
rect 640 285 674 319
rect 812 285 846 319
rect 880 285 914 319
rect 948 285 982 319
rect 1016 285 1050 319
rect 1084 285 1118 319
rect 1152 285 1186 319
rect 1260 285 1294 319
rect 1328 285 1362 319
rect 1396 285 1430 319
rect 1464 285 1498 319
rect 1532 285 1566 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 29 607 88 649
rect 29 573 45 607
rect 79 573 88 607
rect 29 516 88 573
rect 29 482 45 516
rect 79 482 88 516
rect 29 434 88 482
rect 29 400 45 434
rect 79 400 88 434
rect 29 384 88 400
rect 122 599 167 615
rect 122 565 131 599
rect 165 565 167 599
rect 122 516 167 565
rect 122 482 131 516
rect 165 482 167 516
rect 122 434 167 482
rect 201 607 267 649
rect 201 573 217 607
rect 251 573 267 607
rect 201 495 267 573
rect 201 461 217 495
rect 251 461 267 495
rect 201 458 267 461
rect 301 599 353 615
rect 301 565 303 599
rect 337 565 353 599
rect 301 516 353 565
rect 301 482 303 516
rect 337 482 353 516
rect 122 400 131 434
rect 165 424 167 434
rect 301 434 353 482
rect 389 607 455 649
rect 389 573 405 607
rect 439 573 455 607
rect 389 489 455 573
rect 389 455 405 489
rect 439 455 455 489
rect 389 452 455 455
rect 489 599 543 615
rect 489 565 507 599
rect 541 565 543 599
rect 489 516 543 565
rect 489 482 507 516
rect 541 482 543 516
rect 301 424 303 434
rect 165 400 303 424
rect 337 418 353 434
rect 489 434 543 482
rect 577 607 643 649
rect 577 573 593 607
rect 627 573 643 607
rect 577 489 643 573
rect 577 455 593 489
rect 627 455 643 489
rect 577 452 643 455
rect 677 599 715 615
rect 677 565 679 599
rect 713 565 715 599
rect 677 516 715 565
rect 677 482 679 516
rect 713 482 715 516
rect 489 418 507 434
rect 337 400 507 418
rect 541 418 543 434
rect 677 434 715 482
rect 749 607 815 649
rect 749 573 765 607
rect 799 573 815 607
rect 749 489 815 573
rect 749 455 765 489
rect 799 455 815 489
rect 749 452 815 455
rect 849 599 887 615
rect 849 565 851 599
rect 885 565 887 599
rect 849 516 887 565
rect 849 482 851 516
rect 885 482 887 516
rect 677 418 679 434
rect 541 400 679 418
rect 713 418 715 434
rect 849 434 887 482
rect 921 607 987 649
rect 921 573 937 607
rect 971 573 987 607
rect 921 489 987 573
rect 921 455 937 489
rect 971 455 987 489
rect 921 452 987 455
rect 1021 599 1059 615
rect 1021 565 1023 599
rect 1057 565 1059 599
rect 1021 516 1059 565
rect 1021 482 1023 516
rect 1057 482 1059 516
rect 849 418 851 434
rect 713 400 851 418
rect 885 418 887 434
rect 1021 434 1059 482
rect 1093 607 1249 649
rect 1093 573 1109 607
rect 1143 573 1199 607
rect 1233 573 1249 607
rect 1093 489 1249 573
rect 1093 455 1109 489
rect 1143 455 1199 489
rect 1233 455 1249 489
rect 1093 452 1249 455
rect 1283 599 1321 615
rect 1283 565 1285 599
rect 1319 565 1321 599
rect 1283 516 1321 565
rect 1283 482 1285 516
rect 1319 482 1321 516
rect 1021 418 1023 434
rect 885 400 1023 418
rect 1057 418 1059 434
rect 1283 434 1321 482
rect 1355 607 1421 649
rect 1355 573 1371 607
rect 1405 573 1421 607
rect 1355 489 1421 573
rect 1355 455 1371 489
rect 1405 455 1421 489
rect 1355 452 1421 455
rect 1455 599 1493 615
rect 1455 565 1457 599
rect 1491 565 1493 599
rect 1455 516 1493 565
rect 1455 482 1457 516
rect 1491 482 1493 516
rect 1283 418 1285 434
rect 1057 400 1285 418
rect 1319 418 1321 434
rect 1455 434 1493 482
rect 1455 418 1457 434
rect 1319 400 1457 418
rect 1491 400 1493 434
rect 122 384 1493 400
rect 1527 607 1593 649
rect 1527 573 1543 607
rect 1577 573 1593 607
rect 1527 514 1593 573
rect 1527 480 1543 514
rect 1577 480 1593 514
rect 1527 419 1593 480
rect 1527 385 1543 419
rect 1577 385 1593 419
rect 1527 384 1593 385
rect 20 319 353 350
rect 20 285 96 319
rect 130 285 164 319
rect 198 285 232 319
rect 266 285 300 319
rect 334 285 353 319
rect 415 319 690 350
rect 415 285 436 319
rect 470 285 504 319
rect 538 285 572 319
rect 606 285 640 319
rect 674 285 690 319
rect 440 276 690 285
rect 726 251 760 384
rect 796 319 1202 350
rect 796 285 812 319
rect 846 285 880 319
rect 914 285 948 319
rect 982 285 1016 319
rect 1050 285 1084 319
rect 1118 285 1152 319
rect 1186 285 1202 319
rect 1244 319 1601 350
rect 1244 285 1260 319
rect 1294 285 1328 319
rect 1362 285 1396 319
rect 1430 285 1464 319
rect 1498 285 1532 319
rect 1566 285 1601 319
rect 31 221 415 251
rect 31 187 35 221
rect 69 217 207 221
rect 69 187 71 217
rect 31 111 71 187
rect 205 187 207 217
rect 241 217 379 221
rect 241 187 243 217
rect 31 77 35 111
rect 69 77 71 111
rect 31 61 71 77
rect 105 149 121 183
rect 155 149 171 183
rect 105 107 171 149
rect 105 73 121 107
rect 155 73 171 107
rect 105 17 171 73
rect 205 111 243 187
rect 377 187 379 217
rect 413 187 415 221
rect 205 77 207 111
rect 241 77 243 111
rect 205 61 243 77
rect 277 149 293 183
rect 327 149 343 183
rect 277 107 343 149
rect 277 73 293 107
rect 327 73 343 107
rect 277 17 343 73
rect 377 107 415 187
rect 449 225 687 241
rect 449 191 465 225
rect 499 207 637 225
rect 499 191 515 207
rect 449 155 515 191
rect 621 191 637 207
rect 671 191 687 225
rect 726 227 1507 251
rect 726 217 1285 227
rect 621 183 687 191
rect 1269 193 1285 217
rect 1319 217 1457 227
rect 1319 193 1335 217
rect 449 121 465 155
rect 499 121 515 155
rect 549 157 587 173
rect 549 123 551 157
rect 585 123 587 157
rect 377 73 379 107
rect 413 87 415 107
rect 549 87 587 123
rect 621 155 941 183
rect 621 121 637 155
rect 671 149 941 155
rect 975 149 1113 183
rect 1147 149 1163 183
rect 1197 167 1235 183
rect 671 121 687 149
rect 1197 133 1199 167
rect 1233 133 1235 167
rect 1197 115 1235 133
rect 1269 159 1335 193
rect 1441 193 1457 217
rect 1491 193 1507 227
rect 1269 125 1285 159
rect 1319 125 1335 159
rect 1369 167 1407 183
rect 1369 133 1371 167
rect 1405 133 1407 167
rect 723 107 789 113
rect 723 87 739 107
rect 413 73 739 87
rect 773 73 789 107
rect 377 53 789 73
rect 839 109 1235 115
rect 839 75 855 109
rect 889 75 1027 109
rect 1061 89 1235 109
rect 1369 89 1407 133
rect 1441 159 1507 193
rect 1441 125 1457 159
rect 1491 125 1507 159
rect 1541 223 1593 239
rect 1541 189 1543 223
rect 1577 189 1593 223
rect 1541 113 1593 189
rect 1541 89 1543 113
rect 1061 79 1543 89
rect 1577 79 1593 113
rect 1061 75 1593 79
rect 839 55 1593 75
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4622546
string GDS_START 4607944
<< end >>
