magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 112 49 1074 273
rect 0 0 1152 49
<< scnmos >>
rect 191 47 991 247
<< scpmoshvt >>
rect 178 419 978 619
<< ndiff >>
rect 138 229 191 247
rect 138 195 146 229
rect 180 195 191 229
rect 138 161 191 195
rect 138 127 146 161
rect 180 127 191 161
rect 138 93 191 127
rect 138 59 146 93
rect 180 59 191 93
rect 138 47 191 59
rect 991 225 1048 247
rect 991 191 1002 225
rect 1036 191 1048 225
rect 991 157 1048 191
rect 991 123 1002 157
rect 1036 123 1048 157
rect 991 89 1048 123
rect 991 55 1002 89
rect 1036 55 1048 89
rect 991 47 1048 55
<< pdiff >>
rect 123 607 178 619
rect 123 573 131 607
rect 165 573 178 607
rect 123 539 178 573
rect 123 505 131 539
rect 165 505 178 539
rect 123 471 178 505
rect 123 437 131 471
rect 165 437 178 471
rect 123 419 178 437
rect 978 611 1035 619
rect 978 577 989 611
rect 1023 577 1035 611
rect 978 543 1035 577
rect 978 509 989 543
rect 1023 509 1035 543
rect 978 475 1035 509
rect 978 441 989 475
rect 1023 441 1035 475
rect 978 419 1035 441
<< ndiffc >>
rect 146 195 180 229
rect 146 127 180 161
rect 146 59 180 93
rect 1002 191 1036 225
rect 1002 123 1036 157
rect 1002 55 1036 89
<< pdiffc >>
rect 131 573 165 607
rect 131 505 165 539
rect 131 437 165 471
rect 989 577 1023 611
rect 989 509 1023 543
rect 989 441 1023 475
<< poly >>
rect 178 619 978 645
rect 178 387 978 419
rect 174 377 978 387
rect 174 371 516 377
rect 174 337 194 371
rect 228 337 262 371
rect 296 337 330 371
rect 364 337 398 371
rect 432 337 466 371
rect 500 337 516 371
rect 174 321 516 337
rect 585 319 991 335
rect 585 285 601 319
rect 635 285 669 319
rect 703 285 737 319
rect 771 285 805 319
rect 839 285 873 319
rect 907 285 941 319
rect 975 285 991 319
rect 585 273 991 285
rect 191 247 991 273
rect 191 21 991 47
<< polycont >>
rect 194 337 228 371
rect 262 337 296 371
rect 330 337 364 371
rect 398 337 432 371
rect 466 337 500 371
rect 601 285 635 319
rect 669 285 703 319
rect 737 285 771 319
rect 805 285 839 319
rect 873 285 907 319
rect 941 285 975 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 115 607 181 615
rect 115 579 131 607
rect 165 589 181 607
rect 973 611 1039 615
rect 973 589 989 611
rect 165 579 989 589
rect 165 573 187 579
rect 149 545 187 573
rect 221 545 259 579
rect 293 545 331 579
rect 365 545 403 579
rect 437 545 475 579
rect 509 545 547 579
rect 581 545 619 579
rect 653 545 691 579
rect 725 545 770 579
rect 804 545 842 579
rect 876 545 914 579
rect 948 545 986 579
rect 1023 577 1039 611
rect 1020 545 1039 577
rect 115 543 1039 545
rect 115 539 989 543
rect 115 505 131 539
rect 165 535 989 539
rect 165 505 181 535
rect 115 471 181 505
rect 115 437 131 471
rect 165 437 181 471
rect 115 421 181 437
rect 973 509 989 535
rect 1023 509 1039 543
rect 973 475 1039 509
rect 973 441 989 475
rect 1023 441 1039 475
rect 130 371 516 387
rect 130 337 194 371
rect 228 337 262 371
rect 296 337 330 371
rect 364 337 398 371
rect 432 337 466 371
rect 500 337 516 371
rect 130 321 516 337
rect 973 335 1039 441
rect 130 229 196 321
rect 585 319 1039 335
rect 585 285 601 319
rect 635 285 669 319
rect 703 285 737 319
rect 771 285 805 319
rect 839 285 873 319
rect 907 285 941 319
rect 975 285 1039 319
rect 585 268 1039 285
rect 130 195 146 229
rect 180 195 196 229
rect 130 161 196 195
rect 130 127 146 161
rect 180 127 196 161
rect 130 93 196 127
rect 130 59 146 93
rect 180 59 196 93
rect 130 17 196 59
rect 986 191 1002 225
rect 1036 191 1052 225
rect 986 157 1052 191
rect 986 123 1002 157
rect 1036 123 1052 157
rect 986 89 1052 123
rect 986 55 1002 89
rect 1036 55 1052 89
rect 986 17 1052 55
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 115 573 131 579
rect 131 573 149 579
rect 115 545 149 573
rect 187 545 221 579
rect 259 545 293 579
rect 331 545 365 579
rect 403 545 437 579
rect 475 545 509 579
rect 547 545 581 579
rect 619 545 653 579
rect 691 545 725 579
rect 770 545 804 579
rect 842 545 876 579
rect 914 545 948 579
rect 986 577 989 579
rect 989 577 1020 579
rect 986 545 1020 577
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 14 579 1138 589
rect 14 545 115 579
rect 149 545 187 579
rect 221 545 259 579
rect 293 545 331 579
rect 365 545 403 579
rect 437 545 475 579
rect 509 545 547 579
rect 581 545 619 579
rect 653 545 691 579
rect 725 545 770 579
rect 804 545 842 579
rect 876 545 914 579
rect 948 545 986 579
rect 1020 545 1138 579
rect 14 535 1138 545
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 decapkapwr_12
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 14 535 1138 589 0 FreeSans 200 0 0 0 KAPWR
port 1 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE SPACER
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 876342
string GDS_START 870384
<< end >>
