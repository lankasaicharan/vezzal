magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1586 1975
<< nwell >>
rect -38 331 326 704
<< pwell >>
rect 15 49 281 157
rect 0 0 288 49
<< scnmos >>
rect 94 47 124 131
rect 172 47 202 131
<< scpmoshvt >>
rect 86 462 116 590
rect 172 462 202 590
<< ndiff >>
rect 41 106 94 131
rect 41 72 49 106
rect 83 72 94 106
rect 41 47 94 72
rect 124 47 172 131
rect 202 106 255 131
rect 202 72 213 106
rect 247 72 255 106
rect 202 47 255 72
<< pdiff >>
rect 33 578 86 590
rect 33 544 41 578
rect 75 544 86 578
rect 33 508 86 544
rect 33 474 41 508
rect 75 474 86 508
rect 33 462 86 474
rect 116 578 172 590
rect 116 544 127 578
rect 161 544 172 578
rect 116 510 172 544
rect 116 476 127 510
rect 161 476 172 510
rect 116 462 172 476
rect 202 578 255 590
rect 202 544 213 578
rect 247 544 255 578
rect 202 508 255 544
rect 202 474 213 508
rect 247 474 255 508
rect 202 462 255 474
<< ndiffc >>
rect 49 72 83 106
rect 213 72 247 106
<< pdiffc >>
rect 41 544 75 578
rect 41 474 75 508
rect 127 544 161 578
rect 127 476 161 510
rect 213 544 247 578
rect 213 474 247 508
<< poly >>
rect 86 590 116 616
rect 172 590 202 616
rect 86 302 116 462
rect 172 302 202 462
rect 37 286 124 302
rect 37 252 53 286
rect 87 252 124 286
rect 37 218 124 252
rect 37 184 53 218
rect 87 184 124 218
rect 37 168 124 184
rect 94 131 124 168
rect 172 286 247 302
rect 172 252 197 286
rect 231 252 247 286
rect 172 218 247 252
rect 172 184 197 218
rect 231 184 247 218
rect 172 168 247 184
rect 172 131 202 168
rect 94 21 124 47
rect 172 21 202 47
<< polycont >>
rect 53 252 87 286
rect 53 184 87 218
rect 197 252 231 286
rect 197 184 231 218
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 25 578 87 649
rect 25 544 41 578
rect 75 544 87 578
rect 25 508 87 544
rect 25 474 41 508
rect 75 474 87 508
rect 25 458 87 474
rect 121 578 163 594
rect 121 544 127 578
rect 161 544 163 578
rect 121 510 163 544
rect 121 476 127 510
rect 161 476 163 510
rect 17 286 87 424
rect 17 252 53 286
rect 17 218 87 252
rect 17 184 53 218
rect 17 168 87 184
rect 121 122 163 476
rect 197 578 263 649
rect 197 544 213 578
rect 247 544 263 578
rect 197 508 263 544
rect 197 474 213 508
rect 247 474 263 508
rect 197 458 263 474
rect 197 286 271 424
rect 231 252 271 286
rect 197 218 271 252
rect 231 184 271 218
rect 197 168 271 184
rect 33 106 87 122
rect 33 72 49 106
rect 83 72 87 106
rect 33 17 87 72
rect 121 106 263 122
rect 121 72 213 106
rect 247 72 263 106
rect 121 56 263 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
<< metal1 >>
rect 0 683 288 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 0 617 288 649
rect 0 17 288 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
rect 0 -49 288 -17
<< labels >>
flabel pwell s 0 0 288 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 288 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2_0
flabel metal1 s 0 617 288 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 288 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 288 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5785204
string GDS_START 5780196
<< end >>
