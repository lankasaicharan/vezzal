magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 972 229 1246 235
rect 75 157 1246 229
rect 75 49 1535 157
rect 0 0 1536 49
<< scnmos >>
rect 154 119 184 203
rect 240 119 270 203
rect 312 119 342 203
rect 412 119 442 203
rect 484 119 514 203
rect 612 119 642 203
rect 684 119 714 203
rect 770 119 800 203
rect 842 119 872 203
rect 1051 125 1081 209
rect 1137 125 1167 209
rect 1340 47 1370 131
rect 1426 47 1456 131
<< scpmoshvt >>
rect 84 506 114 590
rect 192 506 222 590
rect 264 506 294 590
rect 396 504 426 588
rect 468 504 498 588
rect 583 504 613 588
rect 655 504 685 588
rect 763 504 793 588
rect 835 504 865 588
rect 1045 493 1075 577
rect 1131 493 1161 577
rect 1321 403 1351 487
rect 1426 403 1456 531
<< ndiff >>
rect 101 178 154 203
rect 101 144 109 178
rect 143 144 154 178
rect 101 119 154 144
rect 184 168 240 203
rect 184 134 195 168
rect 229 134 240 168
rect 184 119 240 134
rect 270 119 312 203
rect 342 178 412 203
rect 342 144 367 178
rect 401 144 412 178
rect 342 119 412 144
rect 442 119 484 203
rect 514 178 612 203
rect 514 144 547 178
rect 581 144 612 178
rect 514 119 612 144
rect 642 119 684 203
rect 714 178 770 203
rect 714 144 725 178
rect 759 144 770 178
rect 714 119 770 144
rect 800 119 842 203
rect 872 178 925 203
rect 872 144 883 178
rect 917 144 925 178
rect 872 119 925 144
rect 998 184 1051 209
rect 998 150 1006 184
rect 1040 150 1051 184
rect 998 125 1051 150
rect 1081 184 1137 209
rect 1081 150 1092 184
rect 1126 150 1137 184
rect 1081 125 1137 150
rect 1167 184 1220 209
rect 1167 150 1178 184
rect 1212 150 1220 184
rect 1167 125 1220 150
rect 1287 106 1340 131
rect 1287 72 1295 106
rect 1329 72 1340 106
rect 1287 47 1340 72
rect 1370 106 1426 131
rect 1370 72 1381 106
rect 1415 72 1426 106
rect 1370 47 1426 72
rect 1456 106 1509 131
rect 1456 72 1467 106
rect 1501 72 1509 106
rect 1456 47 1509 72
<< pdiff >>
rect 31 565 84 590
rect 31 531 39 565
rect 73 531 84 565
rect 31 506 84 531
rect 114 578 192 590
rect 114 544 139 578
rect 173 544 192 578
rect 114 506 192 544
rect 222 506 264 590
rect 294 588 374 590
rect 294 545 396 588
rect 294 511 328 545
rect 362 511 396 545
rect 294 506 396 511
rect 316 504 396 506
rect 426 504 468 588
rect 498 578 583 588
rect 498 544 534 578
rect 568 544 583 578
rect 498 504 583 544
rect 613 504 655 588
rect 685 568 763 588
rect 685 534 707 568
rect 741 534 763 568
rect 685 504 763 534
rect 793 504 835 588
rect 865 572 918 588
rect 865 538 876 572
rect 910 538 918 572
rect 865 504 918 538
rect 992 552 1045 577
rect 992 518 1000 552
rect 1034 518 1045 552
rect 316 501 374 504
rect 992 493 1045 518
rect 1075 565 1131 577
rect 1075 531 1086 565
rect 1120 531 1131 565
rect 1075 493 1131 531
rect 1161 542 1214 577
rect 1161 508 1172 542
rect 1206 508 1214 542
rect 1373 519 1426 531
rect 1161 493 1214 508
rect 1373 487 1381 519
rect 1268 462 1321 487
rect 1268 428 1276 462
rect 1310 428 1321 462
rect 1268 403 1321 428
rect 1351 485 1381 487
rect 1415 485 1426 519
rect 1351 449 1426 485
rect 1351 415 1362 449
rect 1396 415 1426 449
rect 1351 403 1426 415
rect 1456 519 1509 531
rect 1456 485 1467 519
rect 1501 485 1509 519
rect 1456 449 1509 485
rect 1456 415 1467 449
rect 1501 415 1509 449
rect 1456 403 1509 415
<< ndiffc >>
rect 109 144 143 178
rect 195 134 229 168
rect 367 144 401 178
rect 547 144 581 178
rect 725 144 759 178
rect 883 144 917 178
rect 1006 150 1040 184
rect 1092 150 1126 184
rect 1178 150 1212 184
rect 1295 72 1329 106
rect 1381 72 1415 106
rect 1467 72 1501 106
<< pdiffc >>
rect 39 531 73 565
rect 139 544 173 578
rect 328 511 362 545
rect 534 544 568 578
rect 707 534 741 568
rect 876 538 910 572
rect 1000 518 1034 552
rect 1086 531 1120 565
rect 1172 508 1206 542
rect 1276 428 1310 462
rect 1381 485 1415 519
rect 1362 415 1396 449
rect 1467 485 1501 519
rect 1467 415 1501 449
<< poly >>
rect 84 590 114 616
rect 192 590 222 616
rect 264 590 294 616
rect 396 588 426 614
rect 468 588 498 614
rect 583 588 613 614
rect 655 588 685 614
rect 763 588 793 614
rect 835 588 865 614
rect 1283 606 1349 622
rect 84 383 114 506
rect 192 461 222 506
rect 186 449 222 461
rect 156 433 222 449
rect 156 399 172 433
rect 206 399 222 433
rect 264 461 294 506
rect 1045 577 1075 603
rect 1131 577 1161 603
rect 264 438 336 461
rect 264 431 286 438
rect 156 383 222 399
rect 270 404 286 431
rect 320 404 336 438
rect 270 388 336 404
rect 78 341 114 383
rect 78 325 144 341
rect 78 291 94 325
rect 128 291 144 325
rect 192 340 222 383
rect 192 310 270 340
rect 396 337 426 504
rect 468 440 498 504
rect 468 424 534 440
rect 468 390 484 424
rect 518 390 534 424
rect 583 404 613 504
rect 655 472 685 504
rect 655 456 721 472
rect 655 422 671 456
rect 705 422 721 456
rect 655 406 721 422
rect 468 374 534 390
rect 78 268 144 291
rect 78 238 184 268
rect 154 203 184 238
rect 240 203 270 310
rect 312 321 426 337
rect 312 287 328 321
rect 362 287 426 321
rect 312 271 426 287
rect 312 203 342 271
rect 412 203 442 229
rect 484 203 514 374
rect 577 364 613 404
rect 576 348 642 364
rect 576 314 592 348
rect 626 314 642 348
rect 576 280 642 314
rect 763 307 793 504
rect 576 246 592 280
rect 626 246 642 280
rect 690 277 793 307
rect 835 322 865 504
rect 1283 572 1299 606
rect 1333 586 1349 606
rect 1333 572 1456 586
rect 1283 556 1456 572
rect 1426 531 1456 556
rect 914 432 981 448
rect 914 398 930 432
rect 964 398 981 432
rect 914 382 981 398
rect 835 292 872 322
rect 690 255 720 277
rect 576 230 642 246
rect 612 203 642 230
rect 684 225 720 255
rect 842 276 909 292
rect 842 242 859 276
rect 893 242 909 276
rect 684 203 714 225
rect 770 203 800 229
rect 842 226 909 242
rect 842 203 872 226
rect 154 51 184 119
rect 240 93 270 119
rect 312 93 342 119
rect 412 51 442 119
rect 484 93 514 119
rect 612 93 642 119
rect 684 51 714 119
rect 154 21 714 51
rect 770 51 800 119
rect 842 93 872 119
rect 951 51 981 382
rect 1045 313 1075 493
rect 1131 385 1161 493
rect 1321 487 1351 513
rect 1131 355 1276 385
rect 1321 365 1351 403
rect 1426 381 1456 403
rect 1210 321 1226 355
rect 1260 321 1276 355
rect 1045 283 1162 313
rect 1210 305 1276 321
rect 1318 349 1384 365
rect 1426 351 1462 381
rect 1318 315 1334 349
rect 1368 315 1384 349
rect 1132 261 1162 283
rect 1318 281 1384 315
rect 1318 261 1334 281
rect 1132 247 1334 261
rect 1368 247 1384 281
rect 1051 209 1081 235
rect 1132 231 1384 247
rect 1137 209 1167 231
rect 1340 131 1370 231
rect 1432 183 1462 351
rect 1426 153 1462 183
rect 1426 131 1456 153
rect 1051 103 1081 125
rect 770 21 981 51
rect 1029 87 1095 103
rect 1137 99 1167 125
rect 1029 53 1045 87
rect 1079 53 1095 87
rect 1029 37 1095 53
rect 1340 21 1370 47
rect 1426 21 1456 47
<< polycont >>
rect 172 399 206 433
rect 286 404 320 438
rect 94 291 128 325
rect 484 390 518 424
rect 671 422 705 456
rect 328 287 362 321
rect 592 314 626 348
rect 592 246 626 280
rect 1299 572 1333 606
rect 930 398 964 432
rect 859 242 893 276
rect 1226 321 1260 355
rect 1334 315 1368 349
rect 1334 247 1368 281
rect 1045 53 1079 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 23 565 89 581
rect 23 531 39 565
rect 73 531 89 565
rect 123 578 189 649
rect 123 544 139 578
rect 173 544 189 578
rect 123 540 189 544
rect 227 581 500 615
rect 23 506 89 531
rect 227 506 261 581
rect 23 472 261 506
rect 312 545 432 547
rect 312 511 328 545
rect 362 511 432 545
rect 312 495 432 511
rect 23 241 60 472
rect 110 433 222 438
rect 110 399 172 433
rect 206 399 222 433
rect 110 386 222 399
rect 258 404 286 438
rect 320 404 336 438
rect 258 388 336 404
rect 258 352 292 388
rect 94 325 292 352
rect 128 316 292 325
rect 326 321 364 337
rect 128 291 258 316
rect 94 275 258 291
rect 326 287 328 321
rect 362 287 364 321
rect 326 273 364 287
rect 297 241 364 273
rect 23 239 364 241
rect 23 207 331 239
rect 23 205 145 207
rect 93 178 145 205
rect 398 203 432 495
rect 466 494 500 581
rect 534 578 584 649
rect 568 544 584 578
rect 534 528 584 544
rect 691 568 775 584
rect 691 534 707 568
rect 741 534 775 568
rect 860 572 926 649
rect 860 538 876 572
rect 910 538 926 572
rect 1084 606 1349 615
rect 1084 581 1299 606
rect 860 534 926 538
rect 984 552 1050 568
rect 691 528 775 534
rect 741 500 775 528
rect 984 518 1000 552
rect 1034 518 1050 552
rect 984 500 1050 518
rect 466 460 707 494
rect 741 466 1050 500
rect 655 456 707 460
rect 468 424 569 426
rect 468 390 484 424
rect 518 390 569 424
rect 468 386 569 390
rect 655 422 671 456
rect 705 432 707 456
rect 705 422 930 432
rect 655 398 930 422
rect 964 398 980 432
rect 655 386 980 398
rect 495 348 737 352
rect 495 314 592 348
rect 626 314 737 348
rect 1016 346 1050 466
rect 495 280 737 314
rect 495 246 592 280
rect 626 246 737 280
rect 495 229 737 246
rect 773 312 1050 346
rect 398 202 465 203
rect 398 194 415 202
rect 93 144 109 178
rect 143 144 145 178
rect 365 178 415 194
rect 93 128 145 144
rect 179 168 245 173
rect 179 134 195 168
rect 229 134 245 168
rect 179 17 245 134
rect 365 144 367 178
rect 401 168 415 178
rect 449 168 465 202
rect 773 194 807 312
rect 843 276 945 278
rect 843 242 859 276
rect 893 242 945 276
rect 843 228 945 242
rect 401 144 465 168
rect 365 128 465 144
rect 531 178 597 194
rect 531 144 547 178
rect 581 144 597 178
rect 531 17 597 144
rect 709 178 807 194
rect 709 144 725 178
rect 759 144 807 178
rect 709 128 807 144
rect 867 178 933 194
rect 867 144 883 178
rect 917 144 933 178
rect 867 17 933 144
rect 990 184 1050 312
rect 990 150 1006 184
rect 1040 150 1050 184
rect 990 134 1050 150
rect 1084 565 1122 581
rect 1084 531 1086 565
rect 1120 531 1122 565
rect 1283 572 1299 581
rect 1333 572 1349 606
rect 1283 556 1349 572
rect 1084 201 1122 531
rect 1156 542 1222 547
rect 1156 508 1172 542
rect 1206 508 1222 542
rect 1383 535 1419 649
rect 1376 523 1419 535
rect 1156 492 1222 508
rect 1360 519 1419 523
rect 1156 269 1190 492
rect 1360 485 1381 519
rect 1415 485 1419 519
rect 1260 462 1326 478
rect 1260 428 1276 462
rect 1310 428 1326 462
rect 1260 412 1326 428
rect 1360 449 1419 485
rect 1360 415 1362 449
rect 1396 415 1419 449
rect 1260 371 1298 412
rect 1360 399 1419 415
rect 1457 519 1517 535
rect 1457 485 1467 519
rect 1501 485 1517 519
rect 1457 449 1517 485
rect 1457 415 1467 449
rect 1501 415 1517 449
rect 1224 355 1298 371
rect 1224 321 1226 355
rect 1260 321 1298 355
rect 1224 305 1298 321
rect 1156 235 1228 269
rect 1162 202 1228 235
rect 1084 184 1128 201
rect 1084 150 1092 184
rect 1126 150 1128 184
rect 1084 134 1128 150
rect 1162 184 1183 202
rect 1162 150 1178 184
rect 1217 168 1228 202
rect 1212 150 1228 168
rect 1162 134 1228 150
rect 1262 122 1298 305
rect 1332 349 1423 365
rect 1332 315 1334 349
rect 1368 315 1423 349
rect 1332 281 1423 315
rect 1332 247 1334 281
rect 1368 247 1423 281
rect 1332 156 1423 247
rect 1262 106 1338 122
rect 1262 100 1295 106
rect 1029 87 1295 100
rect 1029 53 1045 87
rect 1079 72 1295 87
rect 1329 72 1338 106
rect 1079 53 1338 72
rect 1029 51 1338 53
rect 1372 106 1423 122
rect 1372 72 1381 106
rect 1415 72 1423 106
rect 1372 17 1423 72
rect 1457 106 1517 415
rect 1457 72 1467 106
rect 1501 72 1517 106
rect 1457 56 1517 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 415 168 449 202
rect 1183 184 1217 202
rect 1183 168 1212 184
rect 1212 168 1217 184
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 403 202 461 208
rect 403 168 415 202
rect 449 199 461 202
rect 1171 202 1229 208
rect 1171 199 1183 202
rect 449 171 1183 199
rect 449 168 461 171
rect 403 162 461 168
rect 1171 168 1183 171
rect 1217 168 1229 202
rect 1171 162 1229 168
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux4_0
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 1375 168 1409 202 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 1471 94 1505 128 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1471 168 1505 202 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1471 390 1505 424 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1491074
string GDS_START 1477788
<< end >>
