magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 105 233 290 248
rect 671 233 856 277
rect 105 49 856 233
rect 0 0 864 49
<< scpmos >>
rect 177 368 207 592
rect 280 392 310 592
rect 370 392 400 592
rect 564 392 594 592
rect 654 392 684 592
rect 750 392 780 592
<< nmoslvt >>
rect 184 74 214 222
rect 387 79 417 207
rect 459 79 489 207
rect 567 79 597 207
rect 639 79 669 207
rect 747 123 777 251
<< ndiff >>
rect 131 210 184 222
rect 131 176 139 210
rect 173 176 184 210
rect 131 120 184 176
rect 131 86 139 120
rect 173 86 184 120
rect 131 74 184 86
rect 214 207 264 222
rect 697 207 747 251
rect 214 152 387 207
rect 214 118 225 152
rect 259 118 342 152
rect 376 118 387 152
rect 214 79 387 118
rect 417 79 459 207
rect 489 199 567 207
rect 489 165 511 199
rect 545 165 567 199
rect 489 121 567 165
rect 489 87 511 121
rect 545 87 567 121
rect 489 79 567 87
rect 597 79 639 207
rect 669 189 747 207
rect 669 155 684 189
rect 718 155 747 189
rect 669 123 747 155
rect 777 218 830 251
rect 777 184 788 218
rect 822 184 830 218
rect 777 123 830 184
rect 669 121 730 123
rect 669 87 684 121
rect 718 87 730 121
rect 669 79 730 87
rect 214 74 267 79
<< pdiff >>
rect 122 580 177 592
rect 122 546 130 580
rect 164 546 177 580
rect 122 497 177 546
rect 122 463 130 497
rect 164 463 177 497
rect 122 414 177 463
rect 122 380 130 414
rect 164 380 177 414
rect 122 368 177 380
rect 207 580 280 592
rect 207 546 220 580
rect 254 546 280 580
rect 207 510 280 546
rect 207 476 220 510
rect 254 476 280 510
rect 207 440 280 476
rect 207 406 220 440
rect 254 406 280 440
rect 207 392 280 406
rect 310 580 370 592
rect 310 546 323 580
rect 357 546 370 580
rect 310 510 370 546
rect 310 476 323 510
rect 357 476 370 510
rect 310 440 370 476
rect 310 406 323 440
rect 357 406 370 440
rect 310 392 370 406
rect 400 580 455 592
rect 400 546 413 580
rect 447 546 455 580
rect 400 512 455 546
rect 400 478 413 512
rect 447 478 455 512
rect 400 392 455 478
rect 509 580 564 592
rect 509 546 517 580
rect 551 546 564 580
rect 509 512 564 546
rect 509 478 517 512
rect 551 478 564 512
rect 509 392 564 478
rect 594 541 654 592
rect 594 507 607 541
rect 641 507 654 541
rect 594 440 654 507
rect 594 406 607 440
rect 641 406 654 440
rect 594 392 654 406
rect 684 580 750 592
rect 684 546 700 580
rect 734 546 750 580
rect 684 510 750 546
rect 684 476 700 510
rect 734 476 750 510
rect 684 440 750 476
rect 684 406 700 440
rect 734 406 750 440
rect 684 392 750 406
rect 780 580 835 592
rect 780 546 793 580
rect 827 546 835 580
rect 780 509 835 546
rect 780 475 793 509
rect 827 475 835 509
rect 780 438 835 475
rect 780 404 793 438
rect 827 404 835 438
rect 780 392 835 404
rect 207 368 262 392
<< ndiffc >>
rect 139 176 173 210
rect 139 86 173 120
rect 225 118 259 152
rect 342 118 376 152
rect 511 165 545 199
rect 511 87 545 121
rect 684 155 718 189
rect 788 184 822 218
rect 684 87 718 121
<< pdiffc >>
rect 130 546 164 580
rect 130 463 164 497
rect 130 380 164 414
rect 220 546 254 580
rect 220 476 254 510
rect 220 406 254 440
rect 323 546 357 580
rect 323 476 357 510
rect 323 406 357 440
rect 413 546 447 580
rect 413 478 447 512
rect 517 546 551 580
rect 517 478 551 512
rect 607 507 641 541
rect 607 406 641 440
rect 700 546 734 580
rect 700 476 734 510
rect 700 406 734 440
rect 793 546 827 580
rect 793 475 827 509
rect 793 404 827 438
<< poly >>
rect 177 592 207 618
rect 280 592 310 618
rect 370 592 400 618
rect 564 592 594 618
rect 654 592 684 618
rect 750 592 780 618
rect 280 377 310 392
rect 370 377 400 392
rect 564 377 594 392
rect 654 377 684 392
rect 750 377 780 392
rect 177 353 207 368
rect 174 326 210 353
rect 277 336 313 377
rect 367 360 403 377
rect 367 344 489 360
rect 561 356 597 377
rect 651 356 687 377
rect 148 310 214 326
rect 148 276 164 310
rect 198 276 214 310
rect 148 260 214 276
rect 184 222 214 260
rect 259 320 325 336
rect 259 286 275 320
rect 309 286 325 320
rect 367 310 409 344
rect 443 310 489 344
rect 367 294 489 310
rect 259 252 325 286
rect 295 222 417 252
rect 387 207 417 222
rect 459 207 489 294
rect 531 340 597 356
rect 531 306 547 340
rect 581 306 597 340
rect 531 290 597 306
rect 567 207 597 290
rect 639 340 705 356
rect 639 306 655 340
rect 689 306 705 340
rect 639 290 705 306
rect 639 207 669 290
rect 747 266 783 377
rect 747 251 777 266
rect 747 101 777 123
rect 747 85 839 101
rect 184 48 214 74
rect 387 53 417 79
rect 459 53 489 79
rect 567 53 597 79
rect 639 53 669 79
rect 747 51 789 85
rect 823 51 839 85
rect 747 35 839 51
<< polycont >>
rect 164 276 198 310
rect 275 286 309 320
rect 409 310 443 344
rect 547 306 581 340
rect 655 306 689 340
rect 789 51 823 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 25 580 180 596
rect 25 546 130 580
rect 164 546 180 580
rect 25 497 180 546
rect 25 463 130 497
rect 164 463 180 497
rect 25 414 180 463
rect 25 380 130 414
rect 164 380 180 414
rect 220 580 270 649
rect 254 546 270 580
rect 220 510 270 546
rect 254 476 270 510
rect 220 440 270 476
rect 254 406 270 440
rect 220 390 270 406
rect 307 580 357 596
rect 307 546 323 580
rect 307 510 357 546
rect 307 476 323 510
rect 307 440 357 476
rect 397 580 463 649
rect 397 546 413 580
rect 447 546 463 580
rect 397 512 463 546
rect 397 478 413 512
rect 447 478 463 512
rect 397 462 463 478
rect 501 581 737 615
rect 501 580 557 581
rect 501 546 517 580
rect 551 546 557 580
rect 697 580 737 581
rect 501 512 557 546
rect 501 478 517 512
rect 551 478 557 512
rect 501 462 557 478
rect 591 541 657 547
rect 591 507 607 541
rect 641 507 657 541
rect 307 406 323 440
rect 591 440 657 507
rect 591 428 607 440
rect 357 406 607 428
rect 641 406 657 440
rect 307 394 657 406
rect 307 390 357 394
rect 591 390 657 394
rect 697 546 700 580
rect 734 546 737 580
rect 697 510 737 546
rect 697 476 700 510
rect 734 476 737 510
rect 697 440 737 476
rect 697 406 700 440
rect 734 406 737 440
rect 697 390 737 406
rect 777 580 843 596
rect 777 546 793 580
rect 827 546 843 580
rect 777 509 843 546
rect 777 475 793 509
rect 827 475 843 509
rect 777 438 843 475
rect 777 404 793 438
rect 827 404 843 438
rect 25 364 180 380
rect 25 226 100 364
rect 148 310 241 326
rect 148 276 164 310
rect 198 276 241 310
rect 148 260 241 276
rect 275 320 359 356
rect 309 286 359 320
rect 393 344 459 360
rect 393 310 409 344
rect 443 310 459 344
rect 393 294 459 310
rect 505 340 597 356
rect 505 306 547 340
rect 581 306 597 340
rect 505 291 597 306
rect 639 340 743 356
rect 639 306 655 340
rect 689 306 743 340
rect 639 291 743 306
rect 275 270 359 286
rect 207 236 241 260
rect 777 257 843 404
rect 493 236 843 257
rect 25 210 173 226
rect 25 176 139 210
rect 207 223 843 236
rect 207 202 572 223
rect 25 120 173 176
rect 484 199 572 202
rect 25 86 139 120
rect 25 70 173 86
rect 209 152 393 168
rect 209 118 225 152
rect 259 118 342 152
rect 376 118 393 152
rect 209 17 393 118
rect 484 165 511 199
rect 545 165 572 199
rect 772 218 843 223
rect 484 121 572 165
rect 484 87 511 121
rect 545 87 572 121
rect 484 75 572 87
rect 664 155 684 189
rect 718 155 738 189
rect 772 184 788 218
rect 822 184 843 218
rect 772 168 843 184
rect 664 121 738 155
rect 664 87 684 121
rect 718 87 738 121
rect 664 17 738 87
rect 773 85 839 134
rect 773 51 789 85
rect 823 51 839 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a221o_1
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 3996642
string GDS_START 3988170
<< end >>
