magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3122 1975
<< nwell >>
rect -38 331 1862 704
<< pwell >>
rect 1 49 1683 203
rect 0 0 1824 49
<< scnmos >>
rect 80 67 110 177
rect 152 67 182 177
rect 238 67 268 177
rect 310 67 340 177
rect 396 67 426 177
rect 468 67 498 177
rect 554 67 584 177
rect 626 67 656 177
rect 712 67 742 177
rect 784 67 814 177
rect 870 67 900 177
rect 942 67 972 177
rect 1028 67 1058 177
rect 1100 67 1130 177
rect 1186 67 1216 177
rect 1258 67 1288 177
rect 1344 67 1374 177
rect 1416 67 1446 177
rect 1502 67 1532 177
rect 1574 67 1604 177
<< scpmoshvt >>
rect 80 396 130 596
rect 186 396 236 596
rect 292 396 342 596
rect 398 396 448 596
rect 504 396 554 596
rect 610 396 660 596
rect 716 396 766 596
rect 822 396 872 596
rect 928 396 978 596
rect 1034 396 1084 596
rect 1140 396 1190 596
rect 1246 396 1296 596
rect 1352 396 1402 596
rect 1458 396 1508 596
rect 1564 396 1614 596
rect 1670 396 1720 596
<< ndiff >>
rect 27 139 80 177
rect 27 105 35 139
rect 69 105 80 139
rect 27 67 80 105
rect 110 67 152 177
rect 182 126 238 177
rect 182 92 193 126
rect 227 92 238 126
rect 182 67 238 92
rect 268 67 310 177
rect 340 139 396 177
rect 340 105 351 139
rect 385 105 396 139
rect 340 67 396 105
rect 426 67 468 177
rect 498 139 554 177
rect 498 105 509 139
rect 543 105 554 139
rect 498 67 554 105
rect 584 67 626 177
rect 656 139 712 177
rect 656 105 667 139
rect 701 105 712 139
rect 656 67 712 105
rect 742 67 784 177
rect 814 139 870 177
rect 814 105 825 139
rect 859 105 870 139
rect 814 67 870 105
rect 900 67 942 177
rect 972 139 1028 177
rect 972 105 983 139
rect 1017 105 1028 139
rect 972 67 1028 105
rect 1058 67 1100 177
rect 1130 139 1186 177
rect 1130 105 1141 139
rect 1175 105 1186 139
rect 1130 67 1186 105
rect 1216 67 1258 177
rect 1288 139 1344 177
rect 1288 105 1299 139
rect 1333 105 1344 139
rect 1288 67 1344 105
rect 1374 67 1416 177
rect 1446 139 1502 177
rect 1446 105 1457 139
rect 1491 105 1502 139
rect 1446 67 1502 105
rect 1532 67 1574 177
rect 1604 139 1657 177
rect 1604 105 1615 139
rect 1649 105 1657 139
rect 1604 67 1657 105
<< pdiff >>
rect 27 584 80 596
rect 27 550 35 584
rect 69 550 80 584
rect 27 513 80 550
rect 27 479 35 513
rect 69 479 80 513
rect 27 442 80 479
rect 27 408 35 442
rect 69 408 80 442
rect 27 396 80 408
rect 130 584 186 596
rect 130 550 141 584
rect 175 550 186 584
rect 130 513 186 550
rect 130 479 141 513
rect 175 479 186 513
rect 130 442 186 479
rect 130 408 141 442
rect 175 408 186 442
rect 130 396 186 408
rect 236 584 292 596
rect 236 550 247 584
rect 281 550 292 584
rect 236 513 292 550
rect 236 479 247 513
rect 281 479 292 513
rect 236 442 292 479
rect 236 408 247 442
rect 281 408 292 442
rect 236 396 292 408
rect 342 584 398 596
rect 342 550 353 584
rect 387 550 398 584
rect 342 513 398 550
rect 342 479 353 513
rect 387 479 398 513
rect 342 442 398 479
rect 342 408 353 442
rect 387 408 398 442
rect 342 396 398 408
rect 448 584 504 596
rect 448 550 459 584
rect 493 550 504 584
rect 448 513 504 550
rect 448 479 459 513
rect 493 479 504 513
rect 448 442 504 479
rect 448 408 459 442
rect 493 408 504 442
rect 448 396 504 408
rect 554 584 610 596
rect 554 550 565 584
rect 599 550 610 584
rect 554 513 610 550
rect 554 479 565 513
rect 599 479 610 513
rect 554 442 610 479
rect 554 408 565 442
rect 599 408 610 442
rect 554 396 610 408
rect 660 584 716 596
rect 660 550 671 584
rect 705 550 716 584
rect 660 513 716 550
rect 660 479 671 513
rect 705 479 716 513
rect 660 442 716 479
rect 660 408 671 442
rect 705 408 716 442
rect 660 396 716 408
rect 766 584 822 596
rect 766 550 777 584
rect 811 550 822 584
rect 766 513 822 550
rect 766 479 777 513
rect 811 479 822 513
rect 766 442 822 479
rect 766 408 777 442
rect 811 408 822 442
rect 766 396 822 408
rect 872 584 928 596
rect 872 550 883 584
rect 917 550 928 584
rect 872 513 928 550
rect 872 479 883 513
rect 917 479 928 513
rect 872 442 928 479
rect 872 408 883 442
rect 917 408 928 442
rect 872 396 928 408
rect 978 584 1034 596
rect 978 550 989 584
rect 1023 550 1034 584
rect 978 513 1034 550
rect 978 479 989 513
rect 1023 479 1034 513
rect 978 442 1034 479
rect 978 408 989 442
rect 1023 408 1034 442
rect 978 396 1034 408
rect 1084 584 1140 596
rect 1084 550 1095 584
rect 1129 550 1140 584
rect 1084 513 1140 550
rect 1084 479 1095 513
rect 1129 479 1140 513
rect 1084 442 1140 479
rect 1084 408 1095 442
rect 1129 408 1140 442
rect 1084 396 1140 408
rect 1190 584 1246 596
rect 1190 550 1201 584
rect 1235 550 1246 584
rect 1190 513 1246 550
rect 1190 479 1201 513
rect 1235 479 1246 513
rect 1190 442 1246 479
rect 1190 408 1201 442
rect 1235 408 1246 442
rect 1190 396 1246 408
rect 1296 584 1352 596
rect 1296 550 1307 584
rect 1341 550 1352 584
rect 1296 513 1352 550
rect 1296 479 1307 513
rect 1341 479 1352 513
rect 1296 442 1352 479
rect 1296 408 1307 442
rect 1341 408 1352 442
rect 1296 396 1352 408
rect 1402 584 1458 596
rect 1402 550 1413 584
rect 1447 550 1458 584
rect 1402 513 1458 550
rect 1402 479 1413 513
rect 1447 479 1458 513
rect 1402 442 1458 479
rect 1402 408 1413 442
rect 1447 408 1458 442
rect 1402 396 1458 408
rect 1508 584 1564 596
rect 1508 550 1519 584
rect 1553 550 1564 584
rect 1508 513 1564 550
rect 1508 479 1519 513
rect 1553 479 1564 513
rect 1508 442 1564 479
rect 1508 408 1519 442
rect 1553 408 1564 442
rect 1508 396 1564 408
rect 1614 584 1670 596
rect 1614 550 1625 584
rect 1659 550 1670 584
rect 1614 513 1670 550
rect 1614 479 1625 513
rect 1659 479 1670 513
rect 1614 442 1670 479
rect 1614 408 1625 442
rect 1659 408 1670 442
rect 1614 396 1670 408
rect 1720 584 1773 596
rect 1720 550 1731 584
rect 1765 550 1773 584
rect 1720 513 1773 550
rect 1720 479 1731 513
rect 1765 479 1773 513
rect 1720 442 1773 479
rect 1720 408 1731 442
rect 1765 408 1773 442
rect 1720 396 1773 408
<< ndiffc >>
rect 35 105 69 139
rect 193 92 227 126
rect 351 105 385 139
rect 509 105 543 139
rect 667 105 701 139
rect 825 105 859 139
rect 983 105 1017 139
rect 1141 105 1175 139
rect 1299 105 1333 139
rect 1457 105 1491 139
rect 1615 105 1649 139
<< pdiffc >>
rect 35 550 69 584
rect 35 479 69 513
rect 35 408 69 442
rect 141 550 175 584
rect 141 479 175 513
rect 141 408 175 442
rect 247 550 281 584
rect 247 479 281 513
rect 247 408 281 442
rect 353 550 387 584
rect 353 479 387 513
rect 353 408 387 442
rect 459 550 493 584
rect 459 479 493 513
rect 459 408 493 442
rect 565 550 599 584
rect 565 479 599 513
rect 565 408 599 442
rect 671 550 705 584
rect 671 479 705 513
rect 671 408 705 442
rect 777 550 811 584
rect 777 479 811 513
rect 777 408 811 442
rect 883 550 917 584
rect 883 479 917 513
rect 883 408 917 442
rect 989 550 1023 584
rect 989 479 1023 513
rect 989 408 1023 442
rect 1095 550 1129 584
rect 1095 479 1129 513
rect 1095 408 1129 442
rect 1201 550 1235 584
rect 1201 479 1235 513
rect 1201 408 1235 442
rect 1307 550 1341 584
rect 1307 479 1341 513
rect 1307 408 1341 442
rect 1413 550 1447 584
rect 1413 479 1447 513
rect 1413 408 1447 442
rect 1519 550 1553 584
rect 1519 479 1553 513
rect 1519 408 1553 442
rect 1625 550 1659 584
rect 1625 479 1659 513
rect 1625 408 1659 442
rect 1731 550 1765 584
rect 1731 479 1765 513
rect 1731 408 1765 442
<< poly >>
rect 80 596 130 622
rect 186 596 236 622
rect 292 596 342 622
rect 398 596 448 622
rect 504 596 554 622
rect 610 596 660 622
rect 716 596 766 622
rect 822 596 872 622
rect 928 596 978 622
rect 1034 596 1084 622
rect 1140 596 1190 622
rect 1246 596 1296 622
rect 1352 596 1402 622
rect 1458 596 1508 622
rect 1564 596 1614 622
rect 1670 596 1720 622
rect 80 316 130 396
rect 31 313 130 316
rect 186 313 236 396
rect 292 313 342 396
rect 398 313 448 396
rect 504 313 554 396
rect 610 313 660 396
rect 716 313 766 396
rect 822 313 872 396
rect 928 313 978 396
rect 1034 313 1084 396
rect 1140 313 1190 396
rect 1246 313 1296 396
rect 1352 313 1402 396
rect 1458 313 1508 396
rect 1564 313 1614 396
rect 1670 313 1720 396
rect 31 300 1743 313
rect 31 266 47 300
rect 81 297 1743 300
rect 81 266 246 297
rect 31 263 246 266
rect 280 263 314 297
rect 348 263 382 297
rect 416 263 671 297
rect 705 263 947 297
rect 981 263 1026 297
rect 1060 263 1290 297
rect 1324 263 1557 297
rect 1591 263 1625 297
rect 1659 263 1693 297
rect 1727 263 1743 297
rect 31 250 1743 263
rect 80 247 1743 250
rect 80 177 110 247
rect 152 177 182 247
rect 238 177 268 247
rect 310 177 340 247
rect 396 177 426 247
rect 468 177 498 247
rect 554 177 584 247
rect 626 177 656 247
rect 712 177 742 247
rect 784 177 814 247
rect 870 177 900 247
rect 942 177 972 247
rect 1028 177 1058 247
rect 1100 177 1130 247
rect 1186 177 1216 247
rect 1258 177 1288 247
rect 1344 177 1374 247
rect 1416 177 1446 247
rect 1502 177 1532 247
rect 1574 177 1604 247
rect 80 41 110 67
rect 152 41 182 67
rect 238 41 268 67
rect 310 41 340 67
rect 396 41 426 67
rect 468 41 498 67
rect 554 41 584 67
rect 626 41 656 67
rect 712 41 742 67
rect 784 41 814 67
rect 870 41 900 67
rect 942 41 972 67
rect 1028 41 1058 67
rect 1100 41 1130 67
rect 1186 41 1216 67
rect 1258 41 1288 67
rect 1344 41 1374 67
rect 1416 41 1446 67
rect 1502 41 1532 67
rect 1574 41 1604 67
<< polycont >>
rect 47 266 81 300
rect 246 263 280 297
rect 314 263 348 297
rect 382 263 416 297
rect 671 263 705 297
rect 947 263 981 297
rect 1026 263 1060 297
rect 1290 263 1324 297
rect 1557 263 1591 297
rect 1625 263 1659 297
rect 1693 263 1727 297
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 19 584 85 649
rect 19 550 35 584
rect 69 550 85 584
rect 19 513 85 550
rect 19 479 35 513
rect 69 479 85 513
rect 19 442 85 479
rect 19 408 35 442
rect 69 408 85 442
rect 19 392 85 408
rect 125 584 191 600
rect 125 550 141 584
rect 175 550 191 584
rect 125 513 191 550
rect 125 479 141 513
rect 175 479 191 513
rect 125 442 191 479
rect 125 424 141 442
rect 125 390 127 424
rect 175 408 191 442
rect 161 390 191 408
rect 231 584 297 649
rect 231 550 247 584
rect 281 550 297 584
rect 231 513 297 550
rect 231 479 247 513
rect 281 479 297 513
rect 231 442 297 479
rect 231 408 247 442
rect 281 408 297 442
rect 231 392 297 408
rect 337 584 403 600
rect 337 550 353 584
rect 387 550 403 584
rect 337 513 403 550
rect 337 479 353 513
rect 387 479 403 513
rect 337 442 403 479
rect 20 300 91 356
rect 20 276 47 300
rect 20 242 31 276
rect 81 266 91 300
rect 65 242 91 266
rect 20 221 91 242
rect 125 347 191 390
rect 337 390 353 442
rect 387 390 403 442
rect 443 584 509 649
rect 443 550 459 584
rect 493 550 509 584
rect 443 513 509 550
rect 443 479 459 513
rect 493 479 509 513
rect 443 442 509 479
rect 443 408 459 442
rect 493 408 509 442
rect 443 392 509 408
rect 549 584 615 600
rect 549 550 565 584
rect 599 550 615 584
rect 549 513 615 550
rect 549 479 565 513
rect 599 479 615 513
rect 549 442 615 479
rect 337 384 403 390
rect 549 390 565 442
rect 599 390 615 442
rect 655 584 721 649
rect 655 550 671 584
rect 705 550 721 584
rect 655 513 721 550
rect 655 479 671 513
rect 705 479 721 513
rect 655 442 721 479
rect 655 408 671 442
rect 705 408 721 442
rect 655 392 721 408
rect 761 584 827 600
rect 761 550 777 584
rect 811 550 827 584
rect 761 513 827 550
rect 761 479 777 513
rect 811 479 827 513
rect 761 442 827 479
rect 125 202 181 347
rect 549 313 615 390
rect 761 390 777 442
rect 811 390 827 442
rect 867 584 933 649
rect 867 550 883 584
rect 917 550 933 584
rect 867 513 933 550
rect 867 479 883 513
rect 917 479 933 513
rect 867 442 933 479
rect 867 408 883 442
rect 917 408 933 442
rect 867 392 933 408
rect 973 584 1039 600
rect 973 550 989 584
rect 1023 550 1039 584
rect 973 513 1039 550
rect 973 479 989 513
rect 1023 479 1039 513
rect 973 442 1039 479
rect 973 408 989 442
rect 1023 424 1039 442
rect 761 361 827 390
rect 973 390 991 408
rect 1025 390 1039 424
rect 1079 584 1145 649
rect 1079 550 1095 584
rect 1129 550 1145 584
rect 1079 513 1145 550
rect 1079 479 1095 513
rect 1129 479 1145 513
rect 1079 442 1145 479
rect 1079 408 1095 442
rect 1129 408 1145 442
rect 1079 392 1145 408
rect 1179 584 1251 600
rect 1179 550 1201 584
rect 1235 550 1251 584
rect 1179 513 1251 550
rect 1179 479 1201 513
rect 1235 479 1251 513
rect 1179 442 1251 479
rect 1179 424 1201 442
rect 973 384 1039 390
rect 1179 390 1183 424
rect 1235 408 1251 442
rect 1217 390 1251 408
rect 1291 584 1357 649
rect 1291 550 1307 584
rect 1341 550 1357 584
rect 1291 513 1357 550
rect 1291 479 1307 513
rect 1341 479 1357 513
rect 1291 442 1357 479
rect 1291 408 1307 442
rect 1341 408 1357 442
rect 1291 392 1357 408
rect 1397 584 1463 600
rect 1397 550 1413 584
rect 1447 550 1463 584
rect 1397 513 1463 550
rect 1397 479 1413 513
rect 1447 479 1463 513
rect 1397 442 1463 479
rect 776 313 827 361
rect 1179 375 1251 390
rect 1397 390 1413 442
rect 1447 390 1463 442
rect 1503 584 1569 649
rect 1503 550 1519 584
rect 1553 550 1569 584
rect 1503 513 1569 550
rect 1503 479 1519 513
rect 1553 479 1569 513
rect 1503 442 1569 479
rect 1503 408 1519 442
rect 1553 408 1569 442
rect 1503 392 1569 408
rect 1609 584 1675 600
rect 1609 550 1625 584
rect 1659 550 1675 584
rect 1609 513 1675 550
rect 1609 479 1625 513
rect 1659 479 1675 513
rect 1609 442 1675 479
rect 1179 313 1238 375
rect 1397 313 1463 390
rect 1609 390 1625 442
rect 1659 390 1675 442
rect 1715 584 1781 649
rect 1715 550 1731 584
rect 1765 550 1781 584
rect 1715 513 1781 550
rect 1715 479 1731 513
rect 1765 479 1781 513
rect 1715 442 1781 479
rect 1715 408 1731 442
rect 1765 408 1781 442
rect 1715 392 1781 408
rect 1609 384 1675 390
rect 215 297 453 313
rect 215 276 246 297
rect 215 242 223 276
rect 280 263 314 297
rect 348 276 382 297
rect 416 276 453 297
rect 353 263 382 276
rect 257 242 319 263
rect 353 242 415 263
rect 449 242 453 276
rect 215 236 453 242
rect 493 239 615 313
rect 655 297 742 313
rect 655 263 671 297
rect 705 276 742 297
rect 655 242 703 263
rect 737 242 742 276
rect 125 156 191 202
rect 19 139 85 155
rect 19 105 35 139
rect 69 105 85 139
rect 19 17 85 105
rect 125 126 243 156
rect 125 92 193 126
rect 227 92 243 126
rect 125 63 243 92
rect 335 139 401 155
rect 335 105 351 139
rect 385 105 401 139
rect 335 17 401 105
rect 493 139 559 239
rect 655 236 742 242
rect 776 239 875 313
rect 493 105 509 139
rect 543 105 559 139
rect 493 89 559 105
rect 651 139 717 155
rect 651 105 667 139
rect 701 105 717 139
rect 651 17 717 105
rect 809 139 875 239
rect 931 297 1076 313
rect 931 263 947 297
rect 981 276 1026 297
rect 981 263 991 276
rect 931 242 991 263
rect 1025 263 1026 276
rect 1060 263 1076 297
rect 1025 242 1076 263
rect 931 236 1076 242
rect 1125 239 1238 313
rect 1274 297 1340 313
rect 1274 276 1290 297
rect 1274 242 1279 276
rect 1324 263 1340 297
rect 1313 242 1340 263
rect 809 105 825 139
rect 859 105 875 139
rect 809 89 875 105
rect 967 139 1033 155
rect 967 105 983 139
rect 1017 105 1033 139
rect 967 17 1033 105
rect 1125 139 1191 239
rect 1274 236 1340 242
rect 1397 239 1507 313
rect 1125 105 1141 139
rect 1175 105 1191 139
rect 1125 89 1191 105
rect 1283 139 1349 155
rect 1283 105 1299 139
rect 1333 105 1349 139
rect 1283 17 1349 105
rect 1441 139 1507 239
rect 1541 297 1743 313
rect 1541 263 1557 297
rect 1591 276 1625 297
rect 1601 263 1625 276
rect 1659 276 1693 297
rect 1659 263 1663 276
rect 1727 263 1743 297
rect 1541 242 1567 263
rect 1601 242 1663 263
rect 1697 242 1743 263
rect 1541 236 1743 242
rect 1441 105 1457 139
rect 1491 105 1507 139
rect 1441 89 1507 105
rect 1599 139 1665 155
rect 1599 105 1615 139
rect 1649 105 1665 139
rect 1599 17 1665 105
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 127 408 141 424
rect 141 408 161 424
rect 127 390 161 408
rect 31 266 47 276
rect 47 266 65 276
rect 31 242 65 266
rect 353 408 387 424
rect 353 390 387 408
rect 565 408 599 424
rect 565 390 599 408
rect 777 408 811 424
rect 777 390 811 408
rect 991 408 1023 424
rect 1023 408 1025 424
rect 991 390 1025 408
rect 1183 408 1201 424
rect 1201 408 1217 424
rect 1183 390 1217 408
rect 1413 408 1447 424
rect 1413 390 1447 408
rect 1625 408 1659 424
rect 1625 390 1659 408
rect 223 263 246 276
rect 246 263 257 276
rect 319 263 348 276
rect 348 263 353 276
rect 415 263 416 276
rect 416 263 449 276
rect 223 242 257 263
rect 319 242 353 263
rect 415 242 449 263
rect 703 263 705 276
rect 705 263 737 276
rect 703 242 737 263
rect 991 242 1025 276
rect 1279 263 1290 276
rect 1290 263 1313 276
rect 1279 242 1313 263
rect 1567 263 1591 276
rect 1591 263 1601 276
rect 1663 263 1693 276
rect 1693 263 1697 276
rect 1567 242 1601 263
rect 1663 242 1697 263
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 115 424 1671 430
rect 115 390 127 424
rect 161 390 353 424
rect 387 390 565 424
rect 599 390 777 424
rect 811 390 991 424
rect 1025 390 1183 424
rect 1217 390 1413 424
rect 1447 390 1625 424
rect 1659 390 1671 424
rect 115 384 1671 390
rect 15 276 1709 282
rect 15 242 31 276
rect 65 242 223 276
rect 257 242 319 276
rect 353 242 415 276
rect 449 242 703 276
rect 737 242 991 276
rect 1025 242 1279 276
rect 1313 242 1567 276
rect 1601 242 1663 276
rect 1697 242 1709 276
rect 15 236 1709 242
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkinvlp_16
flabel metal1 s 115 384 1671 430 0 FreeSans 400 0 0 0 Y
port 6 nsew signal output
flabel metal1 s 15 236 1709 282 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2218814
string GDS_START 2205984
<< end >>
