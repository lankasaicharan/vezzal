magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 487 159 761 243
rect 46 49 761 159
rect 0 0 768 49
<< scnmos >>
rect 125 49 155 133
rect 197 49 227 133
rect 305 49 335 133
rect 413 49 443 133
rect 566 49 596 217
rect 652 49 682 217
<< scpmoshvt >>
rect 125 367 155 451
rect 211 367 241 451
rect 341 367 371 451
rect 427 367 457 451
rect 566 367 596 619
rect 652 367 682 619
<< ndiff >>
rect 513 133 566 217
rect 72 108 125 133
rect 72 74 80 108
rect 114 74 125 108
rect 72 49 125 74
rect 155 49 197 133
rect 227 49 305 133
rect 335 49 413 133
rect 443 95 566 133
rect 443 61 488 95
rect 522 61 566 95
rect 443 49 566 61
rect 596 205 652 217
rect 596 171 607 205
rect 641 171 652 205
rect 596 101 652 171
rect 596 67 607 101
rect 641 67 652 101
rect 596 49 652 67
rect 682 205 735 217
rect 682 171 693 205
rect 727 171 735 205
rect 682 95 735 171
rect 682 61 693 95
rect 727 61 735 95
rect 682 49 735 61
<< pdiff >>
rect 513 607 566 619
rect 513 573 521 607
rect 555 573 566 607
rect 513 516 566 573
rect 513 482 521 516
rect 555 482 566 516
rect 513 451 566 482
rect 72 426 125 451
rect 72 392 80 426
rect 114 392 125 426
rect 72 367 125 392
rect 155 434 211 451
rect 155 400 166 434
rect 200 400 211 434
rect 155 367 211 400
rect 241 439 341 451
rect 241 405 272 439
rect 306 405 341 439
rect 241 367 341 405
rect 371 426 427 451
rect 371 392 382 426
rect 416 392 427 426
rect 371 367 427 392
rect 457 439 566 451
rect 457 405 468 439
rect 502 405 566 439
rect 457 367 566 405
rect 596 599 652 619
rect 596 565 607 599
rect 641 565 652 599
rect 596 503 652 565
rect 596 469 607 503
rect 641 469 652 503
rect 596 413 652 469
rect 596 379 607 413
rect 641 379 652 413
rect 596 367 652 379
rect 682 607 735 619
rect 682 573 693 607
rect 727 573 735 607
rect 682 507 735 573
rect 682 473 693 507
rect 727 473 735 507
rect 682 413 735 473
rect 682 379 693 413
rect 727 379 735 413
rect 682 367 735 379
<< ndiffc >>
rect 80 74 114 108
rect 488 61 522 95
rect 607 171 641 205
rect 607 67 641 101
rect 693 171 727 205
rect 693 61 727 95
<< pdiffc >>
rect 521 573 555 607
rect 521 482 555 516
rect 80 392 114 426
rect 166 400 200 434
rect 272 405 306 439
rect 382 392 416 426
rect 468 405 502 439
rect 607 565 641 599
rect 607 469 641 503
rect 607 379 641 413
rect 693 573 727 607
rect 693 473 727 507
rect 693 379 727 413
<< poly >>
rect 566 619 596 645
rect 652 619 682 645
rect 125 451 155 477
rect 211 451 241 477
rect 341 451 371 477
rect 427 451 457 477
rect 125 335 155 367
rect 84 319 155 335
rect 211 319 241 367
rect 341 319 371 367
rect 427 319 457 367
rect 566 335 596 367
rect 652 335 682 367
rect 521 319 682 335
rect 84 285 100 319
rect 134 285 155 319
rect 84 251 155 285
rect 84 217 100 251
rect 134 217 155 251
rect 84 201 155 217
rect 125 133 155 201
rect 197 303 263 319
rect 197 269 213 303
rect 247 269 263 303
rect 197 235 263 269
rect 197 201 213 235
rect 247 201 263 235
rect 197 185 263 201
rect 305 303 371 319
rect 305 269 321 303
rect 355 269 371 303
rect 305 235 371 269
rect 305 201 321 235
rect 355 201 371 235
rect 305 185 371 201
rect 413 303 479 319
rect 413 269 429 303
rect 463 269 479 303
rect 521 285 537 319
rect 571 285 682 319
rect 521 269 682 285
rect 413 235 479 269
rect 413 201 429 235
rect 463 201 479 235
rect 566 217 596 269
rect 652 217 682 269
rect 413 185 479 201
rect 197 133 227 185
rect 305 133 335 185
rect 413 133 443 185
rect 125 23 155 49
rect 197 23 227 49
rect 305 23 335 49
rect 413 23 443 49
rect 566 23 596 49
rect 652 23 682 49
<< polycont >>
rect 100 285 134 319
rect 100 217 134 251
rect 213 269 247 303
rect 213 201 247 235
rect 321 269 355 303
rect 321 201 355 235
rect 429 269 463 303
rect 537 285 571 319
rect 429 201 463 235
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 64 426 130 649
rect 64 392 80 426
rect 114 392 130 426
rect 64 384 130 392
rect 164 434 216 452
rect 164 400 166 434
rect 200 400 216 434
rect 256 439 322 649
rect 452 607 571 649
rect 452 573 521 607
rect 555 573 571 607
rect 452 516 571 573
rect 452 482 521 516
rect 555 482 571 516
rect 256 405 272 439
rect 306 405 322 439
rect 366 426 418 442
rect 164 384 216 400
rect 168 371 216 384
rect 366 392 382 426
rect 416 392 418 426
rect 452 439 571 482
rect 452 405 468 439
rect 502 405 571 439
rect 605 599 651 615
rect 605 565 607 599
rect 641 565 651 599
rect 605 503 651 565
rect 605 469 607 503
rect 641 469 651 503
rect 605 413 651 469
rect 366 371 418 392
rect 605 379 607 413
rect 641 379 651 413
rect 17 319 134 350
rect 168 337 571 371
rect 17 285 100 319
rect 521 319 571 337
rect 17 251 134 285
rect 17 217 100 251
rect 17 201 134 217
rect 197 269 213 303
rect 247 269 271 303
rect 197 235 271 269
rect 197 201 213 235
rect 247 201 271 235
rect 305 269 321 303
rect 355 269 371 303
rect 305 235 371 269
rect 305 201 321 235
rect 355 201 371 235
rect 405 269 429 303
rect 463 269 479 303
rect 405 235 479 269
rect 405 201 429 235
rect 463 201 479 235
rect 521 285 537 319
rect 521 167 571 285
rect 64 133 571 167
rect 605 205 651 379
rect 685 607 743 649
rect 685 573 693 607
rect 727 573 743 607
rect 685 507 743 573
rect 685 473 693 507
rect 727 473 743 507
rect 685 413 743 473
rect 685 379 693 413
rect 727 379 743 413
rect 685 363 743 379
rect 605 171 607 205
rect 641 171 651 205
rect 64 108 130 133
rect 64 74 80 108
rect 114 74 130 108
rect 605 101 651 171
rect 64 58 130 74
rect 472 95 538 99
rect 472 61 488 95
rect 522 61 538 95
rect 472 17 538 61
rect 605 67 607 101
rect 641 67 651 101
rect 605 51 651 67
rect 685 205 743 221
rect 685 171 693 205
rect 727 171 743 205
rect 685 95 743 171
rect 685 61 693 95
rect 727 61 743 95
rect 685 17 743 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6278778
string GDS_START 6271606
<< end >>
