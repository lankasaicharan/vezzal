magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3986 1975
<< nwell >>
rect -38 331 2726 704
<< pwell >>
rect 1 254 322 289
rect 626 254 1235 281
rect 1 248 1235 254
rect 1740 273 2045 279
rect 1 241 1351 248
rect 1740 241 2403 273
rect 1 226 2403 241
rect 1 49 2687 226
rect 0 0 2688 49
<< scnmos >>
rect 84 95 114 263
rect 209 135 239 263
rect 413 60 443 228
rect 600 100 630 228
rect 957 127 987 255
rect 1043 127 1073 255
rect 1129 127 1159 255
rect 1238 94 1268 222
rect 1498 47 1528 215
rect 1823 125 1853 253
rect 1909 125 1939 253
rect 2041 119 2071 247
rect 2127 119 2157 247
rect 2236 79 2266 247
rect 2488 72 2518 200
rect 2574 72 2604 200
<< scpmoshvt >>
rect 84 367 114 619
rect 224 419 254 619
rect 528 367 558 619
rect 682 371 712 571
rect 814 436 844 604
rect 1022 414 1052 582
rect 1154 379 1184 547
rect 1287 379 1317 547
rect 1396 367 1426 619
rect 1814 367 1844 535
rect 1900 367 1930 535
rect 2025 367 2055 535
rect 2127 367 2157 535
rect 2229 367 2259 619
rect 2488 409 2518 609
rect 2574 409 2604 609
<< ndiff >>
rect 27 251 84 263
rect 27 217 39 251
rect 73 217 84 251
rect 27 141 84 217
rect 27 107 39 141
rect 73 107 84 141
rect 27 95 84 107
rect 114 135 209 263
rect 239 252 296 263
rect 239 218 250 252
rect 284 218 296 252
rect 239 135 296 218
rect 114 112 194 135
rect 114 95 148 112
rect 136 78 148 95
rect 182 78 194 112
rect 136 66 194 78
rect 652 243 710 255
rect 652 228 664 243
rect 356 112 413 228
rect 356 78 368 112
rect 402 78 413 112
rect 356 60 413 78
rect 443 112 600 228
rect 443 78 454 112
rect 488 100 600 112
rect 630 209 664 228
rect 698 209 710 243
rect 630 100 710 209
rect 878 127 957 255
rect 987 243 1043 255
rect 987 209 998 243
rect 1032 209 1043 243
rect 987 127 1043 209
rect 1073 228 1129 255
rect 1073 194 1084 228
rect 1118 194 1129 228
rect 1073 127 1129 194
rect 1159 222 1209 255
rect 1159 158 1238 222
rect 1159 127 1193 158
rect 488 78 500 100
rect 443 60 500 78
rect 878 87 935 127
rect 878 53 890 87
rect 924 53 935 87
rect 878 41 935 53
rect 1181 124 1193 127
rect 1227 124 1238 158
rect 1181 94 1238 124
rect 1268 191 1325 222
rect 1268 157 1279 191
rect 1313 157 1325 191
rect 1268 94 1325 157
rect 1766 241 1823 253
rect 1441 203 1498 215
rect 1441 169 1453 203
rect 1487 169 1498 203
rect 1441 103 1498 169
rect 1441 69 1453 103
rect 1487 69 1498 103
rect 1441 47 1498 69
rect 1528 109 1585 215
rect 1528 75 1539 109
rect 1573 75 1585 109
rect 1528 47 1585 75
rect 1766 207 1778 241
rect 1812 207 1823 241
rect 1766 173 1823 207
rect 1766 139 1778 173
rect 1812 139 1823 173
rect 1766 125 1823 139
rect 1853 241 1909 253
rect 1853 207 1864 241
rect 1898 207 1909 241
rect 1853 173 1909 207
rect 1853 139 1864 173
rect 1898 139 1909 173
rect 1853 125 1909 139
rect 1939 247 2019 253
rect 1939 182 2041 247
rect 1939 148 1973 182
rect 2007 148 2041 182
rect 1939 125 2041 148
rect 1961 119 2041 125
rect 2071 204 2127 247
rect 2071 170 2082 204
rect 2116 170 2127 204
rect 2071 119 2127 170
rect 2157 204 2236 247
rect 2157 170 2191 204
rect 2225 170 2236 204
rect 2157 119 2236 170
rect 2179 79 2236 119
rect 2266 118 2377 247
rect 2266 84 2331 118
rect 2365 84 2377 118
rect 2266 79 2377 84
rect 2288 72 2377 79
rect 2431 188 2488 200
rect 2431 154 2443 188
rect 2477 154 2488 188
rect 2431 118 2488 154
rect 2431 84 2443 118
rect 2477 84 2488 118
rect 2431 72 2488 84
rect 2518 188 2574 200
rect 2518 154 2529 188
rect 2563 154 2574 188
rect 2518 118 2574 154
rect 2518 84 2529 118
rect 2563 84 2574 118
rect 2518 72 2574 84
rect 2604 188 2661 200
rect 2604 154 2615 188
rect 2649 154 2661 188
rect 2604 118 2661 154
rect 2604 84 2615 118
rect 2649 84 2661 118
rect 2604 72 2661 84
<< pdiff >>
rect 573 627 631 639
rect 573 619 585 627
rect 27 597 84 619
rect 27 563 39 597
rect 73 563 84 597
rect 27 505 84 563
rect 27 471 39 505
rect 73 471 84 505
rect 27 413 84 471
rect 27 379 39 413
rect 73 379 84 413
rect 27 367 84 379
rect 114 607 224 619
rect 114 573 125 607
rect 159 573 224 607
rect 114 526 224 573
rect 114 492 125 526
rect 159 492 224 526
rect 114 419 224 492
rect 254 496 311 619
rect 254 462 265 496
rect 299 462 311 496
rect 254 419 311 462
rect 471 591 528 619
rect 471 557 483 591
rect 517 557 528 591
rect 114 367 164 419
rect 471 367 528 557
rect 558 593 585 619
rect 619 593 631 627
rect 558 571 631 593
rect 734 571 814 604
rect 558 371 682 571
rect 712 436 814 571
rect 844 582 894 604
rect 844 504 1022 582
rect 844 470 855 504
rect 889 470 1022 504
rect 844 436 1022 470
rect 712 417 792 436
rect 712 383 746 417
rect 780 383 792 417
rect 972 414 1022 436
rect 1052 570 1132 582
rect 1052 536 1086 570
rect 1120 547 1132 570
rect 1339 597 1396 619
rect 1339 563 1351 597
rect 1385 563 1396 597
rect 1339 547 1396 563
rect 1120 536 1154 547
rect 1052 414 1154 536
rect 712 371 792 383
rect 558 367 631 371
rect 1074 379 1154 414
rect 1184 521 1287 547
rect 1184 487 1195 521
rect 1229 487 1287 521
rect 1184 379 1287 487
rect 1317 519 1396 547
rect 1317 485 1351 519
rect 1385 485 1396 519
rect 1317 442 1396 485
rect 1317 408 1351 442
rect 1385 408 1396 442
rect 1317 379 1396 408
rect 1339 367 1396 379
rect 1426 607 1483 619
rect 1426 573 1437 607
rect 1471 573 1483 607
rect 2281 622 2370 634
rect 2281 619 2324 622
rect 1426 512 1483 573
rect 1426 478 1437 512
rect 1471 478 1483 512
rect 1426 367 1483 478
rect 1952 570 2010 582
rect 1952 536 1964 570
rect 1998 536 2010 570
rect 1952 535 2010 536
rect 2179 535 2229 619
rect 1741 523 1814 535
rect 1741 489 1753 523
rect 1787 489 1814 523
rect 1741 413 1814 489
rect 1741 379 1753 413
rect 1787 379 1814 413
rect 1741 367 1814 379
rect 1844 426 1900 535
rect 1844 392 1855 426
rect 1889 392 1900 426
rect 1844 367 1900 392
rect 1930 367 2025 535
rect 2055 413 2127 535
rect 2055 379 2066 413
rect 2100 379 2127 413
rect 2055 367 2127 379
rect 2157 463 2229 535
rect 2157 429 2168 463
rect 2202 429 2229 463
rect 2157 367 2229 429
rect 2259 588 2324 619
rect 2358 588 2370 622
rect 2259 367 2370 588
rect 2431 597 2488 609
rect 2431 563 2443 597
rect 2477 563 2488 597
rect 2431 462 2488 563
rect 2431 428 2443 462
rect 2477 428 2488 462
rect 2431 409 2488 428
rect 2518 597 2574 609
rect 2518 563 2529 597
rect 2563 563 2574 597
rect 2518 462 2574 563
rect 2518 428 2529 462
rect 2563 428 2574 462
rect 2518 409 2574 428
rect 2604 597 2661 609
rect 2604 563 2615 597
rect 2649 563 2661 597
rect 2604 526 2661 563
rect 2604 492 2615 526
rect 2649 492 2661 526
rect 2604 455 2661 492
rect 2604 421 2615 455
rect 2649 421 2661 455
rect 2604 409 2661 421
<< ndiffc >>
rect 39 217 73 251
rect 39 107 73 141
rect 250 218 284 252
rect 148 78 182 112
rect 368 78 402 112
rect 454 78 488 112
rect 664 209 698 243
rect 998 209 1032 243
rect 1084 194 1118 228
rect 890 53 924 87
rect 1193 124 1227 158
rect 1279 157 1313 191
rect 1453 169 1487 203
rect 1453 69 1487 103
rect 1539 75 1573 109
rect 1778 207 1812 241
rect 1778 139 1812 173
rect 1864 207 1898 241
rect 1864 139 1898 173
rect 1973 148 2007 182
rect 2082 170 2116 204
rect 2191 170 2225 204
rect 2331 84 2365 118
rect 2443 154 2477 188
rect 2443 84 2477 118
rect 2529 154 2563 188
rect 2529 84 2563 118
rect 2615 154 2649 188
rect 2615 84 2649 118
<< pdiffc >>
rect 39 563 73 597
rect 39 471 73 505
rect 39 379 73 413
rect 125 573 159 607
rect 125 492 159 526
rect 265 462 299 496
rect 483 557 517 591
rect 585 593 619 627
rect 855 470 889 504
rect 746 383 780 417
rect 1086 536 1120 570
rect 1351 563 1385 597
rect 1195 487 1229 521
rect 1351 485 1385 519
rect 1351 408 1385 442
rect 1437 573 1471 607
rect 1437 478 1471 512
rect 1964 536 1998 570
rect 1753 489 1787 523
rect 1753 379 1787 413
rect 1855 392 1889 426
rect 2066 379 2100 413
rect 2168 429 2202 463
rect 2324 588 2358 622
rect 2443 563 2477 597
rect 2443 428 2477 462
rect 2529 563 2563 597
rect 2529 428 2563 462
rect 2615 563 2649 597
rect 2615 492 2649 526
rect 2615 421 2649 455
<< poly >>
rect 84 619 114 645
rect 224 619 254 645
rect 528 619 558 645
rect 224 370 254 419
rect 335 414 439 430
rect 335 380 389 414
rect 423 380 439 414
rect 84 263 114 367
rect 197 354 263 370
rect 197 320 213 354
rect 247 320 263 354
rect 197 304 263 320
rect 335 364 439 380
rect 814 604 844 630
rect 1022 615 1317 645
rect 1396 619 1426 645
rect 682 571 712 597
rect 1022 582 1052 615
rect 814 414 844 436
rect 1154 547 1184 573
rect 1287 547 1317 615
rect 814 384 907 414
rect 209 263 239 304
rect 335 273 365 364
rect 528 316 558 367
rect 311 243 365 273
rect 413 300 558 316
rect 682 336 712 371
rect 682 320 829 336
rect 682 300 779 320
rect 413 266 491 300
rect 525 286 558 300
rect 600 286 779 300
rect 813 286 829 320
rect 525 266 541 286
rect 413 250 541 266
rect 600 270 829 286
rect 877 307 907 384
rect 1022 392 1052 414
rect 1022 364 1059 392
rect 1022 362 1073 364
rect 1029 334 1073 362
rect 1154 347 1184 379
rect 877 277 987 307
rect 84 51 114 95
rect 209 109 239 135
rect 311 51 341 243
rect 413 228 443 250
rect 600 228 630 270
rect 957 255 987 277
rect 1043 255 1073 334
rect 1115 331 1184 347
rect 1287 337 1317 379
rect 1577 609 2157 639
rect 2229 619 2259 645
rect 1577 592 1607 609
rect 1541 576 1607 592
rect 1541 542 1557 576
rect 1591 542 1607 576
rect 1541 508 1607 542
rect 1814 535 1844 561
rect 1900 535 1930 609
rect 2025 535 2055 561
rect 2127 535 2157 609
rect 1541 474 1557 508
rect 1591 474 1607 508
rect 1541 458 1607 474
rect 1115 297 1131 331
rect 1165 297 1184 331
rect 1115 281 1184 297
rect 1129 255 1159 281
rect 1238 267 1317 337
rect 1396 345 1426 367
rect 1541 345 1571 458
rect 2488 609 2518 635
rect 2574 609 2604 635
rect 2488 376 2518 409
rect 1396 315 1571 345
rect 1238 251 1417 267
rect 1238 237 1367 251
rect 1238 222 1268 237
rect 600 74 630 100
rect 84 21 341 51
rect 413 34 443 60
rect 957 53 987 127
rect 1043 101 1073 127
rect 1129 53 1159 127
rect 1351 217 1367 237
rect 1401 217 1417 251
rect 1351 183 1417 217
rect 1498 215 1528 315
rect 1814 305 1844 367
rect 1900 345 1930 367
rect 1900 315 1939 345
rect 1814 275 1853 305
rect 1823 253 1853 275
rect 1909 253 1939 315
rect 2025 299 2055 367
rect 2025 269 2071 299
rect 1351 149 1367 183
rect 1401 149 1417 183
rect 1351 133 1417 149
rect 1238 68 1268 94
rect 957 23 1159 53
rect 1607 196 1673 212
rect 1607 162 1623 196
rect 1657 162 1673 196
rect 1607 128 1673 162
rect 1607 94 1623 128
rect 1657 94 1673 128
rect 2041 247 2071 269
rect 2127 247 2157 367
rect 2229 335 2259 367
rect 2452 360 2518 376
rect 2229 319 2355 335
rect 2229 285 2305 319
rect 2339 285 2355 319
rect 2452 326 2468 360
rect 2502 340 2518 360
rect 2574 340 2604 409
rect 2502 326 2604 340
rect 2452 310 2604 326
rect 2229 269 2355 285
rect 2236 247 2266 269
rect 1607 51 1673 94
rect 1823 51 1853 125
rect 1909 99 1939 125
rect 2041 51 2071 119
rect 2127 93 2157 119
rect 2488 200 2518 310
rect 2574 200 2604 310
rect 2236 53 2266 79
rect 1498 21 1528 47
rect 1607 21 2071 51
rect 2488 46 2518 72
rect 2574 46 2604 72
<< polycont >>
rect 389 380 423 414
rect 213 320 247 354
rect 491 266 525 300
rect 779 286 813 320
rect 1557 542 1591 576
rect 1557 474 1591 508
rect 1131 297 1165 331
rect 1367 217 1401 251
rect 1367 149 1401 183
rect 1623 162 1657 196
rect 1623 94 1657 128
rect 2305 285 2339 319
rect 2468 326 2502 360
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 505 89 563
rect 23 471 39 505
rect 73 471 89 505
rect 125 607 159 649
rect 569 627 635 649
rect 125 526 159 573
rect 125 476 159 492
rect 195 591 517 613
rect 569 593 585 627
rect 619 593 635 627
rect 195 579 483 591
rect 23 413 89 471
rect 195 440 229 579
rect 467 557 483 579
rect 671 579 1315 613
rect 671 557 705 579
rect 23 379 39 413
rect 73 379 89 413
rect 23 251 89 379
rect 23 217 39 251
rect 73 217 89 251
rect 23 141 89 217
rect 127 406 229 440
rect 265 500 333 543
rect 467 536 517 557
rect 553 523 705 557
rect 941 570 1136 579
rect 553 500 587 523
rect 265 496 587 500
rect 299 466 587 496
rect 839 504 905 543
rect 839 487 855 504
rect 623 470 855 487
rect 889 470 905 504
rect 299 462 333 466
rect 265 415 333 462
rect 623 453 905 470
rect 623 430 657 453
rect 839 432 905 453
rect 941 536 1086 570
rect 1120 536 1136 570
rect 127 182 161 406
rect 197 354 263 370
rect 197 320 213 354
rect 247 320 263 354
rect 197 304 263 320
rect 299 268 333 415
rect 234 252 333 268
rect 234 218 250 252
rect 284 218 333 252
rect 373 414 657 430
rect 373 380 389 414
rect 423 396 657 414
rect 423 380 439 396
rect 373 204 439 380
rect 693 383 746 417
rect 780 383 796 417
rect 941 396 975 536
rect 1179 521 1245 543
rect 1179 500 1195 521
rect 693 356 727 383
rect 601 350 727 356
rect 601 316 607 350
rect 641 322 727 350
rect 832 362 975 396
rect 1011 487 1195 500
rect 1229 487 1245 521
rect 1011 466 1245 487
rect 832 336 866 362
rect 641 316 698 322
rect 475 300 541 316
rect 601 310 698 316
rect 475 266 491 300
rect 525 274 541 300
rect 525 266 628 274
rect 475 240 628 266
rect 127 148 337 182
rect 373 170 558 204
rect 23 107 39 141
rect 73 107 89 141
rect 303 134 337 148
rect 303 112 418 134
rect 23 88 89 107
rect 132 78 148 112
rect 182 78 198 112
rect 303 88 368 112
rect 132 17 198 78
rect 352 78 368 88
rect 402 78 418 112
rect 352 56 418 78
rect 454 112 488 134
rect 454 17 488 78
rect 524 87 558 170
rect 594 157 628 240
rect 664 243 698 310
rect 763 320 866 336
rect 763 286 779 320
rect 813 286 866 320
rect 1011 315 1045 466
rect 763 270 866 286
rect 998 281 1045 315
rect 1081 424 1173 430
rect 1281 426 1315 579
rect 1081 390 1087 424
rect 1121 390 1173 424
rect 1081 331 1173 390
rect 1081 297 1131 331
rect 1165 297 1173 331
rect 1081 281 1173 297
rect 1209 392 1315 426
rect 1351 597 1385 613
rect 1351 519 1385 563
rect 1351 442 1385 485
rect 1421 607 1487 649
rect 2324 622 2374 649
rect 1421 573 1437 607
rect 1471 573 1487 607
rect 1421 512 1487 573
rect 1421 478 1437 512
rect 1471 478 1487 512
rect 1421 462 1487 478
rect 1541 576 1607 592
rect 1541 542 1557 576
rect 1591 542 1607 576
rect 1541 508 1607 542
rect 1541 474 1557 508
rect 1591 474 1607 508
rect 1541 458 1607 474
rect 1667 575 2014 609
rect 1385 408 1487 426
rect 1351 392 1487 408
rect 998 259 1032 281
rect 982 243 1032 259
rect 1209 245 1243 392
rect 982 227 998 243
rect 664 193 698 209
rect 734 209 998 227
rect 734 193 1032 209
rect 1068 228 1243 245
rect 1068 194 1084 228
rect 1118 211 1243 228
rect 1279 350 1315 356
rect 1313 316 1315 350
rect 1118 194 1134 211
rect 1068 193 1134 194
rect 734 157 768 193
rect 1279 191 1315 316
rect 1177 158 1243 175
rect 1177 157 1193 158
rect 594 123 768 157
rect 804 124 1193 157
rect 1227 124 1243 158
rect 804 123 1243 124
rect 1313 157 1315 191
rect 1279 123 1315 157
rect 1351 350 1417 356
rect 1351 316 1375 350
rect 1409 316 1417 350
rect 1351 251 1417 316
rect 1351 217 1367 251
rect 1401 217 1417 251
rect 1351 183 1417 217
rect 1351 149 1367 183
rect 1401 149 1417 183
rect 1351 133 1417 149
rect 1453 212 1487 392
rect 1667 282 1701 575
rect 1948 570 2014 575
rect 2358 588 2374 622
rect 2324 572 2374 588
rect 2427 597 2493 613
rect 1737 523 1803 539
rect 1948 536 1964 570
rect 1998 536 2288 570
rect 2427 563 2443 597
rect 2477 563 2493 597
rect 2427 536 2493 563
rect 1737 489 1753 523
rect 1787 500 1803 523
rect 2254 502 2493 536
rect 1787 489 2218 500
rect 1737 466 2218 489
rect 1737 413 1803 466
rect 2152 463 2218 466
rect 1737 379 1753 413
rect 1787 379 1803 413
rect 1839 426 1984 430
rect 1839 390 1855 426
rect 1889 390 1984 426
rect 1839 388 1984 390
rect 1737 352 1803 379
rect 1737 318 1812 352
rect 1667 248 1742 282
rect 1453 203 1672 212
rect 1487 196 1672 203
rect 1487 178 1623 196
rect 804 87 838 123
rect 1453 103 1487 169
rect 1609 162 1623 178
rect 1657 162 1672 196
rect 524 53 838 87
rect 874 53 890 87
rect 924 69 1453 87
rect 924 53 1487 69
rect 1523 109 1573 142
rect 1523 75 1539 109
rect 1609 128 1672 162
rect 1609 94 1623 128
rect 1657 94 1672 128
rect 1609 78 1672 94
rect 1708 87 1742 248
rect 1778 241 1812 318
rect 1778 173 1812 207
rect 1778 123 1812 139
rect 1848 350 1914 352
rect 1848 316 1855 350
rect 1889 316 1914 350
rect 1848 241 1914 316
rect 1950 286 1984 388
rect 2050 413 2116 430
rect 2050 379 2066 413
rect 2100 379 2116 413
rect 2152 429 2168 463
rect 2202 429 2218 463
rect 2152 426 2218 429
rect 2427 462 2493 502
rect 2427 428 2443 462
rect 2477 428 2493 462
rect 2152 392 2253 426
rect 2427 412 2493 428
rect 2529 597 2563 649
rect 2529 462 2563 563
rect 2529 412 2563 428
rect 2599 597 2665 613
rect 2599 563 2615 597
rect 2649 563 2665 597
rect 2599 526 2665 563
rect 2599 492 2615 526
rect 2649 492 2665 526
rect 2599 455 2665 492
rect 2599 421 2615 455
rect 2649 421 2665 455
rect 2050 356 2116 379
rect 2050 350 2183 356
rect 2050 322 2143 350
rect 2137 316 2143 322
rect 2177 316 2183 350
rect 2137 310 2183 316
rect 1950 252 2100 286
rect 2219 274 2253 392
rect 2425 360 2518 376
rect 1848 207 1864 241
rect 1898 207 1914 241
rect 2066 251 2100 252
rect 1848 173 1914 207
rect 1848 139 1864 173
rect 1898 139 1914 173
rect 1848 123 1914 139
rect 1957 182 2023 216
rect 1957 148 1973 182
rect 2007 148 2023 182
rect 1957 87 2023 148
rect 2066 204 2132 251
rect 2066 170 2082 204
rect 2116 170 2132 204
rect 2066 123 2132 170
rect 2175 240 2253 274
rect 2289 319 2355 335
rect 2289 285 2305 319
rect 2339 285 2355 319
rect 2425 326 2468 360
rect 2502 326 2518 360
rect 2425 310 2518 326
rect 2289 274 2355 285
rect 2599 274 2665 421
rect 2289 240 2665 274
rect 2175 204 2225 240
rect 2175 170 2191 204
rect 2175 123 2225 170
rect 2261 188 2493 204
rect 2261 170 2443 188
rect 2261 87 2295 170
rect 2427 154 2443 170
rect 2477 154 2493 188
rect 1523 17 1573 75
rect 1708 53 2295 87
rect 2331 118 2381 134
rect 2365 84 2381 118
rect 2331 17 2381 84
rect 2427 118 2493 154
rect 2427 84 2443 118
rect 2477 84 2493 118
rect 2427 68 2493 84
rect 2529 188 2563 204
rect 2529 118 2563 154
rect 2529 17 2563 84
rect 2599 188 2665 240
rect 2599 154 2615 188
rect 2649 154 2665 188
rect 2599 118 2665 154
rect 2599 84 2615 118
rect 2649 84 2665 118
rect 2599 68 2665 84
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 607 316 641 350
rect 1087 390 1121 424
rect 1279 316 1313 350
rect 1375 316 1409 350
rect 1855 392 1889 424
rect 1855 390 1889 392
rect 1855 316 1889 350
rect 2143 316 2177 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 1843 424 1901 430
rect 1843 421 1855 424
rect 1121 393 1855 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1843 390 1855 393
rect 1889 390 1901 424
rect 1843 384 1901 390
rect 595 350 653 356
rect 595 316 607 350
rect 641 347 653 350
rect 1267 350 1325 356
rect 1267 347 1279 350
rect 641 319 1279 347
rect 641 316 653 319
rect 595 310 653 316
rect 1267 316 1279 319
rect 1313 316 1325 350
rect 1267 310 1325 316
rect 1363 350 1421 356
rect 1363 316 1375 350
rect 1409 347 1421 350
rect 1843 350 1901 356
rect 1843 347 1855 350
rect 1409 319 1855 347
rect 1409 316 1421 319
rect 1363 310 1421 316
rect 1843 316 1855 319
rect 1889 347 1901 350
rect 2131 350 2189 356
rect 2131 347 2143 350
rect 1889 319 2143 347
rect 1889 316 1901 319
rect 1843 310 1901 316
rect 2131 316 2143 319
rect 2177 316 2189 350
rect 2131 310 2189 316
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
flabel pwell s 0 0 2688 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2688 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fah_1
flabel metal1 s 0 617 2688 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2688 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 CI
port 3 nsew signal input
flabel locali s 2431 316 2465 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2688 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6500174
string GDS_START 6481674
<< end >>
