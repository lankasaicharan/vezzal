magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 742 241
rect 0 0 768 49
<< scnmos >>
rect 80 47 110 215
rect 237 47 267 215
rect 336 47 366 215
rect 453 47 483 215
rect 561 47 591 215
rect 633 47 663 215
<< scpmoshvt >>
rect 129 367 159 619
rect 237 367 267 619
rect 326 367 356 619
rect 417 367 447 619
rect 525 367 555 619
rect 633 367 663 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 101 80 169
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 203 237 215
rect 110 169 133 203
rect 167 169 237 203
rect 110 93 237 169
rect 110 59 133 93
rect 167 59 237 93
rect 110 47 237 59
rect 267 187 336 215
rect 267 153 291 187
rect 325 153 336 187
rect 267 101 336 153
rect 267 67 291 101
rect 325 67 336 101
rect 267 47 336 67
rect 366 127 453 215
rect 366 93 393 127
rect 427 93 453 127
rect 366 47 453 93
rect 483 203 561 215
rect 483 169 506 203
rect 540 169 561 203
rect 483 93 561 169
rect 483 59 506 93
rect 540 59 561 93
rect 483 47 561 59
rect 591 47 633 215
rect 663 203 716 215
rect 663 169 674 203
rect 708 169 716 203
rect 663 93 716 169
rect 663 59 674 93
rect 708 59 716 93
rect 663 47 716 59
<< pdiff >>
rect 76 607 129 619
rect 76 573 84 607
rect 118 573 129 607
rect 76 529 129 573
rect 76 495 84 529
rect 118 495 129 529
rect 76 443 129 495
rect 76 409 84 443
rect 118 409 129 443
rect 76 367 129 409
rect 159 607 237 619
rect 159 573 184 607
rect 218 573 237 607
rect 159 529 237 573
rect 159 495 184 529
rect 218 495 237 529
rect 159 443 237 495
rect 159 409 184 443
rect 218 409 237 443
rect 159 367 237 409
rect 267 367 326 619
rect 356 367 417 619
rect 447 599 525 619
rect 447 565 468 599
rect 502 565 525 599
rect 447 507 525 565
rect 447 473 468 507
rect 502 473 525 507
rect 447 413 525 473
rect 447 379 468 413
rect 502 379 525 413
rect 447 367 525 379
rect 555 607 633 619
rect 555 573 576 607
rect 610 573 633 607
rect 555 529 633 573
rect 555 495 576 529
rect 610 495 633 529
rect 555 443 633 495
rect 555 409 576 443
rect 610 409 633 443
rect 555 367 633 409
rect 663 599 722 619
rect 663 565 680 599
rect 714 565 722 599
rect 663 507 722 565
rect 663 473 680 507
rect 714 473 722 507
rect 663 413 722 473
rect 663 379 680 413
rect 714 379 722 413
rect 663 367 722 379
<< ndiffc >>
rect 35 169 69 203
rect 35 67 69 101
rect 133 169 167 203
rect 133 59 167 93
rect 291 153 325 187
rect 291 67 325 101
rect 393 93 427 127
rect 506 169 540 203
rect 506 59 540 93
rect 674 169 708 203
rect 674 59 708 93
<< pdiffc >>
rect 84 573 118 607
rect 84 495 118 529
rect 84 409 118 443
rect 184 573 218 607
rect 184 495 218 529
rect 184 409 218 443
rect 468 565 502 599
rect 468 473 502 507
rect 468 379 502 413
rect 576 573 610 607
rect 576 495 610 529
rect 576 409 610 443
rect 680 565 714 599
rect 680 473 714 507
rect 680 379 714 413
<< poly >>
rect 129 619 159 645
rect 237 619 267 645
rect 326 619 356 645
rect 417 619 447 645
rect 525 619 555 645
rect 633 619 663 645
rect 129 335 159 367
rect 80 319 159 335
rect 80 285 109 319
rect 143 285 159 319
rect 237 303 267 367
rect 326 303 356 367
rect 417 303 447 367
rect 525 303 555 367
rect 633 305 663 367
rect 80 269 159 285
rect 201 287 267 303
rect 80 215 110 269
rect 201 253 217 287
rect 251 253 267 287
rect 201 237 267 253
rect 309 287 375 303
rect 309 253 325 287
rect 359 253 375 287
rect 309 237 375 253
rect 417 287 483 303
rect 417 253 433 287
rect 467 253 483 287
rect 417 237 483 253
rect 525 287 591 303
rect 525 253 541 287
rect 575 253 591 287
rect 525 237 591 253
rect 237 215 267 237
rect 336 215 366 237
rect 453 215 483 237
rect 561 215 591 237
rect 633 289 735 305
rect 633 255 685 289
rect 719 255 735 289
rect 633 239 735 255
rect 633 215 663 239
rect 80 21 110 47
rect 237 21 267 47
rect 336 21 366 47
rect 453 21 483 47
rect 561 21 591 47
rect 633 21 663 47
<< polycont >>
rect 109 285 143 319
rect 217 253 251 287
rect 325 253 359 287
rect 433 253 467 287
rect 541 253 575 287
rect 685 255 719 289
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 19 607 134 615
rect 19 573 84 607
rect 118 573 134 607
rect 19 529 134 573
rect 19 495 84 529
rect 118 495 134 529
rect 19 443 134 495
rect 19 409 84 443
rect 118 409 134 443
rect 168 607 234 649
rect 168 573 184 607
rect 218 573 234 607
rect 168 529 234 573
rect 168 495 184 529
rect 218 495 234 529
rect 168 443 234 495
rect 168 409 184 443
rect 218 409 234 443
rect 452 599 518 615
rect 452 565 468 599
rect 502 565 518 599
rect 452 507 518 565
rect 452 473 468 507
rect 502 473 518 507
rect 452 413 518 473
rect 19 203 73 409
rect 452 379 468 413
rect 502 379 518 413
rect 560 607 626 649
rect 560 573 576 607
rect 610 573 626 607
rect 560 529 626 573
rect 560 495 576 529
rect 610 495 626 529
rect 560 443 626 495
rect 560 409 576 443
rect 610 409 626 443
rect 676 599 730 615
rect 676 565 680 599
rect 714 565 730 599
rect 676 507 730 565
rect 676 473 680 507
rect 714 473 730 507
rect 676 413 730 473
rect 452 375 518 379
rect 676 379 680 413
rect 714 379 730 413
rect 676 375 730 379
rect 107 341 730 375
rect 107 319 159 341
rect 107 285 109 319
rect 143 285 159 319
rect 107 269 159 285
rect 217 287 269 303
rect 409 287 467 303
rect 251 253 269 287
rect 217 237 269 253
rect 303 253 325 287
rect 359 253 375 287
rect 303 237 375 253
rect 409 253 433 287
rect 409 237 467 253
rect 501 287 575 303
rect 501 253 541 287
rect 501 237 575 253
rect 19 169 35 203
rect 69 169 73 203
rect 19 101 73 169
rect 19 67 35 101
rect 69 67 73 101
rect 19 51 73 67
rect 117 203 183 219
rect 117 169 133 203
rect 167 169 183 203
rect 117 93 183 169
rect 117 59 133 93
rect 167 59 183 93
rect 217 76 257 237
rect 615 203 649 341
rect 685 289 750 305
rect 719 255 750 289
rect 685 239 750 255
rect 291 187 506 203
rect 325 169 506 187
rect 540 169 556 203
rect 325 153 335 169
rect 291 101 335 153
rect 117 17 183 59
rect 325 67 335 101
rect 291 51 335 67
rect 377 127 443 135
rect 377 93 393 127
rect 427 93 443 127
rect 377 17 443 93
rect 490 93 556 169
rect 490 59 506 93
rect 540 59 556 93
rect 490 51 556 59
rect 615 169 674 203
rect 708 169 724 203
rect 615 93 724 169
rect 615 59 674 93
rect 708 59 724 93
rect 615 51 724 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o311a_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4406688
string GDS_START 4398958
<< end >>
