magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2218 1852
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 157 292 203
rect 1 21 899 157
rect 27 -17 61 21
<< scnmos >>
rect 84 47 114 177
rect 178 47 208 177
rect 283 47 313 131
rect 389 47 419 131
rect 597 47 627 131
rect 695 47 725 131
rect 790 47 820 131
<< scpmoshvt >>
rect 86 297 122 497
rect 180 297 216 497
rect 285 369 321 497
rect 407 369 443 497
rect 589 369 625 497
rect 687 369 723 497
rect 792 369 828 497
<< ndiff >>
rect 27 159 84 177
rect 27 125 39 159
rect 73 125 84 159
rect 27 91 84 125
rect 27 57 39 91
rect 73 57 84 91
rect 27 47 84 57
rect 114 159 178 177
rect 114 125 134 159
rect 168 125 178 159
rect 114 91 178 125
rect 114 57 134 91
rect 168 57 178 91
rect 114 47 178 57
rect 208 131 266 177
rect 208 122 283 131
rect 208 88 227 122
rect 261 88 283 122
rect 208 47 283 88
rect 313 47 389 131
rect 419 113 479 131
rect 419 79 437 113
rect 471 79 479 113
rect 419 47 479 79
rect 539 114 597 131
rect 539 80 547 114
rect 581 80 597 114
rect 539 47 597 80
rect 627 114 695 131
rect 627 80 641 114
rect 675 80 695 114
rect 627 47 695 80
rect 725 95 790 131
rect 725 61 735 95
rect 769 61 790 95
rect 725 47 790 61
rect 820 104 873 131
rect 820 70 831 104
rect 865 70 873 104
rect 820 47 873 70
<< pdiff >>
rect 27 477 86 497
rect 27 443 39 477
rect 73 443 86 477
rect 27 409 86 443
rect 27 375 39 409
rect 73 375 86 409
rect 27 341 86 375
rect 27 307 39 341
rect 73 307 86 341
rect 27 297 86 307
rect 122 477 180 497
rect 122 443 134 477
rect 168 443 180 477
rect 122 409 180 443
rect 122 375 134 409
rect 168 375 180 409
rect 122 297 180 375
rect 216 481 285 497
rect 216 447 228 481
rect 262 447 285 481
rect 216 369 285 447
rect 321 369 407 497
rect 443 481 589 497
rect 443 447 496 481
rect 530 447 589 481
rect 443 369 589 447
rect 625 485 687 497
rect 625 451 637 485
rect 671 451 687 485
rect 625 417 687 451
rect 625 383 637 417
rect 671 383 687 417
rect 625 369 687 383
rect 723 369 792 497
rect 828 485 884 497
rect 828 451 842 485
rect 876 451 884 485
rect 828 417 884 451
rect 828 383 842 417
rect 876 383 884 417
rect 828 369 884 383
rect 216 297 268 369
rect 340 343 390 369
rect 340 309 348 343
rect 382 309 390 343
rect 340 297 390 309
<< ndiffc >>
rect 39 125 73 159
rect 39 57 73 91
rect 134 125 168 159
rect 134 57 168 91
rect 227 88 261 122
rect 437 79 471 113
rect 547 80 581 114
rect 641 80 675 114
rect 735 61 769 95
rect 831 70 865 104
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 134 443 168 477
rect 134 375 168 409
rect 228 447 262 481
rect 496 447 530 481
rect 637 451 671 485
rect 637 383 671 417
rect 842 451 876 485
rect 842 383 876 417
rect 348 309 382 343
<< poly >>
rect 86 497 122 523
rect 180 497 216 523
rect 285 497 321 523
rect 407 497 443 523
rect 589 497 625 523
rect 687 497 723 523
rect 792 497 828 523
rect 285 354 321 369
rect 86 282 122 297
rect 180 282 216 297
rect 84 265 124 282
rect 178 265 218 282
rect 283 265 323 354
rect 407 354 443 369
rect 589 354 625 369
rect 687 354 723 369
rect 792 354 828 369
rect 84 249 239 265
rect 84 215 185 249
rect 219 215 239 249
rect 84 199 239 215
rect 283 249 347 265
rect 283 215 293 249
rect 327 215 347 249
rect 405 220 445 354
rect 587 337 627 354
rect 488 321 627 337
rect 488 287 498 321
rect 532 287 627 321
rect 488 271 627 287
rect 283 199 347 215
rect 389 204 455 220
rect 84 177 114 199
rect 178 177 208 199
rect 283 131 313 199
rect 389 170 401 204
rect 435 170 455 204
rect 389 154 455 170
rect 389 131 419 154
rect 597 131 627 271
rect 685 265 725 354
rect 790 265 830 354
rect 673 249 737 265
rect 673 215 683 249
rect 717 215 737 249
rect 673 199 737 215
rect 790 249 875 265
rect 790 215 826 249
rect 860 215 875 249
rect 790 199 875 215
rect 695 131 725 199
rect 790 131 820 199
rect 84 21 114 47
rect 178 21 208 47
rect 283 21 313 47
rect 389 21 419 47
rect 597 21 627 47
rect 695 21 725 47
rect 790 21 820 47
<< polycont >>
rect 185 215 219 249
rect 293 215 327 249
rect 498 287 532 321
rect 401 170 435 204
rect 683 215 717 249
rect 826 215 860 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 22 477 73 527
rect 22 443 39 477
rect 22 409 73 443
rect 22 375 39 409
rect 22 341 73 375
rect 22 307 39 341
rect 22 282 73 307
rect 107 477 168 493
rect 107 443 134 477
rect 202 481 278 527
rect 202 447 228 481
rect 262 447 278 481
rect 472 481 553 527
rect 833 485 896 527
rect 472 447 496 481
rect 530 447 553 481
rect 607 451 637 485
rect 671 451 687 485
rect 107 409 168 443
rect 607 417 687 451
rect 607 411 637 417
rect 107 375 134 409
rect 107 359 168 375
rect 240 383 637 411
rect 671 383 687 417
rect 240 377 687 383
rect 22 159 73 182
rect 22 125 39 159
rect 22 91 73 125
rect 22 57 39 91
rect 22 17 73 57
rect 107 165 151 359
rect 240 323 274 377
rect 185 289 274 323
rect 308 309 348 343
rect 382 321 532 343
rect 382 309 498 321
rect 308 299 498 309
rect 185 249 229 289
rect 479 287 498 299
rect 479 271 532 287
rect 566 299 687 377
rect 731 383 799 485
rect 833 451 842 485
rect 876 451 896 485
rect 833 417 896 451
rect 833 383 842 417
rect 876 383 896 417
rect 219 215 229 249
rect 263 249 367 255
rect 263 215 293 249
rect 327 215 367 249
rect 185 199 229 215
rect 401 204 445 220
rect 304 170 401 181
rect 435 170 445 204
rect 107 159 184 165
rect 107 125 134 159
rect 168 125 184 159
rect 107 91 184 125
rect 107 57 134 91
rect 168 57 184 91
rect 107 51 184 57
rect 227 122 261 150
rect 227 17 261 88
rect 304 147 445 170
rect 304 76 377 147
rect 479 113 513 271
rect 566 249 600 299
rect 731 265 765 383
rect 833 363 896 383
rect 562 215 600 249
rect 644 249 765 265
rect 644 215 683 249
rect 717 215 765 249
rect 800 249 893 329
rect 800 215 826 249
rect 860 215 893 249
rect 562 138 596 215
rect 411 79 437 113
rect 471 79 513 113
rect 547 114 596 138
rect 581 80 596 114
rect 547 64 596 80
rect 641 145 881 181
rect 641 114 687 145
rect 675 80 687 114
rect 641 64 687 80
rect 735 95 769 111
rect 803 104 881 145
rect 803 70 831 104
rect 865 70 881 104
rect 803 64 881 70
rect 735 17 769 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 305 219 339 253 0 FreeSans 400 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 122 425 156 459 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 311 85 345 119 0 FreeSans 400 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 675 216 709 250 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 833 221 867 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 761 425 795 459 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 833 289 867 323 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel pwell s 27 -17 61 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 27 527 61 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 27 -17 61 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 27 527 61 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2bb2a_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2547724
string GDS_START 2540152
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
