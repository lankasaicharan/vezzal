magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 22 49 1604 248
rect 0 0 1632 49
<< scpmos >>
rect 97 368 133 592
rect 187 368 223 592
rect 277 368 313 592
rect 367 368 403 592
rect 457 368 493 592
rect 547 368 583 592
rect 637 368 673 592
rect 727 368 763 592
rect 817 368 853 592
rect 907 368 943 592
rect 997 368 1033 592
rect 1133 368 1169 592
rect 1223 368 1259 592
rect 1313 368 1349 592
rect 1403 368 1439 592
rect 1493 368 1529 592
<< nmoslvt >>
rect 101 74 131 222
rect 187 74 217 222
rect 273 74 303 222
rect 359 74 389 222
rect 445 74 475 222
rect 531 74 561 222
rect 617 74 647 222
rect 703 74 733 222
rect 893 74 923 222
rect 979 74 1009 222
rect 1065 74 1095 222
rect 1151 74 1181 222
rect 1237 74 1267 222
rect 1323 74 1353 222
rect 1409 74 1439 222
rect 1495 74 1525 222
<< ndiff >>
rect 48 210 101 222
rect 48 176 56 210
rect 90 176 101 210
rect 48 120 101 176
rect 48 86 56 120
rect 90 86 101 120
rect 48 74 101 86
rect 131 152 187 222
rect 131 118 142 152
rect 176 118 187 152
rect 131 74 187 118
rect 217 210 273 222
rect 217 176 228 210
rect 262 176 273 210
rect 217 120 273 176
rect 217 86 228 120
rect 262 86 273 120
rect 217 74 273 86
rect 303 152 359 222
rect 303 118 314 152
rect 348 118 359 152
rect 303 74 359 118
rect 389 210 445 222
rect 389 176 400 210
rect 434 176 445 210
rect 389 120 445 176
rect 389 86 400 120
rect 434 86 445 120
rect 389 74 445 86
rect 475 169 531 222
rect 475 135 486 169
rect 520 135 531 169
rect 475 74 531 135
rect 561 136 617 222
rect 561 102 572 136
rect 606 102 617 136
rect 561 74 617 102
rect 647 199 703 222
rect 647 165 658 199
rect 692 165 703 199
rect 647 74 703 165
rect 733 120 786 222
rect 733 86 744 120
rect 778 86 786 120
rect 733 74 786 86
rect 840 120 893 222
rect 840 86 848 120
rect 882 86 893 120
rect 840 74 893 86
rect 923 207 979 222
rect 923 173 934 207
rect 968 173 979 207
rect 923 74 979 173
rect 1009 120 1065 222
rect 1009 86 1020 120
rect 1054 86 1065 120
rect 1009 74 1065 86
rect 1095 207 1151 222
rect 1095 173 1106 207
rect 1140 173 1151 207
rect 1095 74 1151 173
rect 1181 210 1237 222
rect 1181 176 1192 210
rect 1226 176 1237 210
rect 1181 120 1237 176
rect 1181 86 1192 120
rect 1226 86 1237 120
rect 1181 74 1237 86
rect 1267 136 1323 222
rect 1267 102 1278 136
rect 1312 102 1323 136
rect 1267 74 1323 102
rect 1353 210 1409 222
rect 1353 176 1364 210
rect 1398 176 1409 210
rect 1353 120 1409 176
rect 1353 86 1364 120
rect 1398 86 1409 120
rect 1353 74 1409 86
rect 1439 136 1495 222
rect 1439 102 1450 136
rect 1484 102 1495 136
rect 1439 74 1495 102
rect 1525 210 1578 222
rect 1525 176 1536 210
rect 1570 176 1578 210
rect 1525 120 1578 176
rect 1525 86 1536 120
rect 1570 86 1578 120
rect 1525 74 1578 86
<< pdiff >>
rect 45 580 97 592
rect 45 546 53 580
rect 87 546 97 580
rect 45 497 97 546
rect 45 463 53 497
rect 87 463 97 497
rect 45 414 97 463
rect 45 380 53 414
rect 87 380 97 414
rect 45 368 97 380
rect 133 531 187 592
rect 133 497 143 531
rect 177 497 187 531
rect 133 424 187 497
rect 133 390 143 424
rect 177 390 187 424
rect 133 368 187 390
rect 223 580 277 592
rect 223 546 233 580
rect 267 546 277 580
rect 223 492 277 546
rect 223 458 233 492
rect 267 458 277 492
rect 223 368 277 458
rect 313 531 367 592
rect 313 497 323 531
rect 357 497 367 531
rect 313 424 367 497
rect 313 390 323 424
rect 357 390 367 424
rect 313 368 367 390
rect 403 580 457 592
rect 403 546 413 580
rect 447 546 457 580
rect 403 492 457 546
rect 403 458 413 492
rect 447 458 457 492
rect 403 368 457 458
rect 493 531 547 592
rect 493 497 503 531
rect 537 497 547 531
rect 493 424 547 497
rect 493 390 503 424
rect 537 390 547 424
rect 493 368 547 390
rect 583 580 637 592
rect 583 546 593 580
rect 627 546 637 580
rect 583 492 637 546
rect 583 458 593 492
rect 627 458 637 492
rect 583 368 637 458
rect 673 531 727 592
rect 673 497 683 531
rect 717 497 727 531
rect 673 440 727 497
rect 673 406 683 440
rect 717 406 727 440
rect 673 368 727 406
rect 763 580 817 592
rect 763 546 773 580
rect 807 546 817 580
rect 763 497 817 546
rect 763 463 773 497
rect 807 463 817 497
rect 763 414 817 463
rect 763 380 773 414
rect 807 380 817 414
rect 763 368 817 380
rect 853 580 907 592
rect 853 546 863 580
rect 897 546 907 580
rect 853 492 907 546
rect 853 458 863 492
rect 897 458 907 492
rect 853 368 907 458
rect 943 580 997 592
rect 943 546 953 580
rect 987 546 997 580
rect 943 500 997 546
rect 943 466 953 500
rect 987 466 997 500
rect 943 424 997 466
rect 943 390 953 424
rect 987 390 997 424
rect 943 368 997 390
rect 1033 580 1133 592
rect 1033 546 1066 580
rect 1100 546 1133 580
rect 1033 492 1133 546
rect 1033 458 1066 492
rect 1100 458 1133 492
rect 1033 368 1133 458
rect 1169 580 1223 592
rect 1169 546 1179 580
rect 1213 546 1223 580
rect 1169 510 1223 546
rect 1169 476 1179 510
rect 1213 476 1223 510
rect 1169 424 1223 476
rect 1169 390 1179 424
rect 1213 390 1223 424
rect 1169 368 1223 390
rect 1259 580 1313 592
rect 1259 546 1269 580
rect 1303 546 1313 580
rect 1259 492 1313 546
rect 1259 458 1269 492
rect 1303 458 1313 492
rect 1259 368 1313 458
rect 1349 580 1403 592
rect 1349 546 1359 580
rect 1393 546 1403 580
rect 1349 510 1403 546
rect 1349 476 1359 510
rect 1393 476 1403 510
rect 1349 424 1403 476
rect 1349 390 1359 424
rect 1393 390 1403 424
rect 1349 368 1403 390
rect 1439 580 1493 592
rect 1439 546 1449 580
rect 1483 546 1493 580
rect 1439 492 1493 546
rect 1439 458 1449 492
rect 1483 458 1493 492
rect 1439 368 1493 458
rect 1529 580 1581 592
rect 1529 546 1539 580
rect 1573 546 1581 580
rect 1529 497 1581 546
rect 1529 463 1539 497
rect 1573 463 1581 497
rect 1529 414 1581 463
rect 1529 380 1539 414
rect 1573 380 1581 414
rect 1529 368 1581 380
<< ndiffc >>
rect 56 176 90 210
rect 56 86 90 120
rect 142 118 176 152
rect 228 176 262 210
rect 228 86 262 120
rect 314 118 348 152
rect 400 176 434 210
rect 400 86 434 120
rect 486 135 520 169
rect 572 102 606 136
rect 658 165 692 199
rect 744 86 778 120
rect 848 86 882 120
rect 934 173 968 207
rect 1020 86 1054 120
rect 1106 173 1140 207
rect 1192 176 1226 210
rect 1192 86 1226 120
rect 1278 102 1312 136
rect 1364 176 1398 210
rect 1364 86 1398 120
rect 1450 102 1484 136
rect 1536 176 1570 210
rect 1536 86 1570 120
<< pdiffc >>
rect 53 546 87 580
rect 53 463 87 497
rect 53 380 87 414
rect 143 497 177 531
rect 143 390 177 424
rect 233 546 267 580
rect 233 458 267 492
rect 323 497 357 531
rect 323 390 357 424
rect 413 546 447 580
rect 413 458 447 492
rect 503 497 537 531
rect 503 390 537 424
rect 593 546 627 580
rect 593 458 627 492
rect 683 497 717 531
rect 683 406 717 440
rect 773 546 807 580
rect 773 463 807 497
rect 773 380 807 414
rect 863 546 897 580
rect 863 458 897 492
rect 953 546 987 580
rect 953 466 987 500
rect 953 390 987 424
rect 1066 546 1100 580
rect 1066 458 1100 492
rect 1179 546 1213 580
rect 1179 476 1213 510
rect 1179 390 1213 424
rect 1269 546 1303 580
rect 1269 458 1303 492
rect 1359 546 1393 580
rect 1359 476 1393 510
rect 1359 390 1393 424
rect 1449 546 1483 580
rect 1449 458 1483 492
rect 1539 546 1573 580
rect 1539 463 1573 497
rect 1539 380 1573 414
<< poly >>
rect 97 592 133 618
rect 187 592 223 618
rect 277 592 313 618
rect 367 592 403 618
rect 457 592 493 618
rect 547 592 583 618
rect 637 592 673 618
rect 727 592 763 618
rect 817 592 853 618
rect 907 592 943 618
rect 997 592 1033 618
rect 1133 592 1169 618
rect 1223 592 1259 618
rect 1313 592 1349 618
rect 1403 592 1439 618
rect 1493 592 1529 618
rect 97 336 133 368
rect 187 336 223 368
rect 277 336 313 368
rect 367 336 403 368
rect 457 336 493 368
rect 547 336 583 368
rect 637 336 673 368
rect 727 336 763 368
rect 101 320 403 336
rect 101 286 137 320
rect 171 286 205 320
rect 239 286 273 320
rect 307 286 341 320
rect 375 286 403 320
rect 453 320 763 336
rect 453 294 469 320
rect 101 270 403 286
rect 445 286 469 294
rect 503 286 537 320
rect 571 286 605 320
rect 639 286 763 320
rect 817 330 853 368
rect 907 336 943 368
rect 997 336 1033 368
rect 1133 336 1169 368
rect 1223 336 1259 368
rect 1313 336 1349 368
rect 1403 336 1439 368
rect 1493 336 1529 368
rect 907 330 1181 336
rect 817 320 1181 330
rect 817 300 929 320
rect 101 222 131 270
rect 187 222 217 270
rect 273 222 303 270
rect 359 222 389 270
rect 445 264 763 286
rect 893 286 929 300
rect 963 286 997 320
rect 1031 286 1065 320
rect 1099 286 1181 320
rect 893 270 1181 286
rect 1223 320 1529 336
rect 1223 286 1239 320
rect 1273 286 1307 320
rect 1341 286 1375 320
rect 1409 286 1443 320
rect 1477 286 1529 320
rect 1223 270 1529 286
rect 445 222 475 264
rect 531 222 561 264
rect 617 222 647 264
rect 703 222 733 264
rect 893 222 923 270
rect 979 222 1009 270
rect 1065 222 1095 270
rect 1151 222 1181 270
rect 1237 222 1267 270
rect 1323 222 1353 270
rect 1409 222 1439 270
rect 1495 222 1525 270
rect 101 48 131 74
rect 187 48 217 74
rect 273 48 303 74
rect 359 48 389 74
rect 445 48 475 74
rect 531 48 561 74
rect 617 48 647 74
rect 703 48 733 74
rect 893 48 923 74
rect 979 48 1009 74
rect 1065 48 1095 74
rect 1151 48 1181 74
rect 1237 48 1267 74
rect 1323 48 1353 74
rect 1409 48 1439 74
rect 1495 48 1525 74
<< polycont >>
rect 137 286 171 320
rect 205 286 239 320
rect 273 286 307 320
rect 341 286 375 320
rect 469 286 503 320
rect 537 286 571 320
rect 605 286 639 320
rect 929 286 963 320
rect 997 286 1031 320
rect 1065 286 1099 320
rect 1239 286 1273 320
rect 1307 286 1341 320
rect 1375 286 1409 320
rect 1443 286 1477 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 37 581 807 615
rect 37 580 87 581
rect 37 546 53 580
rect 217 580 283 581
rect 37 497 87 546
rect 37 463 53 497
rect 37 414 87 463
rect 37 380 53 414
rect 127 531 177 547
rect 127 497 143 531
rect 127 424 177 497
rect 217 546 233 580
rect 267 546 283 580
rect 397 580 463 581
rect 217 492 283 546
rect 217 458 233 492
rect 267 458 283 492
rect 323 531 357 547
rect 323 424 357 497
rect 397 546 413 580
rect 447 546 463 580
rect 577 580 643 581
rect 397 492 463 546
rect 397 458 413 492
rect 447 458 463 492
rect 503 531 537 547
rect 503 424 537 497
rect 577 546 593 580
rect 627 546 643 580
rect 757 580 807 581
rect 577 492 643 546
rect 577 458 593 492
rect 627 458 643 492
rect 683 531 723 547
rect 717 497 723 531
rect 683 440 723 497
rect 127 390 143 424
rect 177 390 323 424
rect 357 390 503 424
rect 537 406 683 424
rect 717 406 723 440
rect 537 390 723 406
rect 37 364 87 380
rect 121 320 391 356
rect 121 286 137 320
rect 171 286 205 320
rect 239 286 273 320
rect 307 286 341 320
rect 375 286 391 320
rect 121 270 391 286
rect 453 320 655 356
rect 453 286 469 320
rect 503 286 537 320
rect 571 286 605 320
rect 639 286 655 320
rect 453 270 655 286
rect 689 304 723 390
rect 757 546 773 580
rect 757 497 807 546
rect 757 463 773 497
rect 757 424 807 463
rect 847 580 913 649
rect 847 546 863 580
rect 897 546 913 580
rect 847 492 913 546
rect 847 458 863 492
rect 897 458 913 492
rect 953 580 1003 596
rect 987 546 1003 580
rect 953 500 1003 546
rect 987 466 1003 500
rect 953 424 1003 466
rect 1037 580 1129 649
rect 1037 546 1066 580
rect 1100 546 1129 580
rect 1037 492 1129 546
rect 1037 458 1066 492
rect 1100 458 1129 492
rect 1163 580 1213 596
rect 1163 546 1179 580
rect 1163 510 1213 546
rect 1163 476 1179 510
rect 1163 424 1213 476
rect 1253 580 1319 649
rect 1253 546 1269 580
rect 1303 546 1319 580
rect 1253 492 1319 546
rect 1253 458 1269 492
rect 1303 458 1319 492
rect 1359 580 1393 596
rect 1359 510 1393 546
rect 1359 424 1393 476
rect 1433 580 1499 649
rect 1433 546 1449 580
rect 1483 546 1499 580
rect 1433 492 1499 546
rect 1433 458 1449 492
rect 1483 458 1499 492
rect 1539 580 1589 596
rect 1573 546 1589 580
rect 1539 497 1589 546
rect 1573 463 1589 497
rect 1539 424 1589 463
rect 757 414 953 424
rect 757 380 773 414
rect 807 390 953 414
rect 987 390 1179 424
rect 1213 390 1359 424
rect 1393 414 1589 424
rect 1393 390 1539 414
rect 757 364 807 380
rect 1573 380 1589 414
rect 1539 364 1589 380
rect 889 320 1127 356
rect 689 236 839 304
rect 889 286 929 320
rect 963 286 997 320
rect 1031 286 1065 320
rect 1099 286 1127 320
rect 889 270 1127 286
rect 1177 320 1493 356
rect 1177 286 1239 320
rect 1273 286 1307 320
rect 1341 286 1375 320
rect 1409 286 1443 320
rect 1477 286 1493 320
rect 1177 270 1493 286
rect 40 210 434 236
rect 40 176 56 210
rect 90 202 228 210
rect 40 120 90 176
rect 212 176 228 202
rect 262 202 400 210
rect 40 86 56 120
rect 40 70 90 86
rect 126 152 176 168
rect 126 118 142 152
rect 126 17 176 118
rect 212 120 262 176
rect 212 86 228 120
rect 212 70 262 86
rect 298 152 364 168
rect 298 118 314 152
rect 348 118 364 152
rect 298 17 364 118
rect 400 120 434 176
rect 470 226 839 236
rect 470 207 1156 226
rect 470 202 934 207
rect 470 169 536 202
rect 470 135 486 169
rect 520 135 536 169
rect 642 199 934 202
rect 470 119 536 135
rect 572 136 606 168
rect 642 165 658 199
rect 692 173 934 199
rect 968 173 1106 207
rect 1140 173 1156 207
rect 692 170 1156 173
rect 692 165 798 170
rect 642 154 798 165
rect 1090 154 1156 170
rect 1192 210 1586 236
rect 1226 202 1364 210
rect 400 85 434 86
rect 832 120 898 136
rect 1192 120 1226 176
rect 1348 176 1364 202
rect 1398 202 1536 210
rect 606 102 744 120
rect 572 86 744 102
rect 778 86 794 120
rect 572 85 794 86
rect 400 51 794 85
rect 832 86 848 120
rect 882 86 1020 120
rect 1054 86 1192 120
rect 832 70 1226 86
rect 1262 136 1312 168
rect 1262 102 1278 136
rect 1262 17 1312 102
rect 1348 120 1398 176
rect 1520 176 1536 202
rect 1570 176 1586 210
rect 1348 86 1364 120
rect 1348 70 1398 86
rect 1434 136 1484 168
rect 1434 102 1450 136
rect 1434 17 1484 102
rect 1520 120 1586 176
rect 1520 86 1536 120
rect 1570 86 1586 120
rect 1520 70 1586 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a22oi_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 352106
string GDS_START 339062
<< end >>
