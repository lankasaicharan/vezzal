magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 3 241 481 259
rect 3 49 1998 241
rect 0 0 2016 49
<< scnmos >>
rect 82 65 112 233
rect 168 65 198 233
rect 270 65 300 233
rect 372 65 402 233
rect 562 47 592 215
rect 648 47 678 215
rect 734 47 764 215
rect 820 47 850 215
rect 906 47 936 215
rect 992 47 1022 215
rect 1078 47 1108 215
rect 1164 47 1194 215
rect 1287 47 1317 215
rect 1373 47 1403 215
rect 1459 47 1489 215
rect 1545 47 1575 215
rect 1631 47 1661 215
rect 1717 47 1747 215
rect 1803 47 1833 215
rect 1889 47 1919 215
<< scpmoshvt >>
rect 218 367 248 619
rect 304 367 334 619
rect 390 367 420 619
rect 476 367 506 619
rect 562 367 592 619
rect 648 367 678 619
rect 734 367 764 619
rect 820 367 850 619
rect 906 367 936 619
rect 992 367 1022 619
rect 1078 367 1108 619
rect 1164 367 1194 619
rect 1287 367 1317 619
rect 1373 367 1403 619
rect 1459 367 1489 619
rect 1545 367 1575 619
rect 1631 367 1661 619
rect 1724 367 1754 619
rect 1810 367 1840 619
rect 1896 367 1926 619
<< ndiff >>
rect 29 221 82 233
rect 29 187 37 221
rect 71 187 82 221
rect 29 111 82 187
rect 29 77 37 111
rect 71 77 82 111
rect 29 65 82 77
rect 112 225 168 233
rect 112 191 123 225
rect 157 191 168 225
rect 112 157 168 191
rect 112 123 123 157
rect 157 123 168 157
rect 112 65 168 123
rect 198 175 270 233
rect 198 141 223 175
rect 257 141 270 175
rect 198 107 270 141
rect 198 73 223 107
rect 257 73 270 107
rect 198 65 270 73
rect 300 225 372 233
rect 300 191 323 225
rect 357 191 372 225
rect 300 157 372 191
rect 300 123 323 157
rect 357 123 372 157
rect 300 65 372 123
rect 402 167 455 233
rect 402 133 413 167
rect 447 133 455 167
rect 402 65 455 133
rect 509 93 562 215
rect 509 59 517 93
rect 551 59 562 93
rect 509 47 562 59
rect 592 181 648 215
rect 592 147 603 181
rect 637 147 648 181
rect 592 47 648 147
rect 678 163 734 215
rect 678 129 689 163
rect 723 129 734 163
rect 678 93 734 129
rect 678 59 689 93
rect 723 59 734 93
rect 678 47 734 59
rect 764 173 820 215
rect 764 139 775 173
rect 809 139 820 173
rect 764 47 820 139
rect 850 105 906 215
rect 850 71 861 105
rect 895 71 906 105
rect 850 47 906 71
rect 936 195 992 215
rect 936 161 947 195
rect 981 161 992 195
rect 936 47 992 161
rect 1022 105 1078 215
rect 1022 71 1033 105
rect 1067 71 1078 105
rect 1022 47 1078 71
rect 1108 183 1164 215
rect 1108 149 1119 183
rect 1153 149 1164 183
rect 1108 47 1164 149
rect 1194 181 1287 215
rect 1194 147 1228 181
rect 1262 147 1287 181
rect 1194 93 1287 147
rect 1194 59 1228 93
rect 1262 59 1287 93
rect 1194 47 1287 59
rect 1317 105 1373 215
rect 1317 71 1328 105
rect 1362 71 1373 105
rect 1317 47 1373 71
rect 1403 181 1459 215
rect 1403 147 1414 181
rect 1448 147 1459 181
rect 1403 101 1459 147
rect 1403 67 1414 101
rect 1448 67 1459 101
rect 1403 47 1459 67
rect 1489 105 1545 215
rect 1489 71 1500 105
rect 1534 71 1545 105
rect 1489 47 1545 71
rect 1575 181 1631 215
rect 1575 147 1586 181
rect 1620 147 1631 181
rect 1575 101 1631 147
rect 1575 67 1586 101
rect 1620 67 1631 101
rect 1575 47 1631 67
rect 1661 105 1717 215
rect 1661 71 1672 105
rect 1706 71 1717 105
rect 1661 47 1717 71
rect 1747 192 1803 215
rect 1747 158 1758 192
rect 1792 158 1803 192
rect 1747 101 1803 158
rect 1747 67 1758 101
rect 1792 67 1803 101
rect 1747 47 1803 67
rect 1833 128 1889 215
rect 1833 94 1844 128
rect 1878 94 1889 128
rect 1833 47 1889 94
rect 1919 192 1972 215
rect 1919 158 1930 192
rect 1964 158 1972 192
rect 1919 101 1972 158
rect 1919 67 1930 101
rect 1964 67 1972 101
rect 1919 47 1972 67
<< pdiff >>
rect 165 607 218 619
rect 165 573 173 607
rect 207 573 218 607
rect 165 511 218 573
rect 165 477 173 511
rect 207 477 218 511
rect 165 418 218 477
rect 165 384 173 418
rect 207 384 218 418
rect 165 367 218 384
rect 248 599 304 619
rect 248 565 259 599
rect 293 565 304 599
rect 248 524 304 565
rect 248 490 259 524
rect 293 490 304 524
rect 248 434 304 490
rect 248 400 259 434
rect 293 400 304 434
rect 248 367 304 400
rect 334 607 390 619
rect 334 573 345 607
rect 379 573 390 607
rect 334 493 390 573
rect 334 459 345 493
rect 379 459 390 493
rect 334 367 390 459
rect 420 599 476 619
rect 420 565 431 599
rect 465 565 476 599
rect 420 513 476 565
rect 420 479 431 513
rect 465 479 476 513
rect 420 418 476 479
rect 420 384 431 418
rect 465 384 476 418
rect 420 367 476 384
rect 506 607 562 619
rect 506 573 517 607
rect 551 573 562 607
rect 506 501 562 573
rect 506 467 517 501
rect 551 467 562 501
rect 506 367 562 467
rect 592 599 648 619
rect 592 565 603 599
rect 637 565 648 599
rect 592 509 648 565
rect 592 475 603 509
rect 637 475 648 509
rect 592 367 648 475
rect 678 567 734 619
rect 678 533 689 567
rect 723 533 734 567
rect 678 367 734 533
rect 764 599 820 619
rect 764 565 775 599
rect 809 565 820 599
rect 764 509 820 565
rect 764 475 775 509
rect 809 475 820 509
rect 764 367 820 475
rect 850 539 906 619
rect 850 505 861 539
rect 895 505 906 539
rect 850 425 906 505
rect 850 391 861 425
rect 895 391 906 425
rect 850 367 906 391
rect 936 599 992 619
rect 936 565 947 599
rect 981 565 992 599
rect 936 513 992 565
rect 936 479 947 513
rect 981 479 992 513
rect 936 367 992 479
rect 1022 539 1078 619
rect 1022 505 1033 539
rect 1067 505 1078 539
rect 1022 425 1078 505
rect 1022 391 1033 425
rect 1067 391 1078 425
rect 1022 367 1078 391
rect 1108 599 1164 619
rect 1108 565 1119 599
rect 1153 565 1164 599
rect 1108 511 1164 565
rect 1108 477 1119 511
rect 1153 477 1164 511
rect 1108 367 1164 477
rect 1194 607 1287 619
rect 1194 573 1226 607
rect 1260 573 1287 607
rect 1194 504 1287 573
rect 1194 470 1226 504
rect 1260 470 1287 504
rect 1194 367 1287 470
rect 1317 599 1373 619
rect 1317 565 1328 599
rect 1362 565 1373 599
rect 1317 511 1373 565
rect 1317 477 1328 511
rect 1362 477 1373 511
rect 1317 367 1373 477
rect 1403 540 1459 619
rect 1403 506 1414 540
rect 1448 506 1459 540
rect 1403 424 1459 506
rect 1403 390 1414 424
rect 1448 390 1459 424
rect 1403 367 1459 390
rect 1489 599 1545 619
rect 1489 565 1500 599
rect 1534 565 1545 599
rect 1489 508 1545 565
rect 1489 474 1500 508
rect 1534 474 1545 508
rect 1489 367 1545 474
rect 1575 540 1631 619
rect 1575 506 1586 540
rect 1620 506 1631 540
rect 1575 424 1631 506
rect 1575 390 1586 424
rect 1620 390 1631 424
rect 1575 367 1631 390
rect 1661 599 1724 619
rect 1661 565 1679 599
rect 1713 565 1724 599
rect 1661 504 1724 565
rect 1661 470 1679 504
rect 1713 470 1724 504
rect 1661 413 1724 470
rect 1661 379 1679 413
rect 1713 379 1724 413
rect 1661 367 1724 379
rect 1754 607 1810 619
rect 1754 573 1765 607
rect 1799 573 1810 607
rect 1754 530 1810 573
rect 1754 496 1765 530
rect 1799 496 1810 530
rect 1754 440 1810 496
rect 1754 406 1765 440
rect 1799 406 1810 440
rect 1754 367 1810 406
rect 1840 599 1896 619
rect 1840 565 1851 599
rect 1885 565 1896 599
rect 1840 504 1896 565
rect 1840 470 1851 504
rect 1885 470 1896 504
rect 1840 413 1896 470
rect 1840 379 1851 413
rect 1885 379 1896 413
rect 1840 367 1896 379
rect 1926 607 1979 619
rect 1926 573 1937 607
rect 1971 573 1979 607
rect 1926 509 1979 573
rect 1926 475 1937 509
rect 1971 475 1979 509
rect 1926 413 1979 475
rect 1926 379 1937 413
rect 1971 379 1979 413
rect 1926 367 1979 379
<< ndiffc >>
rect 37 187 71 221
rect 37 77 71 111
rect 123 191 157 225
rect 123 123 157 157
rect 223 141 257 175
rect 223 73 257 107
rect 323 191 357 225
rect 323 123 357 157
rect 413 133 447 167
rect 517 59 551 93
rect 603 147 637 181
rect 689 129 723 163
rect 689 59 723 93
rect 775 139 809 173
rect 861 71 895 105
rect 947 161 981 195
rect 1033 71 1067 105
rect 1119 149 1153 183
rect 1228 147 1262 181
rect 1228 59 1262 93
rect 1328 71 1362 105
rect 1414 147 1448 181
rect 1414 67 1448 101
rect 1500 71 1534 105
rect 1586 147 1620 181
rect 1586 67 1620 101
rect 1672 71 1706 105
rect 1758 158 1792 192
rect 1758 67 1792 101
rect 1844 94 1878 128
rect 1930 158 1964 192
rect 1930 67 1964 101
<< pdiffc >>
rect 173 573 207 607
rect 173 477 207 511
rect 173 384 207 418
rect 259 565 293 599
rect 259 490 293 524
rect 259 400 293 434
rect 345 573 379 607
rect 345 459 379 493
rect 431 565 465 599
rect 431 479 465 513
rect 431 384 465 418
rect 517 573 551 607
rect 517 467 551 501
rect 603 565 637 599
rect 603 475 637 509
rect 689 533 723 567
rect 775 565 809 599
rect 775 475 809 509
rect 861 505 895 539
rect 861 391 895 425
rect 947 565 981 599
rect 947 479 981 513
rect 1033 505 1067 539
rect 1033 391 1067 425
rect 1119 565 1153 599
rect 1119 477 1153 511
rect 1226 573 1260 607
rect 1226 470 1260 504
rect 1328 565 1362 599
rect 1328 477 1362 511
rect 1414 506 1448 540
rect 1414 390 1448 424
rect 1500 565 1534 599
rect 1500 474 1534 508
rect 1586 506 1620 540
rect 1586 390 1620 424
rect 1679 565 1713 599
rect 1679 470 1713 504
rect 1679 379 1713 413
rect 1765 573 1799 607
rect 1765 496 1799 530
rect 1765 406 1799 440
rect 1851 565 1885 599
rect 1851 470 1885 504
rect 1851 379 1885 413
rect 1937 573 1971 607
rect 1937 475 1971 509
rect 1937 379 1971 413
<< poly >>
rect 218 619 248 645
rect 304 619 334 645
rect 390 619 420 645
rect 476 619 506 645
rect 562 619 592 645
rect 648 619 678 645
rect 734 619 764 645
rect 820 619 850 645
rect 906 619 936 645
rect 992 619 1022 645
rect 1078 619 1108 645
rect 1164 619 1194 645
rect 1287 619 1317 645
rect 1373 619 1403 645
rect 1459 619 1489 645
rect 1545 619 1575 645
rect 1631 619 1661 645
rect 1724 619 1754 645
rect 1810 619 1840 645
rect 1896 619 1926 645
rect 218 335 248 367
rect 304 335 334 367
rect 390 335 420 367
rect 476 335 506 367
rect 50 319 506 335
rect 50 285 66 319
rect 100 285 134 319
rect 168 285 202 319
rect 236 285 270 319
rect 304 285 338 319
rect 372 285 406 319
rect 440 285 506 319
rect 50 269 506 285
rect 562 335 592 367
rect 648 335 678 367
rect 734 335 764 367
rect 562 319 764 335
rect 562 285 578 319
rect 612 285 646 319
rect 680 285 714 319
rect 748 285 764 319
rect 562 269 764 285
rect 82 233 112 269
rect 168 233 198 269
rect 270 233 300 269
rect 372 233 402 269
rect 562 215 592 269
rect 648 215 678 269
rect 734 215 764 269
rect 820 303 850 367
rect 906 303 936 367
rect 992 303 1022 367
rect 1078 303 1108 367
rect 1164 325 1194 367
rect 1157 309 1223 325
rect 820 287 1115 303
rect 820 253 861 287
rect 895 253 929 287
rect 963 253 997 287
rect 1031 253 1065 287
rect 1099 253 1115 287
rect 1157 275 1173 309
rect 1207 275 1223 309
rect 1287 303 1317 367
rect 1373 335 1403 367
rect 1459 335 1489 367
rect 1545 335 1575 367
rect 1631 335 1661 367
rect 1373 319 1661 335
rect 1157 259 1223 275
rect 1265 287 1331 303
rect 820 237 1115 253
rect 820 215 850 237
rect 906 215 936 237
rect 992 215 1022 237
rect 1078 215 1108 237
rect 1164 215 1194 259
rect 1265 253 1281 287
rect 1315 253 1331 287
rect 1265 237 1331 253
rect 1373 285 1389 319
rect 1423 285 1457 319
rect 1491 285 1525 319
rect 1559 285 1593 319
rect 1627 285 1661 319
rect 1724 303 1754 367
rect 1810 303 1840 367
rect 1896 303 1926 367
rect 1373 269 1661 285
rect 1287 215 1317 237
rect 1373 215 1403 269
rect 1459 215 1489 269
rect 1545 215 1575 269
rect 1631 215 1661 269
rect 1717 287 1987 303
rect 1717 253 1733 287
rect 1767 253 1801 287
rect 1835 253 1869 287
rect 1903 253 1937 287
rect 1971 253 1987 287
rect 1717 237 1987 253
rect 1717 215 1747 237
rect 1803 215 1833 237
rect 1889 215 1919 237
rect 82 39 112 65
rect 168 39 198 65
rect 270 39 300 65
rect 372 39 402 65
rect 562 21 592 47
rect 648 21 678 47
rect 734 21 764 47
rect 820 21 850 47
rect 906 21 936 47
rect 992 21 1022 47
rect 1078 21 1108 47
rect 1164 21 1194 47
rect 1287 21 1317 47
rect 1373 21 1403 47
rect 1459 21 1489 47
rect 1545 21 1575 47
rect 1631 21 1661 47
rect 1717 21 1747 47
rect 1803 21 1833 47
rect 1889 21 1919 47
<< polycont >>
rect 66 285 100 319
rect 134 285 168 319
rect 202 285 236 319
rect 270 285 304 319
rect 338 285 372 319
rect 406 285 440 319
rect 578 285 612 319
rect 646 285 680 319
rect 714 285 748 319
rect 861 253 895 287
rect 929 253 963 287
rect 997 253 1031 287
rect 1065 253 1099 287
rect 1173 275 1207 309
rect 1281 253 1315 287
rect 1389 285 1423 319
rect 1457 285 1491 319
rect 1525 285 1559 319
rect 1593 285 1627 319
rect 1733 253 1767 287
rect 1801 253 1835 287
rect 1869 253 1903 287
rect 1937 253 1971 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 157 607 223 649
rect 157 573 173 607
rect 207 573 223 607
rect 157 511 223 573
rect 157 477 173 511
rect 207 477 223 511
rect 157 418 223 477
rect 157 384 173 418
rect 207 384 223 418
rect 257 599 293 615
rect 257 565 259 599
rect 257 524 293 565
rect 257 490 259 524
rect 257 434 293 490
rect 329 607 395 649
rect 329 573 345 607
rect 379 573 395 607
rect 329 493 395 573
rect 329 459 345 493
rect 379 459 395 493
rect 329 452 395 459
rect 429 599 467 615
rect 429 565 431 599
rect 465 565 467 599
rect 429 513 467 565
rect 429 479 431 513
rect 465 479 467 513
rect 257 400 259 434
rect 429 425 467 479
rect 501 607 567 649
rect 501 573 517 607
rect 551 573 567 607
rect 501 501 567 573
rect 501 467 517 501
rect 551 467 567 501
rect 501 459 567 467
rect 601 599 639 615
rect 601 565 603 599
rect 637 565 639 599
rect 601 509 639 565
rect 673 567 739 649
rect 673 533 689 567
rect 723 533 739 567
rect 673 527 739 533
rect 773 599 1169 615
rect 773 565 775 599
rect 809 581 947 599
rect 809 565 811 581
rect 601 475 603 509
rect 637 493 639 509
rect 773 509 811 565
rect 945 565 947 581
rect 981 581 1119 599
rect 981 565 983 581
rect 773 493 775 509
rect 637 475 775 493
rect 809 475 811 509
rect 601 459 811 475
rect 845 539 911 547
rect 845 505 861 539
rect 895 505 911 539
rect 845 427 911 505
rect 945 513 983 565
rect 1117 565 1119 581
rect 1153 565 1169 599
rect 945 479 947 513
rect 981 479 983 513
rect 945 463 983 479
rect 1017 539 1083 547
rect 1017 505 1033 539
rect 1067 505 1083 539
rect 1017 427 1083 505
rect 1117 511 1169 565
rect 1117 477 1119 511
rect 1153 477 1169 511
rect 1117 461 1169 477
rect 1210 607 1276 649
rect 1210 573 1226 607
rect 1260 573 1276 607
rect 1210 504 1276 573
rect 1210 470 1226 504
rect 1260 470 1276 504
rect 1210 461 1276 470
rect 1312 599 1715 615
rect 1312 565 1328 599
rect 1362 581 1500 599
rect 1362 565 1364 581
rect 1312 511 1364 565
rect 1498 565 1500 581
rect 1534 581 1679 599
rect 1534 565 1536 581
rect 1312 477 1328 511
rect 1362 477 1364 511
rect 1312 461 1364 477
rect 1398 540 1464 547
rect 1398 506 1414 540
rect 1448 506 1464 540
rect 1398 427 1464 506
rect 1498 508 1536 565
rect 1677 565 1679 581
rect 1713 565 1715 599
rect 1498 474 1500 508
rect 1534 474 1536 508
rect 1498 458 1536 474
rect 1570 540 1636 547
rect 1570 506 1586 540
rect 1620 506 1636 540
rect 845 425 1464 427
rect 429 418 861 425
rect 293 400 431 418
rect 257 384 431 400
rect 465 391 861 418
rect 895 391 1033 425
rect 1067 424 1464 425
rect 1570 424 1636 506
rect 1067 391 1414 424
rect 465 384 528 391
rect 1279 390 1414 391
rect 1448 390 1586 424
rect 1620 390 1636 424
rect 1677 504 1715 565
rect 1677 470 1679 504
rect 1713 470 1715 504
rect 1677 413 1715 470
rect 17 319 458 350
rect 17 285 66 319
rect 100 285 134 319
rect 168 285 202 319
rect 236 285 270 319
rect 304 285 338 319
rect 372 285 406 319
rect 440 285 458 319
rect 492 251 528 384
rect 1677 379 1679 413
rect 1713 379 1715 413
rect 1749 607 1815 649
rect 1749 573 1765 607
rect 1799 573 1815 607
rect 1749 530 1815 573
rect 1749 496 1765 530
rect 1799 496 1815 530
rect 1749 440 1815 496
rect 1749 406 1765 440
rect 1799 406 1815 440
rect 1849 599 1894 615
rect 1849 565 1851 599
rect 1885 565 1894 599
rect 1849 504 1894 565
rect 1849 470 1851 504
rect 1885 470 1894 504
rect 1849 413 1894 470
rect 1677 372 1715 379
rect 1849 379 1851 413
rect 1885 379 1894 413
rect 1849 372 1894 379
rect 562 323 1229 357
rect 562 319 764 323
rect 562 285 578 319
rect 612 285 646 319
rect 680 285 714 319
rect 748 285 764 319
rect 1163 309 1229 323
rect 562 280 764 285
rect 845 287 1129 289
rect 21 221 73 237
rect 21 187 37 221
rect 71 187 73 221
rect 21 111 73 187
rect 107 225 528 251
rect 845 253 861 287
rect 895 253 929 287
rect 963 253 997 287
rect 1031 253 1065 287
rect 1099 253 1129 287
rect 1163 275 1173 309
rect 1207 275 1229 309
rect 1365 319 1643 350
rect 1677 338 1894 372
rect 1928 607 1987 649
rect 1928 573 1937 607
rect 1971 573 1987 607
rect 1928 509 1987 573
rect 1928 475 1937 509
rect 1971 475 1987 509
rect 1928 413 1987 475
rect 1928 379 1937 413
rect 1971 379 1987 413
rect 1928 363 1987 379
rect 1163 259 1229 275
rect 1281 287 1331 303
rect 107 191 123 225
rect 157 217 323 225
rect 157 191 173 217
rect 107 157 173 191
rect 307 191 323 217
rect 357 217 528 225
rect 357 191 373 217
rect 107 123 123 157
rect 157 123 173 157
rect 107 119 173 123
rect 207 175 273 179
rect 207 141 223 175
rect 257 141 273 175
rect 21 77 37 111
rect 71 85 73 111
rect 207 107 273 141
rect 307 157 373 191
rect 562 205 809 246
rect 845 239 1129 253
rect 1315 253 1331 287
rect 1365 285 1389 319
rect 1423 285 1457 319
rect 1491 285 1525 319
rect 1559 285 1593 319
rect 1627 285 1643 319
rect 1677 287 1998 304
rect 1281 249 1331 253
rect 1677 253 1733 287
rect 1767 253 1801 287
rect 1835 253 1869 287
rect 1903 253 1937 287
rect 1971 253 1998 287
rect 1677 249 1998 253
rect 1281 242 1998 249
rect 1281 215 1718 242
rect 562 201 1169 205
rect 562 183 639 201
rect 307 123 323 157
rect 357 123 373 157
rect 307 119 373 123
rect 407 181 639 183
rect 407 167 603 181
rect 407 133 413 167
rect 447 147 603 167
rect 637 147 639 181
rect 773 195 1169 201
rect 773 173 947 195
rect 447 133 639 147
rect 407 131 639 133
rect 673 163 739 167
rect 207 85 223 107
rect 71 77 223 85
rect 21 73 223 77
rect 257 85 273 107
rect 407 85 463 131
rect 673 129 689 163
rect 723 129 739 163
rect 673 97 739 129
rect 773 139 775 173
rect 809 161 947 173
rect 981 183 1169 195
rect 1752 192 1980 208
rect 981 161 1119 183
rect 809 155 1119 161
rect 809 139 823 155
rect 773 123 823 139
rect 1103 149 1119 155
rect 1153 149 1169 183
rect 1103 133 1169 149
rect 1212 181 1258 189
rect 1752 181 1758 192
rect 1212 147 1228 181
rect 1262 147 1414 181
rect 1448 147 1586 181
rect 1620 158 1758 181
rect 1792 174 1930 192
rect 1792 158 1794 174
rect 1620 147 1794 158
rect 257 73 463 85
rect 21 51 463 73
rect 501 93 739 97
rect 501 59 517 93
rect 551 59 689 93
rect 723 89 739 93
rect 857 105 1071 121
rect 857 89 861 105
rect 723 71 861 89
rect 895 71 1033 105
rect 1067 89 1071 105
rect 1212 93 1278 147
rect 1212 89 1228 93
rect 1067 71 1228 89
rect 723 59 1228 71
rect 1262 59 1278 93
rect 501 51 1278 59
rect 1312 105 1378 113
rect 1312 71 1328 105
rect 1362 71 1378 105
rect 1312 17 1378 71
rect 1412 101 1450 147
rect 1412 67 1414 101
rect 1448 67 1450 101
rect 1412 51 1450 67
rect 1484 105 1550 113
rect 1484 71 1500 105
rect 1534 71 1550 105
rect 1484 17 1550 71
rect 1584 101 1622 147
rect 1584 67 1586 101
rect 1620 67 1622 101
rect 1584 51 1622 67
rect 1656 105 1722 113
rect 1656 71 1672 105
rect 1706 71 1722 105
rect 1656 17 1722 71
rect 1756 101 1794 147
rect 1928 158 1930 174
rect 1964 158 1980 192
rect 1756 67 1758 101
rect 1792 67 1794 101
rect 1756 51 1794 67
rect 1828 128 1894 140
rect 1828 94 1844 128
rect 1878 94 1894 128
rect 1828 17 1894 94
rect 1928 101 1980 158
rect 1928 67 1930 101
rect 1964 67 1980 101
rect 1928 51 1980 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221ai_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1375 390 1409 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5886336
string GDS_START 5869748
<< end >>
