magic
tech sky130A
magscale 1 2
timestamp 1627201166
<< checkpaint >>
rect -1250 -1349 2066 1561
<< pwell >>
rect 10 10 806 230
<< nmoslvt >>
rect 92 36 122 204
rect 178 36 208 204
rect 264 36 294 204
rect 350 36 380 204
rect 436 36 466 204
rect 522 36 552 204
rect 608 36 638 204
rect 694 36 724 204
<< ndiff >>
rect 36 173 92 204
rect 36 139 47 173
rect 81 139 92 173
rect 36 101 92 139
rect 36 67 47 101
rect 81 67 92 101
rect 36 36 92 67
rect 122 173 178 204
rect 122 139 133 173
rect 167 139 178 173
rect 122 101 178 139
rect 122 67 133 101
rect 167 67 178 101
rect 122 36 178 67
rect 208 173 264 204
rect 208 139 219 173
rect 253 139 264 173
rect 208 101 264 139
rect 208 67 219 101
rect 253 67 264 101
rect 208 36 264 67
rect 294 173 350 204
rect 294 139 305 173
rect 339 139 350 173
rect 294 101 350 139
rect 294 67 305 101
rect 339 67 350 101
rect 294 36 350 67
rect 380 173 436 204
rect 380 139 391 173
rect 425 139 436 173
rect 380 101 436 139
rect 380 67 391 101
rect 425 67 436 101
rect 380 36 436 67
rect 466 173 522 204
rect 466 139 477 173
rect 511 139 522 173
rect 466 101 522 139
rect 466 67 477 101
rect 511 67 522 101
rect 466 36 522 67
rect 552 173 608 204
rect 552 139 563 173
rect 597 139 608 173
rect 552 101 608 139
rect 552 67 563 101
rect 597 67 608 101
rect 552 36 608 67
rect 638 173 694 204
rect 638 139 649 173
rect 683 139 694 173
rect 638 101 694 139
rect 638 67 649 101
rect 683 67 694 101
rect 638 36 694 67
rect 724 173 780 204
rect 724 139 735 173
rect 769 139 780 173
rect 724 101 780 139
rect 724 67 735 101
rect 769 67 780 101
rect 724 36 780 67
<< ndiffc >>
rect 47 139 81 173
rect 47 67 81 101
rect 133 139 167 173
rect 133 67 167 101
rect 219 139 253 173
rect 219 67 253 101
rect 305 139 339 173
rect 305 67 339 101
rect 391 139 425 173
rect 391 67 425 101
rect 477 139 511 173
rect 477 67 511 101
rect 563 139 597 173
rect 563 67 597 101
rect 649 139 683 173
rect 649 67 683 101
rect 735 139 769 173
rect 735 67 769 101
<< poly >>
rect 92 285 724 301
rect 92 251 153 285
rect 187 251 221 285
rect 255 251 289 285
rect 323 251 357 285
rect 391 251 425 285
rect 459 251 493 285
rect 527 251 561 285
rect 595 251 629 285
rect 663 251 724 285
rect 92 230 724 251
rect 92 204 122 230
rect 178 204 208 230
rect 264 204 294 230
rect 350 204 380 230
rect 436 204 466 230
rect 522 204 552 230
rect 608 204 638 230
rect 694 204 724 230
rect 92 10 122 36
rect 178 10 208 36
rect 264 10 294 36
rect 350 10 380 36
rect 436 10 466 36
rect 522 10 552 36
rect 608 10 638 36
rect 694 10 724 36
<< polycont >>
rect 153 251 187 285
rect 221 251 255 285
rect 289 251 323 285
rect 357 251 391 285
rect 425 251 459 285
rect 493 251 527 285
rect 561 251 595 285
rect 629 251 663 285
<< locali >>
rect 137 285 679 301
rect 137 251 139 285
rect 187 251 211 285
rect 255 251 283 285
rect 323 251 355 285
rect 391 251 425 285
rect 461 251 493 285
rect 533 251 561 285
rect 605 251 629 285
rect 677 251 679 285
rect 137 235 679 251
rect 47 173 81 189
rect 47 101 81 139
rect 47 51 81 67
rect 133 173 167 189
rect 133 101 167 139
rect 133 51 167 67
rect 219 173 253 189
rect 219 101 253 139
rect 219 51 253 67
rect 305 173 339 189
rect 305 101 339 139
rect 305 51 339 67
rect 391 173 425 189
rect 391 101 425 139
rect 391 51 425 67
rect 477 173 511 189
rect 477 101 511 139
rect 477 51 511 67
rect 563 173 597 189
rect 563 101 597 139
rect 563 51 597 67
rect 649 173 683 189
rect 649 101 683 139
rect 649 51 683 67
rect 735 173 769 189
rect 735 101 769 139
rect 735 51 769 67
<< viali >>
rect 139 251 153 285
rect 153 251 173 285
rect 211 251 221 285
rect 221 251 245 285
rect 283 251 289 285
rect 289 251 317 285
rect 355 251 357 285
rect 357 251 389 285
rect 427 251 459 285
rect 459 251 461 285
rect 499 251 527 285
rect 527 251 533 285
rect 571 251 595 285
rect 595 251 605 285
rect 643 251 663 285
rect 663 251 677 285
rect 47 139 81 173
rect 47 67 81 101
rect 133 139 167 173
rect 133 67 167 101
rect 219 139 253 173
rect 219 67 253 101
rect 305 139 339 173
rect 305 67 339 101
rect 391 139 425 173
rect 391 67 425 101
rect 477 139 511 173
rect 477 67 511 101
rect 563 139 597 173
rect 563 67 597 101
rect 649 139 683 173
rect 649 67 683 101
rect 735 139 769 173
rect 735 67 769 101
<< metal1 >>
rect 127 285 689 297
rect 127 251 139 285
rect 173 251 211 285
rect 245 251 283 285
rect 317 251 355 285
rect 389 251 427 285
rect 461 251 499 285
rect 533 251 571 285
rect 605 251 643 285
rect 677 251 689 285
rect 127 239 689 251
rect 41 173 87 189
rect 41 139 47 173
rect 81 139 87 173
rect 41 101 87 139
rect 41 67 47 101
rect 81 67 87 101
rect 41 -29 87 67
rect 124 178 176 189
rect 124 114 176 126
rect 124 51 176 62
rect 213 173 259 189
rect 213 139 219 173
rect 253 139 259 173
rect 213 101 259 139
rect 213 67 219 101
rect 253 67 259 101
rect 213 -29 259 67
rect 296 176 348 189
rect 296 112 348 124
rect 296 51 348 60
rect 385 173 431 189
rect 385 139 391 173
rect 425 139 431 173
rect 385 101 431 139
rect 385 67 391 101
rect 425 67 431 101
rect 385 -29 431 67
rect 468 176 520 189
rect 468 112 520 124
rect 468 51 520 60
rect 557 173 603 189
rect 557 139 563 173
rect 597 139 603 173
rect 557 101 603 139
rect 557 67 563 101
rect 597 67 603 101
rect 557 -29 603 67
rect 640 176 692 189
rect 640 112 692 124
rect 640 51 692 60
rect 729 173 775 189
rect 729 139 735 173
rect 769 139 775 173
rect 729 101 775 139
rect 729 67 735 101
rect 769 67 775 101
rect 729 -29 775 67
rect 41 -89 775 -29
<< via1 >>
rect 124 173 176 178
rect 124 139 133 173
rect 133 139 167 173
rect 167 139 176 173
rect 124 126 176 139
rect 124 101 176 114
rect 124 67 133 101
rect 133 67 167 101
rect 167 67 176 101
rect 124 62 176 67
rect 296 173 348 176
rect 296 139 305 173
rect 305 139 339 173
rect 339 139 348 173
rect 296 124 348 139
rect 296 101 348 112
rect 296 67 305 101
rect 305 67 339 101
rect 339 67 348 101
rect 296 60 348 67
rect 468 173 520 176
rect 468 139 477 173
rect 477 139 511 173
rect 511 139 520 173
rect 468 124 520 139
rect 468 101 520 112
rect 468 67 477 101
rect 477 67 511 101
rect 511 67 520 101
rect 468 60 520 67
rect 640 173 692 176
rect 640 139 649 173
rect 649 139 683 173
rect 683 139 692 173
rect 640 124 692 139
rect 640 101 692 112
rect 640 67 649 101
rect 649 67 683 101
rect 683 67 692 101
rect 640 60 692 67
<< metal2 >>
rect 117 186 183 195
rect 117 130 122 186
rect 178 130 183 186
rect 117 126 124 130
rect 176 126 183 130
rect 117 114 183 126
rect 117 106 124 114
rect 176 106 183 114
rect 117 50 122 106
rect 178 50 183 106
rect 117 41 183 50
rect 289 186 355 195
rect 289 130 294 186
rect 350 130 355 186
rect 289 124 296 130
rect 348 124 355 130
rect 289 112 355 124
rect 289 106 296 112
rect 348 106 355 112
rect 289 50 294 106
rect 350 50 355 106
rect 289 41 355 50
rect 461 186 527 195
rect 461 130 466 186
rect 522 130 527 186
rect 461 124 468 130
rect 520 124 527 130
rect 461 112 527 124
rect 461 106 468 112
rect 520 106 527 112
rect 461 50 466 106
rect 522 50 527 106
rect 461 41 527 50
rect 633 186 699 195
rect 633 130 638 186
rect 694 130 699 186
rect 633 124 640 130
rect 692 124 699 130
rect 633 112 699 124
rect 633 106 640 112
rect 692 106 699 112
rect 633 50 638 106
rect 694 50 699 106
rect 633 41 699 50
<< via2 >>
rect 122 178 178 186
rect 122 130 124 178
rect 124 130 176 178
rect 176 130 178 178
rect 122 62 124 106
rect 124 62 176 106
rect 176 62 178 106
rect 122 50 178 62
rect 294 176 350 186
rect 294 130 296 176
rect 296 130 348 176
rect 348 130 350 176
rect 294 60 296 106
rect 296 60 348 106
rect 348 60 350 106
rect 294 50 350 60
rect 466 176 522 186
rect 466 130 468 176
rect 468 130 520 176
rect 520 130 522 176
rect 466 60 468 106
rect 468 60 520 106
rect 520 60 522 106
rect 466 50 522 60
rect 638 176 694 186
rect 638 130 640 176
rect 640 130 692 176
rect 692 130 694 176
rect 638 60 640 106
rect 640 60 692 106
rect 692 60 694 106
rect 638 50 694 60
<< metal3 >>
rect 117 186 699 195
rect 117 130 122 186
rect 178 130 294 186
rect 350 130 466 186
rect 522 130 638 186
rect 694 130 699 186
rect 117 129 699 130
rect 117 106 183 129
rect 117 50 122 106
rect 178 50 183 106
rect 117 41 183 50
rect 289 106 355 129
rect 289 50 294 106
rect 350 50 355 106
rect 289 41 355 50
rect 461 106 527 129
rect 461 50 466 106
rect 522 50 527 106
rect 461 41 527 50
rect 633 106 699 129
rect 633 50 638 106
rect 694 50 699 106
rect 633 41 699 50
<< labels >>
flabel metal3 s 117 129 699 195 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 127 239 689 297 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 41 -89 775 -29 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel pwell s 76 211 90 226 0 FreeSans 200 0 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 5963028
string GDS_START 5950406
string path 1.600 4.725 1.600 -2.225 
<< end >>
