magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3602 1975
<< nwell >>
rect -38 332 2342 704
<< pwell >>
rect 1 164 1564 190
rect 1 49 1987 164
rect 0 0 2304 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 263 368 299 592
rect 353 368 389 592
rect 443 368 479 592
rect 533 368 569 592
rect 623 368 659 592
rect 713 368 749 592
rect 803 368 839 592
rect 893 368 929 592
rect 983 368 1019 592
rect 1073 368 1109 592
rect 1173 368 1209 592
rect 1263 368 1299 592
rect 1363 368 1399 592
rect 1465 368 1501 592
rect 1555 368 1591 592
rect 1645 368 1681 592
rect 1735 368 1771 592
rect 1825 368 1861 592
rect 1915 368 1951 592
rect 2005 368 2041 592
rect 2095 368 2131 592
rect 2185 368 2221 592
<< nmoslvt >>
rect 84 80 114 164
rect 170 80 200 164
rect 256 80 286 164
rect 342 80 372 164
rect 442 80 472 164
rect 528 80 558 164
rect 628 80 658 164
rect 714 80 744 164
rect 828 80 858 164
rect 914 80 944 164
rect 1028 80 1058 164
rect 1114 80 1144 164
rect 1200 80 1230 164
rect 1286 80 1316 164
rect 1372 80 1402 164
rect 1458 80 1488 164
<< ndiff >>
rect 27 139 84 164
rect 27 105 39 139
rect 73 105 84 139
rect 27 80 84 105
rect 114 139 170 164
rect 114 105 125 139
rect 159 105 170 139
rect 114 80 170 105
rect 200 139 256 164
rect 200 105 211 139
rect 245 105 256 139
rect 200 80 256 105
rect 286 139 342 164
rect 286 105 297 139
rect 331 105 342 139
rect 286 80 342 105
rect 372 139 442 164
rect 372 105 383 139
rect 417 105 442 139
rect 372 80 442 105
rect 472 139 528 164
rect 472 105 483 139
rect 517 105 528 139
rect 472 80 528 105
rect 558 139 628 164
rect 558 105 569 139
rect 603 105 628 139
rect 558 80 628 105
rect 658 139 714 164
rect 658 105 669 139
rect 703 105 714 139
rect 658 80 714 105
rect 744 139 828 164
rect 744 105 769 139
rect 803 105 828 139
rect 744 80 828 105
rect 858 139 914 164
rect 858 105 869 139
rect 903 105 914 139
rect 858 80 914 105
rect 944 139 1028 164
rect 944 105 969 139
rect 1003 105 1028 139
rect 944 80 1028 105
rect 1058 139 1114 164
rect 1058 105 1069 139
rect 1103 105 1114 139
rect 1058 80 1114 105
rect 1144 139 1200 164
rect 1144 105 1155 139
rect 1189 105 1200 139
rect 1144 80 1200 105
rect 1230 139 1286 164
rect 1230 105 1241 139
rect 1275 105 1286 139
rect 1230 80 1286 105
rect 1316 139 1372 164
rect 1316 105 1327 139
rect 1361 105 1372 139
rect 1316 80 1372 105
rect 1402 139 1458 164
rect 1402 105 1413 139
rect 1447 105 1458 139
rect 1402 80 1458 105
rect 1488 138 1538 164
rect 1488 126 1961 138
rect 1488 92 1513 126
rect 1547 92 1593 126
rect 1627 92 1673 126
rect 1707 92 1755 126
rect 1789 92 1835 126
rect 1869 92 1915 126
rect 1949 92 1961 126
rect 1488 80 1961 92
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 497 173 546
rect 119 463 129 497
rect 163 463 173 497
rect 119 414 173 463
rect 119 380 129 414
rect 163 380 173 414
rect 119 368 173 380
rect 209 580 263 592
rect 209 546 219 580
rect 253 546 263 580
rect 209 497 263 546
rect 209 463 219 497
rect 253 463 263 497
rect 209 414 263 463
rect 209 380 219 414
rect 253 380 263 414
rect 209 368 263 380
rect 299 580 353 592
rect 299 546 309 580
rect 343 546 353 580
rect 299 497 353 546
rect 299 463 309 497
rect 343 463 353 497
rect 299 414 353 463
rect 299 380 309 414
rect 343 380 353 414
rect 299 368 353 380
rect 389 580 443 592
rect 389 546 399 580
rect 433 546 443 580
rect 389 497 443 546
rect 389 463 399 497
rect 433 463 443 497
rect 389 414 443 463
rect 389 380 399 414
rect 433 380 443 414
rect 389 368 443 380
rect 479 580 533 592
rect 479 546 489 580
rect 523 546 533 580
rect 479 497 533 546
rect 479 463 489 497
rect 523 463 533 497
rect 479 414 533 463
rect 479 380 489 414
rect 523 380 533 414
rect 479 368 533 380
rect 569 580 623 592
rect 569 546 579 580
rect 613 546 623 580
rect 569 497 623 546
rect 569 463 579 497
rect 613 463 623 497
rect 569 414 623 463
rect 569 380 579 414
rect 613 380 623 414
rect 569 368 623 380
rect 659 580 713 592
rect 659 546 669 580
rect 703 546 713 580
rect 659 497 713 546
rect 659 463 669 497
rect 703 463 713 497
rect 659 414 713 463
rect 659 380 669 414
rect 703 380 713 414
rect 659 368 713 380
rect 749 580 803 592
rect 749 546 759 580
rect 793 546 803 580
rect 749 497 803 546
rect 749 463 759 497
rect 793 463 803 497
rect 749 414 803 463
rect 749 380 759 414
rect 793 380 803 414
rect 749 368 803 380
rect 839 580 893 592
rect 839 546 849 580
rect 883 546 893 580
rect 839 497 893 546
rect 839 463 849 497
rect 883 463 893 497
rect 839 414 893 463
rect 839 380 849 414
rect 883 380 893 414
rect 839 368 893 380
rect 929 580 983 592
rect 929 546 939 580
rect 973 546 983 580
rect 929 497 983 546
rect 929 463 939 497
rect 973 463 983 497
rect 929 414 983 463
rect 929 380 939 414
rect 973 380 983 414
rect 929 368 983 380
rect 1019 580 1073 592
rect 1019 546 1029 580
rect 1063 546 1073 580
rect 1019 497 1073 546
rect 1019 463 1029 497
rect 1063 463 1073 497
rect 1019 414 1073 463
rect 1019 380 1029 414
rect 1063 380 1073 414
rect 1019 368 1073 380
rect 1109 580 1173 592
rect 1109 546 1119 580
rect 1153 546 1173 580
rect 1109 497 1173 546
rect 1109 463 1119 497
rect 1153 463 1173 497
rect 1109 414 1173 463
rect 1109 380 1119 414
rect 1153 380 1173 414
rect 1109 368 1173 380
rect 1209 580 1263 592
rect 1209 546 1219 580
rect 1253 546 1263 580
rect 1209 497 1263 546
rect 1209 463 1219 497
rect 1253 463 1263 497
rect 1209 414 1263 463
rect 1209 380 1219 414
rect 1253 380 1263 414
rect 1209 368 1263 380
rect 1299 580 1363 592
rect 1299 546 1309 580
rect 1343 546 1363 580
rect 1299 497 1363 546
rect 1299 463 1309 497
rect 1343 463 1363 497
rect 1299 414 1363 463
rect 1299 380 1309 414
rect 1343 380 1363 414
rect 1299 368 1363 380
rect 1399 580 1465 592
rect 1399 546 1415 580
rect 1449 546 1465 580
rect 1399 497 1465 546
rect 1399 463 1415 497
rect 1449 463 1465 497
rect 1399 414 1465 463
rect 1399 380 1415 414
rect 1449 380 1465 414
rect 1399 368 1465 380
rect 1501 580 1555 592
rect 1501 546 1511 580
rect 1545 546 1555 580
rect 1501 497 1555 546
rect 1501 463 1511 497
rect 1545 463 1555 497
rect 1501 414 1555 463
rect 1501 380 1511 414
rect 1545 380 1555 414
rect 1501 368 1555 380
rect 1591 580 1645 592
rect 1591 546 1601 580
rect 1635 546 1645 580
rect 1591 497 1645 546
rect 1591 463 1601 497
rect 1635 463 1645 497
rect 1591 414 1645 463
rect 1591 380 1601 414
rect 1635 380 1645 414
rect 1591 368 1645 380
rect 1681 580 1735 592
rect 1681 546 1691 580
rect 1725 546 1735 580
rect 1681 497 1735 546
rect 1681 463 1691 497
rect 1725 463 1735 497
rect 1681 414 1735 463
rect 1681 380 1691 414
rect 1725 380 1735 414
rect 1681 368 1735 380
rect 1771 580 1825 592
rect 1771 546 1781 580
rect 1815 546 1825 580
rect 1771 497 1825 546
rect 1771 463 1781 497
rect 1815 463 1825 497
rect 1771 414 1825 463
rect 1771 380 1781 414
rect 1815 380 1825 414
rect 1771 368 1825 380
rect 1861 580 1915 592
rect 1861 546 1871 580
rect 1905 546 1915 580
rect 1861 497 1915 546
rect 1861 463 1871 497
rect 1905 463 1915 497
rect 1861 414 1915 463
rect 1861 380 1871 414
rect 1905 380 1915 414
rect 1861 368 1915 380
rect 1951 580 2005 592
rect 1951 546 1961 580
rect 1995 546 2005 580
rect 1951 497 2005 546
rect 1951 463 1961 497
rect 1995 463 2005 497
rect 1951 414 2005 463
rect 1951 380 1961 414
rect 1995 380 2005 414
rect 1951 368 2005 380
rect 2041 580 2095 592
rect 2041 546 2051 580
rect 2085 546 2095 580
rect 2041 497 2095 546
rect 2041 463 2051 497
rect 2085 463 2095 497
rect 2041 414 2095 463
rect 2041 380 2051 414
rect 2085 380 2095 414
rect 2041 368 2095 380
rect 2131 580 2185 592
rect 2131 546 2141 580
rect 2175 546 2185 580
rect 2131 497 2185 546
rect 2131 463 2141 497
rect 2175 463 2185 497
rect 2131 414 2185 463
rect 2131 380 2141 414
rect 2175 380 2185 414
rect 2131 368 2185 380
rect 2221 580 2277 592
rect 2221 546 2231 580
rect 2265 546 2277 580
rect 2221 497 2277 546
rect 2221 463 2231 497
rect 2265 463 2277 497
rect 2221 414 2277 463
rect 2221 380 2231 414
rect 2265 380 2277 414
rect 2221 368 2277 380
<< ndiffc >>
rect 39 105 73 139
rect 125 105 159 139
rect 211 105 245 139
rect 297 105 331 139
rect 383 105 417 139
rect 483 105 517 139
rect 569 105 603 139
rect 669 105 703 139
rect 769 105 803 139
rect 869 105 903 139
rect 969 105 1003 139
rect 1069 105 1103 139
rect 1155 105 1189 139
rect 1241 105 1275 139
rect 1327 105 1361 139
rect 1413 105 1447 139
rect 1513 92 1547 126
rect 1593 92 1627 126
rect 1673 92 1707 126
rect 1755 92 1789 126
rect 1835 92 1869 126
rect 1915 92 1949 126
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 219 546 253 580
rect 219 463 253 497
rect 219 380 253 414
rect 309 546 343 580
rect 309 463 343 497
rect 309 380 343 414
rect 399 546 433 580
rect 399 463 433 497
rect 399 380 433 414
rect 489 546 523 580
rect 489 463 523 497
rect 489 380 523 414
rect 579 546 613 580
rect 579 463 613 497
rect 579 380 613 414
rect 669 546 703 580
rect 669 463 703 497
rect 669 380 703 414
rect 759 546 793 580
rect 759 463 793 497
rect 759 380 793 414
rect 849 546 883 580
rect 849 463 883 497
rect 849 380 883 414
rect 939 546 973 580
rect 939 463 973 497
rect 939 380 973 414
rect 1029 546 1063 580
rect 1029 463 1063 497
rect 1029 380 1063 414
rect 1119 546 1153 580
rect 1119 463 1153 497
rect 1119 380 1153 414
rect 1219 546 1253 580
rect 1219 463 1253 497
rect 1219 380 1253 414
rect 1309 546 1343 580
rect 1309 463 1343 497
rect 1309 380 1343 414
rect 1415 546 1449 580
rect 1415 463 1449 497
rect 1415 380 1449 414
rect 1511 546 1545 580
rect 1511 463 1545 497
rect 1511 380 1545 414
rect 1601 546 1635 580
rect 1601 463 1635 497
rect 1601 380 1635 414
rect 1691 546 1725 580
rect 1691 463 1725 497
rect 1691 380 1725 414
rect 1781 546 1815 580
rect 1781 463 1815 497
rect 1781 380 1815 414
rect 1871 546 1905 580
rect 1871 463 1905 497
rect 1871 380 1905 414
rect 1961 546 1995 580
rect 1961 463 1995 497
rect 1961 380 1995 414
rect 2051 546 2085 580
rect 2051 463 2085 497
rect 2051 380 2085 414
rect 2141 546 2175 580
rect 2141 463 2175 497
rect 2141 380 2175 414
rect 2231 546 2265 580
rect 2231 463 2265 497
rect 2231 380 2265 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 263 592 299 618
rect 353 592 389 618
rect 443 592 479 618
rect 533 592 569 618
rect 623 592 659 618
rect 713 592 749 618
rect 803 592 839 618
rect 893 592 929 618
rect 983 592 1019 618
rect 1073 592 1109 618
rect 1173 592 1209 618
rect 1263 592 1299 618
rect 1363 592 1399 618
rect 1465 592 1501 618
rect 1555 592 1591 618
rect 1645 592 1681 618
rect 1735 592 1771 618
rect 1825 592 1861 618
rect 1915 592 1951 618
rect 2005 592 2041 618
rect 2095 592 2131 618
rect 2185 592 2221 618
rect 83 336 119 368
rect 173 336 209 368
rect 263 336 299 368
rect 353 336 389 368
rect 443 336 479 368
rect 533 336 569 368
rect 623 336 659 368
rect 713 336 749 368
rect 803 336 839 368
rect 893 336 929 368
rect 983 336 1019 368
rect 1073 336 1109 368
rect 1173 336 1209 368
rect 1263 336 1299 368
rect 1363 336 1399 368
rect 1465 336 1501 368
rect 1555 336 1591 368
rect 1645 336 1681 368
rect 1735 336 1771 368
rect 1825 336 1861 368
rect 1915 336 1951 368
rect 2005 336 2041 368
rect 2095 336 2131 368
rect 2185 336 2221 368
rect 83 314 2221 336
rect 83 300 209 314
rect 84 280 209 300
rect 243 280 389 314
rect 423 280 583 314
rect 617 280 769 314
rect 803 280 967 314
rect 1001 280 1135 314
rect 1169 280 1325 314
rect 1359 280 1521 314
rect 1555 280 1589 314
rect 1623 280 1657 314
rect 1691 280 1725 314
rect 1759 280 1793 314
rect 1827 280 1861 314
rect 1895 280 1929 314
rect 1963 280 1997 314
rect 2031 280 2065 314
rect 2099 280 2133 314
rect 2167 280 2221 314
rect 84 264 2221 280
rect 84 164 114 264
rect 170 164 200 264
rect 256 164 286 264
rect 342 164 372 264
rect 442 164 472 264
rect 528 164 558 264
rect 628 164 658 264
rect 714 164 744 264
rect 828 164 858 264
rect 914 164 944 264
rect 1028 164 1058 264
rect 1114 164 1144 264
rect 1200 164 1230 264
rect 1286 164 1316 264
rect 1372 164 1402 264
rect 1458 164 1488 264
rect 84 54 114 80
rect 170 54 200 80
rect 256 54 286 80
rect 342 54 372 80
rect 442 54 472 80
rect 528 54 558 80
rect 628 54 658 80
rect 714 54 744 80
rect 828 54 858 80
rect 914 54 944 80
rect 1028 54 1058 80
rect 1114 54 1144 80
rect 1200 54 1230 80
rect 1286 54 1316 80
rect 1372 54 1402 80
rect 1458 54 1488 80
<< polycont >>
rect 209 280 243 314
rect 389 280 423 314
rect 583 280 617 314
rect 769 280 803 314
rect 967 280 1001 314
rect 1135 280 1169 314
rect 1325 280 1359 314
rect 1521 280 1555 314
rect 1589 280 1623 314
rect 1657 280 1691 314
rect 1725 280 1759 314
rect 1793 280 1827 314
rect 1861 280 1895 314
rect 1929 280 1963 314
rect 1997 280 2031 314
rect 2065 280 2099 314
rect 2133 280 2167 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 497 89 546
rect 23 463 39 497
rect 73 463 89 497
rect 23 414 89 463
rect 23 380 39 414
rect 73 380 89 414
rect 125 580 163 596
rect 125 546 129 580
rect 125 497 163 546
rect 125 463 129 497
rect 125 424 163 463
rect 125 390 127 424
rect 161 414 163 424
rect 125 380 129 390
rect 125 364 163 380
rect 203 580 253 649
rect 203 546 219 580
rect 203 497 253 546
rect 203 463 219 497
rect 203 414 253 463
rect 203 380 219 414
rect 203 364 253 380
rect 293 580 359 596
rect 293 546 309 580
rect 343 546 359 580
rect 293 497 359 546
rect 293 463 309 497
rect 343 463 359 497
rect 293 424 359 463
rect 293 380 309 424
rect 343 380 359 424
rect 293 377 359 380
rect 399 580 433 649
rect 399 497 433 546
rect 399 414 433 463
rect 23 139 89 168
rect 125 155 161 364
rect 195 314 259 330
rect 195 280 209 314
rect 243 280 259 314
rect 195 276 259 280
rect 195 242 209 276
rect 243 242 259 276
rect 195 230 259 242
rect 23 105 39 139
rect 73 105 89 139
rect 23 17 89 105
rect 123 139 161 155
rect 123 105 125 139
rect 159 105 161 139
rect 123 76 161 105
rect 195 139 252 168
rect 293 155 339 377
rect 399 364 433 380
rect 473 580 539 596
rect 473 546 489 580
rect 523 546 539 580
rect 473 497 539 546
rect 473 463 489 497
rect 523 463 539 497
rect 473 424 539 463
rect 473 380 489 424
rect 523 380 539 424
rect 473 377 539 380
rect 579 580 613 649
rect 579 497 613 546
rect 579 414 613 463
rect 373 314 439 330
rect 373 280 389 314
rect 423 280 439 314
rect 373 276 439 280
rect 373 242 389 276
rect 423 242 439 276
rect 373 230 439 242
rect 195 105 211 139
rect 245 105 252 139
rect 195 17 252 105
rect 288 139 340 155
rect 288 105 297 139
rect 331 105 340 139
rect 288 76 340 105
rect 377 139 433 168
rect 473 155 533 377
rect 579 364 613 380
rect 667 580 719 596
rect 667 546 669 580
rect 703 546 719 580
rect 667 497 719 546
rect 667 463 669 497
rect 703 463 719 497
rect 667 424 719 463
rect 667 414 675 424
rect 667 380 669 414
rect 709 390 719 424
rect 703 380 719 390
rect 567 314 633 330
rect 567 280 583 314
rect 617 280 633 314
rect 567 276 633 280
rect 567 242 583 276
rect 617 242 633 276
rect 567 230 633 242
rect 377 105 383 139
rect 417 105 433 139
rect 377 17 433 105
rect 470 139 533 155
rect 470 105 483 139
rect 517 105 533 139
rect 470 76 533 105
rect 569 139 619 168
rect 667 155 719 380
rect 759 580 793 649
rect 759 497 793 546
rect 759 414 793 463
rect 759 364 793 380
rect 833 580 899 596
rect 833 546 849 580
rect 883 546 899 580
rect 833 497 899 546
rect 833 463 849 497
rect 883 463 899 497
rect 833 424 899 463
rect 833 380 849 424
rect 883 380 899 424
rect 939 580 973 649
rect 939 497 973 546
rect 939 414 973 463
rect 833 370 905 380
rect 753 314 819 330
rect 753 280 769 314
rect 803 280 819 314
rect 753 276 819 280
rect 753 242 769 276
rect 803 242 819 276
rect 753 230 819 242
rect 603 105 619 139
rect 569 17 619 105
rect 660 139 719 155
rect 660 105 669 139
rect 703 105 719 139
rect 660 76 719 105
rect 753 139 819 168
rect 753 105 769 139
rect 803 105 819 139
rect 753 17 819 105
rect 853 139 905 370
rect 939 364 973 380
rect 1013 580 1079 596
rect 1013 546 1029 580
rect 1063 546 1079 580
rect 1013 497 1079 546
rect 1013 463 1029 497
rect 1063 463 1079 497
rect 1013 424 1079 463
rect 1013 380 1029 424
rect 1063 402 1079 424
rect 1119 580 1169 649
rect 1153 546 1169 580
rect 1119 497 1169 546
rect 1153 463 1169 497
rect 1119 414 1169 463
rect 1063 380 1085 402
rect 1013 370 1085 380
rect 951 314 1017 330
rect 951 280 967 314
rect 1001 280 1017 314
rect 951 276 1017 280
rect 951 242 967 276
rect 1001 242 1017 276
rect 951 230 1017 242
rect 853 105 869 139
rect 903 105 905 139
rect 853 76 905 105
rect 953 139 1017 168
rect 953 105 969 139
rect 1003 105 1017 139
rect 953 17 1017 105
rect 1051 155 1085 370
rect 1153 380 1169 414
rect 1119 364 1169 380
rect 1203 580 1266 596
rect 1203 546 1219 580
rect 1253 546 1266 580
rect 1203 497 1266 546
rect 1203 463 1219 497
rect 1253 463 1266 497
rect 1203 424 1266 463
rect 1203 380 1219 424
rect 1253 380 1266 424
rect 1203 364 1266 380
rect 1302 580 1359 649
rect 1302 546 1309 580
rect 1343 546 1359 580
rect 1302 497 1359 546
rect 1302 463 1309 497
rect 1343 463 1359 497
rect 1302 414 1359 463
rect 1302 380 1309 414
rect 1343 380 1359 414
rect 1302 364 1359 380
rect 1409 580 1458 596
rect 1409 546 1415 580
rect 1449 546 1458 580
rect 1409 497 1458 546
rect 1409 463 1415 497
rect 1449 463 1458 497
rect 1409 424 1458 463
rect 1409 380 1415 424
rect 1449 380 1458 424
rect 1219 352 1266 364
rect 1119 314 1185 330
rect 1119 280 1135 314
rect 1169 280 1185 314
rect 1119 276 1185 280
rect 1119 242 1135 276
rect 1169 242 1185 276
rect 1119 230 1185 242
rect 1219 202 1268 352
rect 1309 314 1375 330
rect 1309 280 1325 314
rect 1359 280 1375 314
rect 1309 276 1375 280
rect 1309 242 1325 276
rect 1359 242 1375 276
rect 1309 230 1375 242
rect 1051 139 1105 155
rect 1051 105 1069 139
rect 1103 105 1105 139
rect 1051 76 1105 105
rect 1139 139 1196 168
rect 1139 105 1155 139
rect 1189 105 1196 139
rect 1139 17 1196 105
rect 1232 157 1268 202
rect 1232 139 1277 157
rect 1232 105 1241 139
rect 1275 105 1277 139
rect 1232 76 1277 105
rect 1311 139 1375 168
rect 1311 105 1327 139
rect 1361 105 1375 139
rect 1311 17 1375 105
rect 1409 139 1458 380
rect 1495 580 1561 649
rect 1495 546 1511 580
rect 1545 546 1561 580
rect 1495 497 1561 546
rect 1495 463 1511 497
rect 1545 463 1561 497
rect 1495 414 1561 463
rect 1495 380 1511 414
rect 1545 380 1561 414
rect 1495 364 1561 380
rect 1601 580 1635 596
rect 1601 497 1635 546
rect 1601 424 1635 463
rect 1601 364 1635 380
rect 1675 580 1725 649
rect 1675 546 1691 580
rect 1675 497 1725 546
rect 1675 463 1691 497
rect 1675 414 1725 463
rect 1675 380 1691 414
rect 1675 364 1725 380
rect 1781 580 1815 596
rect 1781 497 1815 546
rect 1781 424 1815 463
rect 1781 364 1815 380
rect 1855 580 1921 649
rect 1855 546 1871 580
rect 1905 546 1921 580
rect 1855 497 1921 546
rect 1855 463 1871 497
rect 1905 463 1921 497
rect 1855 414 1921 463
rect 1855 380 1871 414
rect 1905 380 1921 414
rect 1855 364 1921 380
rect 1961 580 1995 596
rect 1961 497 1995 546
rect 1961 424 1995 463
rect 1961 364 1995 380
rect 2035 580 2101 649
rect 2035 546 2051 580
rect 2085 546 2101 580
rect 2035 497 2101 546
rect 2035 463 2051 497
rect 2085 463 2101 497
rect 2035 414 2101 463
rect 2035 380 2051 414
rect 2085 380 2101 414
rect 2035 364 2101 380
rect 2141 580 2175 596
rect 2141 497 2175 546
rect 2141 424 2175 463
rect 2141 364 2175 380
rect 2215 580 2281 649
rect 2215 546 2231 580
rect 2265 546 2281 580
rect 2215 497 2281 546
rect 2215 463 2231 497
rect 2265 463 2281 497
rect 2215 414 2281 463
rect 2215 380 2231 414
rect 2265 380 2281 414
rect 2215 364 2281 380
rect 1505 314 2183 330
rect 1505 280 1521 314
rect 1555 280 1589 314
rect 1623 280 1657 314
rect 1691 280 1725 314
rect 1759 280 1793 314
rect 1827 280 1861 314
rect 1895 280 1929 314
rect 1963 280 1997 314
rect 2031 280 2065 314
rect 2099 280 2133 314
rect 2167 280 2183 314
rect 1505 276 2183 280
rect 1505 242 1549 276
rect 1583 242 1621 276
rect 1655 242 1693 276
rect 1727 242 1765 276
rect 1799 242 1837 276
rect 1871 242 1909 276
rect 1943 242 1981 276
rect 2015 242 2053 276
rect 2087 242 2125 276
rect 2159 242 2183 276
rect 1505 230 2183 242
rect 1409 105 1413 139
rect 1447 105 1458 139
rect 1409 76 1458 105
rect 1497 126 1965 142
rect 1497 92 1513 126
rect 1547 92 1593 126
rect 1627 92 1673 126
rect 1707 92 1755 126
rect 1789 92 1835 126
rect 1869 92 1915 126
rect 1949 92 1965 126
rect 1497 17 1965 92
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 127 414 161 424
rect 127 390 129 414
rect 129 390 161 414
rect 309 414 343 424
rect 309 390 343 414
rect 209 242 243 276
rect 489 414 523 424
rect 489 390 523 414
rect 389 242 423 276
rect 675 414 709 424
rect 675 390 703 414
rect 703 390 709 414
rect 583 242 617 276
rect 849 414 883 424
rect 849 390 883 414
rect 769 242 803 276
rect 1029 414 1063 424
rect 1029 390 1063 414
rect 967 242 1001 276
rect 1219 414 1253 424
rect 1219 390 1253 414
rect 1415 414 1449 424
rect 1415 390 1449 414
rect 1135 242 1169 276
rect 1325 242 1359 276
rect 1601 414 1635 424
rect 1601 390 1635 414
rect 1781 414 1815 424
rect 1781 390 1815 414
rect 1961 414 1995 424
rect 1961 390 1995 414
rect 2141 414 2175 424
rect 2141 390 2175 414
rect 1549 242 1583 276
rect 1621 242 1655 276
rect 1693 242 1727 276
rect 1765 242 1799 276
rect 1837 242 1871 276
rect 1909 242 1943 276
rect 1981 242 2015 276
rect 2053 242 2087 276
rect 2125 242 2159 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 115 424 2187 430
rect 115 390 127 424
rect 161 390 309 424
rect 343 390 489 424
rect 523 390 675 424
rect 709 390 849 424
rect 883 390 1029 424
rect 1063 390 1219 424
rect 1253 390 1415 424
rect 1449 390 1601 424
rect 1635 390 1781 424
rect 1815 390 1961 424
rect 1995 390 2141 424
rect 2175 390 2187 424
rect 115 384 2187 390
rect 197 276 2187 282
rect 197 242 209 276
rect 243 242 389 276
rect 423 242 583 276
rect 617 242 769 276
rect 803 242 967 276
rect 1001 242 1135 276
rect 1169 242 1325 276
rect 1359 242 1549 276
rect 1583 242 1621 276
rect 1655 242 1693 276
rect 1727 242 1765 276
rect 1799 242 1837 276
rect 1871 242 1909 276
rect 1943 242 1981 276
rect 2015 242 2053 276
rect 2087 242 2125 276
rect 2159 242 2187 276
rect 197 236 2187 242
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
flabel pwell s 0 0 2304 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 2304 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkinv_16
flabel metal1 s 0 617 2304 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 2304 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 197 236 2187 282 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel metal1 s 115 384 2187 430 0 FreeSans 400 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2304 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 2675646
string GDS_START 2658066
<< end >>
