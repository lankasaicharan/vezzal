magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 356 1382 704
rect -38 332 232 356
rect 581 332 1382 356
<< pwell >>
rect 337 248 444 294
rect 22 228 539 248
rect 22 184 750 228
rect 932 184 1308 248
rect 22 49 1308 184
rect 0 0 1344 49
<< scpmos >>
rect 86 424 116 592
rect 186 424 216 592
rect 422 392 452 560
rect 538 392 568 592
rect 622 392 652 592
rect 729 508 759 592
rect 860 508 890 592
rect 1012 392 1042 592
rect 1112 392 1142 592
rect 1228 368 1258 592
<< nmoslvt >>
rect 105 112 135 222
rect 222 74 252 222
rect 433 74 463 222
rect 535 74 565 202
rect 613 74 643 202
rect 739 74 769 158
rect 817 74 847 158
rect 1015 74 1045 222
rect 1093 74 1123 222
rect 1195 74 1225 222
<< ndiff >>
rect 363 256 418 268
rect 363 222 375 256
rect 409 222 418 256
rect 48 184 105 222
rect 48 150 60 184
rect 94 150 105 184
rect 48 112 105 150
rect 135 210 222 222
rect 135 176 177 210
rect 211 176 222 210
rect 135 120 222 176
rect 135 112 177 120
rect 165 86 177 112
rect 211 86 222 120
rect 165 74 222 86
rect 252 210 309 222
rect 252 176 263 210
rect 297 176 309 210
rect 252 120 309 176
rect 252 86 263 120
rect 297 86 309 120
rect 252 74 309 86
rect 363 74 433 222
rect 463 202 513 222
rect 463 120 535 202
rect 463 86 480 120
rect 514 86 535 120
rect 463 74 535 86
rect 565 74 613 202
rect 643 169 724 202
rect 643 135 666 169
rect 700 158 724 169
rect 958 210 1015 222
rect 958 176 970 210
rect 1004 176 1015 210
rect 700 135 739 158
rect 643 74 739 135
rect 769 74 817 158
rect 847 133 904 158
rect 847 99 858 133
rect 892 99 904 133
rect 847 74 904 99
rect 958 120 1015 176
rect 958 86 970 120
rect 1004 86 1015 120
rect 958 74 1015 86
rect 1045 74 1093 222
rect 1123 152 1195 222
rect 1123 118 1134 152
rect 1168 118 1195 152
rect 1123 74 1195 118
rect 1225 152 1282 222
rect 1225 118 1236 152
rect 1270 118 1282 152
rect 1225 74 1282 118
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 470 86 546
rect 27 436 39 470
rect 73 436 86 470
rect 27 424 86 436
rect 116 580 186 592
rect 116 546 139 580
rect 173 546 186 580
rect 116 424 186 546
rect 216 444 309 592
rect 470 580 538 592
rect 470 560 486 580
rect 216 424 254 444
rect 234 410 254 424
rect 288 410 309 444
rect 234 398 309 410
rect 363 441 422 560
rect 363 407 375 441
rect 409 407 422 441
rect 363 392 422 407
rect 452 546 486 560
rect 520 546 538 580
rect 452 392 538 546
rect 568 392 622 592
rect 652 531 729 592
rect 652 497 665 531
rect 699 508 729 531
rect 759 508 860 592
rect 890 580 1012 592
rect 890 546 934 580
rect 968 546 1012 580
rect 890 508 1012 546
rect 699 497 711 508
rect 652 392 711 497
rect 959 392 1012 508
rect 1042 580 1112 592
rect 1042 546 1065 580
rect 1099 546 1112 580
rect 1042 510 1112 546
rect 1042 476 1065 510
rect 1099 476 1112 510
rect 1042 440 1112 476
rect 1042 406 1065 440
rect 1099 406 1112 440
rect 1042 392 1112 406
rect 1142 580 1228 592
rect 1142 546 1165 580
rect 1199 546 1228 580
rect 1142 510 1228 546
rect 1142 476 1165 510
rect 1199 476 1228 510
rect 1142 440 1228 476
rect 1142 406 1165 440
rect 1199 406 1228 440
rect 1142 392 1228 406
rect 1175 368 1228 392
rect 1258 580 1317 592
rect 1258 546 1271 580
rect 1305 546 1317 580
rect 1258 497 1317 546
rect 1258 463 1271 497
rect 1305 463 1317 497
rect 1258 414 1317 463
rect 1258 380 1271 414
rect 1305 380 1317 414
rect 1258 368 1317 380
<< ndiffc >>
rect 375 222 409 256
rect 60 150 94 184
rect 177 176 211 210
rect 177 86 211 120
rect 263 176 297 210
rect 263 86 297 120
rect 480 86 514 120
rect 666 135 700 169
rect 970 176 1004 210
rect 858 99 892 133
rect 970 86 1004 120
rect 1134 118 1168 152
rect 1236 118 1270 152
<< pdiffc >>
rect 39 546 73 580
rect 39 436 73 470
rect 139 546 173 580
rect 254 410 288 444
rect 375 407 409 441
rect 486 546 520 580
rect 665 497 699 531
rect 934 546 968 580
rect 1065 546 1099 580
rect 1065 476 1099 510
rect 1065 406 1099 440
rect 1165 546 1199 580
rect 1165 476 1199 510
rect 1165 406 1199 440
rect 1271 546 1305 580
rect 1271 463 1305 497
rect 1271 380 1305 414
<< poly >>
rect 86 592 116 618
rect 186 592 216 618
rect 538 592 568 618
rect 622 592 652 618
rect 729 592 759 618
rect 860 592 890 618
rect 1012 592 1042 618
rect 1112 592 1142 618
rect 1228 592 1258 618
rect 422 560 452 586
rect 86 409 116 424
rect 186 409 216 424
rect 83 338 119 409
rect 183 356 219 409
rect 729 493 759 508
rect 860 493 890 508
rect 726 476 762 493
rect 857 476 893 493
rect 726 460 809 476
rect 726 426 759 460
rect 793 426 809 460
rect 857 460 927 476
rect 857 446 877 460
rect 726 410 809 426
rect 861 426 877 446
rect 911 426 927 460
rect 861 410 927 426
rect 422 377 452 392
rect 538 377 568 392
rect 622 377 652 392
rect 183 340 252 356
rect 83 326 113 338
rect 21 310 113 326
rect 21 276 37 310
rect 71 290 113 310
rect 183 306 202 340
rect 236 306 252 340
rect 183 290 252 306
rect 300 340 366 356
rect 300 306 316 340
rect 350 320 366 340
rect 419 320 455 377
rect 535 360 571 377
rect 505 344 571 360
rect 350 306 463 320
rect 300 290 463 306
rect 505 310 521 344
rect 555 310 571 344
rect 619 368 655 377
rect 619 338 769 368
rect 505 294 571 310
rect 739 311 769 338
rect 739 295 819 311
rect 71 276 135 290
rect 21 260 135 276
rect 105 222 135 260
rect 222 222 252 290
rect 433 222 463 290
rect 105 86 135 112
rect 535 202 565 294
rect 613 274 679 290
rect 613 240 629 274
rect 663 240 679 274
rect 613 224 679 240
rect 739 261 769 295
rect 803 261 819 295
rect 739 245 819 261
rect 613 202 643 224
rect 739 158 769 245
rect 861 203 891 410
rect 1012 377 1042 392
rect 1112 377 1142 392
rect 1009 360 1045 377
rect 933 344 1045 360
rect 933 310 949 344
rect 983 310 1045 344
rect 1109 336 1145 377
rect 1228 353 1258 368
rect 933 294 1045 310
rect 1015 222 1045 294
rect 1087 320 1153 336
rect 1087 286 1103 320
rect 1137 286 1153 320
rect 1225 310 1261 353
rect 1087 270 1153 286
rect 1195 294 1261 310
rect 1093 222 1123 270
rect 1195 260 1211 294
rect 1245 260 1261 294
rect 1195 244 1261 260
rect 1195 222 1225 244
rect 817 173 891 203
rect 817 158 847 173
rect 222 48 252 74
rect 433 48 463 74
rect 535 48 565 74
rect 613 48 643 74
rect 739 48 769 74
rect 817 48 847 74
rect 1015 48 1045 74
rect 1093 48 1123 74
rect 1195 48 1225 74
<< polycont >>
rect 759 426 793 460
rect 877 426 911 460
rect 37 276 71 310
rect 202 306 236 340
rect 316 306 350 340
rect 521 310 555 344
rect 629 240 663 274
rect 769 261 803 295
rect 949 310 983 344
rect 1103 286 1137 320
rect 1211 260 1245 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 123 580 189 649
rect 123 546 139 580
rect 173 546 189 580
rect 466 580 541 649
rect 466 546 486 580
rect 520 546 541 580
rect 581 581 809 615
rect 23 512 89 546
rect 23 478 539 512
rect 23 470 143 478
rect 23 436 39 470
rect 73 436 143 470
rect 23 420 143 436
rect 21 310 75 356
rect 21 276 37 310
rect 71 276 75 310
rect 21 260 75 276
rect 109 226 143 420
rect 230 410 254 444
rect 288 410 325 444
rect 230 394 325 410
rect 359 441 434 444
rect 359 407 375 441
rect 409 407 434 441
rect 359 404 434 407
rect 291 356 325 394
rect 186 340 257 356
rect 186 306 202 340
rect 236 306 257 340
rect 186 290 257 306
rect 291 340 366 356
rect 291 306 316 340
rect 350 306 366 340
rect 291 290 366 306
rect 291 226 325 290
rect 400 256 434 404
rect 505 360 539 478
rect 581 428 615 581
rect 649 531 707 547
rect 649 497 665 531
rect 699 497 707 531
rect 649 481 707 497
rect 581 394 639 428
rect 505 344 571 360
rect 505 310 521 344
rect 555 310 571 344
rect 505 294 571 310
rect 605 290 639 394
rect 673 379 707 481
rect 743 460 809 581
rect 887 580 1015 649
rect 887 546 934 580
rect 968 546 1015 580
rect 887 530 1015 546
rect 1049 580 1115 596
rect 1049 546 1065 580
rect 1099 546 1115 580
rect 1049 510 1115 546
rect 1049 476 1065 510
rect 1099 476 1115 510
rect 743 426 759 460
rect 793 426 809 460
rect 743 413 809 426
rect 861 460 1115 476
rect 861 426 877 460
rect 911 440 1115 460
rect 911 426 1065 440
rect 861 413 1065 426
rect 1019 406 1065 413
rect 1099 406 1115 440
rect 1019 390 1115 406
rect 1149 580 1215 649
rect 1149 546 1165 580
rect 1199 546 1215 580
rect 1149 510 1215 546
rect 1149 476 1165 510
rect 1199 476 1215 510
rect 1149 440 1215 476
rect 1149 406 1165 440
rect 1199 406 1215 440
rect 1149 390 1215 406
rect 1255 580 1327 596
rect 1255 546 1271 580
rect 1305 546 1327 580
rect 1255 497 1327 546
rect 1255 463 1271 497
rect 1305 463 1327 497
rect 1255 414 1327 463
rect 673 345 985 379
rect 605 274 665 290
rect 605 256 629 274
rect 44 184 143 226
rect 44 150 60 184
rect 94 150 143 184
rect 44 108 143 150
rect 177 210 211 226
rect 177 120 211 176
rect 177 17 211 86
rect 247 210 325 226
rect 359 222 375 256
rect 409 240 629 256
rect 663 240 665 274
rect 409 222 665 240
rect 247 176 263 210
rect 297 188 325 210
rect 297 176 604 188
rect 699 185 733 345
rect 933 344 985 345
rect 247 154 604 176
rect 247 120 325 154
rect 247 86 263 120
rect 297 86 325 120
rect 247 70 325 86
rect 459 86 480 120
rect 514 86 536 120
rect 459 17 536 86
rect 570 85 604 154
rect 638 169 733 185
rect 638 135 666 169
rect 700 135 733 169
rect 638 119 733 135
rect 767 295 819 311
rect 767 261 769 295
rect 803 261 819 295
rect 933 310 949 344
rect 983 310 985 344
rect 933 294 985 310
rect 767 245 819 261
rect 767 85 801 245
rect 1019 236 1053 390
rect 1255 380 1271 414
rect 1305 380 1327 414
rect 1255 364 1327 380
rect 1087 320 1153 356
rect 1087 286 1103 320
rect 1137 286 1153 320
rect 1087 270 1153 286
rect 1195 294 1259 310
rect 1195 260 1211 294
rect 1245 260 1259 294
rect 1195 236 1259 260
rect 954 210 1259 236
rect 954 176 970 210
rect 1004 202 1259 210
rect 1004 176 1020 202
rect 570 51 801 85
rect 842 133 908 162
rect 842 99 858 133
rect 892 99 908 133
rect 842 17 908 99
rect 954 120 1020 176
rect 1293 168 1327 364
rect 954 86 970 120
rect 1004 86 1020 120
rect 954 70 1020 86
rect 1118 152 1184 168
rect 1118 118 1134 152
rect 1168 118 1184 152
rect 1118 17 1184 118
rect 1220 152 1327 168
rect 1220 118 1236 152
rect 1270 118 1327 152
rect 1220 70 1327 118
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlrtp_1
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1279 94 1313 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 900494
string GDS_START 890208
<< end >>
