magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 112 49 674 273
rect 0 0 768 49
<< scnmos >>
rect 191 47 591 247
<< scpmoshvt >>
rect 178 419 578 619
<< ndiff >>
rect 138 229 191 247
rect 138 195 146 229
rect 180 195 191 229
rect 138 161 191 195
rect 138 127 146 161
rect 180 127 191 161
rect 138 93 191 127
rect 138 59 146 93
rect 180 59 191 93
rect 138 47 191 59
rect 591 225 648 247
rect 591 191 602 225
rect 636 191 648 225
rect 591 157 648 191
rect 591 123 602 157
rect 636 123 648 157
rect 591 89 648 123
rect 591 55 602 89
rect 636 55 648 89
rect 591 47 648 55
<< pdiff >>
rect 123 607 178 619
rect 123 573 131 607
rect 165 573 178 607
rect 123 539 178 573
rect 123 505 131 539
rect 165 505 178 539
rect 123 471 178 505
rect 123 437 131 471
rect 165 437 178 471
rect 123 419 178 437
rect 578 611 635 619
rect 578 577 589 611
rect 623 577 635 611
rect 578 543 635 577
rect 578 509 589 543
rect 623 509 635 543
rect 578 475 635 509
rect 578 441 589 475
rect 623 441 635 475
rect 578 419 635 441
<< ndiffc >>
rect 146 195 180 229
rect 146 127 180 161
rect 146 59 180 93
rect 602 191 636 225
rect 602 123 636 157
rect 602 55 636 89
<< pdiffc >>
rect 131 573 165 607
rect 131 505 165 539
rect 131 437 165 471
rect 589 577 623 611
rect 589 509 623 543
rect 589 441 623 475
<< poly >>
rect 178 619 578 645
rect 178 387 578 419
rect 174 377 578 387
rect 174 371 312 377
rect 174 337 194 371
rect 228 337 262 371
rect 296 337 312 371
rect 174 321 312 337
rect 391 319 593 335
rect 391 285 407 319
rect 441 285 475 319
rect 509 285 543 319
rect 577 285 593 319
rect 391 273 593 285
rect 191 262 593 273
rect 191 247 591 262
rect 191 21 591 47
<< polycont >>
rect 194 337 228 371
rect 262 337 296 371
rect 407 285 441 319
rect 475 285 509 319
rect 543 285 577 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 115 607 181 649
rect 115 573 131 607
rect 165 573 181 607
rect 115 539 181 573
rect 115 505 131 539
rect 165 505 181 539
rect 115 471 181 505
rect 115 437 131 471
rect 165 437 181 471
rect 115 421 181 437
rect 573 611 639 649
rect 573 577 589 611
rect 623 577 639 611
rect 573 543 639 577
rect 573 509 589 543
rect 623 509 639 543
rect 573 475 639 509
rect 573 441 589 475
rect 623 441 639 475
rect 130 371 312 387
rect 130 337 194 371
rect 228 337 262 371
rect 296 337 312 371
rect 130 321 312 337
rect 573 335 639 441
rect 130 229 196 321
rect 391 319 639 335
rect 391 285 407 319
rect 441 285 475 319
rect 509 285 543 319
rect 577 285 639 319
rect 391 268 639 285
rect 130 195 146 229
rect 180 195 196 229
rect 130 161 196 195
rect 130 127 146 161
rect 180 127 196 161
rect 130 93 196 127
rect 130 59 146 93
rect 180 59 196 93
rect 130 17 196 59
rect 586 191 602 225
rect 636 191 652 225
rect 586 157 652 191
rect 586 123 602 157
rect 636 123 652 157
rect 586 89 652 123
rect 586 55 602 89
rect 636 55 652 89
rect 586 17 652 55
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 2 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 3 nsew power bidirectional
rlabel comment s 0 0 0 0 4 decap_8
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 4 nsew power bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE SPACER
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5968434
string GDS_START 5964420
<< end >>
