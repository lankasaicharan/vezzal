magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 32 49 881 241
rect 0 0 960 49
<< scnmos >>
rect 111 47 141 215
rect 183 47 213 215
rect 291 47 321 215
rect 399 47 429 215
rect 514 47 544 215
rect 600 47 630 215
rect 686 47 716 215
rect 772 47 802 215
<< scpmoshvt >>
rect 111 367 141 619
rect 197 367 227 619
rect 313 367 343 619
rect 399 367 429 619
rect 514 367 544 619
rect 600 367 630 619
rect 686 367 716 619
rect 772 367 802 619
<< ndiff >>
rect 58 190 111 215
rect 58 156 66 190
rect 100 156 111 190
rect 58 122 111 156
rect 58 88 66 122
rect 100 88 111 122
rect 58 47 111 88
rect 141 47 183 215
rect 213 47 291 215
rect 321 47 399 215
rect 429 122 514 215
rect 429 88 452 122
rect 486 88 514 122
rect 429 47 514 88
rect 544 203 600 215
rect 544 169 555 203
rect 589 169 600 203
rect 544 101 600 169
rect 544 67 555 101
rect 589 67 600 101
rect 544 47 600 67
rect 630 177 686 215
rect 630 143 641 177
rect 675 143 686 177
rect 630 93 686 143
rect 630 59 641 93
rect 675 59 686 93
rect 630 47 686 59
rect 716 203 772 215
rect 716 169 727 203
rect 761 169 772 203
rect 716 101 772 169
rect 716 67 727 101
rect 761 67 772 101
rect 716 47 772 67
rect 802 163 855 215
rect 802 129 813 163
rect 847 129 855 163
rect 802 93 855 129
rect 802 59 813 93
rect 847 59 855 93
rect 802 47 855 59
<< pdiff >>
rect 58 607 111 619
rect 58 573 66 607
rect 100 573 111 607
rect 58 508 111 573
rect 58 474 66 508
rect 100 474 111 508
rect 58 418 111 474
rect 58 384 66 418
rect 100 384 111 418
rect 58 367 111 384
rect 141 599 197 619
rect 141 565 152 599
rect 186 565 197 599
rect 141 506 197 565
rect 141 472 152 506
rect 186 472 197 506
rect 141 413 197 472
rect 141 379 152 413
rect 186 379 197 413
rect 141 367 197 379
rect 227 607 313 619
rect 227 573 253 607
rect 287 573 313 607
rect 227 531 313 573
rect 227 497 253 531
rect 287 497 313 531
rect 227 455 313 497
rect 227 421 253 455
rect 287 421 313 455
rect 227 367 313 421
rect 343 599 399 619
rect 343 565 354 599
rect 388 565 399 599
rect 343 506 399 565
rect 343 472 354 506
rect 388 472 399 506
rect 343 413 399 472
rect 343 379 354 413
rect 388 379 399 413
rect 343 367 399 379
rect 429 607 514 619
rect 429 573 452 607
rect 486 573 514 607
rect 429 531 514 573
rect 429 497 452 531
rect 486 497 514 531
rect 429 455 514 497
rect 429 421 452 455
rect 486 421 514 455
rect 429 367 514 421
rect 544 599 600 619
rect 544 565 555 599
rect 589 565 600 599
rect 544 506 600 565
rect 544 472 555 506
rect 589 472 600 506
rect 544 413 600 472
rect 544 379 555 413
rect 589 379 600 413
rect 544 367 600 379
rect 630 611 686 619
rect 630 577 641 611
rect 675 577 686 611
rect 630 535 686 577
rect 630 501 641 535
rect 675 501 686 535
rect 630 457 686 501
rect 630 423 641 457
rect 675 423 686 457
rect 630 367 686 423
rect 716 599 772 619
rect 716 565 727 599
rect 761 565 772 599
rect 716 506 772 565
rect 716 472 727 506
rect 761 472 772 506
rect 716 413 772 472
rect 716 379 727 413
rect 761 379 772 413
rect 716 367 772 379
rect 802 607 855 619
rect 802 573 813 607
rect 847 573 855 607
rect 802 535 855 573
rect 802 501 813 535
rect 847 501 855 535
rect 802 457 855 501
rect 802 423 813 457
rect 847 423 855 457
rect 802 367 855 423
<< ndiffc >>
rect 66 156 100 190
rect 66 88 100 122
rect 452 88 486 122
rect 555 169 589 203
rect 555 67 589 101
rect 641 143 675 177
rect 641 59 675 93
rect 727 169 761 203
rect 727 67 761 101
rect 813 129 847 163
rect 813 59 847 93
<< pdiffc >>
rect 66 573 100 607
rect 66 474 100 508
rect 66 384 100 418
rect 152 565 186 599
rect 152 472 186 506
rect 152 379 186 413
rect 253 573 287 607
rect 253 497 287 531
rect 253 421 287 455
rect 354 565 388 599
rect 354 472 388 506
rect 354 379 388 413
rect 452 573 486 607
rect 452 497 486 531
rect 452 421 486 455
rect 555 565 589 599
rect 555 472 589 506
rect 555 379 589 413
rect 641 577 675 611
rect 641 501 675 535
rect 641 423 675 457
rect 727 565 761 599
rect 727 472 761 506
rect 727 379 761 413
rect 813 573 847 607
rect 813 501 847 535
rect 813 423 847 457
<< poly >>
rect 111 619 141 645
rect 197 619 227 645
rect 313 619 343 645
rect 399 619 429 645
rect 514 619 544 645
rect 600 619 630 645
rect 686 619 716 645
rect 772 619 802 645
rect 111 345 141 367
rect 81 308 141 345
rect 41 292 141 308
rect 197 303 227 367
rect 313 308 343 367
rect 399 308 429 367
rect 514 333 544 367
rect 600 333 630 367
rect 686 333 716 367
rect 772 333 802 367
rect 514 317 852 333
rect 41 258 57 292
rect 91 258 141 292
rect 41 237 141 258
rect 111 215 141 237
rect 183 287 249 303
rect 183 253 199 287
rect 233 253 249 287
rect 183 237 249 253
rect 291 292 357 308
rect 291 258 307 292
rect 341 258 357 292
rect 291 242 357 258
rect 399 292 465 308
rect 399 258 415 292
rect 449 258 465 292
rect 399 242 465 258
rect 514 283 530 317
rect 564 283 598 317
rect 632 283 666 317
rect 700 283 734 317
rect 768 283 802 317
rect 836 283 852 317
rect 514 267 852 283
rect 183 215 213 237
rect 291 215 321 242
rect 399 215 429 242
rect 514 215 544 267
rect 600 215 630 267
rect 686 215 716 267
rect 772 215 802 267
rect 111 21 141 47
rect 183 21 213 47
rect 291 21 321 47
rect 399 21 429 47
rect 514 21 544 47
rect 600 21 630 47
rect 686 21 716 47
rect 772 21 802 47
<< polycont >>
rect 57 258 91 292
rect 199 253 233 287
rect 307 258 341 292
rect 415 258 449 292
rect 530 283 564 317
rect 598 283 632 317
rect 666 283 700 317
rect 734 283 768 317
rect 802 283 836 317
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 50 607 116 649
rect 50 573 66 607
rect 100 573 116 607
rect 50 508 116 573
rect 50 474 66 508
rect 100 474 116 508
rect 50 418 116 474
rect 50 384 66 418
rect 100 384 116 418
rect 150 599 203 615
rect 150 565 152 599
rect 186 565 203 599
rect 150 506 203 565
rect 150 472 152 506
rect 186 472 203 506
rect 150 413 203 472
rect 237 607 303 649
rect 237 573 253 607
rect 287 573 303 607
rect 237 531 303 573
rect 237 497 253 531
rect 287 497 303 531
rect 237 455 303 497
rect 237 421 253 455
rect 287 421 303 455
rect 337 599 402 615
rect 337 565 354 599
rect 388 565 402 599
rect 337 506 402 565
rect 337 472 354 506
rect 388 472 402 506
rect 150 379 152 413
rect 186 385 203 413
rect 337 413 402 472
rect 436 607 502 649
rect 436 573 452 607
rect 486 573 502 607
rect 436 531 502 573
rect 436 497 452 531
rect 486 497 502 531
rect 436 455 502 497
rect 436 421 452 455
rect 486 421 502 455
rect 553 599 591 615
rect 553 565 555 599
rect 589 565 591 599
rect 553 506 591 565
rect 553 472 555 506
rect 589 472 591 506
rect 337 385 354 413
rect 186 379 354 385
rect 388 385 402 413
rect 553 413 591 472
rect 625 611 691 649
rect 625 577 641 611
rect 675 577 691 611
rect 625 535 691 577
rect 625 501 641 535
rect 675 501 691 535
rect 625 457 691 501
rect 625 423 641 457
rect 675 423 691 457
rect 725 599 763 615
rect 725 565 727 599
rect 761 565 763 599
rect 725 506 763 565
rect 725 472 727 506
rect 761 472 763 506
rect 388 379 519 385
rect 150 351 519 379
rect 553 379 555 413
rect 589 389 591 413
rect 725 413 763 472
rect 797 607 863 649
rect 797 573 813 607
rect 847 573 863 607
rect 797 535 863 573
rect 797 501 813 535
rect 847 501 863 535
rect 797 457 863 501
rect 797 423 813 457
rect 847 423 863 457
rect 725 389 727 413
rect 589 379 727 389
rect 761 389 763 413
rect 761 379 940 389
rect 553 355 940 379
rect 20 292 91 350
rect 485 317 519 351
rect 20 258 57 292
rect 20 240 91 258
rect 125 287 267 303
rect 125 253 199 287
rect 233 253 267 287
rect 125 240 267 253
rect 301 292 366 308
rect 301 258 307 292
rect 341 258 366 292
rect 301 240 366 258
rect 400 292 451 308
rect 400 258 415 292
rect 449 258 451 292
rect 400 240 451 258
rect 485 283 530 317
rect 564 283 598 317
rect 632 283 666 317
rect 700 283 734 317
rect 768 283 802 317
rect 836 283 852 317
rect 485 206 519 283
rect 886 247 940 355
rect 62 190 519 206
rect 62 156 66 190
rect 100 172 519 190
rect 555 213 940 247
rect 555 203 591 213
rect 62 122 100 156
rect 589 169 591 203
rect 725 203 773 213
rect 62 88 66 122
rect 62 72 100 88
rect 436 122 502 138
rect 436 88 452 122
rect 486 88 502 122
rect 436 17 502 88
rect 555 101 591 169
rect 589 67 591 101
rect 555 51 591 67
rect 625 177 691 179
rect 625 143 641 177
rect 675 143 691 177
rect 625 93 691 143
rect 625 59 641 93
rect 675 59 691 93
rect 625 17 691 59
rect 725 169 727 203
rect 761 169 773 203
rect 725 101 773 169
rect 725 67 727 101
rect 761 67 773 101
rect 725 51 773 67
rect 807 163 853 179
rect 807 129 813 163
rect 847 129 853 163
rect 807 93 853 129
rect 807 59 813 93
rect 847 59 853 93
rect 887 78 940 213
rect 807 17 853 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4_4
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 895 94 929 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6271550
string GDS_START 6262854
<< end >>
