magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 24 157 298 159
rect 24 49 863 157
rect 0 0 864 49
<< scnmos >>
rect 103 49 133 133
rect 189 49 219 133
rect 379 47 409 131
rect 465 47 495 131
rect 567 47 597 131
rect 653 47 683 131
rect 754 47 784 131
<< scpmoshvt >>
rect 80 530 110 614
rect 166 530 196 614
rect 389 439 419 523
rect 461 439 491 523
rect 563 485 593 569
rect 635 485 665 569
rect 750 485 780 569
<< ndiff >>
rect 50 103 103 133
rect 50 69 58 103
rect 92 69 103 103
rect 50 49 103 69
rect 133 95 189 133
rect 133 61 144 95
rect 178 61 189 95
rect 133 49 189 61
rect 219 121 272 133
rect 219 87 230 121
rect 264 87 272 121
rect 219 49 272 87
rect 326 93 379 131
rect 326 59 334 93
rect 368 59 379 93
rect 326 47 379 59
rect 409 123 465 131
rect 409 89 420 123
rect 454 89 465 123
rect 409 47 465 89
rect 495 89 567 131
rect 495 55 510 89
rect 544 55 567 89
rect 495 47 567 55
rect 597 119 653 131
rect 597 85 608 119
rect 642 85 653 119
rect 597 47 653 85
rect 683 93 754 131
rect 683 59 709 93
rect 743 59 754 93
rect 683 47 754 59
rect 784 119 837 131
rect 784 85 795 119
rect 829 85 837 119
rect 784 47 837 85
<< pdiff >>
rect 27 576 80 614
rect 27 542 35 576
rect 69 542 80 576
rect 27 530 80 542
rect 110 602 166 614
rect 110 568 121 602
rect 155 568 166 602
rect 110 530 166 568
rect 196 589 249 614
rect 196 555 207 589
rect 241 555 249 589
rect 196 530 249 555
rect 513 523 563 569
rect 336 485 389 523
rect 336 451 344 485
rect 378 451 389 485
rect 336 439 389 451
rect 419 439 461 523
rect 491 485 563 523
rect 593 485 635 569
rect 665 557 750 569
rect 665 523 693 557
rect 727 523 750 557
rect 665 485 750 523
rect 780 531 833 569
rect 780 497 791 531
rect 825 497 833 531
rect 780 485 833 497
rect 491 439 541 485
<< ndiffc >>
rect 58 69 92 103
rect 144 61 178 95
rect 230 87 264 121
rect 334 59 368 93
rect 420 89 454 123
rect 510 55 544 89
rect 608 85 642 119
rect 709 59 743 93
rect 795 85 829 119
<< pdiffc >>
rect 35 542 69 576
rect 121 568 155 602
rect 207 555 241 589
rect 344 451 378 485
rect 693 523 727 557
rect 791 497 825 531
<< poly >>
rect 80 614 110 640
rect 166 614 196 640
rect 281 605 347 621
rect 281 571 297 605
rect 331 571 347 605
rect 281 555 347 571
rect 563 569 593 595
rect 635 569 665 595
rect 750 569 780 595
rect 80 289 110 530
rect 166 467 196 530
rect 166 451 232 467
rect 166 417 182 451
rect 216 417 232 451
rect 166 401 232 417
rect 291 417 321 555
rect 389 523 419 549
rect 461 523 491 549
rect 389 417 419 439
rect 75 273 141 289
rect 75 239 91 273
rect 125 239 141 273
rect 75 205 141 239
rect 75 171 91 205
rect 125 171 141 205
rect 75 155 141 171
rect 103 133 133 155
rect 189 133 219 401
rect 291 387 419 417
rect 291 289 321 387
rect 461 339 491 439
rect 425 323 491 339
rect 425 289 441 323
rect 475 303 491 323
rect 563 313 593 485
rect 635 453 665 485
rect 635 437 701 453
rect 635 403 651 437
rect 685 403 701 437
rect 635 387 701 403
rect 475 289 495 303
rect 291 273 357 289
rect 425 273 495 289
rect 291 239 307 273
rect 341 239 357 273
rect 291 205 357 239
rect 291 171 307 205
rect 341 185 357 205
rect 341 171 409 185
rect 291 155 409 171
rect 379 131 409 155
rect 465 131 495 273
rect 537 297 603 313
rect 537 263 553 297
rect 587 263 603 297
rect 537 229 603 263
rect 537 195 553 229
rect 587 195 603 229
rect 537 179 603 195
rect 567 131 597 179
rect 653 131 683 387
rect 750 339 780 485
rect 725 323 791 339
rect 725 289 741 323
rect 775 289 791 323
rect 725 255 791 289
rect 725 221 741 255
rect 775 221 791 255
rect 725 205 791 221
rect 754 131 784 205
rect 103 23 133 49
rect 189 23 219 49
rect 379 21 409 47
rect 465 21 495 47
rect 567 21 597 47
rect 653 21 683 47
rect 754 21 784 47
<< polycont >>
rect 297 571 331 605
rect 182 417 216 451
rect 91 239 125 273
rect 91 171 125 205
rect 441 289 475 323
rect 651 403 685 437
rect 307 239 341 273
rect 307 171 341 205
rect 553 263 587 297
rect 553 195 587 229
rect 741 289 775 323
rect 741 221 775 255
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 117 602 155 649
rect 21 576 73 592
rect 21 542 35 576
rect 69 542 73 576
rect 117 568 121 602
rect 117 552 155 568
rect 203 589 297 605
rect 203 555 207 589
rect 241 571 297 589
rect 331 571 347 605
rect 241 555 347 571
rect 21 359 73 542
rect 203 539 347 555
rect 117 451 232 505
rect 117 417 182 451
rect 216 417 232 451
rect 340 485 571 501
rect 340 451 344 485
rect 378 451 571 485
rect 340 435 571 451
rect 117 401 232 417
rect 537 367 571 435
rect 607 464 641 582
rect 677 557 743 649
rect 677 523 693 557
rect 727 523 743 557
rect 677 519 743 523
rect 787 531 845 582
rect 787 497 791 531
rect 825 497 845 531
rect 787 464 845 497
rect 607 437 701 464
rect 607 403 651 437
rect 685 403 701 437
rect 21 325 475 359
rect 537 333 775 367
rect 21 119 55 325
rect 441 323 475 325
rect 91 273 161 289
rect 125 239 161 273
rect 91 205 161 239
rect 125 171 161 205
rect 307 273 341 289
rect 441 273 475 289
rect 307 205 341 239
rect 91 155 161 171
rect 226 171 307 181
rect 511 263 553 297
rect 587 263 603 297
rect 511 229 603 263
rect 511 195 553 229
rect 587 195 603 229
rect 226 147 341 171
rect 639 159 673 333
rect 741 323 775 333
rect 741 255 775 289
rect 741 205 775 221
rect 226 121 268 147
rect 21 103 96 119
rect 21 69 58 103
rect 92 69 96 103
rect 21 53 96 69
rect 140 95 182 111
rect 140 61 144 95
rect 178 61 182 95
rect 226 87 230 121
rect 264 87 268 121
rect 416 125 673 159
rect 811 135 845 464
rect 416 123 458 125
rect 226 71 268 87
rect 330 93 372 109
rect 140 17 182 61
rect 330 59 334 93
rect 368 59 372 93
rect 416 89 420 123
rect 454 89 458 123
rect 604 119 673 125
rect 416 73 458 89
rect 330 17 372 59
rect 494 55 510 89
rect 544 55 560 89
rect 604 85 608 119
rect 642 85 673 119
rect 791 119 845 135
rect 604 69 673 85
rect 709 93 747 109
rect 494 17 560 55
rect 743 59 747 93
rect 791 85 795 119
rect 829 85 845 119
rect 791 69 845 85
rect 709 17 747 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or4bb_m
flabel comment s 305 406 305 406 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6804974
string GDS_START 6796930
<< end >>
