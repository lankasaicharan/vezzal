magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 15 49 638 162
rect 0 0 672 49
<< scnmos >>
rect 94 52 124 136
rect 241 52 271 136
rect 313 52 343 136
rect 421 52 451 136
rect 529 52 559 136
<< scpmoshvt >>
rect 88 392 118 476
rect 242 392 272 476
rect 328 392 358 476
rect 414 392 444 476
rect 500 392 530 476
<< ndiff >>
rect 41 124 94 136
rect 41 90 49 124
rect 83 90 94 124
rect 41 52 94 90
rect 124 98 241 136
rect 124 64 135 98
rect 169 64 241 98
rect 124 52 241 64
rect 271 52 313 136
rect 343 52 421 136
rect 451 52 529 136
rect 559 124 612 136
rect 559 90 570 124
rect 604 90 612 124
rect 559 52 612 90
<< pdiff >>
rect 35 438 88 476
rect 35 404 43 438
rect 77 404 88 438
rect 35 392 88 404
rect 118 464 242 476
rect 118 430 197 464
rect 231 430 242 464
rect 118 392 242 430
rect 272 438 328 476
rect 272 404 283 438
rect 317 404 328 438
rect 272 392 328 404
rect 358 464 414 476
rect 358 430 369 464
rect 403 430 414 464
rect 358 392 414 430
rect 444 438 500 476
rect 444 404 455 438
rect 489 404 500 438
rect 444 392 500 404
rect 530 464 583 476
rect 530 430 541 464
rect 575 430 583 464
rect 530 392 583 430
<< ndiffc >>
rect 49 90 83 124
rect 135 64 169 98
rect 570 90 604 124
<< pdiffc >>
rect 43 404 77 438
rect 197 430 231 464
rect 283 404 317 438
rect 369 430 403 464
rect 455 404 489 438
rect 541 430 575 464
<< poly >>
rect 111 594 530 610
rect 111 560 127 594
rect 161 580 530 594
rect 161 560 177 580
rect 111 544 177 560
rect 88 476 118 502
rect 242 476 272 502
rect 328 476 358 502
rect 414 476 444 502
rect 500 476 530 580
rect 88 302 118 392
rect 242 370 272 392
rect 241 340 272 370
rect 88 286 163 302
rect 241 292 271 340
rect 328 292 358 392
rect 414 370 444 392
rect 500 370 530 392
rect 414 340 451 370
rect 500 340 559 370
rect 421 292 451 340
rect 88 272 113 286
rect 94 252 113 272
rect 147 252 163 286
rect 94 218 163 252
rect 94 184 113 218
rect 147 184 163 218
rect 94 168 163 184
rect 205 276 271 292
rect 205 242 221 276
rect 255 242 271 276
rect 205 208 271 242
rect 205 174 221 208
rect 255 174 271 208
rect 94 136 124 168
rect 205 158 271 174
rect 241 136 271 158
rect 313 276 379 292
rect 313 242 329 276
rect 363 242 379 276
rect 313 208 379 242
rect 313 174 329 208
rect 363 174 379 208
rect 313 158 379 174
rect 421 276 487 292
rect 421 242 437 276
rect 471 242 487 276
rect 421 208 487 242
rect 421 174 437 208
rect 471 174 487 208
rect 421 158 487 174
rect 313 136 343 158
rect 421 136 451 158
rect 529 136 559 340
rect 94 26 124 52
rect 241 26 271 52
rect 313 26 343 52
rect 421 26 451 52
rect 529 26 559 52
<< polycont >>
rect 127 560 161 594
rect 113 252 147 286
rect 113 184 147 218
rect 221 242 255 276
rect 221 174 255 208
rect 329 242 363 276
rect 329 174 363 208
rect 437 242 471 276
rect 437 174 471 208
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 33 594 161 610
rect 33 560 127 594
rect 33 544 161 560
rect 33 438 77 544
rect 33 404 43 438
rect 33 128 77 404
rect 113 286 161 498
rect 197 464 231 649
rect 369 464 403 649
rect 197 414 231 430
rect 267 438 333 442
rect 267 404 283 438
rect 317 404 333 438
rect 541 464 579 649
rect 369 414 403 430
rect 439 438 505 442
rect 267 350 333 404
rect 439 404 455 438
rect 489 404 505 438
rect 575 430 579 464
rect 541 414 579 430
rect 439 350 505 404
rect 223 316 641 350
rect 147 252 161 286
rect 113 218 161 252
rect 147 184 161 218
rect 113 168 161 184
rect 205 242 221 276
rect 255 242 271 276
rect 205 208 271 242
rect 205 174 221 208
rect 255 174 271 208
rect 33 124 99 128
rect 33 90 49 124
rect 83 90 99 124
rect 33 86 99 90
rect 135 98 169 114
rect 205 94 271 174
rect 313 242 329 276
rect 363 242 379 276
rect 313 208 379 242
rect 313 174 329 208
rect 363 174 379 208
rect 313 94 379 174
rect 415 242 437 276
rect 471 242 487 276
rect 415 208 487 242
rect 415 174 437 208
rect 471 174 487 208
rect 415 94 487 174
rect 607 128 641 316
rect 554 124 641 128
rect 554 90 570 124
rect 604 90 641 124
rect 554 86 641 90
rect 135 17 169 64
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4b_m
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 776028
string GDS_START 768714
<< end >>
