magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 106 159 690 243
rect 1 49 690 159
rect 0 0 768 49
<< scnmos >>
rect 80 49 110 133
rect 198 49 228 217
rect 284 49 314 217
rect 413 133 443 217
rect 521 133 551 217
<< scpmoshvt >>
rect 93 367 123 451
rect 191 367 221 619
rect 277 367 307 619
rect 449 367 479 451
rect 521 367 551 451
<< ndiff >>
rect 132 133 198 217
rect 27 108 80 133
rect 27 74 35 108
rect 69 74 80 108
rect 27 49 80 74
rect 110 69 198 133
rect 110 49 137 69
rect 125 35 137 49
rect 171 49 198 69
rect 228 209 284 217
rect 228 175 239 209
rect 273 175 284 209
rect 228 49 284 175
rect 314 133 413 217
rect 443 209 521 217
rect 443 175 454 209
rect 488 175 521 209
rect 443 133 521 175
rect 551 179 664 217
rect 551 145 622 179
rect 656 145 664 179
rect 551 133 664 145
rect 314 69 387 133
rect 314 49 341 69
rect 171 35 183 49
rect 125 27 183 35
rect 329 35 341 49
rect 375 35 387 69
rect 329 27 387 35
<< pdiff >>
rect 138 607 191 619
rect 138 573 146 607
rect 180 573 191 607
rect 138 539 191 573
rect 138 505 146 539
rect 180 505 191 539
rect 138 461 191 505
rect 138 451 146 461
rect 36 426 93 451
rect 36 392 48 426
rect 82 392 93 426
rect 36 367 93 392
rect 123 427 146 451
rect 180 427 191 461
rect 123 367 191 427
rect 221 599 277 619
rect 221 565 232 599
rect 266 565 277 599
rect 221 505 277 565
rect 221 471 232 505
rect 266 471 277 505
rect 221 409 277 471
rect 221 375 232 409
rect 266 375 277 409
rect 221 367 277 375
rect 307 607 360 619
rect 307 573 318 607
rect 352 573 360 607
rect 307 504 360 573
rect 307 470 318 504
rect 352 470 360 504
rect 307 451 360 470
rect 307 367 449 451
rect 479 367 521 451
rect 551 436 604 451
rect 551 402 562 436
rect 596 402 604 436
rect 551 367 604 402
<< ndiffc >>
rect 35 74 69 108
rect 137 35 171 69
rect 239 175 273 209
rect 454 175 488 209
rect 622 145 656 179
rect 341 35 375 69
<< pdiffc >>
rect 146 573 180 607
rect 146 505 180 539
rect 48 392 82 426
rect 146 427 180 461
rect 232 565 266 599
rect 232 471 266 505
rect 232 375 266 409
rect 318 573 352 607
rect 318 470 352 504
rect 562 402 596 436
<< poly >>
rect 191 619 221 645
rect 277 619 307 645
rect 93 451 123 477
rect 449 451 479 477
rect 521 451 551 477
rect 93 309 123 367
rect 44 293 123 309
rect 44 259 60 293
rect 94 279 123 293
rect 191 305 221 367
rect 277 305 307 367
rect 449 335 479 367
rect 413 319 479 335
rect 191 289 366 305
rect 94 259 110 279
rect 44 225 110 259
rect 191 255 316 289
rect 350 255 366 289
rect 191 254 366 255
rect 44 191 60 225
rect 94 191 110 225
rect 198 239 366 254
rect 413 285 429 319
rect 463 285 479 319
rect 413 269 479 285
rect 521 305 551 367
rect 521 289 727 305
rect 198 217 228 239
rect 284 217 314 239
rect 413 217 443 269
rect 521 255 589 289
rect 623 255 677 289
rect 711 255 727 289
rect 521 239 727 255
rect 521 217 551 239
rect 44 175 110 191
rect 80 133 110 175
rect 80 23 110 49
rect 413 107 443 133
rect 521 107 551 133
rect 198 23 228 49
rect 284 23 314 49
<< polycont >>
rect 60 259 94 293
rect 316 255 350 289
rect 60 191 94 225
rect 429 285 463 319
rect 589 255 623 289
rect 677 255 711 289
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 137 607 182 649
rect 137 573 146 607
rect 180 573 182 607
rect 137 539 182 573
rect 137 505 146 539
rect 180 505 182 539
rect 137 461 182 505
rect 32 426 98 442
rect 32 392 48 426
rect 82 392 98 426
rect 137 427 146 461
rect 180 427 182 461
rect 137 411 182 427
rect 216 599 282 615
rect 216 565 232 599
rect 266 565 282 599
rect 216 505 282 565
rect 216 471 232 505
rect 266 471 282 505
rect 32 377 98 392
rect 216 409 282 471
rect 316 607 368 649
rect 316 573 318 607
rect 352 573 368 607
rect 316 504 368 573
rect 316 470 318 504
rect 352 470 368 504
rect 316 454 368 470
rect 546 436 612 452
rect 546 420 562 436
rect 32 343 164 377
rect 17 293 94 309
rect 17 259 60 293
rect 17 225 94 259
rect 17 191 60 225
rect 17 175 94 191
rect 130 139 164 343
rect 216 375 232 409
rect 266 375 282 409
rect 216 209 282 375
rect 316 402 562 420
rect 596 402 612 436
rect 316 386 612 402
rect 316 289 366 386
rect 350 255 366 289
rect 400 319 555 352
rect 400 285 429 319
rect 463 285 555 319
rect 400 283 555 285
rect 589 289 727 305
rect 316 231 366 255
rect 623 255 677 289
rect 711 255 727 289
rect 589 249 727 255
rect 323 225 366 231
rect 323 209 504 225
rect 216 175 239 209
rect 273 175 289 209
rect 216 173 289 175
rect 323 175 454 209
rect 488 175 504 209
rect 323 173 504 175
rect 538 215 727 249
rect 538 139 572 215
rect 19 108 572 139
rect 19 74 35 108
rect 69 105 572 108
rect 606 179 672 181
rect 606 145 622 179
rect 656 145 672 179
rect 69 74 84 105
rect 19 58 84 74
rect 118 69 187 71
rect 118 35 137 69
rect 171 35 187 69
rect 118 17 187 35
rect 325 69 391 71
rect 325 35 341 69
rect 375 35 391 69
rect 325 17 391 35
rect 606 17 672 145
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or2b_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2265944
string GDS_START 2259690
<< end >>
