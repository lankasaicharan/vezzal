magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 332 614 704
<< pwell >>
rect 4 49 575 184
rect 0 0 576 49
<< scpmos >>
rect 83 368 119 592
rect 173 368 209 592
rect 263 368 299 592
rect 353 368 389 592
rect 453 368 489 592
<< nmoslvt >>
rect 87 74 117 158
rect 173 74 203 158
rect 259 74 289 158
rect 353 74 383 158
rect 459 74 489 158
<< ndiff >>
rect 30 133 87 158
rect 30 99 42 133
rect 76 99 87 133
rect 30 74 87 99
rect 117 133 173 158
rect 117 99 128 133
rect 162 99 173 133
rect 117 74 173 99
rect 203 133 259 158
rect 203 99 214 133
rect 248 99 259 133
rect 203 74 259 99
rect 289 133 353 158
rect 289 99 300 133
rect 334 99 353 133
rect 289 74 353 99
rect 383 133 459 158
rect 383 99 400 133
rect 434 99 459 133
rect 383 74 459 99
rect 489 146 549 158
rect 489 112 501 146
rect 535 112 549 146
rect 489 74 549 112
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 507 173 546
rect 119 473 129 507
rect 163 473 173 507
rect 119 434 173 473
rect 119 400 129 434
rect 163 400 173 434
rect 119 368 173 400
rect 209 580 263 592
rect 209 546 219 580
rect 253 546 263 580
rect 209 502 263 546
rect 209 468 219 502
rect 253 468 263 502
rect 209 368 263 468
rect 299 580 353 592
rect 299 546 309 580
rect 343 546 353 580
rect 299 507 353 546
rect 299 473 309 507
rect 343 473 353 507
rect 299 434 353 473
rect 299 400 309 434
rect 343 400 353 434
rect 299 368 353 400
rect 389 580 453 592
rect 389 546 399 580
rect 433 546 453 580
rect 389 507 453 546
rect 389 473 399 507
rect 433 473 453 507
rect 389 434 453 473
rect 389 400 399 434
rect 433 400 453 434
rect 389 368 453 400
rect 489 580 545 592
rect 489 546 499 580
rect 533 546 545 580
rect 489 497 545 546
rect 489 463 499 497
rect 533 463 545 497
rect 489 414 545 463
rect 489 380 499 414
rect 533 380 545 414
rect 489 368 545 380
<< ndiffc >>
rect 42 99 76 133
rect 128 99 162 133
rect 214 99 248 133
rect 300 99 334 133
rect 400 99 434 133
rect 501 112 535 146
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 473 163 507
rect 129 400 163 434
rect 219 546 253 580
rect 219 468 253 502
rect 309 546 343 580
rect 309 473 343 507
rect 309 400 343 434
rect 399 546 433 580
rect 399 473 433 507
rect 399 400 433 434
rect 499 546 533 580
rect 499 463 533 497
rect 499 380 533 414
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 263 592 299 618
rect 353 592 389 618
rect 453 592 489 618
rect 83 336 119 368
rect 173 336 209 368
rect 263 336 299 368
rect 353 336 389 368
rect 83 320 389 336
rect 83 286 191 320
rect 225 286 259 320
rect 293 286 327 320
rect 361 286 389 320
rect 83 270 389 286
rect 453 282 489 368
rect 87 158 117 270
rect 173 158 203 270
rect 259 158 289 270
rect 353 158 383 270
rect 431 266 497 282
rect 431 232 447 266
rect 481 232 497 266
rect 431 216 497 232
rect 459 158 489 216
rect 87 48 117 74
rect 173 48 203 74
rect 259 48 289 74
rect 353 48 383 74
rect 459 48 489 74
<< polycont >>
rect 191 286 225 320
rect 259 286 293 320
rect 327 286 361 320
rect 447 232 481 266
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 107 580 163 596
rect 107 546 129 580
rect 107 507 163 546
rect 107 473 129 507
rect 107 434 163 473
rect 203 580 253 649
rect 203 546 219 580
rect 203 502 253 546
rect 203 468 219 502
rect 203 452 253 468
rect 293 580 359 596
rect 293 546 309 580
rect 343 546 359 580
rect 293 507 359 546
rect 293 473 309 507
rect 343 473 359 507
rect 107 400 129 434
rect 293 434 359 473
rect 293 418 309 434
rect 163 400 309 418
rect 343 400 359 434
rect 107 384 359 400
rect 399 580 449 649
rect 433 546 449 580
rect 399 507 449 546
rect 433 473 449 507
rect 399 434 449 473
rect 433 400 449 434
rect 399 384 449 400
rect 483 580 559 596
rect 483 546 499 580
rect 533 546 559 580
rect 483 497 559 546
rect 483 463 499 497
rect 533 463 559 497
rect 483 414 559 463
rect 107 230 141 384
rect 483 380 499 414
rect 533 380 559 414
rect 483 350 559 380
rect 175 320 559 350
rect 175 286 191 320
rect 225 286 259 320
rect 293 286 327 320
rect 361 316 559 320
rect 361 286 377 316
rect 175 270 377 286
rect 411 266 491 282
rect 411 232 447 266
rect 481 232 491 266
rect 107 196 350 230
rect 411 216 491 232
rect 26 133 76 162
rect 26 99 42 133
rect 26 17 76 99
rect 112 133 178 196
rect 112 99 128 133
rect 162 99 178 133
rect 112 70 178 99
rect 214 133 248 162
rect 214 17 248 99
rect 284 133 350 196
rect 525 162 559 316
rect 284 99 300 133
rect 334 99 350 133
rect 284 70 350 99
rect 384 133 450 162
rect 384 99 400 133
rect 434 99 450 133
rect 384 17 450 99
rect 484 146 559 162
rect 484 112 501 146
rect 535 112 559 146
rect 484 96 559 112
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkbuf_4
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 786880
string GDS_START 781544
<< end >>
