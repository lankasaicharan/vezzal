magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 337 710 704
rect -38 331 240 337
rect 494 331 710 337
<< pwell >>
rect 302 263 491 295
rect 25 157 491 263
rect 25 49 671 157
rect 0 0 672 49
<< scnmos >>
rect 108 153 138 237
rect 186 153 216 237
rect 283 153 313 237
rect 378 185 408 269
rect 480 47 510 131
rect 558 47 588 131
<< scpmoshvt >>
rect 125 419 175 619
rect 272 419 322 619
rect 378 419 428 619
rect 509 419 559 619
<< ndiff >>
rect 328 237 378 269
rect 51 212 108 237
rect 51 178 63 212
rect 97 178 108 212
rect 51 153 108 178
rect 138 153 186 237
rect 216 199 283 237
rect 216 165 227 199
rect 261 165 283 199
rect 216 153 283 165
rect 313 185 378 237
rect 408 244 465 269
rect 408 210 419 244
rect 453 210 465 244
rect 408 185 465 210
rect 313 153 363 185
rect 423 106 480 131
rect 423 72 435 106
rect 469 72 480 106
rect 423 47 480 72
rect 510 47 558 131
rect 588 106 645 131
rect 588 72 599 106
rect 633 72 645 106
rect 588 47 645 72
<< pdiff >>
rect 68 597 125 619
rect 68 563 80 597
rect 114 563 125 597
rect 68 465 125 563
rect 68 431 80 465
rect 114 431 125 465
rect 68 419 125 431
rect 175 596 272 619
rect 175 562 186 596
rect 220 562 272 596
rect 175 419 272 562
rect 322 597 378 619
rect 322 563 333 597
rect 367 563 378 597
rect 322 516 378 563
rect 322 482 333 516
rect 367 482 378 516
rect 322 419 378 482
rect 428 607 509 619
rect 428 573 439 607
rect 473 573 509 607
rect 428 473 509 573
rect 428 439 439 473
rect 473 439 509 473
rect 428 419 509 439
rect 559 597 616 619
rect 559 563 570 597
rect 604 563 616 597
rect 559 465 616 563
rect 559 431 570 465
rect 604 431 616 465
rect 559 419 616 431
<< ndiffc >>
rect 63 178 97 212
rect 227 165 261 199
rect 419 210 453 244
rect 435 72 469 106
rect 599 72 633 106
<< pdiffc >>
rect 80 563 114 597
rect 80 431 114 465
rect 186 562 220 596
rect 333 563 367 597
rect 333 482 367 516
rect 439 573 473 607
rect 439 439 473 473
rect 570 563 604 597
rect 570 431 604 465
<< poly >>
rect 125 619 175 645
rect 272 619 322 645
rect 378 619 428 645
rect 509 619 559 645
rect 125 325 175 419
rect 272 387 322 419
rect 378 387 428 419
rect 264 371 330 387
rect 264 337 280 371
rect 314 337 330 371
rect 108 309 216 325
rect 264 321 330 337
rect 378 371 461 387
rect 378 337 411 371
rect 445 337 461 371
rect 378 321 461 337
rect 108 275 166 309
rect 200 275 216 309
rect 108 259 216 275
rect 108 237 138 259
rect 186 237 216 259
rect 283 237 313 321
rect 378 269 408 321
rect 509 273 559 419
rect 480 257 588 273
rect 480 223 521 257
rect 555 223 588 257
rect 480 207 588 223
rect 378 159 408 185
rect 108 127 138 153
rect 186 127 216 153
rect 283 127 313 153
rect 480 131 510 207
rect 558 131 588 207
rect 480 21 510 47
rect 558 21 588 47
<< polycont >>
rect 280 337 314 371
rect 411 337 445 371
rect 166 275 200 309
rect 521 223 555 257
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 25 597 114 613
rect 25 563 80 597
rect 25 465 114 563
rect 170 596 236 649
rect 170 562 186 596
rect 220 562 236 596
rect 170 536 236 562
rect 317 597 383 613
rect 317 563 333 597
rect 367 563 383 597
rect 317 516 383 563
rect 317 500 333 516
rect 25 431 80 465
rect 25 212 114 431
rect 150 482 333 500
rect 367 482 383 516
rect 150 466 383 482
rect 423 607 489 649
rect 423 573 439 607
rect 473 573 489 607
rect 423 473 489 573
rect 150 309 216 466
rect 423 439 439 473
rect 473 439 489 473
rect 264 371 359 430
rect 423 423 489 439
rect 554 597 620 613
rect 554 563 570 597
rect 604 563 620 597
rect 554 465 620 563
rect 554 431 570 465
rect 604 431 620 465
rect 554 387 620 431
rect 264 337 280 371
rect 314 337 359 371
rect 264 321 359 337
rect 395 371 649 387
rect 395 337 411 371
rect 445 337 649 371
rect 395 321 649 337
rect 150 275 166 309
rect 200 285 216 309
rect 200 275 469 285
rect 150 251 469 275
rect 403 244 469 251
rect 25 178 63 212
rect 97 178 114 212
rect 25 88 114 178
rect 211 199 277 215
rect 211 165 227 199
rect 261 165 277 199
rect 403 210 419 244
rect 453 210 469 244
rect 403 181 469 210
rect 505 257 571 282
rect 505 223 521 257
rect 555 223 571 257
rect 505 207 571 223
rect 211 17 277 165
rect 615 135 649 321
rect 419 106 485 135
rect 419 72 435 106
rect 469 72 485 106
rect 419 17 485 72
rect 583 106 649 135
rect 583 72 599 106
rect 633 72 649 106
rect 583 59 649 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and2b_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5156618
string GDS_START 5150636
<< end >>
