magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3138 1852
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 1 21 1830 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 287 47 317 177
rect 391 47 421 177
rect 485 47 515 177
rect 579 47 609 177
rect 673 47 703 177
rect 767 47 797 177
rect 861 47 891 177
rect 958 47 988 177
rect 1050 47 1080 177
rect 1144 47 1174 177
rect 1238 47 1268 177
rect 1332 47 1362 177
rect 1426 47 1456 177
rect 1520 47 1550 177
rect 1614 47 1644 177
rect 1718 47 1748 177
<< scpmoshvt >>
rect 81 297 117 497
rect 186 309 222 497
rect 280 309 316 497
rect 374 309 410 497
rect 468 309 504 497
rect 562 309 598 497
rect 656 309 692 497
rect 750 309 786 497
rect 844 309 880 497
rect 1052 297 1088 497
rect 1146 297 1182 497
rect 1240 297 1276 497
rect 1334 297 1370 497
rect 1428 297 1464 497
rect 1522 297 1558 497
rect 1616 297 1652 497
rect 1710 297 1746 497
<< ndiff >>
rect 27 129 89 177
rect 27 95 35 129
rect 69 95 89 129
rect 27 47 89 95
rect 119 93 171 177
rect 119 59 129 93
rect 163 59 171 93
rect 119 47 171 59
rect 235 129 287 177
rect 235 95 243 129
rect 277 95 287 129
rect 235 47 287 95
rect 317 89 391 177
rect 317 55 337 89
rect 371 55 391 89
rect 317 47 391 55
rect 421 129 485 177
rect 421 95 431 129
rect 465 95 485 129
rect 421 47 485 95
rect 515 89 579 177
rect 515 55 525 89
rect 559 55 579 89
rect 515 47 579 55
rect 609 129 673 177
rect 609 95 619 129
rect 653 95 673 129
rect 609 47 673 95
rect 703 89 767 177
rect 703 55 713 89
rect 747 55 767 89
rect 703 47 767 55
rect 797 129 861 177
rect 797 95 807 129
rect 841 95 861 129
rect 797 47 861 95
rect 891 89 958 177
rect 891 55 901 89
rect 935 55 958 89
rect 891 47 958 55
rect 988 129 1050 177
rect 988 95 1001 129
rect 1035 95 1050 129
rect 988 47 1050 95
rect 1080 165 1144 177
rect 1080 131 1100 165
rect 1134 131 1144 165
rect 1080 47 1144 131
rect 1174 90 1238 177
rect 1174 56 1194 90
rect 1228 56 1238 90
rect 1174 47 1238 56
rect 1268 165 1332 177
rect 1268 131 1288 165
rect 1322 131 1332 165
rect 1268 47 1332 131
rect 1362 90 1426 177
rect 1362 56 1382 90
rect 1416 56 1426 90
rect 1362 47 1426 56
rect 1456 165 1520 177
rect 1456 131 1476 165
rect 1510 131 1520 165
rect 1456 47 1520 131
rect 1550 90 1614 177
rect 1550 56 1570 90
rect 1604 56 1614 90
rect 1550 47 1614 56
rect 1644 165 1718 177
rect 1644 131 1664 165
rect 1698 131 1718 165
rect 1644 47 1718 131
rect 1748 90 1804 177
rect 1748 56 1758 90
rect 1792 56 1804 90
rect 1748 47 1804 56
<< pdiff >>
rect 27 448 81 497
rect 27 414 35 448
rect 69 414 81 448
rect 27 380 81 414
rect 27 346 35 380
rect 69 346 81 380
rect 27 297 81 346
rect 117 489 186 497
rect 117 455 129 489
rect 163 455 186 489
rect 117 421 186 455
rect 117 387 129 421
rect 163 387 186 421
rect 117 309 186 387
rect 222 448 280 497
rect 222 414 234 448
rect 268 414 280 448
rect 222 380 280 414
rect 222 346 234 380
rect 268 346 280 380
rect 222 309 280 346
rect 316 489 374 497
rect 316 455 328 489
rect 362 455 374 489
rect 316 421 374 455
rect 316 387 328 421
rect 362 387 374 421
rect 316 309 374 387
rect 410 448 468 497
rect 410 414 422 448
rect 456 414 468 448
rect 410 380 468 414
rect 410 346 422 380
rect 456 346 468 380
rect 410 309 468 346
rect 504 489 562 497
rect 504 455 516 489
rect 550 455 562 489
rect 504 421 562 455
rect 504 387 516 421
rect 550 387 562 421
rect 504 309 562 387
rect 598 448 656 497
rect 598 414 610 448
rect 644 414 656 448
rect 598 380 656 414
rect 598 346 610 380
rect 644 346 656 380
rect 598 309 656 346
rect 692 489 750 497
rect 692 455 704 489
rect 738 455 750 489
rect 692 421 750 455
rect 692 387 704 421
rect 738 387 750 421
rect 692 309 750 387
rect 786 448 844 497
rect 786 414 798 448
rect 832 414 844 448
rect 786 380 844 414
rect 786 346 798 380
rect 832 346 844 380
rect 786 309 844 346
rect 880 485 934 497
rect 880 451 892 485
rect 926 451 934 485
rect 880 417 934 451
rect 880 383 892 417
rect 926 383 934 417
rect 880 309 934 383
rect 998 448 1052 497
rect 998 414 1006 448
rect 1040 414 1052 448
rect 998 380 1052 414
rect 998 346 1006 380
rect 1040 346 1052 380
rect 117 297 169 309
rect 998 297 1052 346
rect 1088 425 1146 497
rect 1088 391 1100 425
rect 1134 391 1146 425
rect 1088 357 1146 391
rect 1088 323 1100 357
rect 1134 323 1146 357
rect 1088 297 1146 323
rect 1182 477 1240 497
rect 1182 443 1194 477
rect 1228 443 1240 477
rect 1182 409 1240 443
rect 1182 375 1194 409
rect 1228 375 1240 409
rect 1182 297 1240 375
rect 1276 425 1334 497
rect 1276 391 1288 425
rect 1322 391 1334 425
rect 1276 357 1334 391
rect 1276 323 1288 357
rect 1322 323 1334 357
rect 1276 297 1334 323
rect 1370 477 1428 497
rect 1370 443 1382 477
rect 1416 443 1428 477
rect 1370 409 1428 443
rect 1370 375 1382 409
rect 1416 375 1428 409
rect 1370 297 1428 375
rect 1464 425 1522 497
rect 1464 391 1476 425
rect 1510 391 1522 425
rect 1464 357 1522 391
rect 1464 323 1476 357
rect 1510 323 1522 357
rect 1464 297 1522 323
rect 1558 477 1616 497
rect 1558 443 1570 477
rect 1604 443 1616 477
rect 1558 409 1616 443
rect 1558 375 1570 409
rect 1604 375 1616 409
rect 1558 297 1616 375
rect 1652 425 1710 497
rect 1652 391 1664 425
rect 1698 391 1710 425
rect 1652 357 1710 391
rect 1652 323 1664 357
rect 1698 323 1710 357
rect 1652 297 1710 323
rect 1746 477 1800 497
rect 1746 443 1758 477
rect 1792 443 1800 477
rect 1746 409 1800 443
rect 1746 375 1758 409
rect 1792 375 1800 409
rect 1746 297 1800 375
<< ndiffc >>
rect 35 95 69 129
rect 129 59 163 93
rect 243 95 277 129
rect 337 55 371 89
rect 431 95 465 129
rect 525 55 559 89
rect 619 95 653 129
rect 713 55 747 89
rect 807 95 841 129
rect 901 55 935 89
rect 1001 95 1035 129
rect 1100 131 1134 165
rect 1194 56 1228 90
rect 1288 131 1322 165
rect 1382 56 1416 90
rect 1476 131 1510 165
rect 1570 56 1604 90
rect 1664 131 1698 165
rect 1758 56 1792 90
<< pdiffc >>
rect 35 414 69 448
rect 35 346 69 380
rect 129 455 163 489
rect 129 387 163 421
rect 234 414 268 448
rect 234 346 268 380
rect 328 455 362 489
rect 328 387 362 421
rect 422 414 456 448
rect 422 346 456 380
rect 516 455 550 489
rect 516 387 550 421
rect 610 414 644 448
rect 610 346 644 380
rect 704 455 738 489
rect 704 387 738 421
rect 798 414 832 448
rect 798 346 832 380
rect 892 451 926 485
rect 892 383 926 417
rect 1006 414 1040 448
rect 1006 346 1040 380
rect 1100 391 1134 425
rect 1100 323 1134 357
rect 1194 443 1228 477
rect 1194 375 1228 409
rect 1288 391 1322 425
rect 1288 323 1322 357
rect 1382 443 1416 477
rect 1382 375 1416 409
rect 1476 391 1510 425
rect 1476 323 1510 357
rect 1570 443 1604 477
rect 1570 375 1604 409
rect 1664 391 1698 425
rect 1664 323 1698 357
rect 1758 443 1792 477
rect 1758 375 1792 409
<< poly >>
rect 81 497 117 523
rect 186 497 222 523
rect 280 497 316 523
rect 374 497 410 523
rect 468 497 504 523
rect 562 497 598 523
rect 656 497 692 523
rect 750 497 786 523
rect 844 497 880 523
rect 1052 497 1088 523
rect 1146 497 1182 523
rect 1240 497 1276 523
rect 1334 497 1370 523
rect 1428 497 1464 523
rect 1522 497 1558 523
rect 1616 497 1652 523
rect 1710 497 1746 523
rect 81 282 117 297
rect 186 294 222 309
rect 280 294 316 309
rect 374 294 410 309
rect 468 294 504 309
rect 562 294 598 309
rect 656 294 692 309
rect 750 294 786 309
rect 844 294 880 309
rect 79 265 119 282
rect 184 265 882 294
rect 1052 282 1088 297
rect 1146 282 1182 297
rect 1240 282 1276 297
rect 1334 282 1370 297
rect 1428 282 1464 297
rect 1522 282 1558 297
rect 1616 282 1652 297
rect 1710 282 1746 297
rect 1050 265 1090 282
rect 1144 265 1184 282
rect 1238 265 1278 282
rect 1332 265 1372 282
rect 1426 265 1466 282
rect 1520 265 1560 282
rect 1614 265 1654 282
rect 1708 265 1748 282
rect 22 264 882 265
rect 22 249 224 264
rect 22 215 32 249
rect 66 235 224 249
rect 924 249 988 265
rect 66 215 119 235
rect 924 222 934 249
rect 22 199 119 215
rect 89 177 119 199
rect 287 215 934 222
rect 968 215 988 249
rect 287 192 988 215
rect 287 177 317 192
rect 391 177 421 192
rect 485 177 515 192
rect 579 177 609 192
rect 673 177 703 192
rect 767 177 797 192
rect 861 177 891 192
rect 958 177 988 192
rect 1050 249 1748 265
rect 1050 215 1066 249
rect 1100 215 1144 249
rect 1178 215 1222 249
rect 1256 215 1300 249
rect 1334 215 1378 249
rect 1412 215 1446 249
rect 1480 215 1524 249
rect 1558 215 1602 249
rect 1636 215 1680 249
rect 1714 215 1748 249
rect 1050 199 1748 215
rect 1050 177 1080 199
rect 1144 177 1174 199
rect 1238 177 1268 199
rect 1332 177 1362 199
rect 1426 177 1456 199
rect 1520 177 1550 199
rect 1614 177 1644 199
rect 1718 177 1748 199
rect 89 21 119 47
rect 287 21 317 47
rect 391 21 421 47
rect 485 21 515 47
rect 579 21 609 47
rect 673 21 703 47
rect 767 21 797 47
rect 861 21 891 47
rect 958 21 988 47
rect 1050 21 1080 47
rect 1144 21 1174 47
rect 1238 21 1268 47
rect 1332 21 1362 47
rect 1426 21 1456 47
rect 1520 21 1550 47
rect 1614 21 1644 47
rect 1718 21 1748 47
<< polycont >>
rect 32 215 66 249
rect 934 215 968 249
rect 1066 215 1100 249
rect 1144 215 1178 249
rect 1222 215 1256 249
rect 1300 215 1334 249
rect 1378 215 1412 249
rect 1446 215 1480 249
rect 1524 215 1558 249
rect 1602 215 1636 249
rect 1680 215 1714 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 18 448 69 493
rect 18 414 35 448
rect 18 380 69 414
rect 18 346 35 380
rect 103 489 179 527
rect 103 455 129 489
rect 163 455 179 489
rect 103 421 179 455
rect 103 387 129 421
rect 163 387 179 421
rect 103 367 179 387
rect 213 448 268 493
rect 213 414 234 448
rect 213 380 268 414
rect 18 333 69 346
rect 213 346 234 380
rect 302 489 378 527
rect 302 455 328 489
rect 362 455 378 489
rect 302 421 378 455
rect 302 387 328 421
rect 362 387 378 421
rect 302 367 378 387
rect 422 448 456 493
rect 422 380 456 414
rect 213 333 268 346
rect 490 489 566 527
rect 490 455 516 489
rect 550 455 566 489
rect 490 421 566 455
rect 490 387 516 421
rect 550 387 566 421
rect 490 367 566 387
rect 610 448 644 493
rect 610 380 644 414
rect 422 333 456 346
rect 678 489 754 527
rect 678 455 704 489
rect 738 455 754 489
rect 678 421 754 455
rect 678 387 704 421
rect 738 387 754 421
rect 678 367 754 387
rect 798 448 832 493
rect 798 380 832 414
rect 610 333 644 346
rect 866 485 946 527
rect 866 451 892 485
rect 926 451 946 485
rect 866 417 946 451
rect 866 383 892 417
rect 926 383 946 417
rect 866 367 946 383
rect 990 477 1819 493
rect 990 459 1194 477
rect 990 448 1040 459
rect 990 414 1006 448
rect 1228 459 1382 477
rect 990 380 1040 414
rect 798 333 832 346
rect 990 346 1006 380
rect 990 333 1040 346
rect 18 299 179 333
rect 213 299 1040 333
rect 1074 391 1100 425
rect 1134 391 1150 425
rect 1074 357 1150 391
rect 1194 409 1228 443
rect 1416 459 1570 477
rect 1194 359 1228 375
rect 1262 391 1288 425
rect 1322 391 1338 425
rect 1074 323 1100 357
rect 1134 325 1150 357
rect 1262 357 1338 391
rect 1382 409 1416 443
rect 1604 459 1758 477
rect 1382 359 1416 375
rect 1450 391 1476 425
rect 1510 391 1526 425
rect 1262 325 1288 357
rect 1134 323 1288 325
rect 1322 325 1338 357
rect 1450 357 1526 391
rect 1570 409 1604 443
rect 1792 443 1819 477
rect 1570 359 1604 375
rect 1638 391 1664 425
rect 1698 391 1714 425
rect 1450 325 1476 357
rect 1322 323 1476 325
rect 1510 325 1526 357
rect 1638 357 1714 391
rect 1758 409 1819 443
rect 1792 375 1819 409
rect 1758 359 1819 375
rect 1638 325 1664 357
rect 1510 323 1664 325
rect 1698 325 1714 357
rect 1698 323 1819 325
rect 103 265 179 299
rect 1074 291 1819 323
rect 18 249 69 265
rect 18 215 32 249
rect 66 215 69 249
rect 18 199 69 215
rect 103 249 995 265
rect 103 215 934 249
rect 968 215 995 249
rect 103 199 995 215
rect 1029 249 1730 257
rect 1029 215 1066 249
rect 1100 215 1144 249
rect 1178 215 1222 249
rect 1256 215 1300 249
rect 1334 215 1378 249
rect 1412 215 1446 249
rect 1480 215 1524 249
rect 1558 215 1602 249
rect 1636 215 1680 249
rect 1714 215 1730 249
rect 1029 199 1730 215
rect 103 165 179 199
rect 1774 165 1819 291
rect 18 131 179 165
rect 213 131 1040 165
rect 18 129 69 131
rect 18 95 35 129
rect 213 129 277 131
rect 18 51 69 95
rect 103 93 179 97
rect 103 59 129 93
rect 163 59 179 93
rect 103 17 179 59
rect 213 95 243 129
rect 431 129 465 131
rect 213 51 277 95
rect 321 89 387 97
rect 321 55 337 89
rect 371 55 387 89
rect 321 17 387 55
rect 619 129 653 131
rect 431 51 465 95
rect 509 89 575 97
rect 509 55 525 89
rect 559 55 575 89
rect 509 17 575 55
rect 807 129 841 131
rect 619 51 653 95
rect 697 89 763 97
rect 697 55 713 89
rect 747 55 763 89
rect 697 17 763 55
rect 997 129 1040 131
rect 807 51 841 95
rect 885 89 953 97
rect 885 55 901 89
rect 935 55 953 89
rect 885 17 953 55
rect 997 95 1001 129
rect 1035 95 1040 129
rect 1074 131 1100 165
rect 1134 131 1288 165
rect 1322 131 1476 165
rect 1510 131 1664 165
rect 1698 131 1819 165
rect 1074 124 1819 131
rect 997 90 1040 95
rect 997 56 1194 90
rect 1228 56 1382 90
rect 1416 56 1570 90
rect 1604 56 1758 90
rect 1792 56 1819 90
rect 997 51 1819 56
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel locali s 1316 221 1350 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 1406 221 1440 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1499 221 1533 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1672 357 1706 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1489 357 1523 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1774 153 1808 187 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1774 221 1808 255 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1593 221 1627 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1050 221 1084 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1223 221 1257 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1685 221 1719 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2060134
string GDS_START 2047226
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
