magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2126 1852
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 3 21 795 203
rect 26 -17 60 21
<< scnmos >>
rect 83 47 113 177
rect 175 47 205 177
rect 383 47 413 177
rect 467 47 497 177
rect 599 47 629 177
rect 687 47 717 177
<< scpmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 375 297 411 497
rect 457 297 493 497
rect 591 297 627 497
rect 673 297 709 497
<< ndiff >>
rect 29 161 83 177
rect 29 127 37 161
rect 71 127 83 161
rect 29 93 83 127
rect 29 59 37 93
rect 71 59 83 93
rect 29 47 83 59
rect 113 136 175 177
rect 113 102 131 136
rect 165 102 175 136
rect 113 47 175 102
rect 205 93 267 177
rect 205 59 225 93
rect 259 59 267 93
rect 205 47 267 59
rect 321 95 383 177
rect 321 61 329 95
rect 363 61 383 95
rect 321 47 383 61
rect 413 163 467 177
rect 413 129 423 163
rect 457 129 467 163
rect 413 47 467 129
rect 497 163 599 177
rect 497 129 534 163
rect 568 129 599 163
rect 497 95 599 129
rect 497 61 534 95
rect 568 61 599 95
rect 497 47 599 61
rect 629 89 687 177
rect 629 55 639 89
rect 673 55 687 89
rect 629 47 687 55
rect 717 163 769 177
rect 717 129 727 163
rect 761 129 769 163
rect 717 95 769 129
rect 717 61 727 95
rect 761 61 769 95
rect 717 47 769 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 341 179 375
rect 121 307 133 341
rect 167 307 179 341
rect 121 297 179 307
rect 215 477 375 497
rect 215 443 235 477
rect 269 443 329 477
rect 363 443 375 477
rect 215 409 375 443
rect 215 375 235 409
rect 269 375 329 409
rect 363 375 375 409
rect 215 297 375 375
rect 411 297 457 497
rect 493 477 591 497
rect 493 443 505 477
rect 539 443 591 477
rect 493 409 591 443
rect 493 375 505 409
rect 539 375 591 409
rect 493 341 591 375
rect 493 307 505 341
rect 539 307 591 341
rect 493 297 591 307
rect 627 297 673 497
rect 709 477 767 497
rect 709 443 721 477
rect 755 443 767 477
rect 709 409 767 443
rect 709 375 721 409
rect 755 375 767 409
rect 709 297 767 375
<< ndiffc >>
rect 37 127 71 161
rect 37 59 71 93
rect 131 102 165 136
rect 225 59 259 93
rect 329 61 363 95
rect 423 129 457 163
rect 534 129 568 163
rect 534 61 568 95
rect 639 55 673 89
rect 727 129 761 163
rect 727 61 761 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 443 167 477
rect 133 375 167 409
rect 133 307 167 341
rect 235 443 269 477
rect 329 443 363 477
rect 235 375 269 409
rect 329 375 363 409
rect 505 443 539 477
rect 505 375 539 409
rect 505 307 539 341
rect 721 443 755 477
rect 721 375 755 409
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 375 497 411 523
rect 457 497 493 523
rect 591 497 627 523
rect 673 497 709 523
rect 85 282 121 297
rect 179 282 215 297
rect 375 282 411 297
rect 457 282 493 297
rect 591 282 627 297
rect 673 282 709 297
rect 83 265 123 282
rect 177 265 217 282
rect 373 265 413 282
rect 83 249 274 265
rect 83 215 230 249
rect 264 215 274 249
rect 83 199 274 215
rect 318 249 413 265
rect 318 215 328 249
rect 362 215 413 249
rect 318 199 413 215
rect 455 265 495 282
rect 589 265 629 282
rect 455 249 519 265
rect 455 215 465 249
rect 499 215 519 249
rect 455 199 519 215
rect 561 249 629 265
rect 561 215 575 249
rect 609 215 629 249
rect 561 199 629 215
rect 671 265 711 282
rect 671 249 749 265
rect 671 215 691 249
rect 725 215 749 249
rect 671 199 749 215
rect 83 177 113 199
rect 175 177 205 199
rect 383 177 413 199
rect 467 177 497 199
rect 599 177 629 199
rect 687 177 717 199
rect 83 21 113 47
rect 175 21 205 47
rect 383 21 413 47
rect 467 21 497 47
rect 599 21 629 47
rect 687 21 717 47
<< polycont >>
rect 230 215 264 249
rect 328 215 362 249
rect 465 215 499 249
rect 575 215 609 249
rect 691 215 725 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 23 477 73 527
rect 23 443 39 477
rect 23 409 73 443
rect 23 375 39 409
rect 23 341 73 375
rect 23 307 39 341
rect 23 289 73 307
rect 121 477 171 493
rect 121 443 133 477
rect 167 443 171 477
rect 121 409 171 443
rect 121 375 133 409
rect 167 375 171 409
rect 219 477 379 527
rect 219 443 235 477
rect 269 443 329 477
rect 363 443 379 477
rect 219 409 379 443
rect 219 375 235 409
rect 269 375 329 409
rect 363 375 379 409
rect 468 477 539 493
rect 468 443 505 477
rect 468 409 539 443
rect 468 375 505 409
rect 121 341 171 375
rect 468 341 539 375
rect 121 307 133 341
rect 167 307 171 341
rect 37 161 71 177
rect 37 93 71 127
rect 121 136 171 307
rect 215 307 505 341
rect 215 291 539 307
rect 215 249 271 291
rect 581 255 635 481
rect 714 477 778 527
rect 714 443 721 477
rect 755 443 778 477
rect 714 409 778 443
rect 714 375 721 409
rect 755 375 778 409
rect 714 359 778 375
rect 215 215 230 249
rect 264 215 271 249
rect 305 249 378 255
rect 305 215 328 249
rect 362 215 378 249
rect 422 249 525 255
rect 422 215 465 249
rect 499 215 525 249
rect 559 249 635 255
rect 559 215 575 249
rect 609 215 635 249
rect 669 249 741 323
rect 669 215 691 249
rect 725 215 741 249
rect 215 179 271 215
rect 215 163 473 179
rect 215 143 423 163
rect 121 102 131 136
rect 165 102 171 136
rect 390 129 423 143
rect 457 129 473 163
rect 518 163 778 173
rect 518 129 534 163
rect 568 139 727 163
rect 568 129 586 139
rect 121 73 171 102
rect 225 93 261 109
rect 518 95 586 129
rect 711 129 727 139
rect 761 129 778 163
rect 37 17 71 59
rect 259 59 261 93
rect 313 61 329 95
rect 363 61 534 95
rect 568 61 586 95
rect 313 59 586 61
rect 639 89 673 105
rect 225 17 261 59
rect 711 95 778 129
rect 711 61 727 95
rect 761 61 778 95
rect 711 56 778 61
rect 639 17 673 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 586 357 620 391 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 128 425 162 459 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 324 221 358 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 422 215 525 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel pwell s 26 -17 60 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 26 527 60 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 26 -17 60 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 26 527 60 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o22a_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 941794
string GDS_START 934944
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
