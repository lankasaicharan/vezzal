magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 383 806 704
rect -38 331 270 383
rect 543 331 806 383
<< pwell >>
rect 312 263 501 303
rect 312 157 767 263
rect 1 49 767 157
rect 0 0 768 49
<< scnmos >>
rect 84 47 114 131
rect 162 47 192 131
rect 395 193 425 277
rect 490 153 520 237
rect 576 153 606 237
rect 654 153 684 237
<< scpmoshvt >>
rect 84 409 134 609
rect 425 419 475 619
rect 523 419 573 619
rect 629 419 679 619
<< ndiff >>
rect 27 111 84 131
rect 27 77 39 111
rect 73 77 84 111
rect 27 47 84 77
rect 114 47 162 131
rect 192 93 273 131
rect 192 59 227 93
rect 261 59 273 93
rect 338 265 395 277
rect 338 231 350 265
rect 384 231 395 265
rect 338 193 395 231
rect 425 237 475 277
rect 425 193 490 237
rect 440 153 490 193
rect 520 199 576 237
rect 520 165 531 199
rect 565 165 576 199
rect 520 153 576 165
rect 606 153 654 237
rect 684 212 741 237
rect 684 178 695 212
rect 729 178 741 212
rect 684 153 741 178
rect 192 47 273 59
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 191 609
rect 134 563 145 597
rect 179 563 191 597
rect 134 526 191 563
rect 134 492 145 526
rect 179 492 191 526
rect 134 455 191 492
rect 368 597 425 619
rect 368 563 380 597
rect 414 563 425 597
rect 134 421 145 455
rect 179 421 191 455
rect 134 409 191 421
rect 368 465 425 563
rect 368 431 380 465
rect 414 431 425 465
rect 368 419 425 431
rect 475 419 523 619
rect 573 607 629 619
rect 573 573 584 607
rect 618 573 629 607
rect 573 516 629 573
rect 573 482 584 516
rect 618 482 629 516
rect 573 419 629 482
rect 679 597 736 619
rect 679 563 690 597
rect 724 563 736 597
rect 679 516 736 563
rect 679 482 690 516
rect 724 482 736 516
rect 679 419 736 482
<< ndiffc >>
rect 39 77 73 111
rect 227 59 261 93
rect 350 231 384 265
rect 531 165 565 199
rect 695 178 729 212
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 492 179 526
rect 380 563 414 597
rect 145 421 179 455
rect 380 431 414 465
rect 584 573 618 607
rect 584 482 618 516
rect 690 563 724 597
rect 690 482 724 516
<< poly >>
rect 84 609 134 635
rect 425 619 475 645
rect 523 619 573 645
rect 629 619 679 645
rect 232 463 298 479
rect 232 429 248 463
rect 282 429 298 463
rect 84 287 134 409
rect 232 395 298 429
rect 232 361 248 395
rect 282 375 298 395
rect 425 375 475 419
rect 282 361 475 375
rect 232 345 475 361
rect 523 387 573 419
rect 629 387 679 419
rect 523 371 679 387
rect 84 271 175 287
rect 84 237 125 271
rect 159 237 175 271
rect 84 203 175 237
rect 232 281 318 297
rect 232 247 248 281
rect 282 247 318 281
rect 395 277 425 345
rect 523 337 539 371
rect 573 351 679 371
rect 573 337 684 351
rect 523 321 684 337
rect 232 231 318 247
rect 84 169 125 203
rect 159 183 175 203
rect 159 169 192 183
rect 84 153 192 169
rect 84 131 114 153
rect 162 131 192 153
rect 288 119 318 231
rect 490 237 520 263
rect 576 237 606 321
rect 654 237 684 321
rect 395 167 425 193
rect 490 119 520 153
rect 576 127 606 153
rect 654 127 684 153
rect 288 89 520 119
rect 84 21 114 47
rect 162 21 192 47
<< polycont >>
rect 248 429 282 463
rect 248 361 282 395
rect 125 237 159 271
rect 248 247 282 281
rect 539 337 573 371
rect 125 169 159 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 526 89 563
rect 23 492 39 526
rect 73 492 89 526
rect 23 455 89 492
rect 23 421 39 455
rect 73 421 89 455
rect 23 369 89 421
rect 129 597 195 649
rect 129 563 145 597
rect 179 563 195 597
rect 129 526 195 563
rect 129 492 145 526
rect 179 492 195 526
rect 129 455 195 492
rect 364 597 455 613
rect 364 563 380 597
rect 414 563 455 597
rect 129 421 145 455
rect 179 421 195 455
rect 129 405 195 421
rect 232 463 298 479
rect 232 429 248 463
rect 282 429 298 463
rect 232 395 298 429
rect 364 465 455 563
rect 568 607 634 649
rect 568 573 584 607
rect 618 573 634 607
rect 568 516 634 573
rect 568 482 584 516
rect 618 482 634 516
rect 568 466 634 482
rect 674 597 745 613
rect 674 563 690 597
rect 724 563 745 597
rect 674 516 745 563
rect 674 482 690 516
rect 724 482 745 516
rect 674 466 745 482
rect 364 431 380 465
rect 414 431 455 465
rect 364 415 455 431
rect 232 369 248 395
rect 23 361 248 369
rect 282 361 298 395
rect 23 335 298 361
rect 409 355 455 415
rect 23 111 73 335
rect 334 321 455 355
rect 505 371 647 430
rect 505 337 539 371
rect 573 337 647 371
rect 505 321 647 337
rect 23 77 39 111
rect 109 271 175 287
rect 109 237 125 271
rect 159 237 175 271
rect 109 203 175 237
rect 109 169 125 203
rect 159 169 175 203
rect 109 88 175 169
rect 232 281 298 297
rect 232 247 248 281
rect 282 247 298 281
rect 232 179 298 247
rect 334 265 400 321
rect 711 285 745 466
rect 334 231 350 265
rect 384 231 400 265
rect 334 215 400 231
rect 436 251 745 285
rect 436 179 470 251
rect 232 145 470 179
rect 515 199 581 215
rect 515 165 531 199
rect 565 165 581 199
rect 211 93 277 109
rect 23 53 73 77
rect 211 59 227 93
rect 261 59 277 93
rect 211 17 277 59
rect 515 17 581 165
rect 679 212 745 251
rect 679 178 695 212
rect 729 178 745 212
rect 679 149 745 178
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ebufn_lp2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3403648
string GDS_START 3397036
<< end >>
