magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4178 1975
<< nwell >>
rect -38 331 2918 704
rect 725 321 1027 331
<< pwell >>
rect 1689 273 2009 279
rect 743 229 1057 241
rect 1388 229 2009 273
rect 743 201 2009 229
rect 743 167 2377 201
rect 2577 167 2875 251
rect 1 157 197 164
rect 743 157 2875 167
rect 1 49 2875 157
rect 0 0 2880 49
<< scnmos >>
rect 84 54 114 138
rect 282 47 312 131
rect 360 47 390 131
rect 456 47 486 131
rect 534 47 564 131
rect 620 47 650 131
rect 826 47 856 215
rect 944 47 974 215
rect 1172 119 1202 203
rect 1289 119 1319 203
rect 1361 119 1391 203
rect 1471 119 1501 247
rect 1549 119 1579 247
rect 1795 125 1825 253
rect 1873 125 1903 253
rect 2005 91 2035 175
rect 2083 91 2113 175
rect 2192 47 2222 175
rect 2264 47 2294 175
rect 2462 57 2492 141
rect 2660 57 2690 225
rect 2762 57 2792 225
<< scpmoshvt >>
rect 132 531 162 615
rect 234 531 264 615
rect 312 531 342 615
rect 398 531 428 615
rect 504 531 534 615
rect 606 531 636 615
rect 818 357 848 609
rect 904 357 934 609
rect 1109 463 1139 547
rect 1195 463 1225 547
rect 1273 463 1303 547
rect 1471 373 1501 541
rect 1603 373 1633 541
rect 1801 373 1831 541
rect 1903 409 1933 577
rect 2012 451 2042 535
rect 2090 451 2120 535
rect 2215 451 2245 619
rect 2301 451 2331 619
rect 2426 451 2456 579
rect 2654 367 2684 619
rect 2756 367 2786 619
<< ndiff >>
rect 27 113 84 138
rect 27 79 39 113
rect 73 79 84 113
rect 27 54 84 79
rect 114 114 171 138
rect 769 184 826 215
rect 769 150 781 184
rect 815 150 826 184
rect 114 80 125 114
rect 159 80 171 114
rect 114 54 171 80
rect 225 106 282 131
rect 225 72 237 106
rect 271 72 282 106
rect 225 47 282 72
rect 312 47 360 131
rect 390 111 456 131
rect 390 77 411 111
rect 445 77 456 111
rect 390 47 456 77
rect 486 47 534 131
rect 564 106 620 131
rect 564 72 575 106
rect 609 72 620 106
rect 564 47 620 72
rect 650 111 707 131
rect 650 77 661 111
rect 695 77 707 111
rect 650 47 707 77
rect 769 103 826 150
rect 769 69 781 103
rect 815 69 826 103
rect 769 47 826 69
rect 856 103 944 215
rect 856 69 883 103
rect 917 69 944 103
rect 856 47 944 69
rect 974 193 1031 215
rect 1414 203 1471 247
rect 974 159 985 193
rect 1019 159 1031 193
rect 974 103 1031 159
rect 1115 178 1172 203
rect 1115 144 1127 178
rect 1161 144 1172 178
rect 1115 119 1172 144
rect 1202 178 1289 203
rect 1202 144 1244 178
rect 1278 144 1289 178
rect 1202 119 1289 144
rect 1319 119 1361 203
rect 1391 194 1471 203
rect 1391 160 1426 194
rect 1460 160 1471 194
rect 1391 119 1471 160
rect 1501 119 1549 247
rect 1579 194 1636 247
rect 1579 160 1590 194
rect 1624 160 1636 194
rect 1579 119 1636 160
rect 1715 197 1795 253
rect 1715 163 1727 197
rect 1761 163 1795 197
rect 1715 125 1795 163
rect 1825 125 1873 253
rect 1903 223 1983 253
rect 1903 189 1937 223
rect 1971 189 1983 223
rect 1903 175 1983 189
rect 1903 137 2005 175
rect 1903 125 1937 137
rect 974 69 985 103
rect 1019 69 1031 103
rect 974 47 1031 69
rect 1925 103 1937 125
rect 1971 103 2005 137
rect 1925 91 2005 103
rect 2035 91 2083 175
rect 2113 119 2192 175
rect 2113 91 2147 119
rect 2135 85 2147 91
rect 2181 85 2192 119
rect 2135 47 2192 85
rect 2222 47 2264 175
rect 2294 133 2351 175
rect 2603 213 2660 225
rect 2603 179 2615 213
rect 2649 179 2660 213
rect 2294 99 2305 133
rect 2339 99 2351 133
rect 2294 47 2351 99
rect 2405 116 2462 141
rect 2405 82 2417 116
rect 2451 82 2462 116
rect 2405 57 2462 82
rect 2492 116 2549 141
rect 2492 82 2503 116
rect 2537 82 2549 116
rect 2492 57 2549 82
rect 2603 103 2660 179
rect 2603 69 2615 103
rect 2649 69 2660 103
rect 2603 57 2660 69
rect 2690 213 2762 225
rect 2690 179 2701 213
rect 2735 179 2762 213
rect 2690 103 2762 179
rect 2690 69 2701 103
rect 2735 69 2762 103
rect 2690 57 2762 69
rect 2792 213 2849 225
rect 2792 179 2803 213
rect 2837 179 2849 213
rect 2792 103 2849 179
rect 2792 69 2803 103
rect 2837 69 2849 103
rect 2792 57 2849 69
<< pdiff >>
rect 75 587 132 615
rect 75 553 87 587
rect 121 553 132 587
rect 75 531 132 553
rect 162 590 234 615
rect 162 556 189 590
rect 223 556 234 590
rect 162 531 234 556
rect 264 531 312 615
rect 342 587 398 615
rect 342 553 353 587
rect 387 553 398 587
rect 342 531 398 553
rect 428 531 504 615
rect 534 603 606 615
rect 534 569 545 603
rect 579 569 606 603
rect 534 531 606 569
rect 636 591 693 615
rect 636 557 647 591
rect 681 557 693 591
rect 636 531 693 557
rect 761 597 818 609
rect 761 563 773 597
rect 807 563 818 597
rect 761 500 818 563
rect 761 466 773 500
rect 807 466 818 500
rect 761 403 818 466
rect 761 369 773 403
rect 807 369 818 403
rect 761 357 818 369
rect 848 597 904 609
rect 848 563 859 597
rect 893 563 904 597
rect 848 528 904 563
rect 848 494 859 528
rect 893 494 904 528
rect 848 459 904 494
rect 848 425 859 459
rect 893 425 904 459
rect 848 357 904 425
rect 934 597 991 609
rect 934 563 945 597
rect 979 563 991 597
rect 934 500 991 563
rect 934 466 945 500
rect 979 466 991 500
rect 934 403 991 466
rect 934 369 945 403
rect 979 369 991 403
rect 934 357 991 369
rect 1523 586 1581 598
rect 1052 522 1109 547
rect 1052 488 1064 522
rect 1098 488 1109 522
rect 1052 463 1109 488
rect 1139 528 1195 547
rect 1139 494 1150 528
rect 1184 494 1195 528
rect 1139 463 1195 494
rect 1225 463 1273 547
rect 1303 522 1360 547
rect 1523 552 1535 586
rect 1569 552 1581 586
rect 2142 596 2215 619
rect 1523 541 1581 552
rect 1853 541 1903 577
rect 1303 488 1314 522
rect 1348 488 1360 522
rect 1303 463 1360 488
rect 1414 529 1471 541
rect 1414 495 1426 529
rect 1460 495 1471 529
rect 1414 427 1471 495
rect 1414 393 1426 427
rect 1460 393 1471 427
rect 1414 373 1471 393
rect 1501 373 1603 541
rect 1633 529 1690 541
rect 1633 495 1644 529
rect 1678 495 1690 529
rect 1633 427 1690 495
rect 1633 393 1644 427
rect 1678 393 1690 427
rect 1633 373 1690 393
rect 1744 529 1801 541
rect 1744 495 1756 529
rect 1790 495 1801 529
rect 1744 427 1801 495
rect 1744 393 1756 427
rect 1790 393 1801 427
rect 1744 373 1801 393
rect 1831 409 1903 541
rect 1933 565 1990 577
rect 1933 531 1944 565
rect 1978 535 1990 565
rect 2142 562 2154 596
rect 2188 562 2215 596
rect 2142 535 2215 562
rect 1978 531 2012 535
rect 1933 455 2012 531
rect 1933 421 1944 455
rect 1978 451 2012 455
rect 2042 451 2090 535
rect 2120 451 2215 535
rect 2245 597 2301 619
rect 2245 563 2256 597
rect 2290 563 2301 597
rect 2245 516 2301 563
rect 2245 482 2256 516
rect 2290 482 2301 516
rect 2245 451 2301 482
rect 2331 607 2404 619
rect 2331 573 2358 607
rect 2392 579 2404 607
rect 2392 573 2426 579
rect 2331 505 2426 573
rect 2331 471 2358 505
rect 2392 471 2426 505
rect 2331 451 2426 471
rect 2456 567 2513 579
rect 2456 533 2467 567
rect 2501 533 2513 567
rect 2456 497 2513 533
rect 2456 463 2467 497
rect 2501 463 2513 497
rect 2456 451 2513 463
rect 1978 421 1990 451
rect 1933 409 1990 421
rect 1831 373 1881 409
rect 2597 413 2654 619
rect 2597 379 2609 413
rect 2643 379 2654 413
rect 2597 367 2654 379
rect 2684 596 2756 619
rect 2684 562 2695 596
rect 2729 562 2756 596
rect 2684 367 2756 562
rect 2786 597 2843 619
rect 2786 563 2797 597
rect 2831 563 2843 597
rect 2786 507 2843 563
rect 2786 473 2797 507
rect 2831 473 2843 507
rect 2786 417 2843 473
rect 2786 383 2797 417
rect 2831 383 2843 417
rect 2786 367 2843 383
<< ndiffc >>
rect 39 79 73 113
rect 781 150 815 184
rect 125 80 159 114
rect 237 72 271 106
rect 411 77 445 111
rect 575 72 609 106
rect 661 77 695 111
rect 781 69 815 103
rect 883 69 917 103
rect 985 159 1019 193
rect 1127 144 1161 178
rect 1244 144 1278 178
rect 1426 160 1460 194
rect 1590 160 1624 194
rect 1727 163 1761 197
rect 1937 189 1971 223
rect 985 69 1019 103
rect 1937 103 1971 137
rect 2147 85 2181 119
rect 2615 179 2649 213
rect 2305 99 2339 133
rect 2417 82 2451 116
rect 2503 82 2537 116
rect 2615 69 2649 103
rect 2701 179 2735 213
rect 2701 69 2735 103
rect 2803 179 2837 213
rect 2803 69 2837 103
<< pdiffc >>
rect 87 553 121 587
rect 189 556 223 590
rect 353 553 387 587
rect 545 569 579 603
rect 647 557 681 591
rect 773 563 807 597
rect 773 466 807 500
rect 773 369 807 403
rect 859 563 893 597
rect 859 494 893 528
rect 859 425 893 459
rect 945 563 979 597
rect 945 466 979 500
rect 945 369 979 403
rect 1064 488 1098 522
rect 1150 494 1184 528
rect 1535 552 1569 586
rect 1314 488 1348 522
rect 1426 495 1460 529
rect 1426 393 1460 427
rect 1644 495 1678 529
rect 1644 393 1678 427
rect 1756 495 1790 529
rect 1756 393 1790 427
rect 1944 531 1978 565
rect 2154 562 2188 596
rect 1944 421 1978 455
rect 2256 563 2290 597
rect 2256 482 2290 516
rect 2358 573 2392 607
rect 2358 471 2392 505
rect 2467 533 2501 567
rect 2467 463 2501 497
rect 2609 379 2643 413
rect 2695 562 2729 596
rect 2797 563 2831 597
rect 2797 473 2831 507
rect 2797 383 2831 417
<< poly >>
rect 132 615 162 641
rect 234 615 264 641
rect 312 615 342 641
rect 398 615 428 641
rect 504 615 534 641
rect 606 615 636 641
rect 818 609 848 635
rect 904 609 934 635
rect 1006 615 1933 645
rect 2215 619 2245 645
rect 2301 619 2331 645
rect 2654 619 2684 645
rect 2756 619 2786 645
rect 132 361 162 531
rect 234 361 264 531
rect 84 345 264 361
rect 84 311 112 345
rect 146 331 264 345
rect 146 311 162 331
rect 84 295 162 311
rect 312 322 342 531
rect 398 463 428 531
rect 390 447 456 463
rect 390 413 406 447
rect 440 413 456 447
rect 390 397 456 413
rect 504 401 534 531
rect 606 499 636 531
rect 606 483 672 499
rect 606 449 622 483
rect 656 463 672 483
rect 656 449 732 463
rect 606 433 732 449
rect 504 371 564 401
rect 534 355 660 371
rect 84 138 114 295
rect 312 275 384 322
rect 162 228 228 244
rect 162 194 178 228
rect 212 194 228 228
rect 312 241 328 275
rect 362 241 384 275
rect 426 307 492 323
rect 426 273 442 307
rect 476 273 492 307
rect 426 257 492 273
rect 534 321 610 355
rect 644 321 660 355
rect 534 287 660 321
rect 312 225 384 241
rect 162 183 228 194
rect 354 209 384 225
rect 162 153 312 183
rect 354 179 390 209
rect 282 131 312 153
rect 360 131 390 179
rect 456 131 486 257
rect 534 253 610 287
rect 644 253 660 287
rect 534 237 660 253
rect 534 131 564 237
rect 702 183 732 433
rect 818 303 848 357
rect 774 287 848 303
rect 774 253 790 287
rect 824 267 848 287
rect 904 311 934 357
rect 1006 311 1036 615
rect 1109 547 1139 573
rect 1195 547 1225 615
rect 1273 547 1303 573
rect 1471 541 1501 567
rect 1903 577 1933 615
rect 1603 541 1633 567
rect 1801 541 1831 567
rect 1109 381 1139 463
rect 1195 437 1225 463
rect 1273 423 1303 463
rect 1273 407 1391 423
rect 1273 393 1332 407
rect 1078 365 1144 381
rect 1078 331 1094 365
rect 1128 345 1144 365
rect 1316 373 1332 393
rect 1366 373 1391 407
rect 2012 535 2042 561
rect 2090 535 2120 561
rect 2426 579 2456 605
rect 1903 383 1933 409
rect 1316 357 1391 373
rect 1128 331 1274 345
rect 1078 315 1274 331
rect 904 295 1036 311
rect 824 253 856 267
rect 774 237 856 253
rect 904 261 920 295
rect 954 267 1036 295
rect 1244 309 1274 315
rect 1244 279 1319 309
rect 954 261 1202 267
rect 904 237 1202 261
rect 826 215 856 237
rect 944 215 974 237
rect 620 153 732 183
rect 620 131 650 153
rect 84 28 114 54
rect 1172 203 1202 237
rect 1289 203 1319 279
rect 1361 203 1391 357
rect 1471 341 1501 373
rect 1603 341 1633 373
rect 1801 341 1831 373
rect 2012 341 2042 451
rect 2090 419 2120 451
rect 1435 325 1501 341
rect 1435 291 1451 325
rect 1485 291 1501 325
rect 1435 275 1501 291
rect 1471 247 1501 275
rect 1549 325 1633 341
rect 1549 291 1565 325
rect 1599 291 1633 325
rect 1549 275 1633 291
rect 1747 325 1831 341
rect 1747 291 1763 325
rect 1797 311 1831 325
rect 1873 325 2042 341
rect 1797 291 1825 311
rect 1747 275 1825 291
rect 1549 247 1579 275
rect 1795 253 1825 275
rect 1873 291 1889 325
rect 1923 311 2042 325
rect 2084 403 2150 419
rect 2084 369 2100 403
rect 2134 369 2150 403
rect 2084 353 2150 369
rect 1923 291 1939 311
rect 1873 275 1939 291
rect 1873 253 1903 275
rect 2084 227 2114 353
rect 2215 305 2245 451
rect 2005 175 2035 201
rect 2083 197 2114 227
rect 2156 275 2245 305
rect 2301 419 2331 451
rect 2301 403 2378 419
rect 2301 369 2317 403
rect 2351 369 2378 403
rect 2301 353 2378 369
rect 2426 357 2456 451
rect 2156 247 2222 275
rect 2156 213 2172 247
rect 2206 213 2222 247
rect 2301 227 2331 353
rect 2420 341 2492 357
rect 2420 307 2436 341
rect 2470 321 2492 341
rect 2654 321 2684 367
rect 2756 331 2786 367
rect 2470 307 2690 321
rect 2420 291 2690 307
rect 2156 197 2222 213
rect 2083 175 2113 197
rect 2192 175 2222 197
rect 2264 197 2331 227
rect 2264 175 2294 197
rect 1172 51 1202 119
rect 1289 93 1319 119
rect 1361 93 1391 119
rect 1471 93 1501 119
rect 1549 93 1579 119
rect 1795 99 1825 125
rect 1873 99 1903 125
rect 2005 51 2035 91
rect 2083 65 2113 91
rect 282 21 312 47
rect 360 21 390 47
rect 456 21 486 47
rect 534 21 564 47
rect 620 21 650 47
rect 826 21 856 47
rect 944 21 974 47
rect 1172 21 2035 51
rect 2462 141 2492 291
rect 2660 225 2690 291
rect 2732 315 2798 331
rect 2732 281 2748 315
rect 2782 281 2798 315
rect 2732 265 2798 281
rect 2762 225 2792 265
rect 2192 21 2222 47
rect 2264 21 2294 47
rect 2462 31 2492 57
rect 2660 31 2690 57
rect 2762 31 2792 57
<< polycont >>
rect 112 311 146 345
rect 406 413 440 447
rect 622 449 656 483
rect 178 194 212 228
rect 328 241 362 275
rect 442 273 476 307
rect 610 321 644 355
rect 610 253 644 287
rect 790 253 824 287
rect 1094 331 1128 365
rect 1332 373 1366 407
rect 920 261 954 295
rect 1451 291 1485 325
rect 1565 291 1599 325
rect 1763 291 1797 325
rect 1889 291 1923 325
rect 2100 369 2134 403
rect 2317 369 2351 403
rect 2172 213 2206 247
rect 2436 307 2470 341
rect 2748 281 2782 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 26 587 137 613
rect 26 553 87 587
rect 121 553 137 587
rect 26 527 137 553
rect 173 590 239 649
rect 173 556 189 590
rect 223 556 239 590
rect 173 527 239 556
rect 337 587 403 613
rect 337 553 353 587
rect 387 553 403 587
rect 529 603 595 649
rect 529 569 545 603
rect 579 569 595 603
rect 631 591 697 613
rect 337 533 403 553
rect 631 557 647 591
rect 681 569 697 591
rect 773 597 807 613
rect 681 557 737 569
rect 631 535 737 557
rect 26 463 60 527
rect 337 499 560 533
rect 526 483 667 499
rect 26 447 456 463
rect 26 413 406 447
rect 440 413 456 447
rect 26 397 456 413
rect 526 449 622 483
rect 656 449 667 483
rect 526 433 667 449
rect 26 244 60 397
rect 96 345 490 361
rect 96 311 112 345
rect 146 327 490 345
rect 146 311 263 327
rect 96 295 263 311
rect 426 307 490 327
rect 312 275 378 291
rect 26 228 228 244
rect 26 194 178 228
rect 212 194 228 228
rect 312 241 328 275
rect 362 241 378 275
rect 426 273 442 307
rect 476 273 490 307
rect 426 257 490 273
rect 312 225 378 241
rect 526 205 560 433
rect 596 355 660 371
rect 596 321 610 355
rect 644 321 660 355
rect 596 287 660 321
rect 596 253 610 287
rect 644 253 660 287
rect 596 236 660 253
rect 26 178 228 194
rect 23 113 73 142
rect 23 79 39 113
rect 23 17 73 79
rect 109 114 175 178
rect 427 171 560 205
rect 427 135 461 171
rect 703 135 737 535
rect 773 500 807 563
rect 773 403 807 466
rect 843 597 909 649
rect 843 563 859 597
rect 893 563 909 597
rect 843 528 909 563
rect 843 494 859 528
rect 893 494 909 528
rect 843 459 909 494
rect 843 425 859 459
rect 893 425 909 459
rect 843 409 909 425
rect 945 597 1006 613
rect 979 563 1006 597
rect 945 500 1006 563
rect 979 466 1006 500
rect 945 403 1006 466
rect 1048 522 1098 551
rect 1048 488 1064 522
rect 1048 451 1098 488
rect 1134 528 1278 551
rect 1134 494 1150 528
rect 1184 494 1278 528
rect 1134 487 1278 494
rect 1048 417 1208 451
rect 807 369 909 373
rect 773 339 909 369
rect 979 381 1006 403
rect 979 369 1138 381
rect 945 365 1138 369
rect 945 350 1094 365
rect 945 347 1087 350
rect 875 311 909 339
rect 1006 316 1087 347
rect 1128 331 1138 365
rect 1121 316 1138 331
rect 774 287 839 303
rect 774 253 790 287
rect 824 253 839 287
rect 774 236 839 253
rect 875 295 970 311
rect 875 261 920 295
rect 954 261 970 295
rect 875 245 970 261
rect 1006 310 1138 316
rect 875 200 909 245
rect 1006 209 1040 310
rect 781 184 909 200
rect 815 166 909 184
rect 969 193 1040 209
rect 1174 207 1208 417
rect 815 150 831 166
rect 109 80 125 114
rect 159 80 175 114
rect 109 53 175 80
rect 221 106 287 135
rect 221 72 237 106
rect 271 72 287 106
rect 221 17 287 72
rect 395 111 461 135
rect 395 77 411 111
rect 445 77 461 111
rect 395 53 461 77
rect 559 106 609 135
rect 559 72 575 106
rect 559 17 609 72
rect 645 128 743 135
rect 645 111 703 128
rect 645 77 661 111
rect 695 94 703 111
rect 737 94 743 128
rect 695 77 743 94
rect 645 53 743 77
rect 781 103 831 150
rect 969 159 985 193
rect 1019 159 1040 193
rect 815 69 831 103
rect 781 53 831 69
rect 867 103 933 130
rect 867 69 883 103
rect 917 69 933 103
rect 867 17 933 69
rect 969 103 1040 159
rect 969 69 985 103
rect 1019 69 1040 103
rect 1081 178 1208 207
rect 1081 144 1127 178
rect 1161 144 1208 178
rect 1081 128 1208 144
rect 1081 94 1087 128
rect 1121 94 1208 128
rect 1244 309 1278 487
rect 1314 522 1364 649
rect 1519 586 1585 649
rect 1519 552 1535 586
rect 1569 552 1585 586
rect 1348 488 1364 522
rect 1314 459 1364 488
rect 1410 529 1476 545
rect 1519 536 1585 552
rect 1410 495 1426 529
rect 1460 500 1476 529
rect 1644 529 1694 545
rect 1460 495 1644 500
rect 1678 495 1694 529
rect 1410 466 1694 495
rect 1410 427 1476 466
rect 1410 423 1426 427
rect 1316 407 1426 423
rect 1316 373 1332 407
rect 1366 393 1426 407
rect 1460 393 1476 427
rect 1366 377 1476 393
rect 1549 424 1607 430
rect 1549 390 1567 424
rect 1601 390 1607 424
rect 1366 373 1382 377
rect 1316 357 1382 373
rect 1549 341 1607 390
rect 1644 427 1694 466
rect 1678 393 1694 427
rect 1644 377 1694 393
rect 1740 529 1806 649
rect 2138 596 2204 649
rect 1740 495 1756 529
rect 1790 495 1806 529
rect 1740 427 1806 495
rect 1740 393 1756 427
rect 1790 393 1806 427
rect 1928 565 1994 581
rect 1928 531 1944 565
rect 1978 531 1994 565
rect 2138 562 2154 596
rect 2188 562 2204 596
rect 2138 536 2204 562
rect 2240 597 2306 613
rect 2240 563 2256 597
rect 2290 563 2306 597
rect 1928 455 1994 531
rect 2240 516 2306 563
rect 2240 500 2256 516
rect 1928 421 1944 455
rect 1978 439 1994 455
rect 2116 482 2256 500
rect 2290 482 2306 516
rect 2116 466 2306 482
rect 2342 607 2408 649
rect 2342 573 2358 607
rect 2392 573 2408 607
rect 2679 596 2745 649
rect 2342 505 2408 573
rect 2342 471 2358 505
rect 2392 471 2408 505
rect 1978 421 2009 439
rect 1928 405 2009 421
rect 2116 419 2150 466
rect 2342 455 2408 471
rect 2451 567 2517 583
rect 2451 533 2467 567
rect 2501 533 2517 567
rect 2679 562 2695 596
rect 2729 562 2745 596
rect 2679 535 2745 562
rect 2781 597 2862 613
rect 2781 563 2797 597
rect 2831 563 2862 597
rect 2451 499 2517 533
rect 2781 507 2862 563
rect 2451 497 2745 499
rect 2451 463 2467 497
rect 2501 465 2745 497
rect 2501 463 2556 465
rect 2451 447 2556 463
rect 1740 377 1806 393
rect 1651 341 1685 377
rect 1849 350 1939 356
rect 1435 325 1501 341
rect 1435 309 1451 325
rect 1244 291 1451 309
rect 1485 291 1501 325
rect 1244 275 1501 291
rect 1549 325 1615 341
rect 1549 291 1565 325
rect 1599 291 1615 325
rect 1549 275 1615 291
rect 1651 325 1813 341
rect 1651 291 1763 325
rect 1797 291 1813 325
rect 1651 275 1813 291
rect 1849 316 1855 350
rect 1889 325 1939 350
rect 1849 291 1889 316
rect 1923 291 1939 325
rect 1849 275 1939 291
rect 1244 178 1294 275
rect 1651 239 1685 275
rect 1975 239 2009 405
rect 2084 403 2150 419
rect 2084 369 2100 403
rect 2134 369 2150 403
rect 2084 353 2150 369
rect 2233 424 2279 430
rect 2233 390 2239 424
rect 2273 419 2279 424
rect 2273 403 2367 419
rect 2273 390 2317 403
rect 2233 369 2317 390
rect 2351 369 2367 403
rect 2233 361 2367 369
rect 2116 325 2150 353
rect 2420 341 2486 357
rect 2420 325 2436 341
rect 2116 307 2436 325
rect 2470 307 2486 341
rect 2116 291 2486 307
rect 2156 247 2222 255
rect 2156 239 2172 247
rect 1278 144 1294 178
rect 1244 115 1294 144
rect 1410 194 1476 239
rect 1410 160 1426 194
rect 1460 160 1476 194
rect 1081 88 1208 94
rect 969 53 1040 69
rect 1410 17 1476 160
rect 1574 194 1685 239
rect 1574 160 1590 194
rect 1624 160 1685 194
rect 1574 115 1685 160
rect 1727 197 1777 239
rect 1761 163 1777 197
rect 1727 17 1777 163
rect 1921 223 2172 239
rect 1921 189 1937 223
rect 1971 213 2172 223
rect 2206 213 2222 247
rect 1971 197 2222 213
rect 1971 189 2009 197
rect 1921 137 2009 189
rect 1921 103 1937 137
rect 1971 103 2009 137
rect 1921 87 2009 103
rect 2131 119 2197 161
rect 2131 85 2147 119
rect 2181 85 2197 119
rect 2131 17 2197 85
rect 2289 133 2355 291
rect 2522 145 2556 447
rect 2289 99 2305 133
rect 2339 99 2355 133
rect 2289 53 2355 99
rect 2401 116 2451 145
rect 2401 82 2417 116
rect 2401 17 2451 82
rect 2487 116 2556 145
rect 2487 82 2503 116
rect 2537 82 2556 116
rect 2487 53 2556 82
rect 2593 413 2665 429
rect 2593 379 2609 413
rect 2643 379 2665 413
rect 2593 276 2665 379
rect 2593 242 2623 276
rect 2657 242 2665 276
rect 2711 331 2745 465
rect 2781 473 2797 507
rect 2831 473 2862 507
rect 2781 424 2862 473
rect 2781 417 2815 424
rect 2781 383 2797 417
rect 2849 390 2862 424
rect 2831 383 2862 390
rect 2781 367 2862 383
rect 2711 315 2792 331
rect 2711 281 2748 315
rect 2782 281 2792 315
rect 2711 265 2792 281
rect 2593 213 2665 242
rect 2828 229 2862 367
rect 2593 179 2615 213
rect 2649 179 2665 213
rect 2593 103 2665 179
rect 2593 69 2615 103
rect 2649 69 2665 103
rect 2593 53 2665 69
rect 2701 213 2751 229
rect 2735 179 2751 213
rect 2701 103 2751 179
rect 2735 69 2751 103
rect 2701 17 2751 69
rect 2787 213 2862 229
rect 2787 179 2803 213
rect 2837 179 2862 213
rect 2787 103 2862 179
rect 2787 69 2803 103
rect 2837 69 2862 103
rect 2787 53 2862 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 1087 331 1094 350
rect 1094 331 1121 350
rect 1087 316 1121 331
rect 703 94 737 128
rect 1087 94 1121 128
rect 1567 390 1601 424
rect 1855 316 1889 350
rect 2239 390 2273 424
rect 2623 242 2657 276
rect 2815 417 2849 424
rect 2815 390 2831 417
rect 2831 390 2849 417
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 1555 424 1613 430
rect 1555 390 1567 424
rect 1601 421 1613 424
rect 2227 424 2285 430
rect 2227 421 2239 424
rect 1601 393 2239 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2227 390 2239 393
rect 2273 390 2285 424
rect 2803 424 2861 430
rect 2227 384 2285 390
rect 2626 393 2753 421
rect 1075 350 1133 356
rect 1075 316 1087 350
rect 1121 347 1133 350
rect 1843 350 1901 356
rect 1843 347 1855 350
rect 1121 319 1855 347
rect 1121 316 1133 319
rect 1075 310 1133 316
rect 1843 316 1855 319
rect 1889 316 1901 350
rect 1843 310 1901 316
rect 2626 282 2654 393
rect 2803 390 2815 424
rect 2849 390 2861 424
rect 2803 384 2861 390
rect 2611 276 2669 282
rect 2611 242 2623 276
rect 2657 242 2669 276
rect 2818 273 2846 384
rect 2719 245 2846 273
rect 2611 236 2669 242
rect 691 128 749 134
rect 691 94 703 128
rect 737 125 749 128
rect 1075 128 1133 134
rect 1075 125 1087 128
rect 737 97 1087 125
rect 737 94 749 97
rect 691 88 749 94
rect 1075 94 1087 97
rect 1121 94 1133 128
rect 1075 88 1133 94
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sregrbp_1
flabel metal1 s 2239 390 2273 424 0 FreeSans 200 0 0 0 ASYNC
port 1 nsew signal input
flabel metal1 s 2719 393 2753 421 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel metal1 s 2719 245 2753 273 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 3 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 2 nsew clock input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2880 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2758424
string GDS_START 2737610
<< end >>
