magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 157 605 261
rect 1 49 765 157
rect 0 0 768 49
<< scnmos >>
rect 80 151 110 235
rect 217 151 247 235
rect 289 151 319 235
rect 397 151 427 235
rect 469 151 499 235
rect 656 47 686 131
<< scpmoshvt >>
rect 93 403 123 487
rect 217 411 247 495
rect 303 411 333 495
rect 397 411 427 495
rect 483 411 513 495
rect 616 411 646 495
<< ndiff >>
rect 27 202 80 235
rect 27 168 35 202
rect 69 168 80 202
rect 27 151 80 168
rect 110 197 217 235
rect 110 163 137 197
rect 171 163 217 197
rect 110 151 217 163
rect 247 151 289 235
rect 319 151 397 235
rect 427 151 469 235
rect 499 227 579 235
rect 499 193 533 227
rect 567 193 579 227
rect 499 185 579 193
rect 499 151 549 185
rect 603 93 656 131
rect 603 59 611 93
rect 645 59 656 93
rect 603 47 656 59
rect 686 115 739 131
rect 686 81 697 115
rect 731 81 739 115
rect 686 47 739 81
<< pdiff >>
rect 145 487 217 495
rect 40 475 93 487
rect 40 441 48 475
rect 82 441 93 475
rect 40 403 93 441
rect 123 483 217 487
rect 123 449 153 483
rect 187 449 217 483
rect 123 411 217 449
rect 247 457 303 495
rect 247 423 258 457
rect 292 423 303 457
rect 247 411 303 423
rect 333 483 397 495
rect 333 449 344 483
rect 378 449 397 483
rect 333 411 397 449
rect 427 483 483 495
rect 427 449 438 483
rect 472 449 483 483
rect 427 411 483 449
rect 513 483 616 495
rect 513 449 524 483
rect 558 449 616 483
rect 513 411 616 449
rect 646 457 699 495
rect 646 423 657 457
rect 691 423 699 457
rect 646 411 699 423
rect 123 403 195 411
<< ndiffc >>
rect 35 168 69 202
rect 137 163 171 197
rect 533 193 567 227
rect 611 59 645 93
rect 697 81 731 115
<< pdiffc >>
rect 48 441 82 475
rect 153 449 187 483
rect 258 423 292 457
rect 344 449 378 483
rect 438 449 472 483
rect 524 449 558 483
rect 657 423 691 457
<< poly >>
rect 82 605 427 621
rect 82 571 98 605
rect 132 591 427 605
rect 132 571 148 591
rect 82 555 148 571
rect 93 487 123 513
rect 217 495 247 521
rect 303 495 333 521
rect 397 495 427 591
rect 483 495 513 521
rect 616 495 646 521
rect 93 323 123 403
rect 217 323 247 411
rect 303 323 333 411
rect 73 307 139 323
rect 73 273 89 307
rect 123 273 139 307
rect 73 257 139 273
rect 181 307 247 323
rect 181 273 197 307
rect 231 273 247 307
rect 181 257 247 273
rect 80 235 110 257
rect 217 235 247 257
rect 289 307 355 323
rect 289 273 305 307
rect 339 273 355 307
rect 289 257 355 273
rect 289 235 319 257
rect 397 235 427 411
rect 483 378 513 411
rect 483 362 558 378
rect 483 328 508 362
rect 542 328 558 362
rect 483 311 558 328
rect 469 281 558 311
rect 616 307 646 411
rect 469 235 499 281
rect 616 277 686 307
rect 656 233 686 277
rect 611 217 686 233
rect 611 183 627 217
rect 661 183 686 217
rect 611 167 686 183
rect 80 125 110 151
rect 217 125 247 151
rect 289 125 319 151
rect 397 125 427 151
rect 469 125 499 151
rect 656 131 686 167
rect 656 21 686 47
<< polycont >>
rect 98 571 132 605
rect 89 273 123 307
rect 197 273 231 307
rect 305 273 339 307
rect 508 328 542 362
rect 627 183 661 217
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 44 605 148 615
rect 44 571 98 605
rect 132 571 148 605
rect 44 555 148 571
rect 44 479 110 555
rect 182 521 220 649
rect 19 475 110 479
rect 19 441 48 475
rect 82 441 110 475
rect 19 437 110 441
rect 149 483 220 521
rect 149 449 153 483
rect 187 479 220 483
rect 344 483 378 649
rect 187 449 191 479
rect 19 206 53 437
rect 149 433 191 449
rect 254 457 296 473
rect 254 423 258 457
rect 292 423 296 457
rect 344 433 378 449
rect 415 483 472 508
rect 415 449 438 483
rect 254 397 296 423
rect 415 397 472 449
rect 508 483 574 649
rect 508 449 524 483
rect 558 449 574 483
rect 508 445 574 449
rect 641 457 707 461
rect 254 363 472 397
rect 641 423 657 457
rect 691 423 707 457
rect 641 378 707 423
rect 89 307 161 350
rect 123 273 161 307
rect 89 242 161 273
rect 197 307 257 323
rect 231 273 257 307
rect 197 257 257 273
rect 19 202 85 206
rect 19 168 35 202
rect 69 168 85 202
rect 19 164 85 168
rect 121 197 187 201
rect 121 163 137 197
rect 171 163 187 197
rect 121 17 187 163
rect 223 84 257 257
rect 305 307 353 323
rect 339 273 353 307
rect 305 84 353 273
rect 415 243 472 363
rect 508 362 735 378
rect 542 328 735 362
rect 508 312 735 328
rect 415 227 571 243
rect 415 209 533 227
rect 529 193 533 209
rect 567 193 571 227
rect 529 177 571 193
rect 607 217 661 276
rect 607 183 627 217
rect 607 158 661 183
rect 697 115 735 312
rect 595 93 661 97
rect 595 59 611 93
rect 645 59 661 93
rect 731 81 735 115
rect 697 65 735 81
rect 595 17 661 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4bb_m
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5675108
string GDS_START 5667942
<< end >>
