magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
rect 727 311 1591 331
rect 1256 297 1591 311
<< pwell >>
rect 777 221 1145 265
rect 1623 221 2015 242
rect 1 211 427 219
rect 777 211 2015 221
rect 1 49 2015 211
rect 0 0 2016 49
<< scnmos >>
rect 84 109 114 193
rect 156 109 186 193
rect 242 109 272 193
rect 314 109 344 193
rect 540 101 570 185
rect 618 101 648 185
rect 930 155 960 239
rect 1032 155 1062 239
rect 1134 111 1164 195
rect 1220 111 1250 195
rect 1318 111 1348 195
rect 1404 111 1434 195
rect 1604 89 1634 173
rect 1699 132 1729 216
rect 1830 132 1860 216
rect 1902 132 1932 216
<< scpmoshvt >>
rect 109 409 159 609
rect 215 409 265 609
rect 597 367 647 567
rect 836 347 886 547
rect 1008 347 1058 547
rect 1114 347 1164 547
rect 1220 347 1270 547
rect 1342 333 1392 533
rect 1448 333 1498 533
rect 1724 401 1774 601
rect 1830 401 1880 601
<< ndiff >>
rect 27 168 84 193
rect 27 134 39 168
rect 73 134 84 168
rect 27 109 84 134
rect 114 109 156 193
rect 186 168 242 193
rect 186 134 197 168
rect 231 134 242 168
rect 186 109 242 134
rect 272 109 314 193
rect 344 177 401 193
rect 344 143 355 177
rect 389 143 401 177
rect 344 109 401 143
rect 483 147 540 185
rect 483 113 495 147
rect 529 113 540 147
rect 483 101 540 113
rect 570 101 618 185
rect 648 173 721 185
rect 648 139 675 173
rect 709 139 721 173
rect 648 101 721 139
rect 803 155 930 239
rect 960 227 1032 239
rect 960 193 971 227
rect 1005 193 1032 227
rect 960 155 1032 193
rect 1062 227 1119 239
rect 1062 193 1073 227
rect 1107 195 1119 227
rect 1107 193 1134 195
rect 1062 155 1134 193
rect 803 127 881 155
rect 803 93 815 127
rect 849 93 881 127
rect 1084 111 1134 155
rect 1164 178 1220 195
rect 1164 144 1175 178
rect 1209 144 1220 178
rect 1164 111 1220 144
rect 1250 170 1318 195
rect 1250 136 1261 170
rect 1295 136 1318 170
rect 1250 111 1318 136
rect 1348 170 1404 195
rect 1348 136 1359 170
rect 1393 136 1404 170
rect 1348 111 1404 136
rect 1434 178 1491 195
rect 1434 144 1445 178
rect 1479 144 1491 178
rect 1649 173 1699 216
rect 1434 111 1491 144
rect 1547 158 1604 173
rect 1547 124 1559 158
rect 1593 124 1604 158
rect 803 81 881 93
rect 1547 89 1604 124
rect 1634 132 1699 173
rect 1729 200 1830 216
rect 1729 166 1785 200
rect 1819 166 1830 200
rect 1729 132 1830 166
rect 1860 132 1902 216
rect 1932 191 1989 216
rect 1932 157 1943 191
rect 1977 157 1989 191
rect 1932 132 1989 157
rect 1634 89 1684 132
<< pdiff >>
rect 52 597 109 609
rect 52 563 64 597
rect 98 563 109 597
rect 52 526 109 563
rect 52 492 64 526
rect 98 492 109 526
rect 52 455 109 492
rect 52 421 64 455
rect 98 421 109 455
rect 52 409 109 421
rect 159 597 215 609
rect 159 563 170 597
rect 204 563 215 597
rect 159 526 215 563
rect 159 492 170 526
rect 204 492 215 526
rect 159 455 215 492
rect 159 421 170 455
rect 204 421 215 455
rect 159 409 215 421
rect 265 597 322 609
rect 265 563 276 597
rect 310 563 322 597
rect 265 526 322 563
rect 265 492 276 526
rect 310 492 322 526
rect 265 455 322 492
rect 265 421 276 455
rect 310 421 322 455
rect 265 409 322 421
rect 524 569 582 581
rect 524 535 536 569
rect 570 567 582 569
rect 570 535 597 567
rect 524 367 597 535
rect 647 413 704 567
rect 647 379 658 413
rect 692 379 704 413
rect 647 367 704 379
rect 763 553 821 565
rect 763 519 775 553
rect 809 547 821 553
rect 809 519 836 547
rect 763 347 836 519
rect 886 527 1008 547
rect 886 493 897 527
rect 931 493 1008 527
rect 886 393 1008 493
rect 886 359 897 393
rect 931 359 1008 393
rect 886 347 1008 359
rect 1058 503 1114 547
rect 1058 469 1069 503
rect 1103 469 1114 503
rect 1058 347 1114 469
rect 1164 393 1220 547
rect 1164 359 1175 393
rect 1209 359 1220 393
rect 1164 347 1220 359
rect 1270 535 1327 547
rect 1270 501 1281 535
rect 1315 533 1327 535
rect 1315 501 1342 533
rect 1270 347 1342 501
rect 1292 333 1342 347
rect 1392 379 1448 533
rect 1392 345 1403 379
rect 1437 345 1448 379
rect 1392 333 1448 345
rect 1498 518 1555 533
rect 1498 484 1509 518
rect 1543 484 1555 518
rect 1498 333 1555 484
rect 1667 589 1724 601
rect 1667 555 1679 589
rect 1713 555 1724 589
rect 1667 518 1724 555
rect 1667 484 1679 518
rect 1713 484 1724 518
rect 1667 447 1724 484
rect 1667 413 1679 447
rect 1713 413 1724 447
rect 1667 401 1724 413
rect 1774 589 1830 601
rect 1774 555 1785 589
rect 1819 555 1830 589
rect 1774 518 1830 555
rect 1774 484 1785 518
rect 1819 484 1830 518
rect 1774 447 1830 484
rect 1774 413 1785 447
rect 1819 413 1830 447
rect 1774 401 1830 413
rect 1880 589 1937 601
rect 1880 555 1891 589
rect 1925 555 1937 589
rect 1880 518 1937 555
rect 1880 484 1891 518
rect 1925 484 1937 518
rect 1880 447 1937 484
rect 1880 413 1891 447
rect 1925 413 1937 447
rect 1880 401 1937 413
<< ndiffc >>
rect 39 134 73 168
rect 197 134 231 168
rect 355 143 389 177
rect 495 113 529 147
rect 675 139 709 173
rect 971 193 1005 227
rect 1073 193 1107 227
rect 815 93 849 127
rect 1175 144 1209 178
rect 1261 136 1295 170
rect 1359 136 1393 170
rect 1445 144 1479 178
rect 1559 124 1593 158
rect 1785 166 1819 200
rect 1943 157 1977 191
<< pdiffc >>
rect 64 563 98 597
rect 64 492 98 526
rect 64 421 98 455
rect 170 563 204 597
rect 170 492 204 526
rect 170 421 204 455
rect 276 563 310 597
rect 276 492 310 526
rect 276 421 310 455
rect 536 535 570 569
rect 658 379 692 413
rect 775 519 809 553
rect 897 493 931 527
rect 897 359 931 393
rect 1069 469 1103 503
rect 1175 359 1209 393
rect 1281 501 1315 535
rect 1403 345 1437 379
rect 1509 484 1543 518
rect 1679 555 1713 589
rect 1679 484 1713 518
rect 1679 413 1713 447
rect 1785 555 1819 589
rect 1785 484 1819 518
rect 1785 413 1819 447
rect 1891 555 1925 589
rect 1891 484 1925 518
rect 1891 413 1925 447
<< poly >>
rect 109 609 159 635
rect 215 609 265 635
rect 597 615 1270 645
rect 597 567 647 615
rect 1008 573 1038 615
rect 109 369 159 409
rect 215 381 265 409
rect 84 353 159 369
rect 84 319 109 353
rect 143 333 159 353
rect 235 367 265 381
rect 836 547 886 573
rect 1008 547 1058 573
rect 1114 547 1164 573
rect 1220 547 1270 615
rect 1342 607 1640 637
rect 235 351 344 367
rect 143 319 186 333
rect 84 303 186 319
rect 84 193 114 303
rect 156 193 186 303
rect 235 317 251 351
rect 285 317 344 351
rect 597 335 647 367
rect 1342 533 1392 607
rect 1448 533 1498 559
rect 235 283 344 317
rect 235 249 251 283
rect 285 249 344 283
rect 235 233 344 249
rect 242 193 272 233
rect 314 193 344 233
rect 540 319 648 335
rect 540 285 556 319
rect 590 285 648 319
rect 836 315 886 347
rect 1008 332 1058 347
rect 540 269 648 285
rect 540 185 570 269
rect 618 185 648 269
rect 700 299 960 315
rect 1008 302 1062 332
rect 700 265 716 299
rect 750 285 960 299
rect 750 265 766 285
rect 700 249 766 265
rect 84 83 114 109
rect 156 83 186 109
rect 242 83 272 109
rect 314 83 344 109
rect 540 75 570 101
rect 618 75 648 101
rect 736 66 766 249
rect 930 239 960 285
rect 1032 239 1062 302
rect 1114 254 1164 347
rect 1134 195 1164 254
rect 1220 302 1270 347
rect 1610 369 1640 607
rect 1724 601 1774 627
rect 1830 601 1880 627
rect 1610 353 1676 369
rect 1342 318 1392 333
rect 1220 195 1250 302
rect 1318 288 1392 318
rect 1318 195 1348 288
rect 1448 240 1498 333
rect 1610 319 1626 353
rect 1660 319 1676 353
rect 1610 303 1676 319
rect 1724 261 1774 401
rect 1546 245 1774 261
rect 1546 240 1562 245
rect 1404 211 1562 240
rect 1596 231 1774 245
rect 1830 290 1880 401
rect 1596 211 1634 231
rect 1699 216 1729 231
rect 1830 216 1860 290
rect 1902 216 1932 242
rect 1404 210 1634 211
rect 1404 195 1434 210
rect 1546 195 1634 210
rect 930 129 960 155
rect 1032 129 1062 155
rect 1604 173 1634 195
rect 1134 66 1164 111
rect 1220 85 1250 111
rect 1318 85 1348 111
rect 1404 85 1434 111
rect 1699 106 1729 132
rect 1830 110 1860 132
rect 1902 110 1932 132
rect 1771 94 1932 110
rect 736 36 1164 66
rect 1604 63 1634 89
rect 1771 60 1787 94
rect 1821 80 1932 94
rect 1821 60 1860 80
rect 1771 44 1860 60
<< polycont >>
rect 109 319 143 353
rect 251 317 285 351
rect 251 249 285 283
rect 556 285 590 319
rect 716 265 750 299
rect 1626 319 1660 353
rect 1562 211 1596 245
rect 1787 60 1821 94
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 597 114 613
rect 23 563 64 597
rect 98 563 114 597
rect 23 526 114 563
rect 23 492 64 526
rect 98 492 114 526
rect 23 455 114 492
rect 23 421 64 455
rect 98 421 114 455
rect 23 405 114 421
rect 154 597 220 649
rect 154 563 170 597
rect 204 563 220 597
rect 154 526 220 563
rect 154 492 170 526
rect 204 492 220 526
rect 154 455 220 492
rect 154 421 170 455
rect 204 421 220 455
rect 154 405 220 421
rect 260 597 326 613
rect 260 563 276 597
rect 310 563 326 597
rect 260 526 326 563
rect 260 492 276 526
rect 310 492 326 526
rect 520 569 586 649
rect 520 535 536 569
rect 570 535 586 569
rect 520 519 586 535
rect 759 579 1613 613
rect 759 553 825 579
rect 759 519 775 553
rect 809 519 825 553
rect 881 527 947 543
rect 260 483 326 492
rect 881 493 897 527
rect 931 493 947 527
rect 881 483 947 493
rect 260 455 947 483
rect 260 421 276 455
rect 310 449 947 455
rect 310 421 373 449
rect 260 405 373 421
rect 23 267 57 405
rect 93 353 167 369
rect 93 319 109 353
rect 143 319 167 353
rect 93 303 167 319
rect 235 351 301 367
rect 235 317 251 351
rect 285 317 301 351
rect 235 283 301 317
rect 235 267 251 283
rect 23 249 251 267
rect 285 249 301 283
rect 23 233 301 249
rect 23 168 89 233
rect 23 134 39 168
rect 73 134 89 168
rect 23 105 89 134
rect 181 168 231 197
rect 181 134 197 168
rect 181 17 231 134
rect 267 87 301 233
rect 339 197 373 405
rect 642 379 658 413
rect 692 379 708 413
rect 642 363 708 379
rect 409 319 606 356
rect 409 285 556 319
rect 590 285 606 319
rect 409 269 606 285
rect 659 315 708 363
rect 881 393 947 449
rect 881 359 897 393
rect 931 359 947 393
rect 983 393 1017 579
rect 1053 503 1119 543
rect 1053 469 1069 503
rect 1103 469 1119 503
rect 1265 535 1331 579
rect 1265 501 1281 535
rect 1315 501 1331 535
rect 1493 518 1543 537
rect 1493 499 1509 518
rect 1053 465 1119 469
rect 1367 484 1509 499
rect 1367 465 1543 484
rect 1053 431 1401 465
rect 1053 429 1119 431
rect 983 359 1123 393
rect 659 299 766 315
rect 659 265 716 299
rect 750 265 766 299
rect 659 249 766 265
rect 881 283 947 359
rect 881 249 1021 283
rect 425 199 615 233
rect 339 177 389 197
rect 339 143 355 177
rect 339 123 389 143
rect 425 87 459 199
rect 267 53 459 87
rect 495 147 545 163
rect 529 113 545 147
rect 495 17 545 113
rect 581 87 615 199
rect 659 173 709 249
rect 955 227 1021 249
rect 659 139 675 173
rect 659 123 709 139
rect 745 179 919 213
rect 955 193 971 227
rect 1005 193 1021 227
rect 1057 227 1123 359
rect 1057 193 1073 227
rect 1107 193 1123 227
rect 1159 359 1175 393
rect 1209 359 1225 393
rect 745 87 779 179
rect 885 157 919 179
rect 1159 178 1225 359
rect 1159 157 1175 178
rect 885 144 1175 157
rect 1209 144 1225 178
rect 581 53 779 87
rect 815 127 849 143
rect 885 123 1225 144
rect 1261 170 1295 431
rect 1579 429 1613 579
rect 1473 395 1613 429
rect 1663 589 1729 605
rect 1663 555 1679 589
rect 1713 555 1729 589
rect 1663 518 1729 555
rect 1663 484 1679 518
rect 1713 484 1729 518
rect 1663 447 1729 484
rect 1663 413 1679 447
rect 1713 413 1729 447
rect 815 87 849 93
rect 1261 87 1295 136
rect 815 53 1295 87
rect 1343 379 1437 395
rect 1343 345 1403 379
rect 1343 329 1437 345
rect 1343 170 1393 329
rect 1473 199 1507 395
rect 1663 359 1729 413
rect 1769 589 1835 649
rect 1769 555 1785 589
rect 1819 555 1835 589
rect 1769 518 1835 555
rect 1769 484 1785 518
rect 1819 484 1835 518
rect 1769 447 1835 484
rect 1769 413 1785 447
rect 1819 413 1835 447
rect 1769 397 1835 413
rect 1875 589 1941 605
rect 1875 555 1891 589
rect 1925 578 1941 589
rect 1925 555 1993 578
rect 1875 518 1993 555
rect 1875 484 1891 518
rect 1925 484 1993 518
rect 1875 447 1993 484
rect 1875 413 1891 447
rect 1925 413 1993 447
rect 1610 353 1729 359
rect 1610 319 1626 353
rect 1660 319 1729 353
rect 1610 312 1729 319
rect 1343 136 1359 170
rect 1343 87 1393 136
rect 1429 178 1507 199
rect 1546 245 1612 276
rect 1546 211 1562 245
rect 1596 211 1612 245
rect 1546 195 1612 211
rect 1429 144 1445 178
rect 1479 144 1507 178
rect 1695 159 1729 312
rect 1875 236 1993 413
rect 1429 123 1507 144
rect 1543 158 1729 159
rect 1543 124 1559 158
rect 1593 124 1729 158
rect 1769 200 1835 220
rect 1769 166 1785 200
rect 1819 180 1835 200
rect 1943 191 1993 236
rect 1819 166 1907 180
rect 1769 146 1907 166
rect 1543 123 1729 124
rect 1771 94 1837 110
rect 1771 87 1787 94
rect 1343 60 1787 87
rect 1821 60 1837 94
rect 1343 53 1837 60
rect 1873 17 1907 146
rect 1977 157 1993 191
rect 1943 128 1993 157
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xnor3_lp
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1951 390 1985 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1951 464 1985 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1951 538 1985 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 746080
string GDS_START 733364
<< end >>
