magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 64 162 661 241
rect 64 49 851 162
rect 0 0 864 49
<< scnmos >>
rect 147 131 177 215
rect 264 47 294 215
rect 336 47 366 215
rect 444 47 474 215
rect 552 47 582 215
rect 742 52 772 136
<< scpmoshvt >>
rect 106 367 136 451
rect 264 367 294 619
rect 350 367 380 619
rect 466 367 496 619
rect 552 367 582 619
rect 692 367 722 451
<< ndiff >>
rect 90 202 147 215
rect 90 168 98 202
rect 132 168 147 202
rect 90 131 147 168
rect 177 131 264 215
rect 211 121 264 131
rect 211 87 219 121
rect 253 87 264 121
rect 211 47 264 87
rect 294 47 336 215
rect 366 47 444 215
rect 474 47 552 215
rect 582 203 635 215
rect 582 169 593 203
rect 627 169 635 203
rect 582 93 635 169
rect 582 59 593 93
rect 627 59 635 93
rect 582 47 635 59
rect 689 111 742 136
rect 689 77 697 111
rect 731 77 742 111
rect 689 52 742 77
rect 772 111 825 136
rect 772 77 783 111
rect 817 77 825 111
rect 772 52 825 77
<< pdiff >>
rect 211 607 264 619
rect 211 573 219 607
rect 253 573 264 607
rect 211 519 264 573
rect 211 485 219 519
rect 253 485 264 519
rect 211 451 264 485
rect 49 426 106 451
rect 49 392 57 426
rect 91 392 106 426
rect 49 367 106 392
rect 136 434 264 451
rect 136 400 199 434
rect 233 400 264 434
rect 136 367 264 400
rect 294 599 350 619
rect 294 565 305 599
rect 339 565 350 599
rect 294 502 350 565
rect 294 468 305 502
rect 339 468 350 502
rect 294 413 350 468
rect 294 379 305 413
rect 339 379 350 413
rect 294 367 350 379
rect 380 607 466 619
rect 380 573 406 607
rect 440 573 466 607
rect 380 524 466 573
rect 380 490 406 524
rect 440 490 466 524
rect 380 440 466 490
rect 380 406 406 440
rect 440 406 466 440
rect 380 367 466 406
rect 496 599 552 619
rect 496 565 507 599
rect 541 565 552 599
rect 496 507 552 565
rect 496 473 507 507
rect 541 473 552 507
rect 496 413 552 473
rect 496 379 507 413
rect 541 379 552 413
rect 496 367 552 379
rect 582 607 646 619
rect 582 573 598 607
rect 632 573 646 607
rect 582 514 646 573
rect 582 480 598 514
rect 632 480 646 514
rect 582 451 646 480
rect 582 430 692 451
rect 582 396 645 430
rect 679 396 692 430
rect 582 367 692 396
rect 722 427 775 451
rect 722 393 733 427
rect 767 393 775 427
rect 722 367 775 393
<< ndiffc >>
rect 98 168 132 202
rect 219 87 253 121
rect 593 169 627 203
rect 593 59 627 93
rect 697 77 731 111
rect 783 77 817 111
<< pdiffc >>
rect 219 573 253 607
rect 219 485 253 519
rect 57 392 91 426
rect 199 400 233 434
rect 305 565 339 599
rect 305 468 339 502
rect 305 379 339 413
rect 406 573 440 607
rect 406 490 440 524
rect 406 406 440 440
rect 507 565 541 599
rect 507 473 541 507
rect 507 379 541 413
rect 598 573 632 607
rect 598 480 632 514
rect 645 396 679 430
rect 733 393 767 427
<< poly >>
rect 264 619 294 645
rect 350 619 380 645
rect 466 619 496 645
rect 552 619 582 645
rect 106 451 136 477
rect 692 451 722 477
rect 106 308 136 367
rect 264 308 294 367
rect 106 292 177 308
rect 106 258 127 292
rect 161 258 177 292
rect 106 242 177 258
rect 219 292 294 308
rect 350 303 380 367
rect 466 304 496 367
rect 552 335 582 367
rect 552 319 650 335
rect 219 258 235 292
rect 269 258 294 292
rect 219 242 294 258
rect 147 215 177 242
rect 264 215 294 242
rect 336 287 402 303
rect 336 253 352 287
rect 386 253 402 287
rect 336 237 402 253
rect 444 288 510 304
rect 444 254 460 288
rect 494 254 510 288
rect 444 238 510 254
rect 552 285 600 319
rect 634 285 650 319
rect 552 269 650 285
rect 692 292 722 367
rect 692 276 772 292
rect 336 215 366 237
rect 444 215 474 238
rect 552 215 582 269
rect 692 262 722 276
rect 706 242 722 262
rect 756 242 772 276
rect 147 105 177 131
rect 706 208 772 242
rect 706 174 722 208
rect 756 174 772 208
rect 706 158 772 174
rect 742 136 772 158
rect 264 21 294 47
rect 336 21 366 47
rect 444 21 474 47
rect 552 21 582 47
rect 742 26 772 52
<< polycont >>
rect 127 258 161 292
rect 235 258 269 292
rect 352 253 386 287
rect 460 254 494 288
rect 600 285 634 319
rect 722 242 756 276
rect 722 174 756 208
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 195 607 269 649
rect 41 426 93 442
rect 41 392 57 426
rect 91 392 93 426
rect 41 206 93 392
rect 127 292 161 595
rect 195 573 219 607
rect 253 573 269 607
rect 195 519 269 573
rect 195 485 219 519
rect 253 485 269 519
rect 195 434 269 485
rect 195 400 199 434
rect 233 400 269 434
rect 195 384 269 400
rect 303 599 355 615
rect 303 565 305 599
rect 339 565 355 599
rect 303 502 355 565
rect 303 468 305 502
rect 339 468 355 502
rect 303 413 355 468
rect 303 379 305 413
rect 339 379 355 413
rect 390 607 456 649
rect 390 573 406 607
rect 440 573 456 607
rect 390 524 456 573
rect 390 490 406 524
rect 440 490 456 524
rect 390 440 456 490
rect 390 406 406 440
rect 440 406 456 440
rect 491 599 564 615
rect 491 565 507 599
rect 541 565 564 599
rect 491 507 564 565
rect 491 473 507 507
rect 541 473 564 507
rect 491 413 564 473
rect 303 372 355 379
rect 491 379 507 413
rect 541 379 564 413
rect 598 607 695 649
rect 632 573 695 607
rect 598 514 695 573
rect 632 480 695 514
rect 598 430 695 480
rect 598 396 645 430
rect 679 396 695 430
rect 598 380 695 396
rect 729 427 783 443
rect 729 393 733 427
rect 767 393 783 427
rect 491 372 564 379
rect 127 240 161 258
rect 201 292 269 350
rect 303 338 564 372
rect 729 346 783 393
rect 201 258 235 292
rect 201 242 269 258
rect 303 287 402 304
rect 303 253 352 287
rect 386 253 402 287
rect 303 240 402 253
rect 444 288 496 304
rect 444 254 460 288
rect 494 254 496 288
rect 444 206 496 254
rect 41 202 496 206
rect 41 168 98 202
rect 132 168 496 202
rect 41 164 496 168
rect 530 222 564 338
rect 598 319 842 346
rect 598 285 600 319
rect 634 312 842 319
rect 634 285 650 312
rect 598 269 650 285
rect 684 276 772 278
rect 684 242 722 276
rect 756 242 772 276
rect 530 203 650 222
rect 530 169 593 203
rect 627 169 650 203
rect 203 121 269 130
rect 203 87 219 121
rect 253 87 269 121
rect 203 17 269 87
rect 530 93 650 169
rect 684 208 772 242
rect 684 174 722 208
rect 756 174 772 208
rect 684 161 772 174
rect 806 127 842 312
rect 530 59 593 93
rect 627 59 650 93
rect 530 51 650 59
rect 684 111 739 127
rect 684 77 697 111
rect 731 77 739 111
rect 684 17 739 77
rect 773 111 842 127
rect 773 77 783 111
rect 817 77 842 111
rect 773 61 842 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4bb_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5682852
string GDS_START 5675166
<< end >>
