magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 332 1478 704
rect 934 327 1148 332
<< pwell >>
rect 1 248 315 256
rect 769 248 1138 249
rect 1 233 562 248
rect 769 233 1439 248
rect 1 49 1439 233
rect 0 0 1440 49
<< scnmos >>
rect 84 120 114 230
rect 202 82 232 230
rect 456 74 486 222
rect 628 79 658 207
rect 706 79 736 207
rect 845 139 875 223
rect 923 139 953 223
rect 1025 75 1055 223
rect 1223 74 1253 222
rect 1321 74 1351 222
<< scpmoshvt >>
rect 116 424 146 592
rect 226 424 256 592
rect 428 392 458 560
rect 555 392 585 592
rect 639 392 669 592
rect 761 503 791 587
rect 845 503 875 587
rect 1023 363 1053 587
rect 1225 368 1255 592
rect 1324 368 1354 592
<< ndiff >>
rect 27 188 84 230
rect 27 154 39 188
rect 73 154 84 188
rect 27 120 84 154
rect 114 120 202 230
rect 129 82 202 120
rect 232 218 289 230
rect 232 184 243 218
rect 277 184 289 218
rect 232 82 289 184
rect 399 189 456 222
rect 399 155 411 189
rect 445 155 456 189
rect 129 48 141 82
rect 175 48 187 82
rect 399 74 456 155
rect 486 207 536 222
rect 795 207 845 223
rect 486 195 628 207
rect 486 161 579 195
rect 613 161 628 195
rect 486 125 628 161
rect 486 91 579 125
rect 613 91 628 125
rect 486 79 628 91
rect 658 79 706 207
rect 736 195 845 207
rect 736 161 773 195
rect 807 161 845 195
rect 736 139 845 161
rect 875 139 923 223
rect 953 195 1025 223
rect 953 161 980 195
rect 1014 161 1025 195
rect 953 139 1025 161
rect 736 79 786 139
rect 968 120 1025 139
rect 486 74 536 79
rect 968 86 980 120
rect 1014 86 1025 120
rect 968 75 1025 86
rect 1055 209 1112 223
rect 1055 175 1066 209
rect 1100 175 1112 209
rect 1055 121 1112 175
rect 1055 87 1066 121
rect 1100 87 1112 121
rect 1055 75 1112 87
rect 1166 209 1223 222
rect 1166 175 1178 209
rect 1212 175 1223 209
rect 1166 120 1223 175
rect 1166 86 1178 120
rect 1212 86 1223 120
rect 1166 74 1223 86
rect 1253 209 1321 222
rect 1253 175 1265 209
rect 1299 175 1321 209
rect 1253 120 1321 175
rect 1253 86 1265 120
rect 1299 86 1321 120
rect 1253 74 1321 86
rect 1351 210 1413 222
rect 1351 176 1367 210
rect 1401 176 1413 210
rect 1351 120 1413 176
rect 1351 86 1367 120
rect 1401 86 1413 120
rect 1351 74 1413 86
rect 129 36 187 48
<< pdiff >>
rect 476 606 537 618
rect 57 580 116 592
rect 57 546 69 580
rect 103 546 116 580
rect 57 470 116 546
rect 57 436 69 470
rect 103 436 116 470
rect 57 424 116 436
rect 146 580 226 592
rect 146 546 169 580
rect 203 546 226 580
rect 146 496 226 546
rect 146 462 169 496
rect 203 462 226 496
rect 146 424 226 462
rect 256 580 315 592
rect 256 546 269 580
rect 303 546 315 580
rect 476 572 489 606
rect 523 592 537 606
rect 523 572 555 592
rect 476 560 555 572
rect 256 470 315 546
rect 256 436 269 470
rect 303 436 315 470
rect 256 424 315 436
rect 369 438 428 560
rect 369 404 381 438
rect 415 404 428 438
rect 369 392 428 404
rect 458 392 555 560
rect 585 392 639 592
rect 669 587 722 592
rect 669 547 761 587
rect 669 513 689 547
rect 723 513 761 547
rect 669 503 761 513
rect 791 503 845 587
rect 875 575 1023 587
rect 875 541 888 575
rect 922 541 975 575
rect 1009 541 1023 575
rect 875 503 1023 541
rect 669 462 743 503
rect 669 428 689 462
rect 723 428 743 462
rect 669 392 743 428
rect 970 363 1023 503
rect 1053 575 1112 587
rect 1053 541 1066 575
rect 1100 541 1112 575
rect 1053 492 1112 541
rect 1053 458 1066 492
rect 1100 458 1112 492
rect 1053 409 1112 458
rect 1053 375 1066 409
rect 1100 375 1112 409
rect 1053 363 1112 375
rect 1166 580 1225 592
rect 1166 546 1178 580
rect 1212 546 1225 580
rect 1166 497 1225 546
rect 1166 463 1178 497
rect 1212 463 1225 497
rect 1166 414 1225 463
rect 1166 380 1178 414
rect 1212 380 1225 414
rect 1166 368 1225 380
rect 1255 434 1324 592
rect 1255 400 1272 434
rect 1306 400 1324 434
rect 1255 368 1324 400
rect 1354 580 1413 592
rect 1354 546 1367 580
rect 1401 546 1413 580
rect 1354 497 1413 546
rect 1354 463 1367 497
rect 1401 463 1413 497
rect 1354 414 1413 463
rect 1354 380 1367 414
rect 1401 380 1413 414
rect 1354 368 1413 380
<< ndiffc >>
rect 39 154 73 188
rect 243 184 277 218
rect 411 155 445 189
rect 141 48 175 82
rect 579 161 613 195
rect 579 91 613 125
rect 773 161 807 195
rect 980 161 1014 195
rect 980 86 1014 120
rect 1066 175 1100 209
rect 1066 87 1100 121
rect 1178 175 1212 209
rect 1178 86 1212 120
rect 1265 175 1299 209
rect 1265 86 1299 120
rect 1367 176 1401 210
rect 1367 86 1401 120
<< pdiffc >>
rect 69 546 103 580
rect 69 436 103 470
rect 169 546 203 580
rect 169 462 203 496
rect 269 546 303 580
rect 489 572 523 606
rect 269 436 303 470
rect 381 404 415 438
rect 689 513 723 547
rect 888 541 922 575
rect 975 541 1009 575
rect 689 428 723 462
rect 1066 541 1100 575
rect 1066 458 1100 492
rect 1066 375 1100 409
rect 1178 546 1212 580
rect 1178 463 1212 497
rect 1178 380 1212 414
rect 1272 400 1306 434
rect 1367 546 1401 580
rect 1367 463 1401 497
rect 1367 380 1401 414
<< poly >>
rect 116 592 146 618
rect 226 592 256 618
rect 428 560 458 586
rect 555 592 585 618
rect 639 592 669 618
rect 116 409 146 424
rect 226 409 256 424
rect 113 326 149 409
rect 223 356 259 409
rect 761 587 791 613
rect 845 587 875 613
rect 1023 587 1053 613
rect 1225 592 1255 618
rect 1324 592 1354 618
rect 761 488 791 503
rect 845 488 875 503
rect 428 377 458 392
rect 555 377 585 392
rect 639 377 669 392
rect 25 310 149 326
rect 25 276 41 310
rect 75 276 149 310
rect 197 340 263 356
rect 197 306 213 340
rect 247 306 263 340
rect 197 290 263 306
rect 311 338 377 354
rect 311 304 327 338
rect 361 304 377 338
rect 25 260 149 276
rect 84 230 114 260
rect 202 230 232 290
rect 311 270 377 304
rect 311 236 327 270
rect 361 267 377 270
rect 425 267 461 377
rect 552 326 588 377
rect 636 360 672 377
rect 758 363 794 488
rect 842 471 878 488
rect 842 455 953 471
rect 842 421 888 455
rect 922 421 953 455
rect 842 405 953 421
rect 636 344 702 360
rect 528 310 594 326
rect 528 276 544 310
rect 578 276 594 310
rect 636 310 652 344
rect 686 310 702 344
rect 636 294 702 310
rect 750 347 870 363
rect 750 313 820 347
rect 854 313 870 347
rect 750 297 870 313
rect 361 237 486 267
rect 528 252 594 276
rect 750 252 780 297
rect 361 236 377 237
rect 84 94 114 120
rect 311 202 377 236
rect 456 222 486 237
rect 564 222 658 252
rect 311 168 327 202
rect 361 168 377 202
rect 311 152 377 168
rect 202 56 232 82
rect 628 207 658 222
rect 706 222 780 252
rect 845 223 875 249
rect 923 223 953 405
rect 1023 348 1053 363
rect 1225 353 1255 368
rect 1324 353 1354 368
rect 1020 325 1056 348
rect 1222 325 1258 353
rect 1321 325 1357 353
rect 1001 309 1067 325
rect 1001 275 1017 309
rect 1051 275 1067 309
rect 1001 259 1067 275
rect 1115 309 1357 325
rect 1115 275 1131 309
rect 1165 275 1199 309
rect 1233 289 1357 309
rect 1233 275 1351 289
rect 1115 259 1351 275
rect 1025 223 1055 259
rect 706 207 736 222
rect 845 117 875 139
rect 809 101 875 117
rect 923 113 953 139
rect 456 48 486 74
rect 628 53 658 79
rect 706 53 736 79
rect 809 67 825 101
rect 859 67 875 101
rect 1223 222 1253 259
rect 1321 222 1351 259
rect 809 51 875 67
rect 1025 49 1055 75
rect 1223 48 1253 74
rect 1321 48 1351 74
<< polycont >>
rect 41 276 75 310
rect 213 306 247 340
rect 327 304 361 338
rect 327 236 361 270
rect 888 421 922 455
rect 544 276 578 310
rect 652 310 686 344
rect 820 313 854 347
rect 327 168 361 202
rect 1017 275 1051 309
rect 1131 275 1165 309
rect 1199 275 1233 309
rect 825 67 859 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 53 580 119 596
rect 53 546 69 580
rect 103 546 119 580
rect 53 470 119 546
rect 53 436 69 470
rect 103 436 119 470
rect 153 580 219 649
rect 472 606 541 649
rect 153 546 169 580
rect 203 546 219 580
rect 153 496 219 546
rect 153 462 169 496
rect 203 462 219 496
rect 153 458 219 462
rect 253 580 331 596
rect 253 546 269 580
rect 303 546 331 580
rect 472 572 489 606
rect 523 572 541 606
rect 472 556 541 572
rect 575 581 838 615
rect 253 522 331 546
rect 575 522 609 581
rect 253 488 609 522
rect 666 513 689 547
rect 723 513 770 547
rect 253 470 331 488
rect 53 424 119 436
rect 253 436 269 470
rect 303 436 331 470
rect 666 462 770 513
rect 53 390 159 424
rect 253 420 331 436
rect 25 310 91 356
rect 25 276 41 310
rect 75 276 91 310
rect 25 260 91 276
rect 125 226 159 390
rect 197 340 263 356
rect 197 306 213 340
rect 247 306 263 340
rect 197 290 263 306
rect 297 354 331 420
rect 365 438 445 454
rect 365 404 381 438
rect 415 404 445 438
rect 666 428 689 462
rect 723 428 770 462
rect 365 394 445 404
rect 365 388 702 394
rect 411 360 702 388
rect 297 338 377 354
rect 297 304 327 338
rect 361 304 377 338
rect 297 270 377 304
rect 297 236 327 270
rect 361 236 377 270
rect 297 234 377 236
rect 23 188 159 226
rect 23 154 39 188
rect 73 154 159 188
rect 227 218 377 234
rect 227 184 243 218
rect 277 202 377 218
rect 277 184 327 202
rect 23 150 159 154
rect 297 168 327 184
rect 361 168 377 202
rect 297 152 377 168
rect 411 189 461 360
rect 636 344 702 360
rect 445 155 461 189
rect 23 116 263 150
rect 411 119 461 155
rect 495 310 594 326
rect 495 276 544 310
rect 578 276 594 310
rect 636 310 652 344
rect 686 310 702 344
rect 636 294 702 310
rect 495 260 594 276
rect 229 85 263 116
rect 495 85 529 260
rect 125 48 141 82
rect 175 48 191 82
rect 229 51 529 85
rect 563 195 629 211
rect 563 161 579 195
rect 613 161 629 195
rect 563 125 629 161
rect 563 91 579 125
rect 613 91 629 125
rect 125 17 191 48
rect 563 17 629 91
rect 663 117 697 294
rect 736 211 770 428
rect 804 363 838 581
rect 872 575 1016 649
rect 872 541 888 575
rect 922 541 975 575
rect 1009 541 1016 575
rect 872 525 1016 541
rect 1050 575 1116 591
rect 1050 541 1066 575
rect 1100 541 1116 575
rect 1050 492 1116 541
rect 1050 471 1066 492
rect 872 458 1066 471
rect 1100 458 1116 492
rect 872 455 1116 458
rect 872 421 888 455
rect 922 421 1116 455
rect 872 409 1116 421
rect 872 405 1066 409
rect 1050 375 1066 405
rect 1100 393 1116 409
rect 1169 580 1212 649
rect 1169 546 1178 580
rect 1367 580 1417 649
rect 1169 497 1212 546
rect 1169 463 1178 497
rect 1169 414 1212 463
rect 1100 375 1135 393
rect 804 347 870 363
rect 1050 359 1135 375
rect 1169 380 1178 414
rect 1252 434 1327 578
rect 1252 400 1272 434
rect 1306 400 1327 434
rect 1252 384 1327 400
rect 1401 546 1417 580
rect 1367 497 1417 546
rect 1401 463 1417 497
rect 1367 414 1417 463
rect 1169 364 1212 380
rect 804 313 820 347
rect 854 313 870 347
rect 1101 325 1135 359
rect 804 297 870 313
rect 998 309 1067 325
rect 998 275 1017 309
rect 1051 275 1067 309
rect 998 263 1067 275
rect 816 259 1067 263
rect 1101 309 1249 325
rect 1101 275 1131 309
rect 1165 275 1199 309
rect 1233 275 1249 309
rect 1101 259 1249 275
rect 816 229 1032 259
rect 816 211 850 229
rect 1101 225 1135 259
rect 1283 225 1317 384
rect 1401 380 1417 414
rect 1367 364 1417 380
rect 731 195 850 211
rect 1066 209 1135 225
rect 731 161 773 195
rect 807 161 850 195
rect 964 161 980 195
rect 1014 161 1030 195
rect 964 120 1030 161
rect 663 101 875 117
rect 663 67 825 101
rect 859 67 875 101
rect 663 51 875 67
rect 964 86 980 120
rect 1014 86 1030 120
rect 964 17 1030 86
rect 1100 191 1135 209
rect 1169 209 1228 225
rect 1100 175 1116 191
rect 1066 121 1116 175
rect 1100 87 1116 121
rect 1066 71 1116 87
rect 1169 175 1178 209
rect 1212 175 1228 209
rect 1169 120 1228 175
rect 1169 86 1178 120
rect 1212 86 1228 120
rect 1169 17 1228 86
rect 1264 209 1317 225
rect 1264 175 1265 209
rect 1299 175 1317 209
rect 1264 120 1317 175
rect 1264 86 1265 120
rect 1299 86 1317 120
rect 1264 70 1317 86
rect 1351 210 1417 226
rect 1351 176 1367 210
rect 1401 176 1417 210
rect 1351 120 1417 176
rect 1351 86 1367 120
rect 1401 86 1417 120
rect 1351 17 1417 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlxtn_2
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 464 1313 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 538 1313 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 784800
string GDS_START 773496
<< end >>
