magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1288 -1260 1541 1360
use sky130_fd_pr__hvdfl1sd2__example_55959141808316  sky130_fd_pr__hvdfl1sd2__example_55959141808316_0
timestamp 1627201311
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808137  sky130_fd_pr__hvdfl1sd__example_55959141808137_0
timestamp 1627201311
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 281 100 281 100 0 FreeSans 300 0 0 0 S
flabel comment s 128 97 128 97 0 FreeSans 300 0 0 0 D
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 23257720
string GDS_START 23256282
<< end >>
