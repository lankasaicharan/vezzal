magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1778 1975
<< nwell >>
rect -38 331 518 704
<< pwell >>
rect 1 49 463 259
rect 0 0 480 49
<< scnmos >>
rect 80 65 110 233
rect 166 65 196 233
rect 252 65 282 233
rect 338 65 368 233
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 252 367 282 619
rect 338 367 368 619
<< ndiff >>
rect 27 221 80 233
rect 27 187 35 221
rect 69 187 80 221
rect 27 111 80 187
rect 27 77 35 111
rect 69 77 80 111
rect 27 65 80 77
rect 110 175 166 233
rect 110 141 121 175
rect 155 141 166 175
rect 110 107 166 141
rect 110 73 121 107
rect 155 73 166 107
rect 110 65 166 73
rect 196 221 252 233
rect 196 187 207 221
rect 241 187 252 221
rect 196 111 252 187
rect 196 77 207 111
rect 241 77 252 111
rect 196 65 252 77
rect 282 225 338 233
rect 282 191 293 225
rect 327 191 338 225
rect 282 155 338 191
rect 282 121 293 155
rect 327 121 338 155
rect 282 65 338 121
rect 368 179 437 233
rect 368 145 395 179
rect 429 145 437 179
rect 368 111 437 145
rect 368 77 395 111
rect 429 77 437 111
rect 368 65 437 77
<< pdiff >>
rect 27 607 80 619
rect 27 573 35 607
rect 69 573 80 607
rect 27 518 80 573
rect 27 484 35 518
rect 69 484 80 518
rect 27 435 80 484
rect 27 401 35 435
rect 69 401 80 435
rect 27 367 80 401
rect 110 599 166 619
rect 110 565 121 599
rect 155 565 166 599
rect 110 519 166 565
rect 110 485 121 519
rect 155 485 166 519
rect 110 434 166 485
rect 110 400 121 434
rect 155 400 166 434
rect 110 367 166 400
rect 196 607 252 619
rect 196 573 207 607
rect 241 573 252 607
rect 196 497 252 573
rect 196 463 207 497
rect 241 463 252 497
rect 196 367 252 463
rect 282 599 338 619
rect 282 565 293 599
rect 327 565 338 599
rect 282 519 338 565
rect 282 485 293 519
rect 327 485 338 519
rect 282 434 338 485
rect 282 400 293 434
rect 327 400 338 434
rect 282 367 338 400
rect 368 607 421 619
rect 368 573 379 607
rect 413 573 421 607
rect 368 497 421 573
rect 368 463 379 497
rect 413 463 421 497
rect 368 367 421 463
<< ndiffc >>
rect 35 187 69 221
rect 35 77 69 111
rect 121 141 155 175
rect 121 73 155 107
rect 207 187 241 221
rect 207 77 241 111
rect 293 191 327 225
rect 293 121 327 155
rect 395 145 429 179
rect 395 77 429 111
<< pdiffc >>
rect 35 573 69 607
rect 35 484 69 518
rect 35 401 69 435
rect 121 565 155 599
rect 121 485 155 519
rect 121 400 155 434
rect 207 573 241 607
rect 207 463 241 497
rect 293 565 327 599
rect 293 485 327 519
rect 293 400 327 434
rect 379 573 413 607
rect 379 463 413 497
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 252 619 282 645
rect 338 619 368 645
rect 80 335 110 367
rect 166 335 196 367
rect 80 319 196 335
rect 80 285 110 319
rect 144 285 196 319
rect 80 269 196 285
rect 80 233 110 269
rect 166 233 196 269
rect 252 335 282 367
rect 338 335 368 367
rect 252 319 368 335
rect 252 285 293 319
rect 327 285 368 319
rect 252 269 368 285
rect 252 233 282 269
rect 338 233 368 269
rect 80 39 110 65
rect 166 39 196 65
rect 252 39 282 65
rect 338 39 368 65
<< polycont >>
rect 110 285 144 319
rect 293 285 327 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 19 607 85 649
rect 19 573 35 607
rect 69 573 85 607
rect 19 518 85 573
rect 19 484 35 518
rect 69 484 85 518
rect 19 435 85 484
rect 19 401 35 435
rect 69 401 85 435
rect 19 385 85 401
rect 119 599 157 615
rect 119 565 121 599
rect 155 565 157 599
rect 119 519 157 565
rect 119 485 121 519
rect 155 485 157 519
rect 119 434 157 485
rect 191 607 257 649
rect 191 573 207 607
rect 241 573 257 607
rect 191 497 257 573
rect 191 463 207 497
rect 241 463 257 497
rect 191 454 257 463
rect 291 599 329 615
rect 291 565 293 599
rect 327 565 329 599
rect 291 519 329 565
rect 291 485 293 519
rect 327 485 329 519
rect 119 400 121 434
rect 155 418 157 434
rect 291 434 329 485
rect 363 607 429 649
rect 363 573 379 607
rect 413 573 429 607
rect 363 497 429 573
rect 363 463 379 497
rect 413 463 429 497
rect 363 452 429 463
rect 291 418 293 434
rect 155 400 293 418
rect 327 418 329 434
rect 327 400 462 418
rect 119 384 462 400
rect 17 319 186 350
rect 17 285 110 319
rect 144 285 186 319
rect 17 283 186 285
rect 220 319 366 350
rect 220 285 293 319
rect 327 285 366 319
rect 220 283 366 285
rect 400 249 462 384
rect 19 221 241 249
rect 19 187 35 221
rect 69 215 207 221
rect 69 187 71 215
rect 19 111 71 187
rect 19 77 35 111
rect 69 77 71 111
rect 19 61 71 77
rect 105 175 171 181
rect 105 141 121 175
rect 155 141 171 175
rect 105 107 171 141
rect 105 73 121 107
rect 155 73 171 107
rect 105 17 171 73
rect 207 111 241 187
rect 277 225 462 249
rect 277 191 293 225
rect 327 215 462 225
rect 327 191 343 215
rect 277 155 343 191
rect 277 121 293 155
rect 327 121 343 155
rect 379 145 395 179
rect 429 145 445 179
rect 379 111 445 145
rect 379 87 395 111
rect 241 77 395 87
rect 429 77 445 111
rect 207 53 445 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2_2
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5794608
string GDS_START 5789484
<< end >>
