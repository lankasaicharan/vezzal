magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4082 1975
<< nwell >>
rect -38 331 2822 704
rect 2182 307 2495 331
<< pwell >>
rect 1089 273 1197 281
rect 1089 241 2070 273
rect 2485 241 2783 247
rect 197 220 672 229
rect 1089 220 2783 241
rect 197 177 2783 220
rect 1 49 2783 177
rect 0 0 2784 49
<< scnmos >>
rect 83 67 113 151
rect 278 119 308 203
rect 457 119 487 203
rect 543 119 573 203
rect 672 110 702 194
rect 786 110 816 194
rect 983 66 1013 194
rect 1070 66 1100 194
rect 1186 66 1216 194
rect 1412 119 1442 247
rect 1514 119 1544 247
rect 1663 163 1693 247
rect 1741 163 1771 247
rect 1866 119 1896 247
rect 1964 119 1994 247
rect 2059 77 2089 205
rect 2268 131 2298 215
rect 2370 47 2400 215
rect 2568 137 2598 221
rect 2670 53 2700 221
<< scpmoshvt >>
rect 84 481 114 609
rect 302 449 332 577
rect 430 449 460 533
rect 516 449 546 533
rect 677 449 707 533
rect 755 449 785 533
rect 998 379 1028 547
rect 1198 379 1228 547
rect 1276 379 1306 547
rect 1406 379 1436 547
rect 1501 428 1531 596
rect 1619 512 1649 596
rect 1778 512 1808 596
rect 1920 451 1950 619
rect 2006 451 2036 619
rect 2078 451 2108 619
rect 2273 343 2303 471
rect 2374 343 2404 595
rect 2568 367 2598 495
rect 2670 367 2700 619
<< ndiff >>
rect 223 176 278 203
rect 27 126 83 151
rect 27 92 38 126
rect 72 92 83 126
rect 27 67 83 92
rect 113 126 169 151
rect 113 92 124 126
rect 158 92 169 126
rect 223 142 233 176
rect 267 142 278 176
rect 223 119 278 142
rect 308 174 457 203
rect 308 140 335 174
rect 369 140 457 174
rect 308 119 457 140
rect 487 178 543 203
rect 487 144 498 178
rect 532 144 543 178
rect 487 119 543 144
rect 573 194 646 203
rect 1115 243 1171 255
rect 1115 209 1126 243
rect 1160 209 1171 243
rect 1115 194 1171 209
rect 573 165 672 194
rect 573 131 600 165
rect 634 131 672 165
rect 573 119 672 131
rect 113 67 169 92
rect 588 110 672 119
rect 702 110 786 194
rect 816 135 983 194
rect 816 110 852 135
rect 840 101 852 110
rect 886 101 983 135
rect 840 66 983 101
rect 1013 169 1070 194
rect 1013 135 1024 169
rect 1058 135 1070 169
rect 1013 66 1070 135
rect 1100 66 1186 194
rect 1216 173 1273 194
rect 1216 139 1227 173
rect 1261 139 1273 173
rect 1216 66 1273 139
rect 1355 165 1412 247
rect 1355 131 1367 165
rect 1401 131 1412 165
rect 1355 119 1412 131
rect 1442 119 1514 247
rect 1544 235 1663 247
rect 1544 201 1602 235
rect 1636 201 1663 235
rect 1544 165 1663 201
rect 1544 131 1602 165
rect 1636 163 1663 165
rect 1693 163 1741 247
rect 1771 171 1866 247
rect 1771 163 1805 171
rect 1636 131 1648 163
rect 1793 137 1805 163
rect 1839 137 1866 171
rect 1544 119 1648 131
rect 1793 119 1866 137
rect 1896 171 1964 247
rect 1896 137 1907 171
rect 1941 137 1964 171
rect 1896 119 1964 137
rect 1994 205 2044 247
rect 1994 175 2059 205
rect 1994 141 2009 175
rect 2043 141 2059 175
rect 1994 119 2059 141
rect 2009 77 2059 119
rect 2089 126 2157 205
rect 2211 180 2268 215
rect 2211 146 2223 180
rect 2257 146 2268 180
rect 2211 131 2268 146
rect 2298 184 2370 215
rect 2298 150 2325 184
rect 2359 150 2370 184
rect 2298 131 2370 150
rect 2089 92 2111 126
rect 2145 92 2157 126
rect 2089 77 2157 92
rect 2313 93 2370 131
rect 2313 59 2325 93
rect 2359 59 2370 93
rect 2313 47 2370 59
rect 2400 185 2457 215
rect 2400 151 2411 185
rect 2445 151 2457 185
rect 2400 103 2457 151
rect 2511 196 2568 221
rect 2511 162 2523 196
rect 2557 162 2568 196
rect 2511 137 2568 162
rect 2598 209 2670 221
rect 2598 175 2625 209
rect 2659 175 2670 209
rect 2598 137 2670 175
rect 2400 69 2411 103
rect 2445 69 2457 103
rect 2400 47 2457 69
rect 2613 99 2670 137
rect 2613 65 2625 99
rect 2659 65 2670 99
rect 2613 53 2670 65
rect 2700 209 2757 221
rect 2700 175 2711 209
rect 2745 175 2757 209
rect 2700 103 2757 175
rect 2700 69 2711 103
rect 2745 69 2757 103
rect 2700 53 2757 69
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 527 84 563
rect 27 493 39 527
rect 73 493 84 527
rect 27 481 84 493
rect 114 597 187 609
rect 114 563 141 597
rect 175 563 187 597
rect 114 527 187 563
rect 114 493 141 527
rect 175 493 187 527
rect 114 481 187 493
rect 245 565 302 577
rect 245 531 257 565
rect 291 531 302 565
rect 245 495 302 531
rect 245 461 257 495
rect 291 461 302 495
rect 245 449 302 461
rect 332 565 405 577
rect 332 531 359 565
rect 393 533 405 565
rect 1847 596 1920 619
rect 925 582 983 594
rect 925 548 937 582
rect 971 548 983 582
rect 925 547 983 548
rect 1451 547 1501 596
rect 925 533 998 547
rect 393 531 430 533
rect 332 495 430 531
rect 332 461 359 495
rect 393 461 430 495
rect 332 449 430 461
rect 460 508 516 533
rect 460 474 471 508
rect 505 474 516 508
rect 460 449 516 474
rect 546 508 677 533
rect 546 474 632 508
rect 666 474 677 508
rect 546 449 677 474
rect 707 449 755 533
rect 785 449 998 533
rect 925 379 998 449
rect 1028 535 1198 547
rect 1028 501 1153 535
rect 1187 501 1198 535
rect 1028 433 1198 501
rect 1028 399 1153 433
rect 1187 399 1198 433
rect 1028 379 1198 399
rect 1228 379 1276 547
rect 1306 535 1406 547
rect 1306 501 1361 535
rect 1395 501 1406 535
rect 1306 425 1406 501
rect 1306 391 1361 425
rect 1395 391 1406 425
rect 1306 379 1406 391
rect 1436 428 1501 547
rect 1531 512 1619 596
rect 1649 512 1778 596
rect 1808 586 1920 596
rect 1808 552 1859 586
rect 1893 552 1920 586
rect 1808 512 1920 552
rect 1531 500 1604 512
rect 1531 466 1558 500
rect 1592 466 1604 500
rect 1531 428 1604 466
rect 1436 379 1486 428
rect 1870 451 1920 512
rect 1950 597 2006 619
rect 1950 563 1961 597
rect 1995 563 2006 597
rect 1950 497 2006 563
rect 1950 463 1961 497
rect 1995 463 2006 497
rect 1950 451 2006 463
rect 2036 451 2078 619
rect 2108 584 2164 619
rect 2613 607 2670 619
rect 2108 550 2119 584
rect 2153 550 2164 584
rect 2108 451 2164 550
rect 2318 572 2374 595
rect 2318 538 2329 572
rect 2363 538 2374 572
rect 2318 471 2374 538
rect 2218 389 2273 471
rect 2218 355 2228 389
rect 2262 355 2273 389
rect 2218 343 2273 355
rect 2303 343 2374 471
rect 2404 583 2459 595
rect 2404 549 2415 583
rect 2449 549 2459 583
rect 2404 486 2459 549
rect 2613 573 2625 607
rect 2659 573 2670 607
rect 2613 510 2670 573
rect 2613 495 2625 510
rect 2404 452 2415 486
rect 2449 452 2459 486
rect 2404 389 2459 452
rect 2404 355 2415 389
rect 2449 355 2459 389
rect 2513 483 2568 495
rect 2513 449 2523 483
rect 2557 449 2568 483
rect 2513 413 2568 449
rect 2513 379 2523 413
rect 2557 379 2568 413
rect 2513 367 2568 379
rect 2598 476 2625 495
rect 2659 476 2670 510
rect 2598 413 2670 476
rect 2598 379 2625 413
rect 2659 379 2670 413
rect 2598 367 2670 379
rect 2700 597 2757 619
rect 2700 563 2711 597
rect 2745 563 2757 597
rect 2700 505 2757 563
rect 2700 471 2711 505
rect 2745 471 2757 505
rect 2700 413 2757 471
rect 2700 379 2711 413
rect 2745 379 2757 413
rect 2700 367 2757 379
rect 2404 343 2459 355
<< ndiffc >>
rect 38 92 72 126
rect 124 92 158 126
rect 233 142 267 176
rect 335 140 369 174
rect 498 144 532 178
rect 1126 209 1160 243
rect 600 131 634 165
rect 852 101 886 135
rect 1024 135 1058 169
rect 1227 139 1261 173
rect 1367 131 1401 165
rect 1602 201 1636 235
rect 1602 131 1636 165
rect 1805 137 1839 171
rect 1907 137 1941 171
rect 2009 141 2043 175
rect 2223 146 2257 180
rect 2325 150 2359 184
rect 2111 92 2145 126
rect 2325 59 2359 93
rect 2411 151 2445 185
rect 2523 162 2557 196
rect 2625 175 2659 209
rect 2411 69 2445 103
rect 2625 65 2659 99
rect 2711 175 2745 209
rect 2711 69 2745 103
<< pdiffc >>
rect 39 563 73 597
rect 39 493 73 527
rect 141 563 175 597
rect 141 493 175 527
rect 257 531 291 565
rect 257 461 291 495
rect 359 531 393 565
rect 937 548 971 582
rect 359 461 393 495
rect 471 474 505 508
rect 632 474 666 508
rect 1153 501 1187 535
rect 1153 399 1187 433
rect 1361 501 1395 535
rect 1361 391 1395 425
rect 1859 552 1893 586
rect 1558 466 1592 500
rect 1961 563 1995 597
rect 1961 463 1995 497
rect 2119 550 2153 584
rect 2329 538 2363 572
rect 2228 355 2262 389
rect 2415 549 2449 583
rect 2625 573 2659 607
rect 2415 452 2449 486
rect 2415 355 2449 389
rect 2523 449 2557 483
rect 2523 379 2557 413
rect 2625 476 2659 510
rect 2625 379 2659 413
rect 2711 563 2745 597
rect 2711 471 2745 505
rect 2711 379 2745 413
<< poly >>
rect 84 609 114 635
rect 302 601 546 631
rect 302 577 332 601
rect 84 325 114 481
rect 430 533 460 559
rect 516 533 546 601
rect 677 615 1531 645
rect 677 533 707 615
rect 1501 596 1531 615
rect 1619 596 1649 622
rect 1778 596 1808 622
rect 1920 619 1950 645
rect 2006 619 2036 645
rect 2078 619 2108 645
rect 755 533 785 559
rect 998 547 1028 573
rect 1198 547 1228 573
rect 1276 547 1306 573
rect 1406 547 1436 573
rect 302 380 332 449
rect 430 434 460 449
rect 23 309 114 325
rect 23 275 39 309
rect 73 275 114 309
rect 23 241 114 275
rect 23 207 39 241
rect 73 207 114 241
rect 156 357 332 380
rect 156 323 172 357
rect 206 350 332 357
rect 380 404 460 434
rect 516 423 546 449
rect 677 434 707 449
rect 594 404 707 434
rect 755 428 785 449
rect 206 323 308 350
rect 156 289 308 323
rect 380 302 410 404
rect 594 362 624 404
rect 755 401 882 428
rect 755 398 832 401
rect 458 346 624 362
rect 786 367 832 398
rect 866 367 882 401
rect 1619 491 1649 512
rect 1619 464 1730 491
rect 1778 480 1808 512
rect 1619 461 1680 464
rect 1664 430 1680 461
rect 1714 430 1730 464
rect 1501 413 1531 428
rect 1501 383 1622 413
rect 786 351 882 367
rect 458 312 474 346
rect 508 332 624 346
rect 672 334 738 350
rect 508 312 573 332
rect 156 255 172 289
rect 206 255 308 289
rect 156 239 308 255
rect 23 191 114 207
rect 278 203 308 239
rect 350 286 416 302
rect 458 296 573 312
rect 350 252 366 286
rect 400 252 416 286
rect 350 248 416 252
rect 350 236 487 248
rect 386 218 487 236
rect 457 203 487 218
rect 543 203 573 296
rect 672 300 688 334
rect 722 300 738 334
rect 672 266 738 300
rect 672 232 688 266
rect 722 232 738 266
rect 672 216 738 232
rect 83 151 113 191
rect 672 194 702 216
rect 786 194 816 351
rect 998 347 1028 379
rect 1198 347 1228 379
rect 962 331 1028 347
rect 962 297 978 331
rect 1012 297 1028 331
rect 1125 331 1228 347
rect 1125 311 1141 331
rect 962 281 1028 297
rect 1070 297 1141 311
rect 1175 297 1228 331
rect 1070 281 1228 297
rect 983 194 1013 281
rect 1070 194 1100 281
rect 1276 239 1306 379
rect 1406 346 1436 379
rect 1370 330 1436 346
rect 1370 296 1386 330
rect 1420 310 1436 330
rect 1484 319 1550 335
rect 1420 296 1442 310
rect 1370 280 1442 296
rect 1412 247 1442 280
rect 1484 285 1500 319
rect 1534 285 1550 319
rect 1484 269 1550 285
rect 1592 292 1622 383
rect 1664 396 1730 430
rect 1664 362 1680 396
rect 1714 362 1730 396
rect 1664 346 1730 362
rect 1772 464 1838 480
rect 1772 430 1788 464
rect 1822 430 1838 464
rect 2374 595 2404 621
rect 2670 619 2700 645
rect 2273 471 2303 497
rect 1920 436 1950 451
rect 1772 414 1838 430
rect 1772 292 1802 414
rect 1886 406 1950 436
rect 1886 366 1916 406
rect 1850 350 1916 366
rect 2006 358 2036 451
rect 2078 436 2108 451
rect 2078 406 2160 436
rect 1850 316 1866 350
rect 1900 316 1916 350
rect 1850 300 1916 316
rect 1958 342 2036 358
rect 1958 308 1974 342
rect 2008 308 2036 342
rect 1514 247 1544 269
rect 1592 262 1693 292
rect 1663 247 1693 262
rect 1741 262 1802 292
rect 1741 247 1771 262
rect 1866 247 1896 300
rect 1958 292 2036 308
rect 2130 303 2160 406
rect 2568 495 2598 521
rect 2273 303 2303 343
rect 2374 303 2404 343
rect 1964 247 1994 292
rect 2130 287 2196 303
rect 2130 253 2146 287
rect 2180 253 2196 287
rect 2130 250 2196 253
rect 1186 209 1306 239
rect 1186 194 1216 209
rect 83 41 113 67
rect 278 51 308 119
rect 457 93 487 119
rect 543 93 573 119
rect 672 51 702 110
rect 786 84 816 110
rect 1663 137 1693 163
rect 1741 137 1771 163
rect 2059 220 2196 250
rect 2238 287 2304 303
rect 2238 253 2254 287
rect 2288 253 2304 287
rect 2238 237 2304 253
rect 2351 287 2417 303
rect 2351 253 2367 287
rect 2401 267 2417 287
rect 2568 267 2598 367
rect 2670 327 2700 367
rect 2401 253 2598 267
rect 2640 311 2706 327
rect 2640 277 2656 311
rect 2690 277 2706 311
rect 2640 261 2706 277
rect 2351 237 2598 253
rect 2059 205 2089 220
rect 2268 215 2298 237
rect 2370 215 2400 237
rect 2568 221 2598 237
rect 2670 221 2700 261
rect 1412 93 1442 119
rect 1514 93 1544 119
rect 1866 93 1896 119
rect 1964 93 1994 119
rect 2268 105 2298 131
rect 278 21 702 51
rect 983 40 1013 66
rect 1070 40 1100 66
rect 1186 51 1216 66
rect 2059 51 2089 77
rect 1186 21 2089 51
rect 2568 111 2598 137
rect 2370 21 2400 47
rect 2670 27 2700 53
<< polycont >>
rect 39 275 73 309
rect 39 207 73 241
rect 172 323 206 357
rect 832 367 866 401
rect 1680 430 1714 464
rect 474 312 508 346
rect 172 255 206 289
rect 366 252 400 286
rect 688 300 722 334
rect 688 232 722 266
rect 978 297 1012 331
rect 1141 297 1175 331
rect 1386 296 1420 330
rect 1500 285 1534 319
rect 1680 362 1714 396
rect 1788 430 1822 464
rect 1866 316 1900 350
rect 1974 308 2008 342
rect 2146 253 2180 287
rect 2254 253 2288 287
rect 2367 253 2401 287
rect 2656 277 2690 311
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 23 597 89 649
rect 23 563 39 597
rect 73 563 89 597
rect 23 527 89 563
rect 23 493 39 527
rect 73 493 89 527
rect 23 477 89 493
rect 125 597 191 613
rect 125 563 141 597
rect 175 563 191 597
rect 125 527 191 563
rect 125 493 141 527
rect 175 493 191 527
rect 23 309 89 430
rect 23 275 39 309
rect 73 275 89 309
rect 23 241 89 275
rect 23 207 39 241
rect 73 207 89 241
rect 23 191 89 207
rect 125 373 191 493
rect 241 565 307 581
rect 241 531 257 565
rect 291 531 307 565
rect 241 495 307 531
rect 241 461 257 495
rect 291 461 307 495
rect 241 409 307 461
rect 343 565 409 649
rect 343 531 359 565
rect 393 531 409 565
rect 921 582 987 649
rect 921 548 937 582
rect 971 548 987 582
rect 343 495 409 531
rect 343 461 359 495
rect 393 461 409 495
rect 455 508 521 537
rect 455 474 471 508
rect 505 495 521 508
rect 616 508 682 537
rect 921 532 987 548
rect 1137 535 1203 551
rect 505 474 580 495
rect 455 461 580 474
rect 343 445 409 461
rect 249 375 510 409
rect 125 357 213 373
rect 125 323 172 357
rect 206 323 213 357
rect 125 289 213 323
rect 125 255 172 289
rect 206 255 213 289
rect 125 239 213 255
rect 125 155 174 239
rect 249 203 283 375
rect 458 346 510 375
rect 458 312 474 346
rect 508 312 510 346
rect 319 286 416 302
rect 458 296 510 312
rect 319 252 366 286
rect 400 252 416 286
rect 546 260 580 461
rect 319 236 416 252
rect 22 126 72 155
rect 22 92 38 126
rect 22 17 72 92
rect 108 126 174 155
rect 108 92 124 126
rect 158 92 174 126
rect 217 176 283 203
rect 482 226 580 260
rect 616 474 632 508
rect 666 479 682 508
rect 1137 501 1153 535
rect 1187 501 1203 535
rect 1137 496 1203 501
rect 666 474 794 479
rect 616 445 794 474
rect 217 142 233 176
rect 267 142 283 176
rect 217 115 283 142
rect 319 174 385 200
rect 319 140 335 174
rect 369 140 385 174
rect 108 63 174 92
rect 319 17 385 140
rect 482 178 548 226
rect 616 190 650 445
rect 686 334 724 350
rect 686 300 688 334
rect 722 300 724 334
rect 686 266 724 300
rect 760 315 794 445
rect 830 462 1203 496
rect 830 401 869 462
rect 1137 433 1203 462
rect 830 367 832 401
rect 866 367 869 401
rect 830 351 869 367
rect 905 392 1101 426
rect 905 315 939 392
rect 760 281 939 315
rect 975 350 1031 356
rect 975 331 991 350
rect 975 297 978 331
rect 1025 316 1031 350
rect 1012 297 1031 316
rect 975 281 1031 297
rect 1067 347 1101 392
rect 1137 399 1153 433
rect 1187 417 1203 433
rect 1345 535 1411 649
rect 1345 501 1361 535
rect 1395 501 1411 535
rect 1345 425 1411 501
rect 1187 399 1309 417
rect 1137 383 1309 399
rect 1067 331 1191 347
rect 1275 339 1309 383
rect 1345 391 1361 425
rect 1395 391 1411 425
rect 1345 375 1411 391
rect 1472 579 1723 613
rect 1067 297 1141 331
rect 1175 297 1191 331
rect 1067 295 1191 297
rect 1227 330 1436 339
rect 1227 296 1386 330
rect 1420 296 1436 330
rect 1227 287 1436 296
rect 1472 335 1506 579
rect 1542 500 1620 543
rect 1542 466 1558 500
rect 1592 466 1620 500
rect 1542 424 1620 466
rect 1472 319 1550 335
rect 686 232 688 266
rect 722 245 724 266
rect 1227 259 1261 287
rect 722 232 972 245
rect 686 211 972 232
rect 482 144 498 178
rect 532 144 548 178
rect 482 115 548 144
rect 584 165 650 190
rect 584 131 600 165
rect 634 131 650 165
rect 584 106 650 131
rect 836 135 902 175
rect 836 101 852 135
rect 886 101 902 135
rect 836 17 902 101
rect 938 87 972 211
rect 1110 243 1261 259
rect 1472 285 1500 319
rect 1534 285 1550 319
rect 1472 269 1550 285
rect 1472 251 1506 269
rect 1110 209 1126 243
rect 1160 225 1261 243
rect 1160 209 1176 225
rect 1008 169 1074 198
rect 1110 193 1176 209
rect 1297 217 1506 251
rect 1586 264 1620 424
rect 1664 464 1723 579
rect 1843 586 1909 649
rect 1843 552 1859 586
rect 1893 552 1909 586
rect 1843 516 1909 552
rect 1945 597 2011 613
rect 1945 563 1961 597
rect 1995 563 2011 597
rect 1945 497 2011 563
rect 2103 584 2169 649
rect 2103 550 2119 584
rect 2153 550 2169 584
rect 2103 511 2169 550
rect 2313 572 2379 649
rect 2609 607 2659 649
rect 2313 538 2329 572
rect 2363 538 2379 572
rect 2313 511 2379 538
rect 2415 583 2487 599
rect 2449 549 2487 583
rect 1945 480 1961 497
rect 1664 430 1680 464
rect 1714 430 1723 464
rect 1664 396 1723 430
rect 1772 464 1961 480
rect 1772 430 1788 464
rect 1822 463 1961 464
rect 1995 475 2011 497
rect 2415 486 2487 549
rect 2609 573 2625 607
rect 2609 510 2659 573
rect 1995 463 2379 475
rect 1822 441 2379 463
rect 1822 430 2011 441
rect 1772 414 2011 430
rect 1664 362 1680 396
rect 1714 362 1723 396
rect 1664 346 1723 362
rect 1759 350 1916 366
rect 1793 316 1866 350
rect 1900 316 1916 350
rect 1759 300 1916 316
rect 1955 342 2024 358
rect 1955 308 1974 342
rect 2008 308 2024 342
rect 1955 292 2024 308
rect 1955 264 1989 292
rect 1586 235 1989 264
rect 1008 135 1024 169
rect 1058 157 1074 169
rect 1227 173 1261 189
rect 1058 139 1227 157
rect 1058 135 1261 139
rect 1008 123 1261 135
rect 1297 87 1331 217
rect 1586 201 1602 235
rect 1636 230 1989 235
rect 1636 201 1652 230
rect 938 53 1331 87
rect 1367 165 1417 181
rect 1401 131 1417 165
rect 1367 17 1417 131
rect 1586 165 1652 201
rect 2060 200 2094 441
rect 2025 194 2094 200
rect 1586 131 1602 165
rect 1636 131 1652 165
rect 1586 115 1652 131
rect 1789 171 1855 194
rect 1789 137 1805 171
rect 1839 137 1855 171
rect 1789 17 1855 137
rect 1891 171 1957 194
rect 1891 137 1907 171
rect 1941 137 1957 171
rect 1891 87 1957 137
rect 1993 175 2094 194
rect 1993 141 2009 175
rect 2043 166 2094 175
rect 2130 389 2278 405
rect 2130 355 2228 389
rect 2262 355 2278 389
rect 2130 339 2278 355
rect 2130 287 2196 339
rect 2345 303 2379 441
rect 2449 452 2487 486
rect 2415 389 2487 452
rect 2449 355 2487 389
rect 2415 339 2487 355
rect 2130 253 2146 287
rect 2180 253 2196 287
rect 2130 200 2196 253
rect 2233 287 2304 303
rect 2233 253 2254 287
rect 2288 253 2304 287
rect 2233 236 2304 253
rect 2345 287 2417 303
rect 2345 253 2367 287
rect 2401 253 2417 287
rect 2345 237 2417 253
rect 2453 201 2487 339
rect 2130 180 2273 200
rect 2130 166 2223 180
rect 2043 141 2059 166
rect 1993 123 2059 141
rect 2207 146 2223 166
rect 2257 146 2273 180
rect 2095 126 2161 130
rect 2207 127 2273 146
rect 2309 184 2359 200
rect 2309 150 2325 184
rect 2095 92 2111 126
rect 2145 92 2161 126
rect 2095 87 2161 92
rect 1891 53 2161 87
rect 2309 93 2359 150
rect 2309 59 2325 93
rect 2309 17 2359 59
rect 2395 185 2487 201
rect 2395 151 2411 185
rect 2445 151 2487 185
rect 2395 103 2487 151
rect 2523 483 2573 499
rect 2557 449 2573 483
rect 2523 413 2573 449
rect 2557 379 2573 413
rect 2523 327 2573 379
rect 2609 476 2625 510
rect 2609 413 2659 476
rect 2609 379 2625 413
rect 2609 363 2659 379
rect 2695 597 2766 613
rect 2695 563 2711 597
rect 2745 563 2766 597
rect 2695 505 2766 563
rect 2695 471 2711 505
rect 2745 471 2766 505
rect 2695 413 2766 471
rect 2695 379 2711 413
rect 2745 379 2766 413
rect 2695 363 2766 379
rect 2523 311 2696 327
rect 2523 277 2656 311
rect 2690 277 2696 311
rect 2523 261 2696 277
rect 2523 196 2573 261
rect 2732 225 2766 363
rect 2557 162 2573 196
rect 2523 133 2573 162
rect 2609 209 2659 225
rect 2609 175 2625 209
rect 2395 69 2411 103
rect 2445 69 2487 103
rect 2395 53 2487 69
rect 2609 99 2659 175
rect 2609 65 2625 99
rect 2609 17 2659 65
rect 2695 209 2766 225
rect 2695 175 2711 209
rect 2745 175 2766 209
rect 2695 103 2766 175
rect 2695 69 2711 103
rect 2745 69 2766 103
rect 2695 53 2766 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 991 331 1025 350
rect 991 316 1012 331
rect 1012 316 1025 331
rect 1759 316 1793 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 979 350 1037 356
rect 979 316 991 350
rect 1025 347 1037 350
rect 1747 350 1805 356
rect 1747 347 1759 350
rect 1025 319 1759 347
rect 1025 316 1037 319
rect 979 310 1037 316
rect 1747 316 1759 319
rect 1793 316 1805 350
rect 1747 310 1805 316
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfbbn_1
flabel comment s 488 40 488 40 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 2431 390 2465 424 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2431 464 2465 498 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2431 538 2465 572 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2239 242 2273 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 SET_B
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2133236
string GDS_START 2113988
<< end >>
