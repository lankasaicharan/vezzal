magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 480 157 668 241
rect 1 49 668 157
rect 0 0 672 49
<< scnmos >>
rect 80 47 110 131
rect 274 47 304 131
rect 346 47 376 131
rect 418 47 448 131
rect 559 47 589 215
<< scpmoshvt >>
rect 80 512 110 596
rect 238 367 268 451
rect 341 367 371 451
rect 434 367 464 451
rect 539 367 569 619
<< ndiff >>
rect 506 203 559 215
rect 506 169 514 203
rect 548 169 559 203
rect 506 131 559 169
rect 27 106 80 131
rect 27 72 35 106
rect 69 72 80 106
rect 27 47 80 72
rect 110 106 163 131
rect 110 72 121 106
rect 155 72 163 106
rect 110 47 163 72
rect 221 106 274 131
rect 221 72 229 106
rect 263 72 274 106
rect 221 47 274 72
rect 304 47 346 131
rect 376 47 418 131
rect 448 93 559 131
rect 448 59 502 93
rect 536 59 559 93
rect 448 47 559 59
rect 589 203 642 215
rect 589 169 600 203
rect 634 169 642 203
rect 589 101 642 169
rect 589 67 600 101
rect 634 67 642 101
rect 589 47 642 67
<< pdiff >>
rect 486 607 539 619
rect 27 571 80 596
rect 27 537 35 571
rect 69 537 80 571
rect 27 512 80 537
rect 110 571 163 596
rect 110 537 121 571
rect 155 537 163 571
rect 110 512 163 537
rect 486 573 494 607
rect 528 573 539 607
rect 486 529 539 573
rect 486 495 494 529
rect 528 495 539 529
rect 486 451 539 495
rect 185 426 238 451
rect 185 392 193 426
rect 227 392 238 426
rect 185 367 238 392
rect 268 443 341 451
rect 268 409 287 443
rect 321 409 341 443
rect 268 367 341 409
rect 371 426 434 451
rect 371 392 386 426
rect 420 392 434 426
rect 371 367 434 392
rect 464 437 539 451
rect 464 403 475 437
rect 509 403 539 437
rect 464 367 539 403
rect 569 599 622 619
rect 569 565 580 599
rect 614 565 622 599
rect 569 508 622 565
rect 569 474 580 508
rect 614 474 622 508
rect 569 420 622 474
rect 569 386 580 420
rect 614 386 622 420
rect 569 367 622 386
<< ndiffc >>
rect 514 169 548 203
rect 35 72 69 106
rect 121 72 155 106
rect 229 72 263 106
rect 502 59 536 93
rect 600 169 634 203
rect 600 67 634 101
<< pdiffc >>
rect 35 537 69 571
rect 121 537 155 571
rect 494 573 528 607
rect 494 495 528 529
rect 193 392 227 426
rect 287 409 321 443
rect 386 392 420 426
rect 475 403 509 437
rect 580 565 614 599
rect 580 474 614 508
rect 580 386 614 420
<< poly >>
rect 80 596 110 622
rect 539 619 569 645
rect 80 302 110 512
rect 238 451 268 477
rect 341 451 371 477
rect 434 451 464 477
rect 21 286 110 302
rect 238 287 268 367
rect 341 297 371 367
rect 21 252 37 286
rect 71 252 110 286
rect 21 218 110 252
rect 21 184 37 218
rect 71 184 110 218
rect 21 168 110 184
rect 80 131 110 168
rect 158 271 268 287
rect 158 237 174 271
rect 208 257 268 271
rect 310 281 376 297
rect 434 287 464 367
rect 539 334 569 367
rect 526 318 592 334
rect 208 237 224 257
rect 158 203 224 237
rect 310 247 326 281
rect 360 247 376 281
rect 310 231 376 247
rect 158 169 174 203
rect 208 183 224 203
rect 208 169 304 183
rect 158 153 304 169
rect 274 131 304 153
rect 346 131 376 231
rect 418 271 484 287
rect 418 237 434 271
rect 468 237 484 271
rect 526 284 542 318
rect 576 284 592 318
rect 526 268 592 284
rect 418 203 484 237
rect 559 215 589 268
rect 418 169 434 203
rect 468 169 484 203
rect 418 153 484 169
rect 418 131 448 153
rect 80 21 110 47
rect 274 21 304 47
rect 346 21 376 47
rect 418 21 448 47
rect 559 21 589 47
<< polycont >>
rect 37 252 71 286
rect 37 184 71 218
rect 174 237 208 271
rect 326 247 360 281
rect 174 169 208 203
rect 434 237 468 271
rect 542 284 576 318
rect 434 169 468 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 19 571 79 649
rect 19 537 35 571
rect 69 537 79 571
rect 19 521 79 537
rect 113 571 171 587
rect 113 537 121 571
rect 155 537 171 571
rect 113 521 171 537
rect 17 286 79 443
rect 17 252 37 286
rect 71 252 79 286
rect 17 218 79 252
rect 17 184 37 218
rect 71 184 79 218
rect 17 162 79 184
rect 113 287 151 521
rect 271 443 337 649
rect 185 426 237 442
rect 185 392 193 426
rect 227 392 237 426
rect 271 409 287 443
rect 321 409 337 443
rect 459 607 532 649
rect 459 573 494 607
rect 528 573 532 607
rect 459 529 532 573
rect 459 495 494 529
rect 528 495 532 529
rect 271 403 337 409
rect 371 426 425 442
rect 185 369 237 392
rect 371 392 386 426
rect 420 392 425 426
rect 459 437 532 495
rect 459 403 475 437
rect 509 403 532 437
rect 576 599 655 615
rect 576 565 580 599
rect 614 565 655 599
rect 576 508 655 565
rect 576 474 580 508
rect 614 474 655 508
rect 576 420 655 474
rect 371 369 425 392
rect 576 386 580 420
rect 614 386 655 420
rect 576 370 655 386
rect 185 335 540 369
rect 113 271 210 287
rect 113 237 174 271
rect 208 237 210 271
rect 113 203 210 237
rect 113 169 174 203
rect 208 169 210 203
rect 113 153 210 169
rect 19 106 79 122
rect 19 72 35 106
rect 69 72 79 106
rect 19 17 79 72
rect 113 106 171 153
rect 244 117 279 335
rect 506 334 540 335
rect 506 318 578 334
rect 113 72 121 106
rect 155 72 171 106
rect 113 56 171 72
rect 213 106 279 117
rect 213 72 229 106
rect 263 72 279 106
rect 313 281 372 297
rect 313 247 326 281
rect 360 247 372 281
rect 313 77 372 247
rect 406 271 468 287
rect 406 237 434 271
rect 506 284 542 318
rect 576 284 578 318
rect 506 268 578 284
rect 406 203 468 237
rect 612 219 655 370
rect 406 169 434 203
rect 406 77 468 169
rect 502 203 564 219
rect 502 169 514 203
rect 548 169 564 203
rect 502 93 564 169
rect 213 56 279 72
rect 536 59 564 93
rect 502 17 564 59
rect 598 203 655 219
rect 598 169 600 203
rect 634 169 655 203
rect 598 101 655 169
rect 598 67 600 101
rect 634 67 655 101
rect 598 51 655 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and3b_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6394724
string GDS_START 6387496
<< end >>
