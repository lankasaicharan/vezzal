magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
<< pwell >>
rect 52 157 707 233
rect 942 175 1485 235
rect 1923 219 2111 271
rect 1732 175 2111 219
rect 942 157 2111 175
rect 52 49 2111 157
rect 0 0 2112 49
<< scnmos >>
rect 131 123 161 207
rect 217 123 247 207
rect 289 123 319 207
rect 434 123 464 207
rect 506 123 536 207
rect 598 123 628 207
rect 793 47 823 131
rect 1021 125 1051 209
rect 1107 125 1137 209
rect 1201 125 1231 209
rect 1357 81 1387 209
rect 1481 65 1511 149
rect 1634 65 1664 149
rect 1706 65 1736 149
rect 1811 65 1841 193
rect 2002 77 2032 245
<< scpmoshvt >>
rect 151 491 181 619
rect 253 491 283 619
rect 325 491 355 619
rect 411 491 441 619
rect 505 491 535 619
rect 598 491 628 619
rect 795 481 825 609
rect 1041 449 1071 533
rect 1127 449 1157 533
rect 1201 449 1231 533
rect 1343 449 1373 617
rect 1429 449 1459 617
rect 1585 495 1615 579
rect 1687 495 1717 579
rect 1812 411 1842 579
rect 2002 367 2032 619
<< ndiff >>
rect 78 177 131 207
rect 78 143 86 177
rect 120 143 131 177
rect 78 123 131 143
rect 161 169 217 207
rect 161 135 172 169
rect 206 135 217 169
rect 161 123 217 135
rect 247 123 289 207
rect 319 187 434 207
rect 319 153 389 187
rect 423 153 434 187
rect 319 123 434 153
rect 464 123 506 207
rect 536 171 598 207
rect 536 137 547 171
rect 581 137 598 171
rect 536 123 598 137
rect 628 185 681 207
rect 628 151 639 185
rect 673 151 681 185
rect 628 123 681 151
rect 968 183 1021 209
rect 968 149 976 183
rect 1010 149 1021 183
rect 740 93 793 131
rect 740 59 748 93
rect 782 59 793 93
rect 740 47 793 59
rect 823 93 876 131
rect 968 125 1021 149
rect 1051 181 1107 209
rect 1051 147 1062 181
rect 1096 147 1107 181
rect 1051 125 1107 147
rect 1137 125 1201 209
rect 1231 127 1357 209
rect 1231 125 1261 127
rect 823 59 834 93
rect 868 59 876 93
rect 823 47 876 59
rect 1253 93 1261 125
rect 1295 93 1357 127
rect 1253 81 1357 93
rect 1387 197 1459 209
rect 1387 163 1415 197
rect 1449 163 1459 197
rect 1387 149 1459 163
rect 1949 233 2002 245
rect 1949 199 1957 233
rect 1991 199 2002 233
rect 1758 179 1811 193
rect 1758 149 1766 179
rect 1387 81 1481 149
rect 1409 65 1481 81
rect 1511 119 1634 149
rect 1511 85 1589 119
rect 1623 85 1634 119
rect 1511 65 1634 85
rect 1664 65 1706 149
rect 1736 145 1766 149
rect 1800 145 1811 179
rect 1736 111 1811 145
rect 1736 77 1766 111
rect 1800 77 1811 111
rect 1736 65 1811 77
rect 1841 181 1894 193
rect 1841 147 1852 181
rect 1886 147 1894 181
rect 1841 113 1894 147
rect 1841 79 1852 113
rect 1886 79 1894 113
rect 1841 65 1894 79
rect 1949 123 2002 199
rect 1949 89 1957 123
rect 1991 89 2002 123
rect 1949 77 2002 89
rect 2032 233 2085 245
rect 2032 199 2043 233
rect 2077 199 2085 233
rect 2032 123 2085 199
rect 2032 89 2043 123
rect 2077 89 2085 123
rect 2032 77 2085 89
<< pdiff >>
rect 98 605 151 619
rect 98 571 106 605
rect 140 571 151 605
rect 98 537 151 571
rect 98 503 106 537
rect 140 503 151 537
rect 98 491 151 503
rect 181 578 253 619
rect 181 544 199 578
rect 233 544 253 578
rect 181 491 253 544
rect 283 491 325 619
rect 355 578 411 619
rect 355 544 366 578
rect 400 544 411 578
rect 355 491 411 544
rect 441 491 505 619
rect 535 582 598 619
rect 535 548 551 582
rect 585 548 598 582
rect 535 491 598 548
rect 628 605 681 619
rect 1270 629 1328 639
rect 628 571 639 605
rect 673 571 681 605
rect 628 537 681 571
rect 628 503 639 537
rect 673 503 681 537
rect 628 491 681 503
rect 735 595 795 609
rect 735 561 743 595
rect 777 561 795 595
rect 735 481 795 561
rect 825 529 925 609
rect 1270 595 1282 629
rect 1316 617 1328 629
rect 1316 595 1343 617
rect 1270 533 1343 595
rect 825 495 883 529
rect 917 495 925 529
rect 825 481 925 495
rect 988 495 1041 533
rect 988 461 996 495
rect 1030 461 1041 495
rect 988 449 1041 461
rect 1071 507 1127 533
rect 1071 473 1082 507
rect 1116 473 1127 507
rect 1071 449 1127 473
rect 1157 449 1201 533
rect 1231 449 1343 533
rect 1373 493 1429 617
rect 1373 459 1384 493
rect 1418 459 1429 493
rect 1373 449 1429 459
rect 1459 579 1509 617
rect 1949 607 2002 619
rect 1459 553 1585 579
rect 1459 519 1538 553
rect 1572 519 1585 553
rect 1459 495 1585 519
rect 1615 495 1687 579
rect 1717 571 1812 579
rect 1717 537 1767 571
rect 1801 537 1812 571
rect 1717 503 1812 537
rect 1717 495 1767 503
rect 1459 449 1509 495
rect 1755 469 1767 495
rect 1801 469 1812 503
rect 1755 411 1812 469
rect 1842 566 1895 579
rect 1842 532 1853 566
rect 1887 532 1895 566
rect 1842 457 1895 532
rect 1842 423 1853 457
rect 1887 423 1895 457
rect 1842 411 1895 423
rect 1949 573 1957 607
rect 1991 573 2002 607
rect 1949 513 2002 573
rect 1949 479 1957 513
rect 1991 479 2002 513
rect 1949 413 2002 479
rect 1949 379 1957 413
rect 1991 379 2002 413
rect 1949 367 2002 379
rect 2032 599 2085 619
rect 2032 565 2043 599
rect 2077 565 2085 599
rect 2032 496 2085 565
rect 2032 462 2043 496
rect 2077 462 2085 496
rect 2032 413 2085 462
rect 2032 379 2043 413
rect 2077 379 2085 413
rect 2032 367 2085 379
<< ndiffc >>
rect 86 143 120 177
rect 172 135 206 169
rect 389 153 423 187
rect 547 137 581 171
rect 639 151 673 185
rect 976 149 1010 183
rect 748 59 782 93
rect 1062 147 1096 181
rect 834 59 868 93
rect 1261 93 1295 127
rect 1415 163 1449 197
rect 1957 199 1991 233
rect 1589 85 1623 119
rect 1766 145 1800 179
rect 1766 77 1800 111
rect 1852 147 1886 181
rect 1852 79 1886 113
rect 1957 89 1991 123
rect 2043 199 2077 233
rect 2043 89 2077 123
<< pdiffc >>
rect 106 571 140 605
rect 106 503 140 537
rect 199 544 233 578
rect 366 544 400 578
rect 551 548 585 582
rect 639 571 673 605
rect 639 503 673 537
rect 743 561 777 595
rect 1282 595 1316 629
rect 883 495 917 529
rect 996 461 1030 495
rect 1082 473 1116 507
rect 1384 459 1418 493
rect 1538 519 1572 553
rect 1767 537 1801 571
rect 1767 469 1801 503
rect 1853 532 1887 566
rect 1853 423 1887 457
rect 1957 573 1991 607
rect 1957 479 1991 513
rect 1957 379 1991 413
rect 2043 565 2077 599
rect 2043 462 2077 496
rect 2043 379 2077 413
<< poly >>
rect 151 619 181 645
rect 253 619 283 645
rect 325 619 355 645
rect 411 619 441 645
rect 505 619 535 645
rect 598 619 628 645
rect 795 609 825 635
rect 151 469 181 491
rect 253 469 283 491
rect 103 439 283 469
rect 103 295 133 439
rect 181 381 247 397
rect 325 391 355 491
rect 411 459 441 491
rect 397 443 463 459
rect 397 409 413 443
rect 447 409 463 443
rect 397 393 463 409
rect 181 347 197 381
rect 231 347 247 381
rect 181 331 247 347
rect 73 279 139 295
rect 211 283 247 331
rect 73 245 89 279
rect 123 259 139 279
rect 123 245 161 259
rect 73 229 161 245
rect 131 207 161 229
rect 217 207 247 283
rect 289 375 355 391
rect 289 341 305 375
rect 339 341 355 375
rect 505 351 535 491
rect 598 376 628 491
rect 1343 617 1373 643
rect 1429 617 1459 643
rect 2002 619 2032 645
rect 1041 533 1071 559
rect 1127 533 1157 559
rect 1201 533 1231 559
rect 598 360 701 376
rect 289 307 355 341
rect 289 273 305 307
rect 339 273 355 307
rect 470 335 536 351
rect 470 301 486 335
rect 520 301 536 335
rect 470 285 536 301
rect 289 257 355 273
rect 289 207 319 257
rect 434 207 464 233
rect 506 207 536 285
rect 598 326 651 360
rect 685 326 701 360
rect 598 292 701 326
rect 598 258 651 292
rect 685 258 701 292
rect 795 287 825 481
rect 1585 579 1615 605
rect 1687 579 1717 605
rect 1812 579 1842 605
rect 1041 427 1071 449
rect 867 411 1071 427
rect 867 377 883 411
rect 917 397 1071 411
rect 917 377 933 397
rect 867 343 933 377
rect 1127 355 1157 449
rect 1201 403 1231 449
rect 1201 387 1272 403
rect 867 309 883 343
rect 917 309 933 343
rect 867 293 933 309
rect 1021 339 1159 355
rect 1021 305 1109 339
rect 1143 305 1159 339
rect 598 242 701 258
rect 757 271 825 287
rect 598 207 628 242
rect 757 237 773 271
rect 807 257 825 271
rect 1021 289 1159 305
rect 1201 353 1222 387
rect 1256 353 1272 387
rect 1201 337 1272 353
rect 807 237 823 257
rect 757 203 823 237
rect 1021 209 1051 289
rect 1107 209 1137 235
rect 1201 209 1231 337
rect 1343 301 1373 449
rect 1429 417 1459 449
rect 1429 401 1520 417
rect 1429 367 1470 401
rect 1504 367 1520 401
rect 1429 351 1520 367
rect 1585 309 1615 495
rect 1687 449 1717 495
rect 1657 433 1736 449
rect 1657 399 1673 433
rect 1707 399 1736 433
rect 1657 383 1736 399
rect 1314 285 1387 301
rect 1314 251 1330 285
rect 1364 251 1387 285
rect 1314 235 1387 251
rect 1357 209 1387 235
rect 1481 279 1615 309
rect 1481 223 1553 279
rect 757 169 773 203
rect 807 169 823 203
rect 757 153 823 169
rect 793 131 823 153
rect 131 55 161 123
rect 217 97 247 123
rect 289 97 319 123
rect 434 55 464 123
rect 506 97 536 123
rect 598 97 628 123
rect 131 25 464 55
rect 1021 99 1051 125
rect 1107 103 1137 125
rect 1093 87 1159 103
rect 1201 99 1231 125
rect 1093 53 1109 87
rect 1143 53 1159 87
rect 1481 189 1503 223
rect 1537 189 1553 223
rect 1481 173 1553 189
rect 1598 221 1664 237
rect 1598 187 1614 221
rect 1648 187 1664 221
rect 1481 149 1511 173
rect 1598 171 1664 187
rect 1634 149 1664 171
rect 1706 149 1736 383
rect 1812 379 1842 411
rect 1778 363 1844 379
rect 1778 329 1794 363
rect 1828 329 1844 363
rect 1778 295 1844 329
rect 1778 261 1794 295
rect 1828 261 1844 295
rect 1890 317 1956 333
rect 1890 283 1906 317
rect 1940 297 1956 317
rect 2002 297 2032 367
rect 1940 283 2032 297
rect 1890 267 2032 283
rect 1778 245 1844 261
rect 2002 245 2032 267
rect 1811 193 1841 245
rect 1357 55 1387 81
rect 793 21 823 47
rect 1093 37 1159 53
rect 1481 39 1511 65
rect 1634 39 1664 65
rect 1706 39 1736 65
rect 1811 39 1841 65
rect 2002 51 2032 77
<< polycont >>
rect 413 409 447 443
rect 197 347 231 381
rect 89 245 123 279
rect 305 341 339 375
rect 305 273 339 307
rect 486 301 520 335
rect 651 326 685 360
rect 651 258 685 292
rect 883 377 917 411
rect 883 309 917 343
rect 1109 305 1143 339
rect 773 237 807 271
rect 1222 353 1256 387
rect 1470 367 1504 401
rect 1673 399 1707 433
rect 1330 251 1364 285
rect 773 169 807 203
rect 1109 53 1143 87
rect 1503 189 1537 223
rect 1614 187 1648 221
rect 1794 329 1828 363
rect 1794 261 1828 295
rect 1906 283 1940 317
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 90 605 156 609
rect 90 571 106 605
rect 140 571 156 605
rect 90 537 156 571
rect 90 503 106 537
rect 140 503 156 537
rect 190 578 249 649
rect 190 544 199 578
rect 233 544 249 578
rect 190 528 249 544
rect 350 578 517 594
rect 350 544 366 578
rect 400 544 517 578
rect 350 528 517 544
rect 551 582 589 649
rect 585 548 589 582
rect 551 532 589 548
rect 623 605 689 609
rect 623 571 639 605
rect 673 571 689 605
rect 623 537 689 571
rect 727 595 779 649
rect 1266 629 1332 649
rect 727 561 743 595
rect 777 561 779 595
rect 727 545 779 561
rect 813 579 1186 613
rect 1266 595 1282 629
rect 1316 595 1332 629
rect 90 494 156 503
rect 483 498 517 528
rect 623 503 639 537
rect 673 511 689 537
rect 813 511 847 579
rect 1152 561 1186 579
rect 1751 571 1817 649
rect 1948 607 1995 649
rect 673 503 847 511
rect 90 460 447 494
rect 90 397 247 460
rect 399 443 447 460
rect 19 381 247 397
rect 19 347 197 381
rect 231 347 247 381
rect 19 331 247 347
rect 291 375 355 426
rect 399 409 413 443
rect 399 393 447 409
rect 483 464 511 498
rect 623 477 847 503
rect 483 441 545 464
rect 483 407 615 441
rect 291 341 305 375
rect 339 341 355 375
rect 19 193 53 331
rect 291 307 355 341
rect 89 279 257 295
rect 123 245 257 279
rect 89 229 257 245
rect 291 273 305 307
rect 339 273 355 307
rect 397 335 547 359
rect 397 301 486 335
rect 520 301 547 335
rect 397 299 547 301
rect 19 177 124 193
rect 19 143 86 177
rect 120 143 124 177
rect 19 127 124 143
rect 168 169 210 185
rect 168 135 172 169
rect 206 135 210 169
rect 168 17 210 135
rect 291 77 355 273
rect 581 265 615 407
rect 389 231 615 265
rect 651 360 739 443
rect 685 326 739 360
rect 651 292 739 326
rect 685 258 739 292
rect 651 235 739 258
rect 773 271 847 477
rect 807 237 847 271
rect 389 187 439 231
rect 773 203 847 237
rect 423 153 439 187
rect 389 137 439 153
rect 531 171 589 187
rect 531 137 547 171
rect 581 137 589 171
rect 623 185 773 197
rect 623 151 639 185
rect 673 169 773 185
rect 807 169 847 203
rect 673 151 847 169
rect 623 143 847 151
rect 881 529 919 545
rect 881 495 883 529
rect 917 495 919 529
rect 1152 527 1504 561
rect 881 411 919 495
rect 881 377 883 411
rect 917 377 919 411
rect 881 343 919 377
rect 881 309 883 343
rect 917 309 919 343
rect 531 17 589 137
rect 732 93 784 109
rect 881 97 919 309
rect 953 498 1034 511
rect 953 464 991 498
rect 1025 495 1034 498
rect 953 461 996 464
rect 1030 461 1034 495
rect 953 445 1034 461
rect 1068 507 1118 523
rect 1068 473 1082 507
rect 1116 473 1118 507
rect 953 199 987 445
rect 1068 409 1118 473
rect 1023 375 1118 409
rect 1023 269 1057 375
rect 1152 341 1186 527
rect 1093 339 1186 341
rect 1093 305 1109 339
rect 1143 305 1186 339
rect 1220 459 1384 493
rect 1418 459 1434 493
rect 1220 387 1434 459
rect 1220 353 1222 387
rect 1256 353 1434 387
rect 1220 337 1434 353
rect 1470 417 1504 527
rect 1538 553 1591 569
rect 1572 519 1591 553
rect 1538 503 1591 519
rect 1470 401 1521 417
rect 1504 367 1521 401
rect 1470 351 1521 367
rect 1093 303 1186 305
rect 1330 285 1364 301
rect 1023 251 1330 269
rect 1023 235 1364 251
rect 1400 267 1434 337
rect 1487 293 1521 351
rect 1557 363 1591 503
rect 1751 537 1767 571
rect 1801 537 1817 571
rect 1751 503 1817 537
rect 1751 469 1767 503
rect 1801 469 1817 503
rect 1853 566 1914 582
rect 1887 532 1914 566
rect 1853 457 1914 532
rect 1657 433 1853 435
rect 1657 399 1673 433
rect 1707 423 1853 433
rect 1887 423 1914 457
rect 1707 399 1914 423
rect 1657 397 1914 399
rect 1557 329 1794 363
rect 1828 329 1844 363
rect 1684 295 1844 329
rect 953 183 1019 199
rect 953 149 976 183
rect 1010 149 1019 183
rect 953 133 1019 149
rect 1053 181 1102 235
rect 1400 233 1453 267
rect 1487 259 1650 293
rect 1415 197 1453 233
rect 1053 147 1062 181
rect 1096 147 1102 181
rect 1053 131 1102 147
rect 1136 163 1381 197
rect 1136 97 1170 163
rect 732 59 748 93
rect 782 59 784 93
rect 732 17 784 59
rect 818 93 1170 97
rect 818 59 834 93
rect 868 87 1170 93
rect 868 59 1109 87
rect 818 53 1109 59
rect 1143 53 1170 87
rect 1245 93 1261 127
rect 1295 93 1311 127
rect 1245 17 1311 93
rect 1347 111 1381 163
rect 1449 163 1453 197
rect 1415 147 1453 163
rect 1487 223 1553 225
rect 1487 189 1503 223
rect 1537 189 1553 223
rect 1487 111 1553 189
rect 1598 221 1650 259
rect 1598 187 1614 221
rect 1648 187 1650 221
rect 1598 171 1650 187
rect 1684 261 1794 295
rect 1828 261 1844 295
rect 1880 329 1914 397
rect 1948 573 1957 607
rect 1991 573 1995 607
rect 1948 513 1995 573
rect 1948 479 1957 513
rect 1991 479 1995 513
rect 1948 413 1995 479
rect 1948 379 1957 413
rect 1991 379 1995 413
rect 1948 363 1995 379
rect 2039 599 2093 615
rect 2039 565 2043 599
rect 2077 565 2093 599
rect 2039 496 2093 565
rect 2039 462 2043 496
rect 2077 462 2093 496
rect 2039 413 2093 462
rect 2039 379 2043 413
rect 2077 379 2093 413
rect 1880 317 1956 329
rect 1880 283 1906 317
rect 1940 283 1956 317
rect 1684 135 1718 261
rect 1880 197 1914 283
rect 1347 77 1553 111
rect 1589 119 1718 135
rect 1623 85 1718 119
rect 1589 69 1718 85
rect 1762 179 1804 195
rect 1762 145 1766 179
rect 1800 145 1804 179
rect 1762 111 1804 145
rect 1762 77 1766 111
rect 1800 77 1804 111
rect 1762 17 1804 77
rect 1848 181 1914 197
rect 1848 147 1852 181
rect 1886 147 1914 181
rect 1848 113 1914 147
rect 1848 79 1852 113
rect 1886 79 1914 113
rect 1848 63 1914 79
rect 1948 233 2005 249
rect 1948 199 1957 233
rect 1991 199 2005 233
rect 1948 123 2005 199
rect 1948 89 1957 123
rect 1991 89 2005 123
rect 1948 17 2005 89
rect 2039 233 2093 379
rect 2039 199 2043 233
rect 2077 199 2093 233
rect 2039 123 2093 199
rect 2039 89 2043 123
rect 2077 89 2093 123
rect 2039 73 2093 89
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 511 464 545 498
rect 991 495 1025 498
rect 991 464 996 495
rect 996 464 1025 495
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 499 498 557 504
rect 499 464 511 498
rect 545 495 557 498
rect 979 498 1037 504
rect 979 495 991 498
rect 545 467 991 495
rect 545 464 557 467
rect 499 458 557 464
rect 979 464 991 467
rect 1025 464 1037 498
rect 979 458 1037 464
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfxtp_1
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2047 94 2081 128 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 168 2081 202 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 464 2081 498 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 538 2081 572 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4036394
string GDS_START 4019508
<< end >>
