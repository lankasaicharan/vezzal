magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 3 49 671 157
rect 0 0 672 49
<< scnmos >>
rect 86 47 116 131
rect 164 47 194 131
rect 242 47 272 131
rect 328 47 358 131
rect 400 47 430 131
rect 486 47 516 131
rect 558 47 588 131
<< scpmoshvt >>
rect 84 409 134 609
rect 190 409 240 609
rect 300 409 350 609
rect 406 409 456 609
rect 512 409 562 609
<< ndiff >>
rect 29 106 86 131
rect 29 72 41 106
rect 75 72 86 106
rect 29 47 86 72
rect 116 47 164 131
rect 194 47 242 131
rect 272 102 328 131
rect 272 68 283 102
rect 317 68 328 102
rect 272 47 328 68
rect 358 47 400 131
rect 430 111 486 131
rect 430 77 441 111
rect 475 77 486 111
rect 430 47 486 77
rect 516 47 558 131
rect 588 101 645 131
rect 588 67 599 101
rect 633 67 645 101
rect 588 47 645 67
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 190 609
rect 134 563 145 597
rect 179 563 190 597
rect 134 526 190 563
rect 134 492 145 526
rect 179 492 190 526
rect 134 455 190 492
rect 134 421 145 455
rect 179 421 190 455
rect 134 409 190 421
rect 240 597 300 609
rect 240 563 251 597
rect 285 563 300 597
rect 240 524 300 563
rect 240 490 251 524
rect 285 490 300 524
rect 240 409 300 490
rect 350 597 406 609
rect 350 563 361 597
rect 395 563 406 597
rect 350 526 406 563
rect 350 492 361 526
rect 395 492 406 526
rect 350 455 406 492
rect 350 421 361 455
rect 395 421 406 455
rect 350 409 406 421
rect 456 409 512 609
rect 562 597 619 609
rect 562 563 573 597
rect 607 563 619 597
rect 562 526 619 563
rect 562 492 573 526
rect 607 492 619 526
rect 562 455 619 492
rect 562 421 573 455
rect 607 421 619 455
rect 562 409 619 421
<< ndiffc >>
rect 41 72 75 106
rect 283 68 317 102
rect 441 77 475 111
rect 599 67 633 101
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 492 179 526
rect 145 421 179 455
rect 251 563 285 597
rect 251 490 285 524
rect 361 563 395 597
rect 361 492 395 526
rect 361 421 395 455
rect 573 563 607 597
rect 573 492 607 526
rect 573 421 607 455
<< poly >>
rect 84 609 134 635
rect 190 609 240 635
rect 300 609 350 635
rect 406 609 456 635
rect 512 609 562 635
rect 84 380 134 409
rect 84 228 114 380
rect 190 368 240 409
rect 300 368 350 409
rect 406 368 456 409
rect 512 383 562 409
rect 176 352 242 368
rect 176 332 192 352
rect 164 318 192 332
rect 226 318 242 352
rect 164 302 242 318
rect 284 352 350 368
rect 284 318 300 352
rect 334 318 350 352
rect 50 212 116 228
rect 50 178 66 212
rect 100 178 116 212
rect 50 162 116 178
rect 86 131 116 162
rect 164 131 194 302
rect 284 284 350 318
rect 284 254 300 284
rect 242 250 300 254
rect 334 250 350 284
rect 242 224 350 250
rect 398 352 464 368
rect 398 318 414 352
rect 448 318 464 352
rect 398 284 464 318
rect 398 250 414 284
rect 448 250 464 284
rect 398 234 464 250
rect 512 335 542 383
rect 512 319 578 335
rect 512 285 528 319
rect 562 285 578 319
rect 512 269 578 285
rect 242 131 272 224
rect 400 176 430 234
rect 512 186 542 269
rect 328 146 430 176
rect 328 131 358 146
rect 400 131 430 146
rect 486 156 588 186
rect 486 131 516 156
rect 558 131 588 156
rect 86 21 116 47
rect 164 21 194 47
rect 242 21 272 47
rect 328 21 358 47
rect 400 21 430 47
rect 486 21 516 47
rect 558 21 588 47
<< polycont >>
rect 192 318 226 352
rect 300 318 334 352
rect 66 178 100 212
rect 300 250 334 284
rect 414 318 448 352
rect 414 250 448 284
rect 528 285 562 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 597 89 649
rect 23 563 39 597
rect 73 563 89 597
rect 23 526 89 563
rect 23 492 39 526
rect 73 492 89 526
rect 23 455 89 492
rect 23 421 39 455
rect 73 421 89 455
rect 23 405 89 421
rect 129 597 195 613
rect 129 563 145 597
rect 179 563 195 597
rect 129 526 195 563
rect 129 492 145 526
rect 179 492 195 526
rect 129 455 195 492
rect 235 597 301 649
rect 235 563 251 597
rect 285 563 301 597
rect 235 524 301 563
rect 235 490 251 524
rect 285 490 301 524
rect 235 474 301 490
rect 345 597 411 613
rect 345 563 361 597
rect 395 563 411 597
rect 345 526 411 563
rect 345 492 361 526
rect 395 492 411 526
rect 129 421 145 455
rect 179 438 195 455
rect 345 455 411 492
rect 345 438 361 455
rect 179 421 361 438
rect 395 421 411 455
rect 129 404 411 421
rect 557 597 648 613
rect 557 563 573 597
rect 607 563 648 597
rect 557 526 648 563
rect 557 492 573 526
rect 607 492 648 526
rect 557 455 648 492
rect 557 421 573 455
rect 607 421 648 455
rect 557 405 648 421
rect 25 352 242 368
rect 25 318 192 352
rect 226 318 242 352
rect 25 302 242 318
rect 284 352 359 368
rect 284 318 300 352
rect 334 318 359 352
rect 284 284 359 318
rect 284 250 300 284
rect 334 250 359 284
rect 284 234 359 250
rect 398 352 464 368
rect 398 318 414 352
rect 448 318 464 352
rect 398 284 464 318
rect 398 250 414 284
rect 448 250 464 284
rect 505 319 578 356
rect 505 285 528 319
rect 562 285 578 319
rect 505 269 578 285
rect 398 234 464 250
rect 25 212 116 228
rect 25 178 66 212
rect 100 178 116 212
rect 614 208 648 405
rect 601 198 648 208
rect 25 162 116 178
rect 152 164 648 198
rect 152 126 186 164
rect 25 106 186 126
rect 25 72 41 106
rect 75 92 186 106
rect 267 102 333 128
rect 75 72 91 92
rect 25 53 91 72
rect 267 68 283 102
rect 317 68 333 102
rect 267 17 333 68
rect 425 111 491 164
rect 601 162 648 164
rect 425 77 441 111
rect 475 77 491 111
rect 425 53 491 77
rect 583 101 649 126
rect 583 67 599 101
rect 633 67 649 101
rect 583 17 649 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a311oi_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3268360
string GDS_START 3261626
<< end >>
