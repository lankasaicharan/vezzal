magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 159 228 606 248
rect 159 49 1630 228
rect 0 0 1632 49
<< scpmos >>
rect 140 368 170 592
rect 230 368 260 592
rect 320 368 350 592
rect 410 368 440 592
rect 604 392 634 592
rect 694 392 724 592
rect 784 392 814 592
rect 874 392 904 592
rect 1068 392 1098 592
rect 1158 392 1188 592
rect 1248 392 1278 592
rect 1338 392 1368 592
rect 1428 392 1458 592
rect 1518 392 1548 592
<< nmoslvt >>
rect 242 74 272 222
rect 328 74 358 222
rect 414 74 444 222
rect 500 74 530 222
rect 595 74 625 202
rect 681 74 711 202
rect 769 74 799 202
rect 855 74 885 202
rect 943 74 973 202
rect 1029 74 1059 202
rect 1263 74 1293 202
rect 1349 74 1379 202
rect 1435 74 1465 202
rect 1521 74 1551 202
<< ndiff >>
rect 185 142 242 222
rect 185 108 197 142
rect 231 108 242 142
rect 185 74 242 108
rect 272 210 328 222
rect 272 176 283 210
rect 317 176 328 210
rect 272 120 328 176
rect 272 86 283 120
rect 317 86 328 120
rect 272 74 328 86
rect 358 142 414 222
rect 358 108 369 142
rect 403 108 414 142
rect 358 74 414 108
rect 444 210 500 222
rect 444 176 455 210
rect 489 176 500 210
rect 444 120 500 176
rect 444 86 455 120
rect 489 86 500 120
rect 444 74 500 86
rect 530 202 580 222
rect 530 190 595 202
rect 530 156 541 190
rect 575 156 595 190
rect 530 120 595 156
rect 530 86 541 120
rect 575 86 595 120
rect 530 74 595 86
rect 625 190 681 202
rect 625 156 636 190
rect 670 156 681 190
rect 625 120 681 156
rect 625 86 636 120
rect 670 86 681 120
rect 625 74 681 86
rect 711 127 769 202
rect 711 93 723 127
rect 757 93 769 127
rect 711 74 769 93
rect 799 190 855 202
rect 799 156 810 190
rect 844 156 855 190
rect 799 120 855 156
rect 799 86 810 120
rect 844 86 855 120
rect 799 74 855 86
rect 885 188 943 202
rect 885 154 897 188
rect 931 154 943 188
rect 885 116 943 154
rect 885 82 897 116
rect 931 82 943 116
rect 885 74 943 82
rect 973 190 1029 202
rect 973 156 984 190
rect 1018 156 1029 190
rect 973 120 1029 156
rect 973 86 984 120
rect 1018 86 1029 120
rect 973 74 1029 86
rect 1059 188 1112 202
rect 1059 154 1070 188
rect 1104 154 1112 188
rect 1059 120 1112 154
rect 1059 86 1070 120
rect 1104 86 1112 120
rect 1059 74 1112 86
rect 1210 188 1263 202
rect 1210 154 1218 188
rect 1252 154 1263 188
rect 1210 120 1263 154
rect 1210 86 1218 120
rect 1252 86 1263 120
rect 1210 74 1263 86
rect 1293 175 1349 202
rect 1293 141 1304 175
rect 1338 141 1349 175
rect 1293 74 1349 141
rect 1379 190 1435 202
rect 1379 156 1390 190
rect 1424 156 1435 190
rect 1379 120 1435 156
rect 1379 86 1390 120
rect 1424 86 1435 120
rect 1379 74 1435 86
rect 1465 134 1521 202
rect 1465 100 1476 134
rect 1510 100 1521 134
rect 1465 74 1521 100
rect 1551 190 1604 202
rect 1551 156 1562 190
rect 1596 156 1604 190
rect 1551 120 1604 156
rect 1551 86 1562 120
rect 1596 86 1604 120
rect 1551 74 1604 86
<< pdiff >>
rect 85 580 140 592
rect 85 546 93 580
rect 127 546 140 580
rect 85 478 140 546
rect 85 444 93 478
rect 127 444 140 478
rect 85 368 140 444
rect 170 580 230 592
rect 170 546 183 580
rect 217 546 230 580
rect 170 497 230 546
rect 170 463 183 497
rect 217 463 230 497
rect 170 414 230 463
rect 170 380 183 414
rect 217 380 230 414
rect 170 368 230 380
rect 260 580 320 592
rect 260 546 273 580
rect 307 546 320 580
rect 260 478 320 546
rect 260 444 273 478
rect 307 444 320 478
rect 260 368 320 444
rect 350 580 410 592
rect 350 546 363 580
rect 397 546 410 580
rect 350 497 410 546
rect 350 463 363 497
rect 397 463 410 497
rect 350 414 410 463
rect 350 380 363 414
rect 397 380 410 414
rect 350 368 410 380
rect 440 580 495 592
rect 440 546 453 580
rect 487 546 495 580
rect 440 497 495 546
rect 440 463 453 497
rect 487 463 495 497
rect 440 414 495 463
rect 440 380 453 414
rect 487 380 495 414
rect 549 580 604 592
rect 549 546 557 580
rect 591 546 604 580
rect 549 508 604 546
rect 549 474 557 508
rect 591 474 604 508
rect 549 392 604 474
rect 634 531 694 592
rect 634 497 647 531
rect 681 497 694 531
rect 634 440 694 497
rect 634 406 647 440
rect 681 406 694 440
rect 634 392 694 406
rect 724 580 784 592
rect 724 546 737 580
rect 771 546 784 580
rect 724 510 784 546
rect 724 476 737 510
rect 771 476 784 510
rect 724 440 784 476
rect 724 406 737 440
rect 771 406 784 440
rect 724 392 784 406
rect 814 531 874 592
rect 814 497 827 531
rect 861 497 874 531
rect 814 440 874 497
rect 814 406 827 440
rect 861 406 874 440
rect 814 392 874 406
rect 904 580 959 592
rect 904 546 917 580
rect 951 546 959 580
rect 904 508 959 546
rect 904 474 917 508
rect 951 474 959 508
rect 904 392 959 474
rect 1013 580 1068 592
rect 1013 546 1021 580
rect 1055 546 1068 580
rect 1013 508 1068 546
rect 1013 474 1021 508
rect 1055 474 1068 508
rect 1013 392 1068 474
rect 1098 544 1158 592
rect 1098 510 1111 544
rect 1145 510 1158 544
rect 1098 440 1158 510
rect 1098 406 1111 440
rect 1145 406 1158 440
rect 1098 392 1158 406
rect 1188 580 1248 592
rect 1188 546 1201 580
rect 1235 546 1248 580
rect 1188 510 1248 546
rect 1188 476 1201 510
rect 1235 476 1248 510
rect 1188 440 1248 476
rect 1188 406 1201 440
rect 1235 406 1248 440
rect 1188 392 1248 406
rect 1278 580 1338 592
rect 1278 546 1291 580
rect 1325 546 1338 580
rect 1278 497 1338 546
rect 1278 463 1291 497
rect 1325 463 1338 497
rect 1278 392 1338 463
rect 1368 580 1428 592
rect 1368 546 1381 580
rect 1415 546 1428 580
rect 1368 510 1428 546
rect 1368 476 1381 510
rect 1415 476 1428 510
rect 1368 440 1428 476
rect 1368 406 1381 440
rect 1415 406 1428 440
rect 1368 392 1428 406
rect 1458 580 1518 592
rect 1458 546 1471 580
rect 1505 546 1518 580
rect 1458 508 1518 546
rect 1458 474 1471 508
rect 1505 474 1518 508
rect 1458 392 1518 474
rect 1548 580 1603 592
rect 1548 546 1561 580
rect 1595 546 1603 580
rect 1548 510 1603 546
rect 1548 476 1561 510
rect 1595 476 1603 510
rect 1548 440 1603 476
rect 1548 406 1561 440
rect 1595 406 1603 440
rect 1548 392 1603 406
rect 440 368 495 380
<< ndiffc >>
rect 197 108 231 142
rect 283 176 317 210
rect 283 86 317 120
rect 369 108 403 142
rect 455 176 489 210
rect 455 86 489 120
rect 541 156 575 190
rect 541 86 575 120
rect 636 156 670 190
rect 636 86 670 120
rect 723 93 757 127
rect 810 156 844 190
rect 810 86 844 120
rect 897 154 931 188
rect 897 82 931 116
rect 984 156 1018 190
rect 984 86 1018 120
rect 1070 154 1104 188
rect 1070 86 1104 120
rect 1218 154 1252 188
rect 1218 86 1252 120
rect 1304 141 1338 175
rect 1390 156 1424 190
rect 1390 86 1424 120
rect 1476 100 1510 134
rect 1562 156 1596 190
rect 1562 86 1596 120
<< pdiffc >>
rect 93 546 127 580
rect 93 444 127 478
rect 183 546 217 580
rect 183 463 217 497
rect 183 380 217 414
rect 273 546 307 580
rect 273 444 307 478
rect 363 546 397 580
rect 363 463 397 497
rect 363 380 397 414
rect 453 546 487 580
rect 453 463 487 497
rect 453 380 487 414
rect 557 546 591 580
rect 557 474 591 508
rect 647 497 681 531
rect 647 406 681 440
rect 737 546 771 580
rect 737 476 771 510
rect 737 406 771 440
rect 827 497 861 531
rect 827 406 861 440
rect 917 546 951 580
rect 917 474 951 508
rect 1021 546 1055 580
rect 1021 474 1055 508
rect 1111 510 1145 544
rect 1111 406 1145 440
rect 1201 546 1235 580
rect 1201 476 1235 510
rect 1201 406 1235 440
rect 1291 546 1325 580
rect 1291 463 1325 497
rect 1381 546 1415 580
rect 1381 476 1415 510
rect 1381 406 1415 440
rect 1471 546 1505 580
rect 1471 474 1505 508
rect 1561 546 1595 580
rect 1561 476 1595 510
rect 1561 406 1595 440
<< poly >>
rect 140 592 170 618
rect 230 592 260 618
rect 320 592 350 618
rect 410 592 440 618
rect 604 592 634 618
rect 694 592 724 618
rect 784 592 814 618
rect 874 592 904 618
rect 1068 592 1098 618
rect 1158 592 1188 618
rect 1248 592 1278 618
rect 1338 592 1368 618
rect 1428 592 1458 618
rect 1518 592 1548 618
rect 604 377 634 392
rect 694 377 724 392
rect 784 377 814 392
rect 874 377 904 392
rect 1068 377 1098 392
rect 1158 377 1188 392
rect 1248 377 1278 392
rect 1338 377 1368 392
rect 1428 377 1458 392
rect 1518 377 1548 392
rect 140 353 170 368
rect 230 353 260 368
rect 320 353 350 368
rect 410 353 440 368
rect 137 326 173 353
rect 227 326 263 353
rect 317 326 353 353
rect 407 326 443 353
rect 137 310 530 326
rect 137 276 190 310
rect 224 276 258 310
rect 292 276 326 310
rect 360 276 394 310
rect 428 276 480 310
rect 514 276 530 310
rect 601 318 637 377
rect 691 318 727 377
rect 781 356 817 377
rect 871 356 907 377
rect 1065 356 1101 377
rect 1155 356 1188 377
rect 1245 356 1281 377
rect 1335 356 1371 377
rect 781 340 925 356
rect 781 320 807 340
rect 601 302 727 318
rect 601 282 677 302
rect 137 260 530 276
rect 242 222 272 260
rect 328 222 358 260
rect 414 222 444 260
rect 500 222 530 260
rect 595 268 677 282
rect 711 268 727 302
rect 595 252 727 268
rect 769 306 807 320
rect 841 306 875 340
rect 909 306 925 340
rect 769 290 925 306
rect 1065 340 1185 356
rect 1065 306 1097 340
rect 1131 306 1185 340
rect 595 202 625 252
rect 681 202 711 252
rect 769 202 799 290
rect 859 247 889 290
rect 1065 248 1185 306
rect 1245 340 1371 356
rect 1245 306 1273 340
rect 1307 320 1371 340
rect 1307 306 1379 320
rect 1245 290 1379 306
rect 855 217 889 247
rect 943 218 1185 248
rect 855 202 885 217
rect 943 202 973 218
rect 1029 202 1059 218
rect 1263 202 1293 290
rect 1349 202 1379 290
rect 1425 318 1461 377
rect 1515 318 1551 377
rect 1425 302 1551 318
rect 1425 268 1465 302
rect 1499 268 1551 302
rect 1425 252 1551 268
rect 1435 202 1465 252
rect 1521 202 1551 252
rect 242 48 272 74
rect 328 48 358 74
rect 414 48 444 74
rect 500 48 530 74
rect 595 48 625 74
rect 681 48 711 74
rect 769 48 799 74
rect 855 48 885 74
rect 943 48 973 74
rect 1029 48 1059 74
rect 1263 48 1293 74
rect 1349 48 1379 74
rect 1435 48 1465 74
rect 1521 48 1551 74
<< polycont >>
rect 190 276 224 310
rect 258 276 292 310
rect 326 276 360 310
rect 394 276 428 310
rect 480 276 514 310
rect 677 268 711 302
rect 807 306 841 340
rect 875 306 909 340
rect 1097 306 1131 340
rect 1273 306 1307 340
rect 1465 268 1499 302
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 77 580 127 649
rect 77 546 93 580
rect 77 478 127 546
rect 77 444 93 478
rect 77 428 127 444
rect 167 580 233 596
rect 167 546 183 580
rect 217 546 233 580
rect 167 497 233 546
rect 167 463 183 497
rect 217 463 233 497
rect 167 414 233 463
rect 273 580 307 649
rect 273 478 307 546
rect 273 428 307 444
rect 347 580 413 596
rect 347 546 363 580
rect 397 546 413 580
rect 347 497 413 546
rect 347 463 363 497
rect 397 463 413 497
rect 167 394 183 414
rect 25 380 183 394
rect 217 394 233 414
rect 347 414 413 463
rect 347 394 363 414
rect 217 380 363 394
rect 397 380 413 414
rect 25 360 413 380
rect 453 580 503 649
rect 487 546 503 580
rect 453 497 503 546
rect 487 463 503 497
rect 453 414 503 463
rect 541 581 967 615
rect 541 580 607 581
rect 541 546 557 580
rect 591 546 607 580
rect 721 580 787 581
rect 541 508 607 546
rect 541 474 557 508
rect 591 474 607 508
rect 541 458 607 474
rect 647 531 681 547
rect 647 440 681 497
rect 487 380 503 414
rect 453 364 503 380
rect 609 406 647 424
rect 609 390 681 406
rect 721 546 737 580
rect 771 546 787 580
rect 901 580 967 581
rect 721 510 787 546
rect 721 476 737 510
rect 771 476 787 510
rect 721 440 787 476
rect 721 406 737 440
rect 771 406 787 440
rect 721 390 787 406
rect 827 531 861 547
rect 827 440 861 497
rect 901 546 917 580
rect 951 546 967 580
rect 901 508 967 546
rect 901 474 917 508
rect 951 474 967 508
rect 901 458 967 474
rect 1005 581 1235 615
rect 1005 580 1061 581
rect 1005 546 1021 580
rect 1055 546 1061 580
rect 1201 580 1235 581
rect 1005 508 1061 546
rect 1005 474 1021 508
rect 1055 474 1061 508
rect 1005 458 1061 474
rect 1095 544 1161 547
rect 1095 510 1111 544
rect 1145 510 1161 544
rect 1095 440 1161 510
rect 1095 424 1111 440
rect 861 406 1111 424
rect 1145 406 1161 440
rect 827 390 1161 406
rect 1201 510 1235 546
rect 1201 440 1235 476
rect 1275 580 1341 649
rect 1275 546 1291 580
rect 1325 546 1341 580
rect 1275 497 1341 546
rect 1275 463 1291 497
rect 1325 463 1341 497
rect 1275 458 1341 463
rect 1381 580 1415 596
rect 1381 510 1415 546
rect 1381 440 1415 476
rect 1455 580 1505 649
rect 1455 546 1471 580
rect 1455 508 1505 546
rect 1455 474 1471 508
rect 1455 458 1505 474
rect 1545 580 1611 596
rect 1545 546 1561 580
rect 1595 546 1611 580
rect 1545 510 1611 546
rect 1545 476 1561 510
rect 1595 476 1611 510
rect 1235 406 1381 424
rect 1545 440 1611 476
rect 1545 424 1561 440
rect 1415 406 1561 424
rect 1595 406 1611 440
rect 1201 390 1611 406
rect 25 226 130 360
rect 609 326 643 390
rect 174 310 643 326
rect 174 276 190 310
rect 224 276 258 310
rect 292 276 326 310
rect 360 276 394 310
rect 428 276 480 310
rect 514 276 643 310
rect 174 260 643 276
rect 25 210 489 226
rect 25 192 283 210
rect 317 192 455 210
rect 317 176 333 192
rect 181 142 247 158
rect 181 108 197 142
rect 231 108 247 142
rect 181 17 247 108
rect 283 120 333 176
rect 439 176 455 192
rect 609 218 643 260
rect 677 302 743 356
rect 711 268 743 302
rect 793 340 1031 356
rect 793 306 807 340
rect 841 306 875 340
rect 909 306 1031 340
rect 793 290 1031 306
rect 1081 340 1223 356
rect 1081 306 1097 340
rect 1131 306 1223 340
rect 1081 290 1223 306
rect 1257 340 1415 356
rect 1257 306 1273 340
rect 1307 306 1415 340
rect 1257 290 1415 306
rect 1449 302 1607 356
rect 677 252 743 268
rect 1449 268 1465 302
rect 1499 268 1607 302
rect 810 222 1354 256
rect 1449 252 1607 268
rect 810 218 844 222
rect 317 86 333 120
rect 283 70 333 86
rect 369 142 403 158
rect 369 17 403 108
rect 439 120 489 176
rect 439 86 455 120
rect 439 70 489 86
rect 525 190 575 206
rect 525 156 541 190
rect 525 120 575 156
rect 525 86 541 120
rect 525 17 575 86
rect 609 190 844 218
rect 609 156 636 190
rect 670 184 810 190
rect 609 120 670 156
rect 984 190 1018 222
rect 609 86 636 120
rect 609 70 670 86
rect 706 127 774 150
rect 706 93 723 127
rect 757 93 774 127
rect 706 17 774 93
rect 810 120 844 156
rect 810 70 844 86
rect 880 154 897 188
rect 931 154 948 188
rect 880 116 948 154
rect 880 82 897 116
rect 931 82 948 116
rect 880 17 948 82
rect 984 120 1018 156
rect 984 70 1018 86
rect 1054 154 1070 188
rect 1104 154 1120 188
rect 1054 120 1120 154
rect 1054 86 1070 120
rect 1104 86 1120 120
rect 1054 17 1120 86
rect 1202 154 1218 188
rect 1252 154 1268 188
rect 1202 120 1268 154
rect 1302 175 1354 222
rect 1302 141 1304 175
rect 1338 141 1354 175
rect 1302 125 1354 141
rect 1390 190 1612 218
rect 1424 184 1562 190
rect 1202 86 1218 120
rect 1252 91 1268 120
rect 1390 120 1424 156
rect 1596 156 1612 190
rect 1252 86 1390 91
rect 1202 57 1424 86
rect 1460 134 1526 150
rect 1460 100 1476 134
rect 1510 100 1526 134
rect 1460 17 1526 100
rect 1562 120 1612 156
rect 1596 86 1612 120
rect 1562 70 1612 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a2111o_4
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 75440
string GDS_START 61610
<< end >>
