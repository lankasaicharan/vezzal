magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 112 49 767 157
rect 0 0 768 49
<< scnmos >>
rect 195 47 225 131
rect 273 47 303 131
rect 359 47 389 131
rect 473 47 503 131
rect 576 47 606 131
rect 654 47 684 131
<< scpmoshvt >>
rect 87 409 137 609
rect 193 409 243 609
rect 360 409 410 609
rect 466 409 516 609
rect 618 409 668 609
<< ndiff >>
rect 138 106 195 131
rect 138 72 150 106
rect 184 72 195 106
rect 138 47 195 72
rect 225 47 273 131
rect 303 106 359 131
rect 303 72 314 106
rect 348 72 359 106
rect 303 47 359 72
rect 389 47 473 131
rect 503 98 576 131
rect 503 64 531 98
rect 565 64 576 98
rect 503 47 576 64
rect 606 47 654 131
rect 684 103 741 131
rect 684 69 695 103
rect 729 69 741 103
rect 684 47 741 69
<< pdiff >>
rect 30 597 87 609
rect 30 563 42 597
rect 76 563 87 597
rect 30 526 87 563
rect 30 492 42 526
rect 76 492 87 526
rect 30 455 87 492
rect 30 421 42 455
rect 76 421 87 455
rect 30 409 87 421
rect 137 597 193 609
rect 137 563 148 597
rect 182 563 193 597
rect 137 529 193 563
rect 137 495 148 529
rect 182 495 193 529
rect 137 461 193 495
rect 137 427 148 461
rect 182 427 193 461
rect 137 409 193 427
rect 243 527 360 609
rect 243 493 315 527
rect 349 493 360 527
rect 243 455 360 493
rect 243 421 315 455
rect 349 421 360 455
rect 243 409 360 421
rect 410 597 466 609
rect 410 563 421 597
rect 455 563 466 597
rect 410 515 466 563
rect 410 481 421 515
rect 455 481 466 515
rect 410 409 466 481
rect 516 597 618 609
rect 516 563 527 597
rect 561 563 618 597
rect 516 515 618 563
rect 516 481 527 515
rect 561 481 618 515
rect 516 409 618 481
rect 668 597 725 609
rect 668 563 679 597
rect 713 563 725 597
rect 668 526 725 563
rect 668 492 679 526
rect 713 492 725 526
rect 668 455 725 492
rect 668 421 679 455
rect 713 421 725 455
rect 668 409 725 421
<< ndiffc >>
rect 150 72 184 106
rect 314 72 348 106
rect 531 64 565 98
rect 695 69 729 103
<< pdiffc >>
rect 42 563 76 597
rect 42 492 76 526
rect 42 421 76 455
rect 148 563 182 597
rect 148 495 182 529
rect 148 427 182 461
rect 315 493 349 527
rect 315 421 349 455
rect 421 563 455 597
rect 421 481 455 515
rect 527 563 561 597
rect 527 481 561 515
rect 679 563 713 597
rect 679 492 713 526
rect 679 421 713 455
<< poly >>
rect 87 609 137 635
rect 193 609 243 635
rect 360 609 410 635
rect 466 609 516 635
rect 618 609 668 635
rect 87 358 137 409
rect 193 375 243 409
rect 179 359 245 375
rect 51 342 117 358
rect 51 308 67 342
rect 101 308 117 342
rect 51 274 117 308
rect 51 240 67 274
rect 101 240 117 274
rect 179 325 195 359
rect 229 325 245 359
rect 360 356 410 409
rect 466 359 516 409
rect 179 291 245 325
rect 324 340 390 356
rect 324 320 340 340
rect 179 257 195 291
rect 229 257 245 291
rect 179 241 245 257
rect 287 306 340 320
rect 374 306 390 340
rect 287 290 390 306
rect 473 343 557 359
rect 473 309 507 343
rect 541 309 557 343
rect 51 224 117 240
rect 195 131 225 241
rect 287 176 317 290
rect 473 275 557 309
rect 618 289 668 409
rect 473 241 507 275
rect 541 241 557 275
rect 273 146 317 176
rect 359 221 425 237
rect 359 187 375 221
rect 409 187 425 221
rect 359 171 425 187
rect 473 225 557 241
rect 609 273 684 289
rect 609 239 625 273
rect 659 239 684 273
rect 273 131 303 146
rect 359 131 389 171
rect 473 131 503 225
rect 609 205 684 239
rect 609 177 625 205
rect 576 171 625 177
rect 659 171 684 205
rect 576 147 684 171
rect 576 131 606 147
rect 654 131 684 147
rect 195 21 225 47
rect 273 21 303 47
rect 359 21 389 47
rect 473 21 503 47
rect 576 21 606 47
rect 654 21 684 47
<< polycont >>
rect 67 308 101 342
rect 67 240 101 274
rect 195 325 229 359
rect 195 257 229 291
rect 340 306 374 340
rect 507 309 541 343
rect 507 241 541 275
rect 375 187 409 221
rect 625 239 659 273
rect 625 171 659 205
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 26 597 92 649
rect 26 563 42 597
rect 76 563 92 597
rect 26 526 92 563
rect 26 492 42 526
rect 76 492 92 526
rect 26 455 92 492
rect 26 421 42 455
rect 76 421 92 455
rect 26 405 92 421
rect 132 597 471 613
rect 132 563 148 597
rect 182 579 421 597
rect 182 563 198 579
rect 132 529 198 563
rect 405 563 421 579
rect 455 563 471 597
rect 132 495 148 529
rect 182 495 198 529
rect 132 461 198 495
rect 132 427 148 461
rect 182 427 198 461
rect 132 411 198 427
rect 299 527 365 543
rect 299 493 315 527
rect 349 493 365 527
rect 299 455 365 493
rect 405 515 471 563
rect 405 481 421 515
rect 455 481 471 515
rect 405 465 471 481
rect 511 597 577 649
rect 511 563 527 597
rect 561 563 577 597
rect 511 515 577 563
rect 511 481 527 515
rect 561 481 577 515
rect 511 465 577 481
rect 663 597 745 613
rect 663 563 679 597
rect 713 563 745 597
rect 663 526 745 563
rect 663 492 679 526
rect 713 492 745 526
rect 299 421 315 455
rect 349 429 365 455
rect 663 455 745 492
rect 349 421 627 429
rect 299 395 627 421
rect 663 421 679 455
rect 713 421 745 455
rect 663 405 745 421
rect 179 359 263 375
rect 25 342 117 358
rect 25 308 67 342
rect 101 308 117 342
rect 25 274 117 308
rect 25 240 67 274
rect 101 240 117 274
rect 179 325 195 359
rect 229 325 263 359
rect 179 291 263 325
rect 179 257 195 291
rect 229 257 263 291
rect 313 340 455 356
rect 313 306 340 340
rect 374 306 455 340
rect 313 290 455 306
rect 491 343 557 359
rect 491 309 507 343
rect 541 309 557 343
rect 179 241 263 257
rect 491 275 557 309
rect 491 241 507 275
rect 541 241 557 275
rect 25 224 117 240
rect 83 205 117 224
rect 359 221 425 237
rect 491 225 557 241
rect 593 289 627 395
rect 697 384 745 405
rect 593 273 675 289
rect 593 239 625 273
rect 659 239 675 273
rect 359 205 375 221
rect 83 187 375 205
rect 409 187 425 221
rect 593 205 675 239
rect 593 189 625 205
rect 83 171 425 187
rect 461 171 625 189
rect 659 171 675 205
rect 461 155 675 171
rect 461 135 495 155
rect 134 106 200 135
rect 134 72 150 106
rect 184 72 200 106
rect 134 17 200 72
rect 298 106 495 135
rect 711 119 745 384
rect 298 72 314 106
rect 348 101 495 106
rect 348 72 364 101
rect 298 59 364 72
rect 531 98 581 119
rect 565 64 581 98
rect 531 17 581 64
rect 679 103 745 119
rect 679 69 695 103
rect 729 69 745 103
rect 679 53 745 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a22o_lp
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1119928
string GDS_START 1112590
<< end >>
