magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 2 49 931 167
rect 0 0 960 49
<< scnmos >>
rect 85 57 115 141
rect 157 57 187 141
rect 319 57 349 141
rect 397 57 427 141
rect 560 57 590 141
rect 660 57 690 141
rect 746 57 776 141
rect 818 57 848 141
<< scpmoshvt >>
rect 84 401 134 601
rect 256 401 306 601
rect 354 401 404 601
rect 468 401 518 601
rect 566 401 616 601
rect 672 401 722 601
<< ndiff >>
rect 28 116 85 141
rect 28 82 40 116
rect 74 82 85 116
rect 28 57 85 82
rect 115 57 157 141
rect 187 116 319 141
rect 187 82 198 116
rect 232 82 319 116
rect 187 57 319 82
rect 349 57 397 141
rect 427 116 560 141
rect 427 82 515 116
rect 549 82 560 116
rect 427 57 560 82
rect 590 57 660 141
rect 690 116 746 141
rect 690 82 701 116
rect 735 82 746 116
rect 690 57 746 82
rect 776 57 818 141
rect 848 116 905 141
rect 848 82 859 116
rect 893 82 905 116
rect 848 57 905 82
<< pdiff >>
rect 27 589 84 601
rect 27 555 39 589
rect 73 555 84 589
rect 27 518 84 555
rect 27 484 39 518
rect 73 484 84 518
rect 27 447 84 484
rect 27 413 39 447
rect 73 413 84 447
rect 27 401 84 413
rect 134 588 256 601
rect 134 554 145 588
rect 179 554 256 588
rect 134 401 256 554
rect 306 401 354 601
rect 404 447 468 601
rect 404 413 415 447
rect 449 413 468 447
rect 404 401 468 413
rect 518 401 566 601
rect 616 588 672 601
rect 616 554 627 588
rect 661 554 672 588
rect 616 401 672 554
rect 722 589 779 601
rect 722 555 733 589
rect 767 555 779 589
rect 722 518 779 555
rect 722 484 733 518
rect 767 484 779 518
rect 722 447 779 484
rect 722 413 733 447
rect 767 413 779 447
rect 722 401 779 413
<< ndiffc >>
rect 40 82 74 116
rect 198 82 232 116
rect 515 82 549 116
rect 701 82 735 116
rect 859 82 893 116
<< pdiffc >>
rect 39 555 73 589
rect 39 484 73 518
rect 39 413 73 447
rect 145 554 179 588
rect 415 413 449 447
rect 627 554 661 588
rect 733 555 767 589
rect 733 484 767 518
rect 733 413 767 447
<< poly >>
rect 84 601 134 627
rect 256 601 306 627
rect 354 601 404 627
rect 468 601 518 627
rect 566 601 616 627
rect 672 601 722 627
rect 84 259 134 401
rect 256 369 306 401
rect 182 353 306 369
rect 182 319 198 353
rect 232 319 306 353
rect 182 303 306 319
rect 354 369 404 401
rect 354 353 420 369
rect 354 319 370 353
rect 404 319 420 353
rect 354 303 420 319
rect 104 247 134 259
rect 104 231 192 247
rect 104 211 142 231
rect 85 197 142 211
rect 176 197 192 231
rect 85 181 192 197
rect 276 186 306 303
rect 468 295 518 401
rect 566 361 616 401
rect 672 361 722 401
rect 566 345 848 361
rect 566 311 585 345
rect 619 311 653 345
rect 687 311 721 345
rect 755 311 789 345
rect 823 311 848 345
rect 566 295 848 311
rect 468 229 498 295
rect 397 213 498 229
rect 85 141 115 181
rect 157 141 187 181
rect 276 156 349 186
rect 319 141 349 156
rect 397 179 413 213
rect 447 199 498 213
rect 546 231 612 247
rect 447 179 463 199
rect 546 197 562 231
rect 596 197 612 231
rect 546 181 612 197
rect 397 163 463 179
rect 397 141 427 163
rect 560 141 590 181
rect 660 141 690 295
rect 746 141 776 295
rect 818 141 848 295
rect 85 31 115 57
rect 157 31 187 57
rect 319 31 349 57
rect 397 31 427 57
rect 560 31 590 57
rect 660 31 690 57
rect 746 31 776 57
rect 818 31 848 57
<< polycont >>
rect 198 319 232 353
rect 370 319 404 353
rect 142 197 176 231
rect 585 311 619 345
rect 653 311 687 345
rect 721 311 755 345
rect 789 311 823 345
rect 413 179 447 213
rect 562 197 596 231
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 589 89 605
rect 23 555 39 589
rect 73 555 89 589
rect 23 518 89 555
rect 129 588 195 649
rect 129 554 145 588
rect 179 554 195 588
rect 129 553 195 554
rect 611 588 677 649
rect 611 554 627 588
rect 661 554 677 588
rect 611 553 677 554
rect 717 589 783 605
rect 717 555 733 589
rect 767 555 783 589
rect 23 484 39 518
rect 73 504 89 518
rect 717 518 783 555
rect 717 517 733 518
rect 73 484 90 504
rect 23 447 90 484
rect 23 413 39 447
rect 73 413 90 447
rect 23 116 90 413
rect 182 484 733 517
rect 767 484 783 518
rect 182 483 783 484
rect 182 353 248 483
rect 717 447 783 483
rect 182 319 198 353
rect 232 319 248 353
rect 182 303 248 319
rect 284 413 415 447
rect 449 413 465 447
rect 717 413 733 447
rect 767 431 783 447
rect 767 413 909 431
rect 284 247 318 413
rect 717 397 909 413
rect 354 353 533 369
rect 354 319 370 353
rect 404 319 533 353
rect 354 303 533 319
rect 126 231 318 247
rect 126 197 142 231
rect 176 197 318 231
rect 499 247 533 303
rect 569 345 839 361
rect 569 311 585 345
rect 619 311 653 345
rect 687 311 721 345
rect 755 311 789 345
rect 823 311 839 345
rect 569 295 839 311
rect 499 231 647 247
rect 126 181 318 197
rect 23 82 40 116
rect 74 82 90 116
rect 23 53 90 82
rect 182 116 248 145
rect 182 82 198 116
rect 232 82 248 116
rect 182 17 248 82
rect 284 103 318 181
rect 397 213 463 229
rect 397 179 413 213
rect 447 179 463 213
rect 499 197 562 231
rect 596 197 647 231
rect 499 181 647 197
rect 397 162 463 179
rect 499 116 565 145
rect 499 103 515 116
rect 284 82 515 103
rect 549 82 565 116
rect 601 88 647 181
rect 875 145 909 397
rect 685 116 751 145
rect 284 69 565 82
rect 685 82 701 116
rect 735 82 751 116
rect 685 17 751 82
rect 843 116 909 145
rect 843 82 859 116
rect 893 82 909 116
rect 843 53 909 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2_lp2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1663568
string GDS_START 1656026
<< end >>
