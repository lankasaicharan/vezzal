magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3794 1975
<< nwell >>
rect -38 331 2534 704
<< pwell >>
rect 2 229 198 266
rect 855 261 1220 279
rect 855 229 1546 261
rect 2190 229 2495 250
rect 2 181 1546 229
rect 1810 181 2495 229
rect 2 49 2495 181
rect 0 0 2496 49
<< scnmos >>
rect 81 156 111 240
rect 302 119 332 203
rect 464 119 494 203
rect 550 119 580 203
rect 636 119 666 203
rect 708 119 738 203
rect 934 169 964 253
rect 1006 169 1036 253
rect 1111 125 1141 253
rect 1301 151 1331 235
rect 1410 107 1440 235
rect 1627 71 1657 155
rect 1699 71 1729 155
rect 1889 119 1919 203
rect 1975 119 2005 203
rect 2269 56 2299 224
rect 2386 56 2416 224
<< scpmoshvt >>
rect 81 456 111 584
rect 348 465 378 593
rect 485 533 515 617
rect 571 533 601 617
rect 657 533 687 617
rect 729 533 759 617
rect 1034 533 1064 617
rect 1120 533 1150 617
rect 1229 449 1259 617
rect 1337 449 1367 617
rect 1442 449 1472 533
rect 1535 449 1565 533
rect 1621 449 1651 533
rect 1875 431 1905 515
rect 1984 431 2014 559
rect 2263 367 2293 619
rect 2349 367 2379 619
<< ndiff >>
rect 28 204 81 240
rect 28 170 36 204
rect 70 170 81 204
rect 28 156 81 170
rect 111 216 172 240
rect 111 182 130 216
rect 164 182 172 216
rect 111 156 172 182
rect 881 241 934 253
rect 881 207 889 241
rect 923 207 934 241
rect 249 173 302 203
rect 249 139 257 173
rect 291 139 302 173
rect 249 119 302 139
rect 332 164 464 203
rect 332 130 345 164
rect 379 130 464 164
rect 332 119 464 130
rect 494 179 550 203
rect 494 145 505 179
rect 539 145 550 179
rect 494 119 550 145
rect 580 179 636 203
rect 580 145 591 179
rect 625 145 636 179
rect 580 119 636 145
rect 666 119 708 203
rect 738 165 795 203
rect 881 169 934 207
rect 964 169 1006 253
rect 1036 199 1111 253
rect 1036 169 1066 199
rect 738 131 749 165
rect 783 131 795 165
rect 1058 165 1066 169
rect 1100 165 1111 199
rect 738 119 795 131
rect 1058 125 1111 165
rect 1141 199 1194 253
rect 1141 165 1152 199
rect 1186 165 1194 199
rect 1141 125 1194 165
rect 1248 209 1301 235
rect 1248 175 1256 209
rect 1290 175 1301 209
rect 1248 151 1301 175
rect 1331 227 1410 235
rect 1331 193 1356 227
rect 1390 193 1410 227
rect 1331 151 1410 193
rect 1353 107 1410 151
rect 1440 107 1520 235
rect 1836 178 1889 203
rect 1462 87 1520 107
rect 1462 53 1474 87
rect 1508 53 1520 87
rect 1574 130 1627 155
rect 1574 96 1582 130
rect 1616 96 1627 130
rect 1574 71 1627 96
rect 1657 71 1699 155
rect 1729 130 1782 155
rect 1729 96 1740 130
rect 1774 96 1782 130
rect 1836 144 1844 178
rect 1878 144 1889 178
rect 1836 119 1889 144
rect 1919 178 1975 203
rect 1919 144 1930 178
rect 1964 144 1975 178
rect 1919 119 1975 144
rect 2005 178 2058 203
rect 2216 212 2269 224
rect 2005 144 2016 178
rect 2050 144 2058 178
rect 2005 119 2058 144
rect 2216 178 2224 212
rect 2258 178 2269 212
rect 2216 144 2269 178
rect 1729 71 1782 96
rect 2216 110 2224 144
rect 2258 110 2269 144
rect 1462 45 1520 53
rect 2216 56 2269 110
rect 2299 208 2386 224
rect 2299 174 2332 208
rect 2366 174 2386 208
rect 2299 102 2386 174
rect 2299 68 2332 102
rect 2366 68 2386 102
rect 2299 56 2386 68
rect 2416 212 2469 224
rect 2416 178 2427 212
rect 2461 178 2469 212
rect 2416 102 2469 178
rect 2416 68 2427 102
rect 2461 68 2469 102
rect 2416 56 2469 68
<< pdiff >>
rect 28 572 81 584
rect 28 538 36 572
rect 70 538 81 572
rect 28 456 81 538
rect 111 570 164 584
rect 111 536 122 570
rect 156 536 164 570
rect 421 593 485 617
rect 295 579 348 593
rect 111 502 164 536
rect 111 468 122 502
rect 156 468 164 502
rect 111 456 164 468
rect 295 545 303 579
rect 337 545 348 579
rect 295 511 348 545
rect 295 477 303 511
rect 337 477 348 511
rect 295 465 348 477
rect 378 585 485 593
rect 378 551 416 585
rect 450 551 485 585
rect 378 533 485 551
rect 515 594 571 617
rect 515 560 526 594
rect 560 560 571 594
rect 515 533 571 560
rect 601 594 657 617
rect 601 560 612 594
rect 646 560 657 594
rect 601 533 657 560
rect 687 533 729 617
rect 759 603 1034 617
rect 759 569 770 603
rect 804 569 1034 603
rect 759 533 1034 569
rect 1064 587 1120 617
rect 1064 553 1075 587
rect 1109 553 1120 587
rect 1064 533 1120 553
rect 1150 582 1229 617
rect 1150 548 1180 582
rect 1214 548 1229 582
rect 1150 533 1229 548
rect 378 465 428 533
rect 1172 449 1229 533
rect 1259 449 1337 617
rect 1367 533 1420 617
rect 1927 551 1984 559
rect 1367 519 1442 533
rect 1367 485 1378 519
rect 1412 485 1442 519
rect 1367 449 1442 485
rect 1472 449 1535 533
rect 1565 506 1621 533
rect 1565 472 1576 506
rect 1610 472 1621 506
rect 1565 449 1621 472
rect 1651 495 1704 533
rect 1927 517 1939 551
rect 1973 517 1984 551
rect 1927 515 1984 517
rect 1651 461 1662 495
rect 1696 461 1704 495
rect 1651 449 1704 461
rect 1822 490 1875 515
rect 1822 456 1830 490
rect 1864 456 1875 490
rect 1822 431 1875 456
rect 1905 481 1984 515
rect 1905 447 1916 481
rect 1950 447 1984 481
rect 1905 431 1984 447
rect 2014 545 2067 559
rect 2014 511 2025 545
rect 2059 511 2067 545
rect 2014 477 2067 511
rect 2014 443 2025 477
rect 2059 443 2067 477
rect 2014 431 2067 443
rect 2210 429 2263 619
rect 2210 395 2218 429
rect 2252 395 2263 429
rect 2210 367 2263 395
rect 2293 597 2349 619
rect 2293 563 2304 597
rect 2338 563 2349 597
rect 2293 367 2349 563
rect 2379 599 2432 619
rect 2379 565 2390 599
rect 2424 565 2432 599
rect 2379 503 2432 565
rect 2379 469 2390 503
rect 2424 469 2432 503
rect 2379 413 2432 469
rect 2379 379 2390 413
rect 2424 379 2432 413
rect 2379 367 2432 379
<< ndiffc >>
rect 36 170 70 204
rect 130 182 164 216
rect 889 207 923 241
rect 257 139 291 173
rect 345 130 379 164
rect 505 145 539 179
rect 591 145 625 179
rect 749 131 783 165
rect 1066 165 1100 199
rect 1152 165 1186 199
rect 1256 175 1290 209
rect 1356 193 1390 227
rect 1474 53 1508 87
rect 1582 96 1616 130
rect 1740 96 1774 130
rect 1844 144 1878 178
rect 1930 144 1964 178
rect 2016 144 2050 178
rect 2224 178 2258 212
rect 2224 110 2258 144
rect 2332 174 2366 208
rect 2332 68 2366 102
rect 2427 178 2461 212
rect 2427 68 2461 102
<< pdiffc >>
rect 36 538 70 572
rect 122 536 156 570
rect 122 468 156 502
rect 303 545 337 579
rect 303 477 337 511
rect 416 551 450 585
rect 526 560 560 594
rect 612 560 646 594
rect 770 569 804 603
rect 1075 553 1109 587
rect 1180 548 1214 582
rect 1378 485 1412 519
rect 1576 472 1610 506
rect 1939 517 1973 551
rect 1662 461 1696 495
rect 1830 456 1864 490
rect 1916 447 1950 481
rect 2025 511 2059 545
rect 2025 443 2059 477
rect 2218 395 2252 429
rect 2304 563 2338 597
rect 2390 565 2424 599
rect 2390 469 2424 503
rect 2390 379 2424 413
<< poly >>
rect 197 615 378 645
rect 485 617 515 643
rect 571 617 601 643
rect 657 617 687 643
rect 729 617 759 643
rect 1034 617 1064 643
rect 1120 617 1150 643
rect 1229 617 1259 643
rect 1337 617 1367 643
rect 81 584 111 610
rect 197 605 263 615
rect 197 571 213 605
rect 247 571 263 605
rect 348 593 378 615
rect 197 555 263 571
rect 485 501 515 533
rect 460 485 529 501
rect 81 396 111 456
rect 348 439 378 465
rect 460 451 476 485
rect 510 451 529 485
rect 460 435 529 451
rect 44 380 111 396
rect 44 346 60 380
rect 94 346 111 380
rect 44 312 111 346
rect 44 278 60 312
rect 94 278 111 312
rect 44 262 111 278
rect 81 240 111 262
rect 197 413 270 429
rect 197 379 220 413
rect 254 393 270 413
rect 571 393 601 533
rect 657 433 687 533
rect 729 511 759 533
rect 1034 511 1064 533
rect 729 485 877 511
rect 729 481 827 485
rect 811 451 827 481
rect 861 451 877 485
rect 811 435 877 451
rect 919 485 1064 511
rect 919 451 935 485
rect 969 481 1064 485
rect 969 451 985 481
rect 254 379 601 393
rect 197 363 601 379
rect 643 417 732 433
rect 643 383 682 417
rect 716 383 732 417
rect 81 130 111 156
rect 197 103 227 363
rect 643 349 732 383
rect 643 321 682 349
rect 419 305 494 321
rect 302 275 377 291
rect 302 241 327 275
rect 361 241 377 275
rect 419 271 435 305
rect 469 271 494 305
rect 419 255 494 271
rect 302 225 377 241
rect 302 203 332 225
rect 464 203 494 255
rect 550 315 682 321
rect 716 315 732 349
rect 811 333 841 435
rect 919 417 985 451
rect 1120 439 1150 533
rect 1535 607 1827 637
rect 2263 619 2293 645
rect 2349 619 2379 645
rect 1442 533 1472 559
rect 1535 533 1565 607
rect 1761 597 1827 607
rect 1761 563 1777 597
rect 1811 563 1827 597
rect 1621 533 1651 559
rect 1761 547 1827 563
rect 1984 559 2014 585
rect 1875 515 1905 541
rect 919 383 935 417
rect 969 383 985 417
rect 919 367 985 383
rect 1033 423 1150 439
rect 1033 389 1049 423
rect 1083 409 1150 423
rect 1083 389 1099 409
rect 1229 403 1259 449
rect 1033 373 1099 389
rect 1193 387 1259 403
rect 1337 401 1367 449
rect 550 299 732 315
rect 780 317 846 333
rect 550 291 673 299
rect 550 203 580 291
rect 780 283 796 317
rect 830 283 846 317
rect 780 257 846 283
rect 636 203 666 229
rect 708 227 846 257
rect 934 253 964 367
rect 1033 319 1063 373
rect 1193 353 1209 387
rect 1243 353 1259 387
rect 1193 325 1259 353
rect 1006 289 1063 319
rect 1111 295 1259 325
rect 1301 385 1367 401
rect 1301 351 1317 385
rect 1351 351 1367 385
rect 1301 317 1367 351
rect 1006 253 1036 289
rect 1111 253 1141 295
rect 1301 283 1317 317
rect 1351 283 1367 317
rect 1442 287 1472 449
rect 1301 267 1367 283
rect 708 203 738 227
rect 934 143 964 169
rect 1006 143 1036 169
rect 1301 235 1331 267
rect 1410 257 1472 287
rect 1410 235 1440 257
rect 1535 243 1565 449
rect 1621 409 1651 449
rect 1875 409 1905 431
rect 1984 409 2014 431
rect 1621 393 1729 409
rect 1875 397 2014 409
rect 1621 359 1637 393
rect 1671 359 1729 393
rect 1621 343 1729 359
rect 1301 125 1331 151
rect 161 87 227 103
rect 302 93 332 119
rect 464 93 494 119
rect 550 93 580 119
rect 161 53 177 87
rect 211 53 227 87
rect 161 51 227 53
rect 636 51 666 119
rect 708 93 738 119
rect 1111 99 1141 125
rect 1535 227 1657 243
rect 1535 193 1577 227
rect 1611 193 1657 227
rect 1535 177 1657 193
rect 1627 155 1657 177
rect 1699 155 1729 343
rect 1853 381 2014 397
rect 1853 347 1869 381
rect 1903 379 2014 381
rect 2056 383 2122 399
rect 1903 347 1919 379
rect 1853 313 1919 347
rect 2056 349 2072 383
rect 2106 349 2122 383
rect 2056 333 2122 349
rect 1853 279 1869 313
rect 1903 279 1919 313
rect 1853 255 1919 279
rect 2080 327 2122 333
rect 2263 327 2293 367
rect 2080 297 2299 327
rect 2349 312 2379 367
rect 1889 225 2005 255
rect 1889 203 1919 225
rect 1975 203 2005 225
rect 2080 231 2146 297
rect 1410 51 1440 107
rect 161 21 1440 51
rect 2080 197 2096 231
rect 2130 197 2146 231
rect 2269 224 2299 297
rect 2341 296 2416 312
rect 2341 262 2357 296
rect 2391 262 2416 296
rect 2341 246 2416 262
rect 2386 224 2416 246
rect 2080 181 2146 197
rect 1889 93 1919 119
rect 1975 93 2005 119
rect 1627 45 1657 71
rect 1699 45 1729 71
rect 2269 30 2299 56
rect 2386 30 2416 56
<< polycont >>
rect 213 571 247 605
rect 476 451 510 485
rect 60 346 94 380
rect 60 278 94 312
rect 220 379 254 413
rect 827 451 861 485
rect 935 451 969 485
rect 682 383 716 417
rect 327 241 361 275
rect 435 271 469 305
rect 682 315 716 349
rect 1777 563 1811 597
rect 935 383 969 417
rect 1049 389 1083 423
rect 796 283 830 317
rect 1209 353 1243 387
rect 1317 351 1351 385
rect 1317 283 1351 317
rect 1637 359 1671 393
rect 177 53 211 87
rect 1577 193 1611 227
rect 1869 347 1903 381
rect 2072 349 2106 383
rect 1869 279 1903 313
rect 2096 197 2130 231
rect 2357 262 2391 296
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 20 572 86 649
rect 193 605 263 615
rect 193 586 213 605
rect 20 538 36 572
rect 70 538 86 572
rect 20 532 86 538
rect 120 571 213 586
rect 247 571 263 605
rect 120 570 263 571
rect 120 536 122 570
rect 156 536 263 570
rect 120 502 263 536
rect 17 418 86 498
rect 120 468 122 502
rect 156 468 263 502
rect 120 452 263 468
rect 297 579 353 595
rect 297 545 303 579
rect 337 545 353 579
rect 297 511 353 545
rect 400 585 466 649
rect 400 551 416 585
rect 450 551 466 585
rect 400 535 466 551
rect 510 594 578 610
rect 510 560 526 594
rect 560 560 578 594
rect 510 544 578 560
rect 297 477 303 511
rect 337 477 353 511
rect 17 380 94 418
rect 17 346 60 380
rect 17 312 94 346
rect 17 278 60 312
rect 17 242 94 278
rect 128 291 168 452
rect 297 418 353 477
rect 204 413 353 418
rect 204 379 220 413
rect 254 379 353 413
rect 204 363 353 379
rect 400 485 510 501
rect 400 451 476 485
rect 400 435 510 451
rect 400 305 485 435
rect 544 387 578 544
rect 128 275 366 291
rect 128 257 327 275
rect 128 216 180 257
rect 20 204 86 208
rect 20 170 36 204
rect 70 170 86 204
rect 20 17 86 170
rect 128 182 130 216
rect 164 182 180 216
rect 361 241 366 275
rect 400 271 435 305
rect 469 271 485 305
rect 521 353 578 387
rect 612 594 662 610
rect 646 560 662 594
rect 754 603 820 649
rect 754 569 770 603
rect 804 569 820 603
rect 754 565 820 569
rect 856 587 1113 603
rect 612 531 662 560
rect 856 553 1075 587
rect 1109 553 1113 587
rect 856 537 1113 553
rect 1164 582 1230 649
rect 1164 548 1180 582
rect 1214 548 1230 582
rect 612 497 791 531
rect 856 501 890 537
rect 1164 532 1230 548
rect 1266 569 1536 615
rect 327 237 366 241
rect 327 203 463 237
rect 128 166 180 182
rect 241 173 293 189
rect 241 139 257 173
rect 291 139 293 173
rect 241 103 293 139
rect 161 87 293 103
rect 161 53 177 87
rect 211 53 293 87
rect 329 164 395 169
rect 329 130 345 164
rect 379 130 395 164
rect 329 17 395 130
rect 429 94 463 203
rect 521 195 555 353
rect 612 317 646 497
rect 497 179 555 195
rect 497 145 505 179
rect 539 145 555 179
rect 497 129 555 145
rect 589 283 646 317
rect 680 417 723 433
rect 680 383 682 417
rect 716 383 723 417
rect 680 349 723 383
rect 757 387 791 497
rect 827 485 890 501
rect 861 451 890 485
rect 827 435 890 451
rect 935 485 997 501
rect 1266 498 1300 569
rect 969 451 997 485
rect 935 417 997 451
rect 757 383 935 387
rect 969 383 997 417
rect 1033 449 1300 498
rect 1362 519 1428 535
rect 1362 485 1378 519
rect 1412 485 1428 519
rect 1362 457 1428 485
rect 1033 423 1099 449
rect 1033 389 1049 423
rect 1083 389 1099 423
rect 757 353 997 383
rect 1135 387 1243 403
rect 1135 353 1209 387
rect 680 315 682 349
rect 716 315 723 349
rect 963 337 1243 353
rect 1301 385 1353 401
rect 1301 351 1317 385
rect 1351 351 1353 385
rect 963 319 1169 337
rect 1301 317 1353 351
rect 589 179 631 283
rect 680 249 723 315
rect 780 283 796 317
rect 830 283 927 317
rect 1301 301 1317 317
rect 1254 283 1317 301
rect 1351 283 1353 317
rect 680 247 853 249
rect 589 145 591 179
rect 625 145 631 179
rect 589 129 631 145
rect 665 215 853 247
rect 665 94 699 215
rect 429 60 699 94
rect 745 165 785 181
rect 745 131 749 165
rect 783 131 785 165
rect 745 17 785 131
rect 819 155 853 215
rect 889 241 927 283
rect 923 207 927 241
rect 889 191 927 207
rect 963 267 1353 283
rect 1387 297 1428 457
rect 1502 409 1536 569
rect 1570 506 1618 649
rect 1775 597 1826 613
rect 1775 563 1777 597
rect 1811 563 1826 597
rect 1570 472 1576 506
rect 1610 472 1618 506
rect 1570 456 1618 472
rect 1658 495 1741 511
rect 1658 461 1662 495
rect 1696 461 1741 495
rect 1658 445 1741 461
rect 1502 393 1673 409
rect 1502 359 1637 393
rect 1671 359 1673 393
rect 1502 343 1673 359
rect 1707 297 1741 445
rect 1775 506 1826 563
rect 1914 551 1977 649
rect 2288 597 2354 649
rect 2288 563 2304 597
rect 2338 563 2354 597
rect 1914 517 1939 551
rect 1973 517 1977 551
rect 1775 490 1880 506
rect 1775 456 1830 490
rect 1864 456 1880 490
rect 1775 440 1880 456
rect 1914 481 1977 517
rect 1914 447 1916 481
rect 1950 447 1977 481
rect 1914 431 1977 447
rect 2011 545 2068 561
rect 2288 547 2354 563
rect 2388 599 2479 615
rect 2388 565 2390 599
rect 2424 565 2479 599
rect 2011 511 2025 545
rect 2059 511 2068 545
rect 2011 477 2068 511
rect 2011 443 2025 477
rect 2059 443 2068 477
rect 2011 431 2068 443
rect 2140 479 2350 513
rect 2011 397 2106 431
rect 1853 381 1919 397
rect 1853 347 1869 381
rect 1903 347 1919 381
rect 1853 313 1919 347
rect 2056 383 2106 397
rect 2056 349 2072 383
rect 2056 333 2106 349
rect 1853 297 1869 313
rect 1387 279 1869 297
rect 1903 299 1919 313
rect 2140 299 2174 479
rect 1903 279 2174 299
rect 963 249 1306 267
rect 1387 265 2174 279
rect 2208 429 2282 445
rect 2208 395 2218 429
rect 2252 395 2282 429
rect 1387 263 1919 265
rect 963 155 997 249
rect 1387 233 1421 263
rect 1340 227 1421 233
rect 819 121 997 155
rect 1050 199 1104 215
rect 1050 165 1066 199
rect 1100 165 1104 199
rect 1050 17 1104 165
rect 1148 199 1202 215
rect 1148 165 1152 199
rect 1186 165 1202 199
rect 1148 89 1202 165
rect 1240 209 1306 215
rect 1240 175 1256 209
rect 1290 175 1306 209
rect 1340 193 1356 227
rect 1390 193 1421 227
rect 1340 191 1421 193
rect 1561 227 1887 229
rect 1561 193 1577 227
rect 1611 193 1887 227
rect 2007 197 2096 231
rect 2130 197 2146 231
rect 1561 191 1887 193
rect 1240 157 1306 175
rect 1828 178 1887 191
rect 1240 130 1620 157
rect 1240 123 1582 130
rect 1566 96 1582 123
rect 1616 96 1620 130
rect 1148 87 1524 89
rect 1148 53 1474 87
rect 1508 53 1524 87
rect 1566 80 1620 96
rect 1724 130 1790 146
rect 1724 96 1740 130
rect 1774 96 1790 130
rect 1828 144 1844 178
rect 1878 144 1887 178
rect 1828 128 1887 144
rect 1921 178 1973 194
rect 1921 144 1930 178
rect 1964 144 1973 178
rect 1724 17 1790 96
rect 1921 17 1973 144
rect 2007 178 2146 197
rect 2007 144 2016 178
rect 2050 144 2146 178
rect 2007 128 2146 144
rect 2208 212 2282 395
rect 2316 312 2350 479
rect 2388 503 2479 565
rect 2388 469 2390 503
rect 2424 469 2479 503
rect 2388 413 2479 469
rect 2388 379 2390 413
rect 2424 379 2479 413
rect 2388 348 2479 379
rect 2316 296 2391 312
rect 2316 262 2357 296
rect 2316 246 2391 262
rect 2425 212 2479 348
rect 2208 178 2224 212
rect 2258 178 2282 212
rect 2208 144 2282 178
rect 2208 110 2224 144
rect 2258 110 2282 144
rect 2208 94 2282 110
rect 2316 208 2382 212
rect 2316 174 2332 208
rect 2366 174 2382 208
rect 2316 102 2382 174
rect 2316 68 2332 102
rect 2366 68 2382 102
rect 2316 17 2382 68
rect 2425 178 2427 212
rect 2461 178 2479 212
rect 2425 102 2479 178
rect 2425 68 2427 102
rect 2461 68 2479 102
rect 2425 52 2479 68
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 683 2496 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 0 617 2496 649
rect 0 17 2496 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
rect 0 -49 2496 -17
<< labels >>
flabel pwell s 0 0 2496 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2496 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel comment s 2098 305 2098 305 0 FreeSans 200 90 0 0 no_jumper_check
flabel comment s 1542 328 1542 328 0 FreeSans 200 90 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfsbp_1
flabel comment s 208 233 208 233 0 FreeSans 200 90 0 0 no_jumper_check
flabel comment s 821 379 821 379 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 2496 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2496 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1183 464 1217 498 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2239 94 2273 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 168 2273 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 242 2273 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 316 2273 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 390 2273 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2431 94 2465 128 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2431 168 2465 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2431 242 2465 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2431 316 2465 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2431 390 2465 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2431 464 2465 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2431 538 2465 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2496 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2344728
string GDS_START 2325736
<< end >>
