magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 331 1478 704
<< pwell >>
rect 3 241 629 259
rect 3 49 1433 241
rect 0 0 1440 49
<< scnmos >>
rect 82 65 112 233
rect 168 65 198 233
rect 254 65 284 233
rect 348 65 378 233
rect 434 65 464 233
rect 520 65 550 233
rect 710 47 740 215
rect 796 47 826 215
rect 882 47 912 215
rect 968 47 998 215
rect 1062 47 1092 215
rect 1148 47 1178 215
rect 1234 47 1264 215
rect 1320 47 1350 215
<< scpmoshvt >>
rect 82 367 112 619
rect 168 367 198 619
rect 262 367 292 619
rect 348 367 378 619
rect 434 367 464 619
rect 520 367 550 619
rect 696 367 726 619
rect 782 367 812 619
rect 868 367 898 619
rect 954 367 984 619
rect 1069 367 1099 619
rect 1155 367 1185 619
rect 1241 367 1271 619
rect 1327 367 1357 619
<< ndiff >>
rect 29 192 82 233
rect 29 158 37 192
rect 71 158 82 192
rect 29 111 82 158
rect 29 77 37 111
rect 71 77 82 111
rect 29 65 82 77
rect 112 225 168 233
rect 112 191 123 225
rect 157 191 168 225
rect 112 153 168 191
rect 112 119 123 153
rect 157 119 168 153
rect 112 65 168 119
rect 198 179 254 233
rect 198 145 209 179
rect 243 145 254 179
rect 198 111 254 145
rect 198 77 209 111
rect 243 77 254 111
rect 198 65 254 77
rect 284 178 348 233
rect 284 144 303 178
rect 337 144 348 178
rect 284 65 348 144
rect 378 107 434 233
rect 378 73 389 107
rect 423 73 434 107
rect 378 65 434 73
rect 464 178 520 233
rect 464 144 475 178
rect 509 144 520 178
rect 464 65 520 144
rect 550 111 603 233
rect 550 77 561 111
rect 595 77 603 111
rect 550 65 603 77
rect 657 100 710 215
rect 657 66 665 100
rect 699 66 710 100
rect 657 47 710 66
rect 740 178 796 215
rect 740 144 751 178
rect 785 144 796 178
rect 740 47 796 144
rect 826 100 882 215
rect 826 66 837 100
rect 871 66 882 100
rect 826 47 882 66
rect 912 178 968 215
rect 912 144 923 178
rect 957 144 968 178
rect 912 47 968 144
rect 998 165 1062 215
rect 998 131 1013 165
rect 1047 131 1062 165
rect 998 97 1062 131
rect 998 63 1013 97
rect 1047 63 1062 97
rect 998 47 1062 63
rect 1092 203 1148 215
rect 1092 169 1103 203
rect 1137 169 1148 203
rect 1092 101 1148 169
rect 1092 67 1103 101
rect 1137 67 1148 101
rect 1092 47 1148 67
rect 1178 171 1234 215
rect 1178 137 1189 171
rect 1223 137 1234 171
rect 1178 89 1234 137
rect 1178 55 1189 89
rect 1223 55 1234 89
rect 1178 47 1234 55
rect 1264 203 1320 215
rect 1264 169 1275 203
rect 1309 169 1320 203
rect 1264 101 1320 169
rect 1264 67 1275 101
rect 1309 67 1320 101
rect 1264 47 1320 67
rect 1350 171 1407 215
rect 1350 137 1361 171
rect 1395 137 1407 171
rect 1350 89 1407 137
rect 1350 55 1361 89
rect 1395 55 1407 89
rect 1350 47 1407 55
<< pdiff >>
rect 29 607 82 619
rect 29 573 37 607
rect 71 573 82 607
rect 29 513 82 573
rect 29 479 37 513
rect 71 479 82 513
rect 29 425 82 479
rect 29 391 37 425
rect 71 391 82 425
rect 29 367 82 391
rect 112 599 168 619
rect 112 565 123 599
rect 157 565 168 599
rect 112 512 168 565
rect 112 478 123 512
rect 157 478 168 512
rect 112 413 168 478
rect 112 379 123 413
rect 157 379 168 413
rect 112 367 168 379
rect 198 607 262 619
rect 198 573 213 607
rect 247 573 262 607
rect 198 494 262 573
rect 198 460 213 494
rect 247 460 262 494
rect 198 367 262 460
rect 292 599 348 619
rect 292 565 303 599
rect 337 565 348 599
rect 292 504 348 565
rect 292 470 303 504
rect 337 470 348 504
rect 292 367 348 470
rect 378 536 434 619
rect 378 502 389 536
rect 423 502 434 536
rect 378 436 434 502
rect 378 402 389 436
rect 423 402 434 436
rect 378 367 434 402
rect 464 599 520 619
rect 464 565 475 599
rect 509 565 520 599
rect 464 504 520 565
rect 464 470 475 504
rect 509 470 520 504
rect 464 367 520 470
rect 550 607 696 619
rect 550 573 561 607
rect 595 573 651 607
rect 685 573 696 607
rect 550 494 696 573
rect 550 460 561 494
rect 595 460 651 494
rect 685 460 696 494
rect 550 367 696 460
rect 726 599 782 619
rect 726 565 737 599
rect 771 565 782 599
rect 726 504 782 565
rect 726 470 737 504
rect 771 470 782 504
rect 726 367 782 470
rect 812 538 868 619
rect 812 504 823 538
rect 857 504 868 538
rect 812 436 868 504
rect 812 402 823 436
rect 857 402 868 436
rect 812 367 868 402
rect 898 599 954 619
rect 898 565 909 599
rect 943 565 954 599
rect 898 506 954 565
rect 898 472 909 506
rect 943 472 954 506
rect 898 367 954 472
rect 984 607 1069 619
rect 984 573 1010 607
rect 1044 573 1069 607
rect 984 495 1069 573
rect 984 461 1010 495
rect 1044 461 1069 495
rect 984 367 1069 461
rect 1099 599 1155 619
rect 1099 565 1110 599
rect 1144 565 1155 599
rect 1099 503 1155 565
rect 1099 469 1110 503
rect 1144 469 1155 503
rect 1099 413 1155 469
rect 1099 379 1110 413
rect 1144 379 1155 413
rect 1099 367 1155 379
rect 1185 607 1241 619
rect 1185 573 1196 607
rect 1230 573 1241 607
rect 1185 526 1241 573
rect 1185 492 1196 526
rect 1230 492 1241 526
rect 1185 455 1241 492
rect 1185 421 1196 455
rect 1230 421 1241 455
rect 1185 367 1241 421
rect 1271 599 1327 619
rect 1271 565 1282 599
rect 1316 565 1327 599
rect 1271 503 1327 565
rect 1271 469 1282 503
rect 1316 469 1327 503
rect 1271 413 1327 469
rect 1271 379 1282 413
rect 1316 379 1327 413
rect 1271 367 1327 379
rect 1357 607 1410 619
rect 1357 573 1368 607
rect 1402 573 1410 607
rect 1357 526 1410 573
rect 1357 492 1368 526
rect 1402 492 1410 526
rect 1357 455 1410 492
rect 1357 421 1368 455
rect 1402 421 1410 455
rect 1357 367 1410 421
<< ndiffc >>
rect 37 158 71 192
rect 37 77 71 111
rect 123 191 157 225
rect 123 119 157 153
rect 209 145 243 179
rect 209 77 243 111
rect 303 144 337 178
rect 389 73 423 107
rect 475 144 509 178
rect 561 77 595 111
rect 665 66 699 100
rect 751 144 785 178
rect 837 66 871 100
rect 923 144 957 178
rect 1013 131 1047 165
rect 1013 63 1047 97
rect 1103 169 1137 203
rect 1103 67 1137 101
rect 1189 137 1223 171
rect 1189 55 1223 89
rect 1275 169 1309 203
rect 1275 67 1309 101
rect 1361 137 1395 171
rect 1361 55 1395 89
<< pdiffc >>
rect 37 573 71 607
rect 37 479 71 513
rect 37 391 71 425
rect 123 565 157 599
rect 123 478 157 512
rect 123 379 157 413
rect 213 573 247 607
rect 213 460 247 494
rect 303 565 337 599
rect 303 470 337 504
rect 389 502 423 536
rect 389 402 423 436
rect 475 565 509 599
rect 475 470 509 504
rect 561 573 595 607
rect 651 573 685 607
rect 561 460 595 494
rect 651 460 685 494
rect 737 565 771 599
rect 737 470 771 504
rect 823 504 857 538
rect 823 402 857 436
rect 909 565 943 599
rect 909 472 943 506
rect 1010 573 1044 607
rect 1010 461 1044 495
rect 1110 565 1144 599
rect 1110 469 1144 503
rect 1110 379 1144 413
rect 1196 573 1230 607
rect 1196 492 1230 526
rect 1196 421 1230 455
rect 1282 565 1316 599
rect 1282 469 1316 503
rect 1282 379 1316 413
rect 1368 573 1402 607
rect 1368 492 1402 526
rect 1368 421 1402 455
<< poly >>
rect 82 619 112 645
rect 168 619 198 645
rect 262 619 292 645
rect 348 619 378 645
rect 434 619 464 645
rect 520 619 550 645
rect 696 619 726 645
rect 782 619 812 645
rect 868 619 898 645
rect 954 619 984 645
rect 1069 619 1099 645
rect 1155 619 1185 645
rect 1241 619 1271 645
rect 1327 619 1357 645
rect 82 321 112 367
rect 168 321 198 367
rect 262 321 292 367
rect 348 335 378 367
rect 434 335 464 367
rect 21 305 198 321
rect 21 271 37 305
rect 71 271 198 305
rect 21 255 198 271
rect 240 305 306 321
rect 240 271 256 305
rect 290 271 306 305
rect 240 255 306 271
rect 348 319 464 335
rect 348 285 414 319
rect 448 285 464 319
rect 348 269 464 285
rect 82 233 112 255
rect 168 233 198 255
rect 254 233 284 255
rect 348 233 378 269
rect 434 233 464 269
rect 520 321 550 367
rect 520 305 631 321
rect 520 271 581 305
rect 615 271 631 305
rect 696 303 726 367
rect 782 335 812 367
rect 868 335 898 367
rect 782 319 898 335
rect 782 305 809 319
rect 520 255 631 271
rect 674 287 740 303
rect 520 233 550 255
rect 674 253 690 287
rect 724 253 740 287
rect 793 285 809 305
rect 843 299 898 319
rect 954 303 984 367
rect 1069 331 1099 367
rect 1155 331 1185 367
rect 1241 331 1271 367
rect 1327 331 1357 367
rect 1069 315 1357 331
rect 843 285 912 299
rect 793 269 912 285
rect 674 237 740 253
rect 710 215 740 237
rect 796 215 826 269
rect 882 215 912 269
rect 954 287 1020 303
rect 1069 295 1085 315
rect 954 253 970 287
rect 1004 253 1020 287
rect 954 237 1020 253
rect 1062 281 1085 295
rect 1119 281 1153 315
rect 1187 281 1221 315
rect 1255 281 1289 315
rect 1323 281 1357 315
rect 1062 265 1357 281
rect 968 215 998 237
rect 1062 215 1092 265
rect 1148 215 1178 265
rect 1234 215 1264 265
rect 1320 215 1350 265
rect 82 39 112 65
rect 168 39 198 65
rect 254 39 284 65
rect 348 39 378 65
rect 434 39 464 65
rect 520 39 550 65
rect 710 21 740 47
rect 796 21 826 47
rect 882 21 912 47
rect 968 21 998 47
rect 1062 21 1092 47
rect 1148 21 1178 47
rect 1234 21 1264 47
rect 1320 21 1350 47
<< polycont >>
rect 37 271 71 305
rect 256 271 290 305
rect 414 285 448 319
rect 581 271 615 305
rect 690 253 724 287
rect 809 285 843 319
rect 970 253 1004 287
rect 1085 281 1119 315
rect 1153 281 1187 315
rect 1221 281 1255 315
rect 1289 281 1323 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 21 607 87 649
rect 21 573 37 607
rect 71 573 87 607
rect 21 513 87 573
rect 21 479 37 513
rect 71 479 87 513
rect 21 425 87 479
rect 21 391 37 425
rect 71 391 87 425
rect 121 599 163 615
rect 121 565 123 599
rect 157 565 163 599
rect 121 512 163 565
rect 121 478 123 512
rect 157 478 163 512
rect 121 420 163 478
rect 197 607 263 649
rect 197 573 213 607
rect 247 573 263 607
rect 197 494 263 573
rect 197 460 213 494
rect 247 460 263 494
rect 197 454 263 460
rect 297 599 511 615
rect 297 565 303 599
rect 337 581 475 599
rect 337 565 339 581
rect 297 504 339 565
rect 473 565 475 581
rect 509 565 511 599
rect 297 470 303 504
rect 337 470 339 504
rect 297 454 339 470
rect 373 536 439 547
rect 373 502 389 536
rect 423 502 439 536
rect 373 436 439 502
rect 473 504 511 565
rect 473 470 475 504
rect 509 470 511 504
rect 473 454 511 470
rect 545 607 701 649
rect 545 573 561 607
rect 595 573 651 607
rect 685 573 701 607
rect 545 494 701 573
rect 545 460 561 494
rect 595 460 651 494
rect 685 460 701 494
rect 545 454 701 460
rect 735 599 959 615
rect 735 565 737 599
rect 771 581 909 599
rect 771 565 773 581
rect 735 504 773 565
rect 907 565 909 581
rect 943 565 959 599
rect 735 470 737 504
rect 771 470 773 504
rect 735 454 773 470
rect 807 538 873 547
rect 807 504 823 538
rect 857 504 873 538
rect 373 420 389 436
rect 121 413 389 420
rect 121 379 123 413
rect 157 402 389 413
rect 423 420 439 436
rect 807 436 873 504
rect 907 506 959 565
rect 907 472 909 506
rect 943 472 959 506
rect 907 456 959 472
rect 994 607 1060 649
rect 994 573 1010 607
rect 1044 573 1060 607
rect 994 495 1060 573
rect 994 461 1010 495
rect 1044 461 1060 495
rect 994 454 1060 461
rect 1108 599 1146 615
rect 1108 565 1110 599
rect 1144 565 1146 599
rect 1108 503 1146 565
rect 1108 469 1110 503
rect 1144 469 1146 503
rect 807 420 823 436
rect 423 402 823 420
rect 857 420 873 436
rect 857 402 1074 420
rect 157 386 1074 402
rect 157 379 173 386
rect 17 305 87 357
rect 17 271 37 305
rect 71 271 87 305
rect 17 270 87 271
rect 17 242 70 270
rect 121 229 173 379
rect 207 305 364 321
rect 207 271 256 305
rect 290 271 364 305
rect 398 319 547 352
rect 398 285 414 319
rect 448 285 547 319
rect 581 305 631 321
rect 207 249 364 271
rect 615 271 631 305
rect 772 319 859 352
rect 581 249 631 271
rect 207 242 631 249
rect 107 225 173 229
rect 21 192 73 208
rect 21 158 37 192
rect 71 158 73 192
rect 21 111 73 158
rect 107 191 123 225
rect 157 191 173 225
rect 319 215 631 242
rect 674 287 738 303
rect 674 253 690 287
rect 724 253 738 287
rect 772 285 809 319
rect 843 285 859 319
rect 1040 317 1074 386
rect 1108 413 1146 469
rect 1180 607 1246 649
rect 1180 573 1196 607
rect 1230 573 1246 607
rect 1180 526 1246 573
rect 1180 492 1196 526
rect 1230 492 1246 526
rect 1180 455 1246 492
rect 1180 421 1196 455
rect 1230 421 1246 455
rect 1280 599 1318 615
rect 1280 565 1282 599
rect 1316 565 1318 599
rect 1280 503 1318 565
rect 1280 469 1282 503
rect 1316 469 1318 503
rect 1108 379 1110 413
rect 1144 385 1146 413
rect 1280 413 1318 469
rect 1352 607 1418 649
rect 1352 573 1368 607
rect 1402 573 1418 607
rect 1352 526 1418 573
rect 1352 492 1368 526
rect 1402 492 1418 526
rect 1352 455 1418 492
rect 1352 421 1368 455
rect 1402 421 1418 455
rect 1280 385 1282 413
rect 1144 379 1282 385
rect 1316 385 1318 413
rect 1316 379 1423 385
rect 1108 351 1423 379
rect 1040 315 1339 317
rect 893 287 1006 303
rect 674 249 738 253
rect 893 253 970 287
rect 1004 253 1006 287
rect 1040 281 1085 315
rect 1119 281 1153 315
rect 1187 281 1221 315
rect 1255 281 1289 315
rect 1323 281 1339 315
rect 1040 277 1339 281
rect 893 249 1006 253
rect 674 215 1006 249
rect 1373 243 1423 351
rect 1093 209 1423 243
rect 1093 203 1139 209
rect 107 153 173 191
rect 107 119 123 153
rect 157 119 173 153
rect 207 179 253 195
rect 207 145 209 179
rect 243 145 253 179
rect 21 77 37 111
rect 71 85 73 111
rect 207 111 253 145
rect 287 178 973 181
rect 287 144 303 178
rect 337 144 475 178
rect 509 145 751 178
rect 509 144 529 145
rect 287 142 529 144
rect 627 144 751 145
rect 785 144 923 178
rect 957 144 973 178
rect 627 142 973 144
rect 1007 165 1059 181
rect 1007 131 1013 165
rect 1047 131 1059 165
rect 207 85 209 111
rect 71 77 209 85
rect 243 108 253 111
rect 545 108 561 111
rect 243 107 561 108
rect 243 77 389 107
rect 21 73 389 77
rect 423 77 561 107
rect 595 77 611 111
rect 423 73 611 77
rect 21 51 611 73
rect 649 100 715 108
rect 649 66 665 100
rect 699 66 715 100
rect 649 17 715 66
rect 821 100 887 108
rect 821 66 837 100
rect 871 66 887 100
rect 821 17 887 66
rect 1007 97 1059 131
rect 1007 63 1013 97
rect 1047 63 1059 97
rect 1007 17 1059 63
rect 1093 169 1103 203
rect 1137 169 1139 203
rect 1273 203 1311 209
rect 1093 101 1139 169
rect 1093 67 1103 101
rect 1137 67 1139 101
rect 1093 51 1139 67
rect 1173 171 1239 173
rect 1173 137 1189 171
rect 1223 137 1239 171
rect 1173 89 1239 137
rect 1173 55 1189 89
rect 1223 55 1239 89
rect 1173 17 1239 55
rect 1273 169 1275 203
rect 1309 169 1311 203
rect 1273 101 1311 169
rect 1273 67 1275 101
rect 1309 67 1311 101
rect 1273 51 1311 67
rect 1345 171 1411 175
rect 1345 137 1361 171
rect 1395 137 1411 171
rect 1345 89 1411 137
rect 1345 55 1361 89
rect 1395 55 1411 89
rect 1345 17 1411 55
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221a_4
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4920872
string GDS_START 4908574
<< end >>
