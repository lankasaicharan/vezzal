magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 27 49 651 167
rect 0 0 672 49
<< scnmos >>
rect 110 57 140 141
rect 188 57 218 141
rect 302 57 332 141
rect 374 57 404 141
rect 460 57 490 141
rect 538 57 568 141
<< scpmoshvt >>
rect 90 409 140 609
rect 196 409 246 609
rect 302 409 352 609
rect 538 396 588 596
<< ndiff >>
rect 53 116 110 141
rect 53 82 65 116
rect 99 82 110 116
rect 53 57 110 82
rect 140 57 188 141
rect 218 116 302 141
rect 218 82 257 116
rect 291 82 302 116
rect 218 57 302 82
rect 332 57 374 141
rect 404 103 460 141
rect 404 69 415 103
rect 449 69 460 103
rect 404 57 460 69
rect 490 57 538 141
rect 568 116 625 141
rect 568 82 579 116
rect 613 82 625 116
rect 568 57 625 82
<< pdiff >>
rect 33 597 90 609
rect 33 563 45 597
rect 79 563 90 597
rect 33 526 90 563
rect 33 492 45 526
rect 79 492 90 526
rect 33 455 90 492
rect 33 421 45 455
rect 79 421 90 455
rect 33 409 90 421
rect 140 597 196 609
rect 140 563 151 597
rect 185 563 196 597
rect 140 515 196 563
rect 140 481 151 515
rect 185 481 196 515
rect 140 409 196 481
rect 246 597 302 609
rect 246 563 257 597
rect 291 563 302 597
rect 246 526 302 563
rect 246 492 257 526
rect 291 492 302 526
rect 246 455 302 492
rect 246 421 257 455
rect 291 421 302 455
rect 246 409 302 421
rect 352 597 409 609
rect 352 563 363 597
rect 397 563 409 597
rect 352 526 409 563
rect 352 492 363 526
rect 397 492 409 526
rect 352 455 409 492
rect 352 421 363 455
rect 397 421 409 455
rect 352 409 409 421
rect 481 584 538 596
rect 481 550 493 584
rect 527 550 538 584
rect 481 513 538 550
rect 481 479 493 513
rect 527 479 538 513
rect 481 442 538 479
rect 481 408 493 442
rect 527 408 538 442
rect 481 396 538 408
rect 588 584 645 596
rect 588 550 599 584
rect 633 550 645 584
rect 588 513 645 550
rect 588 479 599 513
rect 633 479 645 513
rect 588 442 645 479
rect 588 408 599 442
rect 633 408 645 442
rect 588 396 645 408
<< ndiffc >>
rect 65 82 99 116
rect 257 82 291 116
rect 415 69 449 103
rect 579 82 613 116
<< pdiffc >>
rect 45 563 79 597
rect 45 492 79 526
rect 45 421 79 455
rect 151 563 185 597
rect 151 481 185 515
rect 257 563 291 597
rect 257 492 291 526
rect 257 421 291 455
rect 363 563 397 597
rect 363 492 397 526
rect 363 421 397 455
rect 493 550 527 584
rect 493 479 527 513
rect 493 408 527 442
rect 599 550 633 584
rect 599 479 633 513
rect 599 408 633 442
<< poly >>
rect 90 609 140 635
rect 196 609 246 635
rect 302 609 352 635
rect 538 596 588 622
rect 90 356 140 409
rect 196 359 246 409
rect 302 359 352 409
rect 44 340 140 356
rect 44 306 60 340
rect 94 306 140 340
rect 44 272 140 306
rect 44 238 60 272
rect 94 238 140 272
rect 44 222 140 238
rect 110 141 140 222
rect 188 343 254 359
rect 188 309 204 343
rect 238 309 254 343
rect 188 275 254 309
rect 188 241 204 275
rect 238 241 254 275
rect 188 225 254 241
rect 302 343 368 359
rect 302 309 318 343
rect 352 309 368 343
rect 302 275 368 309
rect 538 297 588 396
rect 302 241 318 275
rect 352 255 368 275
rect 460 281 588 297
rect 352 241 404 255
rect 302 225 404 241
rect 188 141 218 225
rect 302 141 332 225
rect 374 141 404 225
rect 460 247 476 281
rect 510 247 588 281
rect 460 225 588 247
rect 460 213 568 225
rect 460 179 476 213
rect 510 179 568 213
rect 460 163 568 179
rect 460 141 490 163
rect 538 141 568 163
rect 110 31 140 57
rect 188 31 218 57
rect 302 31 332 57
rect 374 31 404 57
rect 460 31 490 57
rect 538 31 568 57
<< polycont >>
rect 60 306 94 340
rect 60 238 94 272
rect 204 309 238 343
rect 204 241 238 275
rect 318 309 352 343
rect 318 241 352 275
rect 476 247 510 281
rect 476 179 510 213
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 29 597 95 613
rect 29 563 45 597
rect 79 563 95 597
rect 29 526 95 563
rect 29 492 45 526
rect 79 492 95 526
rect 29 455 95 492
rect 135 597 201 649
rect 135 563 151 597
rect 185 563 201 597
rect 135 515 201 563
rect 135 481 151 515
rect 185 481 201 515
rect 135 465 201 481
rect 241 597 307 613
rect 241 563 257 597
rect 291 563 307 597
rect 241 526 307 563
rect 241 492 257 526
rect 291 492 307 526
rect 29 421 45 455
rect 79 429 95 455
rect 241 455 307 492
rect 241 429 257 455
rect 79 421 257 429
rect 291 421 307 455
rect 29 395 307 421
rect 347 597 438 613
rect 347 563 363 597
rect 397 563 438 597
rect 347 526 438 563
rect 347 492 363 526
rect 397 492 438 526
rect 347 455 438 492
rect 347 421 363 455
rect 397 421 438 455
rect 347 405 438 421
rect 25 340 110 356
rect 25 306 60 340
rect 94 306 110 340
rect 25 272 110 306
rect 25 238 60 272
rect 94 238 110 272
rect 25 222 110 238
rect 188 343 263 359
rect 188 309 204 343
rect 238 309 263 343
rect 188 275 263 309
rect 188 241 204 275
rect 238 241 263 275
rect 188 225 263 241
rect 302 343 368 359
rect 302 309 318 343
rect 352 309 368 343
rect 302 275 368 309
rect 302 241 318 275
rect 352 241 368 275
rect 302 225 368 241
rect 404 297 438 405
rect 477 584 543 649
rect 477 550 493 584
rect 527 550 543 584
rect 477 513 543 550
rect 477 479 493 513
rect 527 479 543 513
rect 477 442 543 479
rect 477 408 493 442
rect 527 408 543 442
rect 477 392 543 408
rect 583 584 649 600
rect 583 550 599 584
rect 633 550 649 584
rect 583 513 649 550
rect 583 479 599 513
rect 633 479 649 513
rect 583 442 649 479
rect 583 408 599 442
rect 633 408 649 442
rect 583 356 649 408
rect 404 281 526 297
rect 404 247 476 281
rect 510 247 526 281
rect 404 213 526 247
rect 404 189 476 213
rect 241 179 476 189
rect 510 179 526 213
rect 241 155 526 179
rect 49 116 115 145
rect 49 82 65 116
rect 99 82 115 116
rect 49 17 115 82
rect 241 116 307 155
rect 241 82 257 116
rect 291 82 307 116
rect 241 53 307 82
rect 399 103 465 119
rect 399 69 415 103
rect 449 69 465 103
rect 399 17 465 69
rect 563 116 649 356
rect 563 82 579 116
rect 613 82 649 116
rect 563 53 649 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21o_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2597026
string GDS_START 2590312
<< end >>
