magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 6290 1975
<< nwell >>
rect -38 331 5030 704
rect 2346 269 4196 331
<< pwell >>
rect 314 241 424 267
rect 1 201 556 241
rect 1 49 3204 201
rect 4282 49 4800 241
rect 0 0 4992 49
<< scnmos >>
rect 84 47 114 215
rect 170 47 200 215
rect 288 47 318 215
rect 420 47 450 215
rect 641 47 671 175
rect 743 47 773 175
rect 829 47 859 175
rect 915 47 945 175
rect 1001 47 1031 175
rect 1103 47 1133 175
rect 1189 47 1219 175
rect 1307 47 1337 175
rect 1393 47 1423 175
rect 1479 47 1509 175
rect 1565 47 1595 175
rect 1651 47 1681 175
rect 1737 47 1767 175
rect 1823 47 1853 175
rect 1909 47 1939 175
rect 2011 47 2041 175
rect 2113 47 2143 175
rect 2215 47 2245 175
rect 2301 47 2331 175
rect 2387 47 2417 175
rect 2473 47 2503 175
rect 2559 47 2589 175
rect 2645 47 2675 175
rect 2731 47 2761 175
rect 2817 47 2847 175
rect 2903 47 2933 175
rect 2989 47 3019 175
rect 3075 47 3105 175
rect 4366 47 4396 215
rect 4467 47 4497 215
rect 4585 47 4615 215
rect 4671 47 4701 215
<< scpmos >>
rect 84 367 114 619
rect 170 367 200 619
rect 256 367 286 619
rect 342 367 372 619
rect 428 367 458 619
rect 514 367 544 619
rect 600 367 630 619
rect 686 367 716 619
rect 772 367 802 619
rect 858 367 888 619
rect 944 367 974 619
rect 1030 367 1060 619
rect 1116 367 1146 619
rect 1202 367 1232 619
rect 1288 367 1318 619
rect 1374 367 1404 619
rect 1460 367 1490 619
rect 1546 367 1576 619
rect 1636 367 1666 619
rect 1722 367 1752 619
rect 1808 367 1838 619
rect 1894 367 1924 619
rect 1980 367 2010 619
rect 2066 367 2096 619
rect 2152 367 2182 619
rect 2238 367 2268 619
rect 2439 305 2469 557
rect 2525 305 2555 557
rect 2611 305 2641 557
rect 2697 305 2727 557
rect 2783 305 2813 557
rect 2869 305 2899 557
rect 2955 305 2985 557
rect 3041 305 3071 557
rect 3127 305 3157 557
rect 3213 305 3243 557
rect 3299 305 3329 557
rect 3385 305 3415 557
rect 3471 305 3501 557
rect 3557 305 3587 557
rect 3643 305 3673 557
rect 3729 305 3759 557
rect 3815 305 3845 557
rect 3901 305 3931 557
rect 3987 305 4017 557
rect 4073 305 4103 557
rect 4271 367 4301 619
rect 4357 367 4387 619
rect 4443 367 4473 619
rect 4529 367 4559 619
rect 4615 367 4645 619
rect 4701 367 4731 619
rect 4792 367 4822 619
rect 4878 367 4908 619
<< ndiff >>
rect 340 229 398 241
rect 340 215 352 229
rect 27 184 84 215
rect 27 150 39 184
rect 73 150 84 184
rect 27 93 84 150
rect 27 59 39 93
rect 73 59 84 93
rect 27 47 84 59
rect 114 203 170 215
rect 114 169 125 203
rect 159 169 170 203
rect 114 103 170 169
rect 114 69 125 103
rect 159 69 170 103
rect 114 47 170 69
rect 200 89 288 215
rect 200 55 227 89
rect 261 55 288 89
rect 200 47 288 55
rect 318 195 352 215
rect 386 215 398 229
rect 386 195 420 215
rect 318 47 420 195
rect 450 73 530 215
rect 450 47 484 73
rect 215 43 273 47
rect 472 39 484 47
rect 518 39 530 73
rect 584 126 641 175
rect 584 92 596 126
rect 630 92 641 126
rect 584 47 641 92
rect 671 94 743 175
rect 671 60 698 94
rect 732 60 743 94
rect 671 47 743 60
rect 773 126 829 175
rect 773 92 784 126
rect 818 92 829 126
rect 773 47 829 92
rect 859 94 915 175
rect 859 60 870 94
rect 904 60 915 94
rect 859 47 915 60
rect 945 126 1001 175
rect 945 92 956 126
rect 990 92 1001 126
rect 945 47 1001 92
rect 1031 94 1103 175
rect 1031 60 1042 94
rect 1076 60 1103 94
rect 1031 47 1103 60
rect 1133 126 1189 175
rect 1133 92 1144 126
rect 1178 92 1189 126
rect 1133 47 1189 92
rect 1219 94 1307 175
rect 1219 60 1246 94
rect 1280 60 1307 94
rect 1219 47 1307 60
rect 1337 133 1393 175
rect 1337 99 1348 133
rect 1382 99 1393 133
rect 1337 47 1393 99
rect 1423 120 1479 175
rect 1423 86 1434 120
rect 1468 86 1479 120
rect 1423 47 1479 86
rect 1509 133 1565 175
rect 1509 99 1520 133
rect 1554 99 1565 133
rect 1509 47 1565 99
rect 1595 120 1651 175
rect 1595 86 1606 120
rect 1640 86 1651 120
rect 1595 47 1651 86
rect 1681 133 1737 175
rect 1681 99 1692 133
rect 1726 99 1737 133
rect 1681 47 1737 99
rect 1767 120 1823 175
rect 1767 86 1778 120
rect 1812 86 1823 120
rect 1767 47 1823 86
rect 1853 133 1909 175
rect 1853 99 1864 133
rect 1898 99 1909 133
rect 1853 47 1909 99
rect 1939 167 2011 175
rect 1939 133 1966 167
rect 2000 133 2011 167
rect 1939 47 2011 133
rect 2041 93 2113 175
rect 2041 59 2068 93
rect 2102 59 2113 93
rect 2041 47 2113 59
rect 2143 167 2215 175
rect 2143 133 2170 167
rect 2204 133 2215 167
rect 2143 47 2215 133
rect 2245 93 2301 175
rect 2245 59 2256 93
rect 2290 59 2301 93
rect 2245 47 2301 59
rect 2331 163 2387 175
rect 2331 129 2342 163
rect 2376 129 2387 163
rect 2331 47 2387 129
rect 2417 93 2473 175
rect 2417 59 2428 93
rect 2462 59 2473 93
rect 2417 47 2473 59
rect 2503 163 2559 175
rect 2503 129 2514 163
rect 2548 129 2559 163
rect 2503 47 2559 129
rect 2589 93 2645 175
rect 2589 59 2600 93
rect 2634 59 2645 93
rect 2589 47 2645 59
rect 2675 163 2731 175
rect 2675 129 2686 163
rect 2720 129 2731 163
rect 2675 47 2731 129
rect 2761 93 2817 175
rect 2761 59 2772 93
rect 2806 59 2817 93
rect 2761 47 2817 59
rect 2847 163 2903 175
rect 2847 129 2858 163
rect 2892 129 2903 163
rect 2847 47 2903 129
rect 2933 93 2989 175
rect 2933 59 2944 93
rect 2978 59 2989 93
rect 2933 47 2989 59
rect 3019 163 3075 175
rect 3019 129 3030 163
rect 3064 129 3075 163
rect 3019 47 3075 129
rect 3105 124 3178 175
rect 3105 90 3132 124
rect 3166 90 3178 124
rect 3105 47 3178 90
rect 4308 103 4366 215
rect 4308 69 4320 103
rect 4354 69 4366 103
rect 4308 47 4366 69
rect 4396 184 4467 215
rect 4396 150 4422 184
rect 4456 150 4467 184
rect 4396 93 4467 150
rect 4396 59 4422 93
rect 4456 59 4467 93
rect 4396 47 4467 59
rect 4497 103 4585 215
rect 4497 69 4524 103
rect 4558 69 4585 103
rect 4497 47 4585 69
rect 4615 184 4671 215
rect 4615 150 4626 184
rect 4660 150 4671 184
rect 4615 103 4671 150
rect 4615 69 4626 103
rect 4660 69 4671 103
rect 4615 47 4671 69
rect 4701 184 4774 215
rect 4701 150 4728 184
rect 4762 150 4774 184
rect 4701 93 4774 150
rect 4701 59 4728 93
rect 4762 59 4774 93
rect 4701 47 4774 59
rect 472 27 530 39
<< pdiff >>
rect 27 607 84 619
rect 27 573 39 607
rect 73 573 84 607
rect 27 510 84 573
rect 27 476 39 510
rect 73 476 84 510
rect 27 413 84 476
rect 27 379 39 413
rect 73 379 84 413
rect 27 367 84 379
rect 114 597 170 619
rect 114 563 125 597
rect 159 563 170 597
rect 114 505 170 563
rect 114 471 125 505
rect 159 471 170 505
rect 114 413 170 471
rect 114 379 125 413
rect 159 379 170 413
rect 114 367 170 379
rect 200 607 256 619
rect 200 573 211 607
rect 245 573 256 607
rect 200 510 256 573
rect 200 476 211 510
rect 245 476 256 510
rect 200 413 256 476
rect 200 379 211 413
rect 245 379 256 413
rect 200 367 256 379
rect 286 597 342 619
rect 286 563 297 597
rect 331 563 342 597
rect 286 505 342 563
rect 286 471 297 505
rect 331 471 342 505
rect 286 413 342 471
rect 286 379 297 413
rect 331 379 342 413
rect 286 367 342 379
rect 372 607 428 619
rect 372 573 383 607
rect 417 573 428 607
rect 372 483 428 573
rect 372 449 383 483
rect 417 449 428 483
rect 372 367 428 449
rect 458 597 514 619
rect 458 563 469 597
rect 503 563 514 597
rect 458 505 514 563
rect 458 471 469 505
rect 503 471 514 505
rect 458 413 514 471
rect 458 379 469 413
rect 503 379 514 413
rect 458 367 514 379
rect 544 607 600 619
rect 544 573 555 607
rect 589 573 600 607
rect 544 514 600 573
rect 544 480 555 514
rect 589 480 600 514
rect 544 421 600 480
rect 544 387 555 421
rect 589 387 600 421
rect 544 367 600 387
rect 630 537 686 619
rect 630 503 641 537
rect 675 503 686 537
rect 630 423 686 503
rect 630 389 641 423
rect 675 389 686 423
rect 630 367 686 389
rect 716 611 772 619
rect 716 577 727 611
rect 761 577 772 611
rect 716 491 772 577
rect 716 457 727 491
rect 761 457 772 491
rect 716 367 772 457
rect 802 537 858 619
rect 802 503 813 537
rect 847 503 858 537
rect 802 423 858 503
rect 802 389 813 423
rect 847 389 858 423
rect 802 367 858 389
rect 888 611 944 619
rect 888 577 899 611
rect 933 577 944 611
rect 888 491 944 577
rect 888 457 899 491
rect 933 457 944 491
rect 888 367 944 457
rect 974 537 1030 619
rect 974 503 985 537
rect 1019 503 1030 537
rect 974 423 1030 503
rect 974 389 985 423
rect 1019 389 1030 423
rect 974 367 1030 389
rect 1060 611 1116 619
rect 1060 577 1071 611
rect 1105 577 1116 611
rect 1060 491 1116 577
rect 1060 457 1071 491
rect 1105 457 1116 491
rect 1060 367 1116 457
rect 1146 537 1202 619
rect 1146 503 1157 537
rect 1191 503 1202 537
rect 1146 423 1202 503
rect 1146 389 1157 423
rect 1191 389 1202 423
rect 1146 367 1202 389
rect 1232 611 1288 619
rect 1232 577 1243 611
rect 1277 577 1288 611
rect 1232 491 1288 577
rect 1232 457 1243 491
rect 1277 457 1288 491
rect 1232 367 1288 457
rect 1318 537 1374 619
rect 1318 503 1329 537
rect 1363 503 1374 537
rect 1318 423 1374 503
rect 1318 389 1329 423
rect 1363 389 1374 423
rect 1318 367 1374 389
rect 1404 611 1460 619
rect 1404 577 1415 611
rect 1449 577 1460 611
rect 1404 491 1460 577
rect 1404 457 1415 491
rect 1449 457 1460 491
rect 1404 367 1460 457
rect 1490 537 1546 619
rect 1490 503 1501 537
rect 1535 503 1546 537
rect 1490 423 1546 503
rect 1490 389 1501 423
rect 1535 389 1546 423
rect 1490 367 1546 389
rect 1576 611 1636 619
rect 1576 577 1587 611
rect 1621 577 1636 611
rect 1576 491 1636 577
rect 1576 457 1587 491
rect 1621 457 1636 491
rect 1576 367 1636 457
rect 1666 537 1722 619
rect 1666 503 1677 537
rect 1711 503 1722 537
rect 1666 423 1722 503
rect 1666 389 1677 423
rect 1711 389 1722 423
rect 1666 367 1722 389
rect 1752 611 1808 619
rect 1752 577 1763 611
rect 1797 577 1808 611
rect 1752 491 1808 577
rect 1752 457 1763 491
rect 1797 457 1808 491
rect 1752 367 1808 457
rect 1838 537 1894 619
rect 1838 503 1849 537
rect 1883 503 1894 537
rect 1838 423 1894 503
rect 1838 389 1849 423
rect 1883 389 1894 423
rect 1838 367 1894 389
rect 1924 611 1980 619
rect 1924 577 1935 611
rect 1969 577 1980 611
rect 1924 491 1980 577
rect 1924 457 1935 491
rect 1969 457 1980 491
rect 1924 367 1980 457
rect 2010 597 2066 619
rect 2010 563 2021 597
rect 2055 563 2066 597
rect 2010 505 2066 563
rect 2010 471 2021 505
rect 2055 471 2066 505
rect 2010 413 2066 471
rect 2010 379 2021 413
rect 2055 379 2066 413
rect 2010 367 2066 379
rect 2096 607 2152 619
rect 2096 573 2107 607
rect 2141 573 2152 607
rect 2096 510 2152 573
rect 2096 476 2107 510
rect 2141 476 2152 510
rect 2096 413 2152 476
rect 2096 379 2107 413
rect 2141 379 2152 413
rect 2096 367 2152 379
rect 2182 597 2238 619
rect 2182 563 2193 597
rect 2227 563 2238 597
rect 2182 505 2238 563
rect 2182 471 2193 505
rect 2227 471 2238 505
rect 2182 413 2238 471
rect 2182 379 2193 413
rect 2227 379 2238 413
rect 2182 367 2238 379
rect 2268 607 2325 619
rect 2268 573 2279 607
rect 2313 573 2325 607
rect 4214 607 4271 619
rect 2268 523 2325 573
rect 4214 573 4226 607
rect 4260 573 4271 607
rect 2268 489 2279 523
rect 2313 489 2325 523
rect 2268 367 2325 489
rect 2382 351 2439 557
rect 2382 317 2394 351
rect 2428 317 2439 351
rect 2382 305 2439 317
rect 2469 545 2525 557
rect 2469 511 2480 545
rect 2514 511 2525 545
rect 2469 442 2525 511
rect 2469 408 2480 442
rect 2514 408 2525 442
rect 2469 305 2525 408
rect 2555 527 2611 557
rect 2555 493 2566 527
rect 2600 493 2611 527
rect 2555 439 2611 493
rect 2555 405 2566 439
rect 2600 405 2611 439
rect 2555 351 2611 405
rect 2555 317 2566 351
rect 2600 317 2611 351
rect 2555 305 2611 317
rect 2641 549 2697 557
rect 2641 515 2652 549
rect 2686 515 2697 549
rect 2641 481 2697 515
rect 2641 447 2652 481
rect 2686 447 2697 481
rect 2641 413 2697 447
rect 2641 379 2652 413
rect 2686 379 2697 413
rect 2641 305 2697 379
rect 2727 527 2783 557
rect 2727 493 2738 527
rect 2772 493 2783 527
rect 2727 439 2783 493
rect 2727 405 2738 439
rect 2772 405 2783 439
rect 2727 351 2783 405
rect 2727 317 2738 351
rect 2772 317 2783 351
rect 2727 305 2783 317
rect 2813 549 2869 557
rect 2813 515 2824 549
rect 2858 515 2869 549
rect 2813 481 2869 515
rect 2813 447 2824 481
rect 2858 447 2869 481
rect 2813 413 2869 447
rect 2813 379 2824 413
rect 2858 379 2869 413
rect 2813 305 2869 379
rect 2899 527 2955 557
rect 2899 493 2910 527
rect 2944 493 2955 527
rect 2899 439 2955 493
rect 2899 405 2910 439
rect 2944 405 2955 439
rect 2899 351 2955 405
rect 2899 317 2910 351
rect 2944 317 2955 351
rect 2899 305 2955 317
rect 2985 549 3041 557
rect 2985 515 2996 549
rect 3030 515 3041 549
rect 2985 481 3041 515
rect 2985 447 2996 481
rect 3030 447 3041 481
rect 2985 413 3041 447
rect 2985 379 2996 413
rect 3030 379 3041 413
rect 2985 305 3041 379
rect 3071 527 3127 557
rect 3071 493 3082 527
rect 3116 493 3127 527
rect 3071 439 3127 493
rect 3071 405 3082 439
rect 3116 405 3127 439
rect 3071 351 3127 405
rect 3071 317 3082 351
rect 3116 317 3127 351
rect 3071 305 3127 317
rect 3157 549 3213 557
rect 3157 515 3168 549
rect 3202 515 3213 549
rect 3157 481 3213 515
rect 3157 447 3168 481
rect 3202 447 3213 481
rect 3157 413 3213 447
rect 3157 379 3168 413
rect 3202 379 3213 413
rect 3157 305 3213 379
rect 3243 527 3299 557
rect 3243 493 3254 527
rect 3288 493 3299 527
rect 3243 439 3299 493
rect 3243 405 3254 439
rect 3288 405 3299 439
rect 3243 351 3299 405
rect 3243 317 3254 351
rect 3288 317 3299 351
rect 3243 305 3299 317
rect 3329 549 3385 557
rect 3329 515 3340 549
rect 3374 515 3385 549
rect 3329 481 3385 515
rect 3329 447 3340 481
rect 3374 447 3385 481
rect 3329 413 3385 447
rect 3329 379 3340 413
rect 3374 379 3385 413
rect 3329 305 3385 379
rect 3415 527 3471 557
rect 3415 493 3426 527
rect 3460 493 3471 527
rect 3415 439 3471 493
rect 3415 405 3426 439
rect 3460 405 3471 439
rect 3415 351 3471 405
rect 3415 317 3426 351
rect 3460 317 3471 351
rect 3415 305 3471 317
rect 3501 549 3557 557
rect 3501 515 3512 549
rect 3546 515 3557 549
rect 3501 481 3557 515
rect 3501 447 3512 481
rect 3546 447 3557 481
rect 3501 413 3557 447
rect 3501 379 3512 413
rect 3546 379 3557 413
rect 3501 305 3557 379
rect 3587 527 3643 557
rect 3587 493 3598 527
rect 3632 493 3643 527
rect 3587 439 3643 493
rect 3587 405 3598 439
rect 3632 405 3643 439
rect 3587 351 3643 405
rect 3587 317 3598 351
rect 3632 317 3643 351
rect 3587 305 3643 317
rect 3673 549 3729 557
rect 3673 515 3684 549
rect 3718 515 3729 549
rect 3673 481 3729 515
rect 3673 447 3684 481
rect 3718 447 3729 481
rect 3673 413 3729 447
rect 3673 379 3684 413
rect 3718 379 3729 413
rect 3673 305 3729 379
rect 3759 527 3815 557
rect 3759 493 3770 527
rect 3804 493 3815 527
rect 3759 439 3815 493
rect 3759 405 3770 439
rect 3804 405 3815 439
rect 3759 351 3815 405
rect 3759 317 3770 351
rect 3804 317 3815 351
rect 3759 305 3815 317
rect 3845 549 3901 557
rect 3845 515 3856 549
rect 3890 515 3901 549
rect 3845 481 3901 515
rect 3845 447 3856 481
rect 3890 447 3901 481
rect 3845 413 3901 447
rect 3845 379 3856 413
rect 3890 379 3901 413
rect 3845 305 3901 379
rect 3931 527 3987 557
rect 3931 493 3942 527
rect 3976 493 3987 527
rect 3931 439 3987 493
rect 3931 405 3942 439
rect 3976 405 3987 439
rect 3931 351 3987 405
rect 3931 317 3942 351
rect 3976 317 3987 351
rect 3931 305 3987 317
rect 4017 549 4073 557
rect 4017 515 4028 549
rect 4062 515 4073 549
rect 4017 481 4073 515
rect 4017 447 4028 481
rect 4062 447 4073 481
rect 4017 413 4073 447
rect 4017 379 4028 413
rect 4062 379 4073 413
rect 4017 305 4073 379
rect 4103 545 4160 557
rect 4103 511 4114 545
rect 4148 511 4160 545
rect 4103 448 4160 511
rect 4103 414 4114 448
rect 4148 414 4160 448
rect 4103 351 4160 414
rect 4214 510 4271 573
rect 4214 476 4226 510
rect 4260 476 4271 510
rect 4214 413 4271 476
rect 4214 379 4226 413
rect 4260 379 4271 413
rect 4214 367 4271 379
rect 4301 597 4357 619
rect 4301 563 4312 597
rect 4346 563 4357 597
rect 4301 505 4357 563
rect 4301 471 4312 505
rect 4346 471 4357 505
rect 4301 413 4357 471
rect 4301 379 4312 413
rect 4346 379 4357 413
rect 4301 367 4357 379
rect 4387 607 4443 619
rect 4387 573 4398 607
rect 4432 573 4443 607
rect 4387 483 4443 573
rect 4387 449 4398 483
rect 4432 449 4443 483
rect 4387 367 4443 449
rect 4473 597 4529 619
rect 4473 563 4484 597
rect 4518 563 4529 597
rect 4473 505 4529 563
rect 4473 471 4484 505
rect 4518 471 4529 505
rect 4473 413 4529 471
rect 4473 379 4484 413
rect 4518 379 4529 413
rect 4473 367 4529 379
rect 4559 607 4615 619
rect 4559 573 4570 607
rect 4604 573 4615 607
rect 4559 533 4615 573
rect 4559 499 4570 533
rect 4604 499 4615 533
rect 4559 459 4615 499
rect 4559 425 4570 459
rect 4604 425 4615 459
rect 4559 367 4615 425
rect 4645 597 4701 619
rect 4645 563 4656 597
rect 4690 563 4701 597
rect 4645 505 4701 563
rect 4645 471 4656 505
rect 4690 471 4701 505
rect 4645 413 4701 471
rect 4645 379 4656 413
rect 4690 379 4701 413
rect 4645 367 4701 379
rect 4731 607 4792 619
rect 4731 573 4742 607
rect 4776 573 4792 607
rect 4731 533 4792 573
rect 4731 499 4742 533
rect 4776 499 4792 533
rect 4731 459 4792 499
rect 4731 425 4742 459
rect 4776 425 4792 459
rect 4731 367 4792 425
rect 4822 597 4878 619
rect 4822 563 4833 597
rect 4867 563 4878 597
rect 4822 505 4878 563
rect 4822 471 4833 505
rect 4867 471 4878 505
rect 4822 413 4878 471
rect 4822 379 4833 413
rect 4867 379 4878 413
rect 4822 367 4878 379
rect 4908 607 4965 619
rect 4908 573 4919 607
rect 4953 573 4965 607
rect 4908 510 4965 573
rect 4908 476 4919 510
rect 4953 476 4965 510
rect 4908 413 4965 476
rect 4908 379 4919 413
rect 4953 379 4965 413
rect 4908 367 4965 379
rect 4103 317 4114 351
rect 4148 317 4160 351
rect 4103 305 4160 317
<< ndiffc >>
rect 39 150 73 184
rect 39 59 73 93
rect 125 169 159 203
rect 125 69 159 103
rect 227 55 261 89
rect 352 195 386 229
rect 484 39 518 73
rect 596 92 630 126
rect 698 60 732 94
rect 784 92 818 126
rect 870 60 904 94
rect 956 92 990 126
rect 1042 60 1076 94
rect 1144 92 1178 126
rect 1246 60 1280 94
rect 1348 99 1382 133
rect 1434 86 1468 120
rect 1520 99 1554 133
rect 1606 86 1640 120
rect 1692 99 1726 133
rect 1778 86 1812 120
rect 1864 99 1898 133
rect 1966 133 2000 167
rect 2068 59 2102 93
rect 2170 133 2204 167
rect 2256 59 2290 93
rect 2342 129 2376 163
rect 2428 59 2462 93
rect 2514 129 2548 163
rect 2600 59 2634 93
rect 2686 129 2720 163
rect 2772 59 2806 93
rect 2858 129 2892 163
rect 2944 59 2978 93
rect 3030 129 3064 163
rect 3132 90 3166 124
rect 4320 69 4354 103
rect 4422 150 4456 184
rect 4422 59 4456 93
rect 4524 69 4558 103
rect 4626 150 4660 184
rect 4626 69 4660 103
rect 4728 150 4762 184
rect 4728 59 4762 93
<< pdiffc >>
rect 39 573 73 607
rect 39 476 73 510
rect 39 379 73 413
rect 125 563 159 597
rect 125 471 159 505
rect 125 379 159 413
rect 211 573 245 607
rect 211 476 245 510
rect 211 379 245 413
rect 297 563 331 597
rect 297 471 331 505
rect 297 379 331 413
rect 383 573 417 607
rect 383 449 417 483
rect 469 563 503 597
rect 469 471 503 505
rect 469 379 503 413
rect 555 573 589 607
rect 555 480 589 514
rect 555 387 589 421
rect 641 503 675 537
rect 641 389 675 423
rect 727 577 761 611
rect 727 457 761 491
rect 813 503 847 537
rect 813 389 847 423
rect 899 577 933 611
rect 899 457 933 491
rect 985 503 1019 537
rect 985 389 1019 423
rect 1071 577 1105 611
rect 1071 457 1105 491
rect 1157 503 1191 537
rect 1157 389 1191 423
rect 1243 577 1277 611
rect 1243 457 1277 491
rect 1329 503 1363 537
rect 1329 389 1363 423
rect 1415 577 1449 611
rect 1415 457 1449 491
rect 1501 503 1535 537
rect 1501 389 1535 423
rect 1587 577 1621 611
rect 1587 457 1621 491
rect 1677 503 1711 537
rect 1677 389 1711 423
rect 1763 577 1797 611
rect 1763 457 1797 491
rect 1849 503 1883 537
rect 1849 389 1883 423
rect 1935 577 1969 611
rect 1935 457 1969 491
rect 2021 563 2055 597
rect 2021 471 2055 505
rect 2021 379 2055 413
rect 2107 573 2141 607
rect 2107 476 2141 510
rect 2107 379 2141 413
rect 2193 563 2227 597
rect 2193 471 2227 505
rect 2193 379 2227 413
rect 2279 573 2313 607
rect 4226 573 4260 607
rect 2279 489 2313 523
rect 2394 317 2428 351
rect 2480 511 2514 545
rect 2480 408 2514 442
rect 2566 493 2600 527
rect 2566 405 2600 439
rect 2566 317 2600 351
rect 2652 515 2686 549
rect 2652 447 2686 481
rect 2652 379 2686 413
rect 2738 493 2772 527
rect 2738 405 2772 439
rect 2738 317 2772 351
rect 2824 515 2858 549
rect 2824 447 2858 481
rect 2824 379 2858 413
rect 2910 493 2944 527
rect 2910 405 2944 439
rect 2910 317 2944 351
rect 2996 515 3030 549
rect 2996 447 3030 481
rect 2996 379 3030 413
rect 3082 493 3116 527
rect 3082 405 3116 439
rect 3082 317 3116 351
rect 3168 515 3202 549
rect 3168 447 3202 481
rect 3168 379 3202 413
rect 3254 493 3288 527
rect 3254 405 3288 439
rect 3254 317 3288 351
rect 3340 515 3374 549
rect 3340 447 3374 481
rect 3340 379 3374 413
rect 3426 493 3460 527
rect 3426 405 3460 439
rect 3426 317 3460 351
rect 3512 515 3546 549
rect 3512 447 3546 481
rect 3512 379 3546 413
rect 3598 493 3632 527
rect 3598 405 3632 439
rect 3598 317 3632 351
rect 3684 515 3718 549
rect 3684 447 3718 481
rect 3684 379 3718 413
rect 3770 493 3804 527
rect 3770 405 3804 439
rect 3770 317 3804 351
rect 3856 515 3890 549
rect 3856 447 3890 481
rect 3856 379 3890 413
rect 3942 493 3976 527
rect 3942 405 3976 439
rect 3942 317 3976 351
rect 4028 515 4062 549
rect 4028 447 4062 481
rect 4028 379 4062 413
rect 4114 511 4148 545
rect 4114 414 4148 448
rect 4226 476 4260 510
rect 4226 379 4260 413
rect 4312 563 4346 597
rect 4312 471 4346 505
rect 4312 379 4346 413
rect 4398 573 4432 607
rect 4398 449 4432 483
rect 4484 563 4518 597
rect 4484 471 4518 505
rect 4484 379 4518 413
rect 4570 573 4604 607
rect 4570 499 4604 533
rect 4570 425 4604 459
rect 4656 563 4690 597
rect 4656 471 4690 505
rect 4656 379 4690 413
rect 4742 573 4776 607
rect 4742 499 4776 533
rect 4742 425 4776 459
rect 4833 563 4867 597
rect 4833 471 4867 505
rect 4833 379 4867 413
rect 4919 573 4953 607
rect 4919 476 4953 510
rect 4919 379 4953 413
rect 4114 317 4148 351
<< poly >>
rect 84 619 114 645
rect 170 619 200 645
rect 256 619 286 645
rect 342 619 372 645
rect 428 619 458 645
rect 514 619 544 645
rect 600 619 630 645
rect 686 619 716 645
rect 772 619 802 645
rect 858 619 888 645
rect 944 619 974 645
rect 1030 619 1060 645
rect 1116 619 1146 645
rect 1202 619 1232 645
rect 1288 619 1318 645
rect 1374 619 1404 645
rect 1460 619 1490 645
rect 1546 619 1576 645
rect 1636 619 1666 645
rect 1722 619 1752 645
rect 1808 619 1838 645
rect 1894 619 1924 645
rect 1980 619 2010 645
rect 2066 619 2096 645
rect 2152 619 2182 645
rect 2238 619 2268 645
rect 4271 619 4301 645
rect 4357 619 4387 645
rect 4443 619 4473 645
rect 4529 619 4559 645
rect 4615 619 4645 645
rect 4701 619 4731 645
rect 4792 619 4822 645
rect 4878 619 4908 645
rect 2439 557 2469 583
rect 2525 557 2555 583
rect 2611 557 2641 583
rect 2697 557 2727 583
rect 2783 557 2813 583
rect 2869 557 2899 583
rect 2955 557 2985 583
rect 3041 557 3071 583
rect 3127 557 3157 583
rect 3213 557 3243 583
rect 3299 557 3329 583
rect 3385 557 3415 583
rect 3471 557 3501 583
rect 3557 557 3587 583
rect 3643 557 3673 583
rect 3729 557 3759 583
rect 3815 557 3845 583
rect 3901 557 3931 583
rect 3987 557 4017 583
rect 4073 557 4103 583
rect 84 303 114 367
rect 23 287 114 303
rect 23 253 39 287
rect 73 267 114 287
rect 170 267 200 367
rect 256 297 286 367
rect 342 297 372 367
rect 428 297 458 367
rect 514 297 544 367
rect 600 345 630 367
rect 686 345 716 367
rect 772 345 802 367
rect 858 345 888 367
rect 944 345 974 367
rect 1030 345 1060 367
rect 1116 345 1146 367
rect 1202 345 1232 367
rect 1288 345 1318 367
rect 1374 345 1404 367
rect 1460 345 1490 367
rect 1546 345 1576 367
rect 1636 345 1666 367
rect 1722 345 1752 367
rect 1808 345 1838 367
rect 1894 345 1924 367
rect 1980 345 2010 367
rect 2066 345 2096 367
rect 2152 345 2182 367
rect 2238 345 2268 367
rect 600 319 2268 345
rect 600 315 1294 319
rect 256 267 544 297
rect 1278 285 1294 315
rect 1328 285 1362 319
rect 1396 285 1430 319
rect 1464 285 1498 319
rect 1532 285 1566 319
rect 1600 285 1634 319
rect 1668 285 1702 319
rect 1736 285 1770 319
rect 1804 285 1838 319
rect 1872 285 1906 319
rect 1940 315 2268 319
rect 1940 285 1956 315
rect 4271 341 4301 367
rect 4357 341 4387 367
rect 4271 311 4387 341
rect 1278 269 1956 285
rect 73 253 200 267
rect 23 237 200 253
rect 84 215 114 237
rect 170 215 200 237
rect 288 215 318 267
rect 420 215 450 267
rect 514 251 1230 267
rect 2439 265 2469 305
rect 2525 265 2555 305
rect 2611 265 2641 305
rect 2697 265 2727 305
rect 2783 265 2813 305
rect 2869 265 2899 305
rect 2955 265 2985 305
rect 3041 265 3071 305
rect 3127 265 3157 305
rect 3213 265 3243 305
rect 3299 265 3329 305
rect 3385 265 3415 305
rect 3471 265 3501 305
rect 3557 265 3587 305
rect 3643 265 3673 305
rect 3729 265 3759 305
rect 514 237 568 251
rect 552 217 568 237
rect 602 217 636 251
rect 670 217 704 251
rect 738 217 772 251
rect 806 217 840 251
rect 874 217 908 251
rect 942 217 976 251
rect 1010 217 1044 251
rect 1078 217 1112 251
rect 1146 217 1180 251
rect 1214 227 1230 251
rect 2387 263 3759 265
rect 3815 263 3845 305
rect 3901 263 3931 305
rect 3987 263 4017 305
rect 4073 263 4103 305
rect 4357 303 4387 311
rect 4443 303 4473 367
rect 4529 303 4559 367
rect 4615 303 4645 367
rect 4701 303 4731 367
rect 4792 303 4822 367
rect 4878 303 4908 367
rect 4357 287 4908 303
rect 4357 273 4382 287
rect 2387 249 4286 263
rect 2387 235 2497 249
rect 2387 227 2417 235
rect 1214 217 1853 227
rect 552 197 1853 217
rect 641 175 671 197
rect 743 175 773 197
rect 829 175 859 197
rect 915 175 945 197
rect 1001 175 1031 197
rect 1103 175 1133 197
rect 1189 175 1219 197
rect 1307 175 1337 197
rect 1393 175 1423 197
rect 1479 175 1509 197
rect 1565 175 1595 197
rect 1651 175 1681 197
rect 1737 175 1767 197
rect 1823 175 1853 197
rect 1909 197 2417 227
rect 2469 215 2497 235
rect 2531 215 2565 249
rect 2599 215 2633 249
rect 2667 215 2701 249
rect 2735 215 2769 249
rect 2803 215 2837 249
rect 2871 215 2905 249
rect 2939 215 2973 249
rect 3007 215 3041 249
rect 3075 247 4286 249
rect 3075 215 3148 247
rect 2469 213 3148 215
rect 3182 213 3216 247
rect 3250 213 3284 247
rect 3318 213 3352 247
rect 3386 213 3420 247
rect 3454 213 3488 247
rect 3522 213 3556 247
rect 3590 213 3624 247
rect 3658 213 3692 247
rect 3726 213 3760 247
rect 3794 213 3828 247
rect 3862 213 3896 247
rect 3930 213 3964 247
rect 3998 213 4032 247
rect 4066 213 4100 247
rect 4134 213 4168 247
rect 4202 213 4236 247
rect 4270 213 4286 247
rect 4366 253 4382 273
rect 4416 253 4450 287
rect 4484 253 4518 287
rect 4552 253 4586 287
rect 4620 253 4654 287
rect 4688 253 4722 287
rect 4756 253 4790 287
rect 4824 253 4858 287
rect 4892 253 4908 287
rect 4366 237 4908 253
rect 4366 215 4396 237
rect 4467 215 4497 237
rect 4585 215 4615 237
rect 4671 215 4701 237
rect 2469 197 4286 213
rect 1909 175 1939 197
rect 2011 175 2041 197
rect 2113 175 2143 197
rect 2215 175 2245 197
rect 2301 175 2331 197
rect 2387 175 2417 197
rect 2473 175 2503 197
rect 2559 175 2589 197
rect 2645 175 2675 197
rect 2731 175 2761 197
rect 2817 175 2847 197
rect 2903 175 2933 197
rect 2989 175 3019 197
rect 3075 175 3105 197
rect 84 21 114 47
rect 170 21 200 47
rect 288 21 318 47
rect 420 21 450 47
rect 641 21 671 47
rect 743 21 773 47
rect 829 21 859 47
rect 915 21 945 47
rect 1001 21 1031 47
rect 1103 21 1133 47
rect 1189 21 1219 47
rect 1307 21 1337 47
rect 1393 21 1423 47
rect 1479 21 1509 47
rect 1565 21 1595 47
rect 1651 21 1681 47
rect 1737 21 1767 47
rect 1823 21 1853 47
rect 1909 21 1939 47
rect 2011 21 2041 47
rect 2113 21 2143 47
rect 2215 21 2245 47
rect 2301 21 2331 47
rect 2387 21 2417 47
rect 2473 21 2503 47
rect 2559 21 2589 47
rect 2645 21 2675 47
rect 2731 21 2761 47
rect 2817 21 2847 47
rect 2903 21 2933 47
rect 2989 21 3019 47
rect 3075 21 3105 47
rect 4366 21 4396 47
rect 4467 21 4497 47
rect 4585 21 4615 47
rect 4671 21 4701 47
<< polycont >>
rect 39 253 73 287
rect 1294 285 1328 319
rect 1362 285 1396 319
rect 1430 285 1464 319
rect 1498 285 1532 319
rect 1566 285 1600 319
rect 1634 285 1668 319
rect 1702 285 1736 319
rect 1770 285 1804 319
rect 1838 285 1872 319
rect 1906 285 1940 319
rect 568 217 602 251
rect 636 217 670 251
rect 704 217 738 251
rect 772 217 806 251
rect 840 217 874 251
rect 908 217 942 251
rect 976 217 1010 251
rect 1044 217 1078 251
rect 1112 217 1146 251
rect 1180 217 1214 251
rect 2497 215 2531 249
rect 2565 215 2599 249
rect 2633 215 2667 249
rect 2701 215 2735 249
rect 2769 215 2803 249
rect 2837 215 2871 249
rect 2905 215 2939 249
rect 2973 215 3007 249
rect 3041 215 3075 249
rect 3148 213 3182 247
rect 3216 213 3250 247
rect 3284 213 3318 247
rect 3352 213 3386 247
rect 3420 213 3454 247
rect 3488 213 3522 247
rect 3556 213 3590 247
rect 3624 213 3658 247
rect 3692 213 3726 247
rect 3760 213 3794 247
rect 3828 213 3862 247
rect 3896 213 3930 247
rect 3964 213 3998 247
rect 4032 213 4066 247
rect 4100 213 4134 247
rect 4168 213 4202 247
rect 4236 213 4270 247
rect 4382 253 4416 287
rect 4450 253 4484 287
rect 4518 253 4552 287
rect 4586 253 4620 287
rect 4654 253 4688 287
rect 4722 253 4756 287
rect 4790 253 4824 287
rect 4858 253 4892 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3775 683
rect 3809 649 3871 683
rect 3905 649 3967 683
rect 4001 649 4063 683
rect 4097 649 4159 683
rect 4193 649 4255 683
rect 4289 649 4351 683
rect 4385 649 4447 683
rect 4481 649 4543 683
rect 4577 649 4639 683
rect 4673 649 4735 683
rect 4769 649 4831 683
rect 4865 649 4927 683
rect 4961 649 4992 683
rect 23 607 89 649
rect 23 573 39 607
rect 73 573 89 607
rect 23 510 89 573
rect 23 476 39 510
rect 73 476 89 510
rect 23 413 89 476
rect 23 379 39 413
rect 73 379 89 413
rect 23 363 89 379
rect 125 597 159 613
rect 125 505 159 563
rect 125 413 159 471
rect 23 287 89 303
rect 23 253 39 287
rect 73 253 89 287
rect 23 236 89 253
rect 125 203 159 379
rect 195 607 245 649
rect 195 573 211 607
rect 195 510 245 573
rect 195 476 211 510
rect 195 413 245 476
rect 195 379 211 413
rect 195 363 245 379
rect 281 597 347 613
rect 281 563 297 597
rect 331 563 347 597
rect 281 505 347 563
rect 281 471 297 505
rect 331 471 347 505
rect 281 413 347 471
rect 383 607 417 649
rect 383 483 417 573
rect 383 433 417 449
rect 453 597 519 613
rect 453 563 469 597
rect 503 563 519 597
rect 453 505 519 563
rect 453 471 469 505
rect 503 471 519 505
rect 281 379 297 413
rect 331 397 347 413
rect 453 413 519 471
rect 453 397 469 413
rect 331 379 469 397
rect 503 379 519 413
rect 281 363 519 379
rect 555 607 589 649
rect 555 514 589 573
rect 725 611 763 649
rect 725 577 727 611
rect 761 577 763 611
rect 555 421 589 480
rect 555 371 589 387
rect 625 537 691 553
rect 625 503 641 537
rect 675 503 691 537
rect 625 423 691 503
rect 725 491 763 577
rect 897 611 935 649
rect 897 577 899 611
rect 933 577 935 611
rect 725 457 727 491
rect 761 457 763 491
rect 725 441 763 457
rect 797 537 863 553
rect 797 503 813 537
rect 847 503 863 537
rect 625 389 641 423
rect 675 407 691 423
rect 797 423 863 503
rect 897 491 935 577
rect 1069 611 1107 649
rect 1069 577 1071 611
rect 1105 577 1107 611
rect 897 457 899 491
rect 933 457 935 491
rect 897 441 935 457
rect 969 537 1035 553
rect 969 503 985 537
rect 1019 503 1035 537
rect 797 407 813 423
rect 675 389 813 407
rect 847 407 863 423
rect 969 423 1035 503
rect 1069 491 1107 577
rect 1241 611 1279 649
rect 1241 577 1243 611
rect 1277 577 1279 611
rect 1069 457 1071 491
rect 1105 457 1107 491
rect 1069 441 1107 457
rect 1141 537 1207 553
rect 1141 503 1157 537
rect 1191 503 1207 537
rect 969 407 985 423
rect 847 389 985 407
rect 1019 407 1035 423
rect 1141 423 1207 503
rect 1241 491 1279 577
rect 1413 611 1451 649
rect 1413 577 1415 611
rect 1449 577 1451 611
rect 1241 457 1243 491
rect 1277 457 1279 491
rect 1241 441 1279 457
rect 1313 537 1379 553
rect 1313 503 1329 537
rect 1363 503 1379 537
rect 1141 407 1157 423
rect 1019 389 1157 407
rect 1191 407 1207 423
rect 1313 423 1379 503
rect 1413 491 1451 577
rect 1585 611 1623 649
rect 1585 577 1587 611
rect 1621 577 1623 611
rect 1413 457 1415 491
rect 1449 457 1451 491
rect 1413 441 1451 457
rect 1485 537 1551 553
rect 1485 503 1501 537
rect 1535 503 1551 537
rect 1313 407 1329 423
rect 1191 389 1329 407
rect 1363 407 1379 423
rect 1485 423 1551 503
rect 1585 491 1623 577
rect 1761 611 1799 649
rect 1761 577 1763 611
rect 1797 577 1799 611
rect 1585 457 1587 491
rect 1621 457 1623 491
rect 1585 441 1623 457
rect 1661 537 1727 553
rect 1661 503 1677 537
rect 1711 503 1727 537
rect 1485 407 1501 423
rect 1363 389 1501 407
rect 1535 407 1551 423
rect 1661 423 1727 503
rect 1761 491 1799 577
rect 1933 611 1971 649
rect 1933 577 1935 611
rect 1969 577 1971 611
rect 1761 457 1763 491
rect 1797 457 1799 491
rect 1761 441 1799 457
rect 1833 537 1899 553
rect 1833 503 1849 537
rect 1883 503 1899 537
rect 1661 407 1677 423
rect 1535 389 1677 407
rect 1711 407 1727 423
rect 1833 423 1899 503
rect 1933 491 1971 577
rect 1933 457 1935 491
rect 1969 457 1971 491
rect 1933 441 1971 457
rect 2005 597 2071 613
rect 2005 563 2021 597
rect 2055 563 2071 597
rect 2005 505 2071 563
rect 2005 471 2021 505
rect 2055 471 2071 505
rect 1833 407 1849 423
rect 1711 389 1849 407
rect 1883 407 1899 423
rect 2005 413 2071 471
rect 2005 407 2021 413
rect 1883 389 2021 407
rect 625 379 2021 389
rect 2055 379 2071 413
rect 625 373 2071 379
rect 23 184 89 200
rect 23 150 39 184
rect 73 150 89 184
rect 23 93 89 150
rect 23 59 39 93
rect 73 59 89 93
rect 23 17 89 59
rect 336 229 402 363
rect 453 337 519 363
rect 453 319 1956 337
rect 453 303 1294 319
rect 1278 285 1294 303
rect 1328 285 1362 319
rect 1396 285 1430 319
rect 1464 285 1498 319
rect 1532 285 1566 319
rect 1600 285 1634 319
rect 1668 285 1702 319
rect 1736 285 1770 319
rect 1804 285 1838 319
rect 1872 285 1906 319
rect 1940 285 1956 319
rect 2005 327 2071 373
rect 2107 607 2141 649
rect 2107 510 2141 573
rect 2107 413 2141 476
rect 2107 363 2141 379
rect 2177 597 2227 613
rect 2177 563 2193 597
rect 2177 505 2227 563
rect 2177 471 2193 505
rect 2263 607 2329 649
rect 2263 573 2279 607
rect 2313 573 2329 607
rect 2263 523 2329 573
rect 2263 489 2279 523
rect 2313 489 2329 523
rect 2263 473 2329 489
rect 2464 577 4078 613
rect 2464 545 2530 577
rect 2464 511 2480 545
rect 2514 511 2530 545
rect 2636 549 2702 577
rect 2177 437 2227 471
rect 2464 442 2530 511
rect 2464 437 2480 442
rect 2177 413 2480 437
rect 2177 379 2193 413
rect 2227 408 2480 413
rect 2514 408 2530 442
rect 2227 392 2530 408
rect 2564 527 2602 543
rect 2564 493 2566 527
rect 2600 493 2602 527
rect 2564 439 2602 493
rect 2564 405 2566 439
rect 2600 405 2602 439
rect 2177 327 2227 379
rect 2564 356 2602 405
rect 2636 515 2652 549
rect 2686 515 2702 549
rect 2808 549 2874 577
rect 2636 481 2702 515
rect 2636 447 2652 481
rect 2686 447 2702 481
rect 2636 413 2702 447
rect 2636 379 2652 413
rect 2686 379 2702 413
rect 2736 527 2774 543
rect 2736 493 2738 527
rect 2772 493 2774 527
rect 2736 439 2774 493
rect 2736 405 2738 439
rect 2772 405 2774 439
rect 2005 293 2227 327
rect 2261 351 2602 356
rect 2261 317 2394 351
rect 2428 317 2566 351
rect 2600 345 2602 351
rect 2736 351 2774 405
rect 2808 515 2824 549
rect 2858 515 2874 549
rect 2980 549 3046 577
rect 2808 481 2874 515
rect 2808 447 2824 481
rect 2858 447 2874 481
rect 2808 413 2874 447
rect 2808 379 2824 413
rect 2858 379 2874 413
rect 2908 527 2946 543
rect 2908 493 2910 527
rect 2944 493 2946 527
rect 2908 439 2946 493
rect 2908 405 2910 439
rect 2944 405 2946 439
rect 2736 345 2738 351
rect 2600 317 2738 345
rect 2772 345 2774 351
rect 2908 351 2946 405
rect 2980 515 2996 549
rect 3030 515 3046 549
rect 3152 549 3218 577
rect 2980 481 3046 515
rect 2980 447 2996 481
rect 3030 447 3046 481
rect 2980 413 3046 447
rect 2980 379 2996 413
rect 3030 379 3046 413
rect 3080 527 3118 543
rect 3080 493 3082 527
rect 3116 493 3118 527
rect 3080 439 3118 493
rect 3080 405 3082 439
rect 3116 405 3118 439
rect 2908 345 2910 351
rect 2772 317 2910 345
rect 2944 345 2946 351
rect 3080 351 3118 405
rect 3152 515 3168 549
rect 3202 515 3218 549
rect 3324 549 3390 577
rect 3152 481 3218 515
rect 3152 447 3168 481
rect 3202 447 3218 481
rect 3152 413 3218 447
rect 3152 379 3168 413
rect 3202 379 3218 413
rect 3252 527 3290 543
rect 3252 493 3254 527
rect 3288 493 3290 527
rect 3252 439 3290 493
rect 3252 405 3254 439
rect 3288 405 3290 439
rect 3080 345 3082 351
rect 2944 317 3082 345
rect 3116 345 3118 351
rect 3252 351 3290 405
rect 3324 515 3340 549
rect 3374 515 3390 549
rect 3496 549 3562 577
rect 3324 481 3390 515
rect 3324 447 3340 481
rect 3374 447 3390 481
rect 3324 413 3390 447
rect 3324 379 3340 413
rect 3374 379 3390 413
rect 3424 527 3462 543
rect 3424 493 3426 527
rect 3460 493 3462 527
rect 3424 439 3462 493
rect 3424 405 3426 439
rect 3460 405 3462 439
rect 3252 345 3254 351
rect 3116 317 3254 345
rect 3288 345 3290 351
rect 3424 351 3462 405
rect 3496 515 3512 549
rect 3546 515 3562 549
rect 3668 549 3734 577
rect 3496 481 3562 515
rect 3496 447 3512 481
rect 3546 447 3562 481
rect 3496 413 3562 447
rect 3496 379 3512 413
rect 3546 379 3562 413
rect 3596 527 3634 543
rect 3596 493 3598 527
rect 3632 493 3634 527
rect 3596 439 3634 493
rect 3596 405 3598 439
rect 3632 405 3634 439
rect 3424 345 3426 351
rect 3288 317 3426 345
rect 3460 345 3462 351
rect 3596 351 3634 405
rect 3668 515 3684 549
rect 3718 515 3734 549
rect 3840 549 3906 577
rect 3668 481 3734 515
rect 3668 447 3684 481
rect 3718 447 3734 481
rect 3668 413 3734 447
rect 3668 379 3684 413
rect 3718 379 3734 413
rect 3768 527 3806 543
rect 3768 493 3770 527
rect 3804 493 3806 527
rect 3768 439 3806 493
rect 3768 405 3770 439
rect 3804 405 3806 439
rect 3596 345 3598 351
rect 3460 317 3598 345
rect 3632 345 3634 351
rect 3768 351 3806 405
rect 3840 515 3856 549
rect 3890 515 3906 549
rect 4012 549 4078 577
rect 4210 607 4260 649
rect 4210 573 4226 607
rect 3840 481 3906 515
rect 3840 447 3856 481
rect 3890 447 3906 481
rect 3840 413 3906 447
rect 3840 379 3856 413
rect 3890 379 3906 413
rect 3940 527 3978 543
rect 3940 493 3942 527
rect 3976 493 3978 527
rect 3940 439 3978 493
rect 3940 405 3942 439
rect 3976 405 3978 439
rect 3768 345 3770 351
rect 3632 317 3770 345
rect 3804 345 3806 351
rect 3940 351 3978 405
rect 4012 515 4028 549
rect 4062 515 4078 549
rect 4012 481 4078 515
rect 4012 447 4028 481
rect 4062 447 4078 481
rect 4012 413 4078 447
rect 4012 379 4028 413
rect 4062 379 4078 413
rect 4114 545 4164 561
rect 4148 511 4164 545
rect 4114 448 4164 511
rect 4148 414 4164 448
rect 3940 345 3942 351
rect 3804 317 3942 345
rect 3976 345 3978 351
rect 4114 351 4164 414
rect 4210 510 4260 573
rect 4210 476 4226 510
rect 4210 413 4260 476
rect 4210 379 4226 413
rect 4210 363 4260 379
rect 4296 597 4362 613
rect 4296 563 4312 597
rect 4346 563 4362 597
rect 4296 505 4362 563
rect 4296 471 4312 505
rect 4346 471 4362 505
rect 4296 413 4362 471
rect 4398 607 4432 649
rect 4398 483 4432 573
rect 4398 433 4432 449
rect 4468 597 4534 613
rect 4468 563 4484 597
rect 4518 563 4534 597
rect 4468 505 4534 563
rect 4468 471 4484 505
rect 4518 471 4534 505
rect 4296 379 4312 413
rect 4346 379 4362 413
rect 4296 373 4362 379
rect 4468 413 4534 471
rect 4468 379 4484 413
rect 4518 379 4534 413
rect 4570 607 4604 649
rect 4570 533 4604 573
rect 4570 459 4604 499
rect 4570 409 4604 425
rect 4640 597 4706 613
rect 4640 563 4656 597
rect 4690 563 4706 597
rect 4640 505 4706 563
rect 4640 471 4656 505
rect 4690 471 4706 505
rect 4640 413 4706 471
rect 4468 373 4534 379
rect 4640 379 4656 413
rect 4690 379 4706 413
rect 4742 607 4776 649
rect 4742 533 4776 573
rect 4742 459 4776 499
rect 4742 409 4776 425
rect 4817 597 4883 613
rect 4817 563 4833 597
rect 4867 563 4883 597
rect 4817 505 4883 563
rect 4817 471 4833 505
rect 4867 471 4883 505
rect 4817 413 4883 471
rect 4640 373 4706 379
rect 4817 379 4833 413
rect 4867 379 4883 413
rect 4817 373 4883 379
rect 3976 317 4114 345
rect 4148 317 4164 351
rect 2261 301 4164 317
rect 1278 269 1956 285
rect 336 195 352 229
rect 386 195 402 229
rect 438 251 1230 267
rect 438 217 568 251
rect 602 217 636 251
rect 670 217 704 251
rect 738 217 772 251
rect 806 217 840 251
rect 874 217 908 251
rect 942 217 976 251
rect 1010 217 1044 251
rect 1078 217 1112 251
rect 1146 217 1180 251
rect 1214 217 1230 251
rect 438 201 1230 217
rect 125 159 159 169
rect 438 159 472 201
rect 1332 199 1914 233
rect 1332 165 1398 199
rect 125 125 472 159
rect 580 133 1398 165
rect 580 131 1348 133
rect 580 126 646 131
rect 125 103 159 125
rect 580 92 596 126
rect 630 92 646 126
rect 784 126 818 131
rect 125 53 159 69
rect 211 55 227 89
rect 261 55 277 89
rect 211 17 277 55
rect 468 73 534 89
rect 468 39 484 73
rect 518 39 534 73
rect 580 53 646 92
rect 682 94 748 95
rect 682 60 698 94
rect 732 60 748 94
rect 468 17 534 39
rect 682 17 748 60
rect 956 126 990 131
rect 784 53 818 92
rect 854 94 920 95
rect 854 60 870 94
rect 904 60 920 94
rect 854 17 920 60
rect 1128 126 1194 131
rect 956 53 990 92
rect 1026 94 1092 95
rect 1026 60 1042 94
rect 1076 60 1092 94
rect 1026 17 1092 60
rect 1128 92 1144 126
rect 1178 92 1194 126
rect 1332 99 1348 131
rect 1382 99 1398 133
rect 1128 53 1194 92
rect 1230 94 1296 95
rect 1230 60 1246 94
rect 1280 60 1296 94
rect 1230 17 1296 60
rect 1332 53 1398 99
rect 1434 120 1468 163
rect 1434 17 1468 86
rect 1504 133 1570 199
rect 1504 99 1520 133
rect 1554 99 1570 133
rect 1504 53 1570 99
rect 1606 120 1640 163
rect 1606 17 1640 86
rect 1676 133 1742 199
rect 1676 99 1692 133
rect 1726 99 1742 133
rect 1676 53 1742 99
rect 1778 120 1812 163
rect 1778 17 1812 86
rect 1848 133 1914 199
rect 2261 179 2447 301
rect 3254 299 4164 301
rect 4296 339 4883 373
rect 4919 607 4969 649
rect 4953 573 4969 607
rect 4919 510 4969 573
rect 4953 476 4969 510
rect 4919 413 4969 476
rect 4953 379 4969 413
rect 4919 363 4969 379
rect 2481 263 3091 265
rect 4296 263 4330 339
rect 2481 249 4330 263
rect 2481 215 2497 249
rect 2531 215 2565 249
rect 2599 215 2633 249
rect 2667 215 2701 249
rect 2735 215 2769 249
rect 2803 215 2837 249
rect 2871 215 2905 249
rect 2939 215 2973 249
rect 3007 215 3041 249
rect 3075 247 4330 249
rect 3075 215 3148 247
rect 3132 213 3148 215
rect 3182 213 3216 247
rect 3250 213 3284 247
rect 3318 213 3352 247
rect 3386 213 3420 247
rect 3454 213 3488 247
rect 3522 213 3556 247
rect 3590 213 3624 247
rect 3658 213 3692 247
rect 3726 213 3760 247
rect 3794 213 3828 247
rect 3862 213 3896 247
rect 3930 213 3964 247
rect 3998 213 4032 247
rect 4066 213 4100 247
rect 4134 213 4168 247
rect 4202 213 4236 247
rect 4270 213 4330 247
rect 4366 287 4967 303
rect 4366 253 4382 287
rect 4416 253 4450 287
rect 4484 253 4518 287
rect 4552 253 4586 287
rect 4620 253 4654 287
rect 4688 253 4722 287
rect 4756 253 4790 287
rect 4824 253 4858 287
rect 4892 253 4967 287
rect 4366 236 4967 253
rect 3132 200 4330 213
rect 3132 197 4676 200
rect 4296 184 4676 197
rect 1848 99 1864 133
rect 1898 99 1914 133
rect 1950 167 3080 179
rect 1950 133 1966 167
rect 2000 133 2170 167
rect 2204 163 3080 167
rect 4296 166 4422 184
rect 2204 133 2342 163
rect 1950 129 2342 133
rect 2376 129 2514 163
rect 2548 129 2686 163
rect 2720 129 2858 163
rect 2892 129 3030 163
rect 3064 129 3080 163
rect 1848 95 1914 99
rect 3116 124 3182 161
rect 4406 150 4422 166
rect 4456 166 4626 184
rect 4456 150 4472 166
rect 3116 95 3132 124
rect 1848 93 3132 95
rect 1848 59 2068 93
rect 2102 59 2256 93
rect 2290 59 2428 93
rect 2462 59 2600 93
rect 2634 59 2772 93
rect 2806 59 2944 93
rect 2978 90 3132 93
rect 3166 90 3182 124
rect 2978 59 3182 90
rect 1848 53 3182 59
rect 4304 103 4370 130
rect 4304 69 4320 103
rect 4354 69 4370 103
rect 4304 17 4370 69
rect 4406 93 4472 150
rect 4610 150 4626 166
rect 4660 150 4676 184
rect 4406 59 4422 93
rect 4456 59 4472 93
rect 4508 103 4574 130
rect 4508 69 4524 103
rect 4558 69 4574 103
rect 4508 17 4574 69
rect 4610 103 4676 150
rect 4610 69 4626 103
rect 4660 69 4676 103
rect 4610 53 4676 69
rect 4712 184 4778 200
rect 4712 150 4728 184
rect 4762 150 4778 184
rect 4712 93 4778 150
rect 4712 59 4728 93
rect 4762 59 4778 93
rect 4712 17 4778 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 4992 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 3583 649 3617 683
rect 3679 649 3713 683
rect 3775 649 3809 683
rect 3871 649 3905 683
rect 3967 649 4001 683
rect 4063 649 4097 683
rect 4159 649 4193 683
rect 4255 649 4289 683
rect 4351 649 4385 683
rect 4447 649 4481 683
rect 4543 649 4577 683
rect 4639 649 4673 683
rect 4735 649 4769 683
rect 4831 649 4865 683
rect 4927 649 4961 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
rect 4063 -17 4097 17
rect 4159 -17 4193 17
rect 4255 -17 4289 17
rect 4351 -17 4385 17
rect 4447 -17 4481 17
rect 4543 -17 4577 17
rect 4639 -17 4673 17
rect 4735 -17 4769 17
rect 4831 -17 4865 17
rect 4927 -17 4961 17
<< metal1 >>
rect 0 683 4992 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3775 683
rect 3809 649 3871 683
rect 3905 649 3967 683
rect 4001 649 4063 683
rect 4097 649 4159 683
rect 4193 649 4255 683
rect 4289 649 4351 683
rect 4385 649 4447 683
rect 4481 649 4543 683
rect 4577 649 4639 683
rect 4673 649 4735 683
rect 4769 649 4831 683
rect 4865 649 4927 683
rect 4961 649 4992 683
rect 0 617 4992 649
rect 0 17 4992 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 4992 17
rect 0 -49 4992 -17
<< labels >>
flabel pwell s 0 0 4992 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 4992 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 busdriver_20
flabel metal1 s 0 617 4992 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 4992 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 2335 316 2369 350 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 4447 242 4481 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 4543 242 4577 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 4639 242 4673 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 4735 242 4769 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 4831 242 4865 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 4927 242 4961 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 2335 242 2369 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 2335 168 2369 202 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 4992 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y
string GDS_END 5729378
string GDS_START 5697026
<< end >>
