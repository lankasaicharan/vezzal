magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 5 49 1505 241
rect 0 0 1536 49
<< scnmos >>
rect 84 47 114 215
rect 170 47 200 215
rect 256 47 286 215
rect 342 47 372 215
rect 428 47 458 215
rect 514 47 544 215
rect 600 47 630 215
rect 686 47 716 215
rect 794 47 824 215
rect 880 47 910 215
rect 966 47 996 215
rect 1052 47 1082 215
rect 1138 47 1168 215
rect 1224 47 1254 215
rect 1310 47 1340 215
rect 1396 47 1426 215
<< scpmoshvt >>
rect 98 367 128 619
rect 184 367 214 619
rect 270 367 300 619
rect 356 367 386 619
rect 442 367 472 619
rect 528 367 558 619
rect 614 367 644 619
rect 710 367 740 619
rect 796 367 826 619
rect 882 367 912 619
rect 968 367 998 619
rect 1054 367 1084 619
rect 1140 367 1170 619
rect 1226 367 1256 619
rect 1312 367 1342 619
rect 1398 367 1428 619
<< ndiff >>
rect 31 203 84 215
rect 31 169 39 203
rect 73 169 84 203
rect 31 93 84 169
rect 31 59 39 93
rect 73 59 84 93
rect 31 47 84 59
rect 114 203 170 215
rect 114 169 125 203
rect 159 169 170 203
rect 114 101 170 169
rect 114 67 125 101
rect 159 67 170 101
rect 114 47 170 67
rect 200 164 256 215
rect 200 130 211 164
rect 245 130 256 164
rect 200 93 256 130
rect 200 59 211 93
rect 245 59 256 93
rect 200 47 256 59
rect 286 207 342 215
rect 286 173 297 207
rect 331 173 342 207
rect 286 101 342 173
rect 286 67 297 101
rect 331 67 342 101
rect 286 47 342 67
rect 372 194 428 215
rect 372 160 383 194
rect 417 160 428 194
rect 372 47 428 160
rect 458 101 514 215
rect 458 67 469 101
rect 503 67 514 101
rect 458 47 514 67
rect 544 194 600 215
rect 544 160 555 194
rect 589 160 600 194
rect 544 47 600 160
rect 630 101 686 215
rect 630 67 641 101
rect 675 67 686 101
rect 630 47 686 67
rect 716 107 794 215
rect 716 73 727 107
rect 761 73 794 107
rect 716 47 794 73
rect 824 186 880 215
rect 824 152 835 186
rect 869 152 880 186
rect 824 101 880 152
rect 824 67 835 101
rect 869 67 880 101
rect 824 47 880 67
rect 910 95 966 215
rect 910 61 921 95
rect 955 61 966 95
rect 910 47 966 61
rect 996 175 1052 215
rect 996 141 1007 175
rect 1041 141 1052 175
rect 996 91 1052 141
rect 996 57 1007 91
rect 1041 57 1052 91
rect 996 47 1052 57
rect 1082 99 1138 215
rect 1082 65 1093 99
rect 1127 65 1138 99
rect 1082 47 1138 65
rect 1168 175 1224 215
rect 1168 141 1179 175
rect 1213 141 1224 175
rect 1168 91 1224 141
rect 1168 57 1179 91
rect 1213 57 1224 91
rect 1168 47 1224 57
rect 1254 95 1310 215
rect 1254 61 1265 95
rect 1299 61 1310 95
rect 1254 47 1310 61
rect 1340 175 1396 215
rect 1340 141 1351 175
rect 1385 141 1396 175
rect 1340 91 1396 141
rect 1340 57 1351 91
rect 1385 57 1396 91
rect 1340 47 1396 57
rect 1426 99 1479 215
rect 1426 65 1437 99
rect 1471 65 1479 99
rect 1426 47 1479 65
<< pdiff >>
rect 45 599 98 619
rect 45 565 53 599
rect 87 565 98 599
rect 45 525 98 565
rect 45 491 53 525
rect 87 491 98 525
rect 45 441 98 491
rect 45 407 53 441
rect 87 407 98 441
rect 45 367 98 407
rect 128 607 184 619
rect 128 573 139 607
rect 173 573 184 607
rect 128 497 184 573
rect 128 463 139 497
rect 173 463 184 497
rect 128 367 184 463
rect 214 599 270 619
rect 214 565 225 599
rect 259 565 270 599
rect 214 525 270 565
rect 214 491 225 525
rect 259 491 270 525
rect 214 441 270 491
rect 214 407 225 441
rect 259 407 270 441
rect 214 367 270 407
rect 300 607 356 619
rect 300 573 311 607
rect 345 573 356 607
rect 300 497 356 573
rect 300 463 311 497
rect 345 463 356 497
rect 300 367 356 463
rect 386 599 442 619
rect 386 565 397 599
rect 431 565 442 599
rect 386 525 442 565
rect 386 491 397 525
rect 431 491 442 525
rect 386 441 442 491
rect 386 407 397 441
rect 431 407 442 441
rect 386 367 442 407
rect 472 611 528 619
rect 472 577 483 611
rect 517 577 528 611
rect 472 499 528 577
rect 472 465 483 499
rect 517 465 528 499
rect 472 367 528 465
rect 558 597 614 619
rect 558 563 569 597
rect 603 563 614 597
rect 558 525 614 563
rect 558 491 569 525
rect 603 491 614 525
rect 558 441 614 491
rect 558 407 569 441
rect 603 407 614 441
rect 558 367 614 407
rect 644 611 710 619
rect 644 577 655 611
rect 689 577 710 611
rect 644 499 710 577
rect 644 465 655 499
rect 689 465 710 499
rect 644 367 710 465
rect 740 599 796 619
rect 740 565 751 599
rect 785 565 796 599
rect 740 507 796 565
rect 740 473 751 507
rect 785 473 796 507
rect 740 413 796 473
rect 740 379 751 413
rect 785 379 796 413
rect 740 367 796 379
rect 826 599 882 619
rect 826 565 837 599
rect 871 565 882 599
rect 826 529 882 565
rect 826 495 837 529
rect 871 495 882 529
rect 826 459 882 495
rect 826 425 837 459
rect 871 425 882 459
rect 826 367 882 425
rect 912 481 968 619
rect 912 447 923 481
rect 957 447 968 481
rect 912 413 968 447
rect 912 379 923 413
rect 957 379 968 413
rect 912 367 968 379
rect 998 599 1054 619
rect 998 565 1009 599
rect 1043 565 1054 599
rect 998 367 1054 565
rect 1084 425 1140 619
rect 1084 391 1095 425
rect 1129 391 1140 425
rect 1084 367 1140 391
rect 1170 599 1226 619
rect 1170 565 1181 599
rect 1215 565 1226 599
rect 1170 367 1226 565
rect 1256 413 1312 619
rect 1256 379 1267 413
rect 1301 379 1312 413
rect 1256 367 1312 379
rect 1342 599 1398 619
rect 1342 565 1353 599
rect 1387 565 1398 599
rect 1342 367 1398 565
rect 1428 607 1485 619
rect 1428 573 1443 607
rect 1477 573 1485 607
rect 1428 537 1485 573
rect 1428 503 1443 537
rect 1477 503 1485 537
rect 1428 467 1485 503
rect 1428 433 1443 467
rect 1477 433 1485 467
rect 1428 367 1485 433
<< ndiffc >>
rect 39 169 73 203
rect 39 59 73 93
rect 125 169 159 203
rect 125 67 159 101
rect 211 130 245 164
rect 211 59 245 93
rect 297 173 331 207
rect 297 67 331 101
rect 383 160 417 194
rect 469 67 503 101
rect 555 160 589 194
rect 641 67 675 101
rect 727 73 761 107
rect 835 152 869 186
rect 835 67 869 101
rect 921 61 955 95
rect 1007 141 1041 175
rect 1007 57 1041 91
rect 1093 65 1127 99
rect 1179 141 1213 175
rect 1179 57 1213 91
rect 1265 61 1299 95
rect 1351 141 1385 175
rect 1351 57 1385 91
rect 1437 65 1471 99
<< pdiffc >>
rect 53 565 87 599
rect 53 491 87 525
rect 53 407 87 441
rect 139 573 173 607
rect 139 463 173 497
rect 225 565 259 599
rect 225 491 259 525
rect 225 407 259 441
rect 311 573 345 607
rect 311 463 345 497
rect 397 565 431 599
rect 397 491 431 525
rect 397 407 431 441
rect 483 577 517 611
rect 483 465 517 499
rect 569 563 603 597
rect 569 491 603 525
rect 569 407 603 441
rect 655 577 689 611
rect 655 465 689 499
rect 751 565 785 599
rect 751 473 785 507
rect 751 379 785 413
rect 837 565 871 599
rect 837 495 871 529
rect 837 425 871 459
rect 923 447 957 481
rect 923 379 957 413
rect 1009 565 1043 599
rect 1095 391 1129 425
rect 1181 565 1215 599
rect 1267 379 1301 413
rect 1353 565 1387 599
rect 1443 573 1477 607
rect 1443 503 1477 537
rect 1443 433 1477 467
<< poly >>
rect 98 619 128 645
rect 184 619 214 645
rect 270 619 300 645
rect 356 619 386 645
rect 442 619 472 645
rect 528 619 558 645
rect 614 619 644 645
rect 710 619 740 645
rect 796 619 826 645
rect 882 619 912 645
rect 968 619 998 645
rect 1054 619 1084 645
rect 1140 619 1170 645
rect 1226 619 1256 645
rect 1312 619 1342 645
rect 1398 619 1428 645
rect 98 345 128 367
rect 184 345 214 367
rect 270 345 300 367
rect 24 315 300 345
rect 24 309 294 315
rect 24 275 40 309
rect 74 275 108 309
rect 142 275 176 309
rect 210 275 244 309
rect 278 275 294 309
rect 24 259 294 275
rect 356 303 386 367
rect 442 303 472 367
rect 528 303 558 367
rect 614 303 644 367
rect 710 321 740 367
rect 356 287 644 303
rect 356 267 383 287
rect 84 215 114 259
rect 170 215 200 259
rect 256 215 286 259
rect 342 253 383 267
rect 417 253 451 287
rect 485 253 519 287
rect 553 253 587 287
rect 621 273 644 287
rect 686 305 752 321
rect 621 253 637 273
rect 342 237 637 253
rect 686 271 702 305
rect 736 271 752 305
rect 686 255 752 271
rect 796 303 826 367
rect 882 303 912 367
rect 968 303 998 367
rect 1054 335 1084 367
rect 1140 335 1170 367
rect 1226 335 1256 367
rect 1312 335 1342 367
rect 796 287 998 303
rect 796 267 812 287
rect 342 215 372 237
rect 428 215 458 237
rect 514 215 544 237
rect 600 215 630 237
rect 686 215 716 255
rect 794 253 812 267
rect 846 253 880 287
rect 914 253 948 287
rect 982 253 998 287
rect 794 237 998 253
rect 1052 319 1342 335
rect 1052 285 1086 319
rect 1120 285 1154 319
rect 1188 285 1222 319
rect 1256 285 1290 319
rect 1324 285 1342 319
rect 1398 303 1428 367
rect 1052 269 1342 285
rect 1396 287 1462 303
rect 794 215 824 237
rect 880 215 910 237
rect 966 215 996 237
rect 1052 215 1082 269
rect 1138 215 1168 269
rect 1224 215 1254 269
rect 1310 215 1340 269
rect 1396 253 1412 287
rect 1446 253 1462 287
rect 1396 237 1462 253
rect 1396 215 1426 237
rect 84 21 114 47
rect 170 21 200 47
rect 256 21 286 47
rect 342 21 372 47
rect 428 21 458 47
rect 514 21 544 47
rect 600 21 630 47
rect 686 21 716 47
rect 794 21 824 47
rect 880 21 910 47
rect 966 21 996 47
rect 1052 21 1082 47
rect 1138 21 1168 47
rect 1224 21 1254 47
rect 1310 21 1340 47
rect 1396 21 1426 47
<< polycont >>
rect 40 275 74 309
rect 108 275 142 309
rect 176 275 210 309
rect 244 275 278 309
rect 383 253 417 287
rect 451 253 485 287
rect 519 253 553 287
rect 587 253 621 287
rect 702 271 736 305
rect 812 253 846 287
rect 880 253 914 287
rect 948 253 982 287
rect 1086 285 1120 319
rect 1154 285 1188 319
rect 1222 285 1256 319
rect 1290 285 1324 319
rect 1412 253 1446 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 37 599 89 615
rect 37 565 53 599
rect 87 565 89 599
rect 37 525 89 565
rect 37 491 53 525
rect 87 491 89 525
rect 37 441 89 491
rect 123 607 189 649
rect 123 573 139 607
rect 173 573 189 607
rect 123 497 189 573
rect 123 463 139 497
rect 173 463 189 497
rect 123 459 189 463
rect 223 599 261 615
rect 223 565 225 599
rect 259 565 261 599
rect 223 525 261 565
rect 223 491 225 525
rect 259 491 261 525
rect 37 407 53 441
rect 87 425 89 441
rect 223 441 261 491
rect 295 607 361 649
rect 295 573 311 607
rect 345 573 361 607
rect 295 497 361 573
rect 295 463 311 497
rect 345 463 361 497
rect 295 459 361 463
rect 395 599 433 615
rect 395 565 397 599
rect 431 565 433 599
rect 395 525 433 565
rect 395 491 397 525
rect 431 491 433 525
rect 223 425 225 441
rect 87 407 225 425
rect 259 425 261 441
rect 395 441 433 491
rect 467 611 533 649
rect 467 577 483 611
rect 517 577 533 611
rect 467 499 533 577
rect 467 465 483 499
rect 517 465 533 499
rect 467 459 533 465
rect 567 597 605 615
rect 567 563 569 597
rect 603 563 605 597
rect 567 525 605 563
rect 567 491 569 525
rect 603 491 605 525
rect 395 425 397 441
rect 259 407 397 425
rect 431 425 433 441
rect 567 441 605 491
rect 639 611 705 649
rect 639 577 655 611
rect 689 577 705 611
rect 639 499 705 577
rect 639 465 655 499
rect 689 465 705 499
rect 639 459 705 465
rect 739 599 789 615
rect 739 565 751 599
rect 785 565 789 599
rect 739 507 789 565
rect 739 473 751 507
rect 785 473 789 507
rect 567 425 569 441
rect 431 407 569 425
rect 603 425 605 441
rect 739 425 789 473
rect 603 413 789 425
rect 603 407 751 413
rect 37 391 751 407
rect 747 379 751 391
rect 785 379 789 413
rect 833 599 1393 615
rect 833 565 837 599
rect 871 565 1009 599
rect 1043 565 1181 599
rect 1215 565 1353 599
rect 1387 565 1393 599
rect 833 549 1393 565
rect 1427 607 1493 611
rect 1427 573 1443 607
rect 1477 573 1493 607
rect 833 529 875 549
rect 833 495 837 529
rect 871 495 875 529
rect 1427 537 1493 573
rect 1427 515 1443 537
rect 833 459 875 495
rect 833 425 837 459
rect 871 425 875 459
rect 833 409 875 425
rect 919 503 1443 515
rect 1477 503 1493 537
rect 919 481 1493 503
rect 919 447 923 481
rect 957 467 1493 481
rect 957 465 1443 467
rect 957 447 961 465
rect 919 413 961 447
rect 1427 433 1443 465
rect 1477 433 1493 467
rect 747 375 789 379
rect 919 379 923 413
rect 957 379 961 413
rect 1079 425 1323 429
rect 1079 391 1095 425
rect 1129 413 1323 425
rect 1129 391 1267 413
rect 1079 387 1267 391
rect 919 375 961 379
rect 24 323 711 357
rect 747 341 961 375
rect 1263 379 1267 387
rect 1301 397 1323 413
rect 1301 379 1516 397
rect 1263 363 1516 379
rect 24 309 329 323
rect 24 275 40 309
rect 74 275 108 309
rect 142 275 176 309
rect 210 275 244 309
rect 278 275 329 309
rect 677 307 711 323
rect 1070 329 1229 353
rect 1070 319 1342 329
rect 677 305 752 307
rect 24 269 329 275
rect 367 287 641 289
rect 367 253 383 287
rect 417 253 451 287
rect 485 253 519 287
rect 553 253 587 287
rect 621 253 641 287
rect 677 271 702 305
rect 736 271 752 305
rect 677 254 752 271
rect 796 287 1036 303
rect 367 236 641 253
rect 796 253 812 287
rect 846 253 880 287
rect 914 253 948 287
rect 982 253 1036 287
rect 1070 285 1086 319
rect 1120 285 1154 319
rect 1188 285 1222 319
rect 1256 285 1290 319
rect 1324 285 1342 319
rect 1396 287 1448 303
rect 796 251 1036 253
rect 1396 253 1412 287
rect 1446 253 1448 287
rect 1396 251 1448 253
rect 796 242 1448 251
rect 23 203 83 219
rect 23 169 39 203
rect 73 169 83 203
rect 23 93 83 169
rect 23 59 39 93
rect 73 59 83 93
rect 23 17 83 59
rect 117 207 333 235
rect 979 217 1448 242
rect 117 203 297 207
rect 117 169 125 203
rect 159 201 297 203
rect 159 169 161 201
rect 117 101 161 169
rect 295 173 297 201
rect 331 173 333 207
rect 117 67 125 101
rect 159 67 161 101
rect 117 51 161 67
rect 195 164 261 167
rect 195 130 211 164
rect 245 130 261 164
rect 195 93 261 130
rect 195 59 211 93
rect 245 59 261 93
rect 195 17 261 59
rect 295 117 333 173
rect 367 194 945 202
rect 367 160 383 194
rect 417 160 555 194
rect 589 186 945 194
rect 589 160 835 186
rect 367 152 835 160
rect 869 183 945 186
rect 1482 183 1516 363
rect 869 175 1516 183
rect 869 152 1007 175
rect 367 151 1007 152
rect 811 145 1007 151
rect 295 101 677 117
rect 295 67 297 101
rect 331 67 469 101
rect 503 67 641 101
rect 675 67 677 101
rect 295 51 677 67
rect 711 107 777 117
rect 711 73 727 107
rect 761 73 777 107
rect 711 17 777 73
rect 811 101 871 145
rect 991 141 1007 145
rect 1041 149 1179 175
rect 1041 141 1057 149
rect 811 67 835 101
rect 869 67 871 101
rect 811 51 871 67
rect 905 95 957 111
rect 905 61 921 95
rect 955 61 957 95
rect 905 17 957 61
rect 991 91 1057 141
rect 1163 141 1179 149
rect 1213 149 1351 175
rect 1213 141 1229 149
rect 991 57 1007 91
rect 1041 57 1057 91
rect 991 51 1057 57
rect 1091 99 1129 115
rect 1091 65 1093 99
rect 1127 65 1129 99
rect 1091 17 1129 65
rect 1163 91 1229 141
rect 1335 141 1351 149
rect 1385 149 1516 175
rect 1385 141 1401 149
rect 1163 57 1179 91
rect 1213 57 1229 91
rect 1163 51 1229 57
rect 1263 95 1301 115
rect 1263 61 1265 95
rect 1299 61 1301 95
rect 1263 17 1301 61
rect 1335 91 1401 141
rect 1335 57 1351 91
rect 1385 57 1401 91
rect 1335 51 1401 57
rect 1435 99 1487 115
rect 1435 65 1437 99
rect 1471 65 1487 99
rect 1435 17 1487 65
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a211oi_4
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 199518
string GDS_START 186522
<< end >>
