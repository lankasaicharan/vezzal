magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1299 -1308 2586 1852
<< nwell >>
rect -39 261 1326 582
<< pwell >>
rect 1 21 1287 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 267 47 297 177
rect 371 47 401 177
rect 559 47 589 177
rect 643 47 673 177
rect 727 47 757 177
rect 821 47 851 177
rect 1065 47 1095 177
rect 1179 47 1209 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 635 297 671 497
rect 729 297 765 497
rect 891 297 927 497
rect 987 297 1023 497
rect 1171 297 1207 497
<< ndiff >>
rect 27 161 89 177
rect 27 127 35 161
rect 69 127 89 161
rect 27 93 89 127
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 93 183 177
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 161 267 177
rect 213 127 223 161
rect 257 127 267 161
rect 213 93 267 127
rect 213 59 223 93
rect 257 59 267 93
rect 213 47 267 59
rect 297 165 371 177
rect 297 131 317 165
rect 351 131 371 165
rect 297 47 371 131
rect 401 93 453 177
rect 401 59 411 93
rect 445 59 453 93
rect 401 47 453 59
rect 507 93 559 177
rect 507 59 515 93
rect 549 59 559 93
rect 507 47 559 59
rect 589 165 643 177
rect 589 131 599 165
rect 633 131 643 165
rect 589 47 643 131
rect 673 93 727 177
rect 673 59 683 93
rect 717 59 727 93
rect 673 47 727 59
rect 757 161 821 177
rect 757 127 767 161
rect 801 127 821 161
rect 757 47 821 127
rect 851 93 903 177
rect 851 59 861 93
rect 895 59 903 93
rect 851 47 903 59
rect 982 93 1065 177
rect 982 59 990 93
rect 1024 59 1065 93
rect 982 47 1065 59
rect 1095 161 1179 177
rect 1095 127 1110 161
rect 1144 127 1179 161
rect 1095 89 1179 127
rect 1095 55 1110 89
rect 1144 55 1179 89
rect 1095 47 1179 55
rect 1209 161 1261 177
rect 1209 127 1219 161
rect 1253 127 1261 161
rect 1209 93 1261 127
rect 1209 59 1219 93
rect 1253 59 1261 93
rect 1209 47 1261 59
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 297 81 375
rect 117 425 175 497
rect 117 391 129 425
rect 163 391 175 425
rect 117 357 175 391
rect 117 323 129 357
rect 163 323 175 357
rect 117 297 175 323
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 409 269 443
rect 211 375 223 409
rect 257 375 269 409
rect 211 297 269 375
rect 305 409 363 497
rect 305 375 317 409
rect 351 375 363 409
rect 305 297 363 375
rect 399 477 457 497
rect 399 443 411 477
rect 445 443 457 477
rect 399 409 457 443
rect 399 375 411 409
rect 445 375 457 409
rect 399 297 457 375
rect 493 485 635 497
rect 493 451 512 485
rect 546 451 580 485
rect 614 451 635 485
rect 493 297 635 451
rect 671 477 729 497
rect 671 443 683 477
rect 717 443 729 477
rect 671 409 729 443
rect 671 375 683 409
rect 717 375 729 409
rect 671 297 729 375
rect 765 485 891 497
rect 765 451 777 485
rect 811 451 845 485
rect 879 451 891 485
rect 765 297 891 451
rect 927 477 987 497
rect 927 443 939 477
rect 973 443 987 477
rect 927 409 987 443
rect 927 375 939 409
rect 973 375 987 409
rect 927 297 987 375
rect 1023 485 1171 497
rect 1023 451 1041 485
rect 1075 451 1119 485
rect 1153 451 1171 485
rect 1023 297 1171 451
rect 1207 477 1261 497
rect 1207 443 1219 477
rect 1253 443 1261 477
rect 1207 409 1261 443
rect 1207 375 1219 409
rect 1253 375 1261 409
rect 1207 297 1261 375
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 59 163 93
rect 223 127 257 161
rect 223 59 257 93
rect 317 131 351 165
rect 411 59 445 93
rect 515 59 549 93
rect 599 131 633 165
rect 683 59 717 93
rect 767 127 801 161
rect 861 59 895 93
rect 990 59 1024 93
rect 1110 127 1144 161
rect 1110 55 1144 89
rect 1219 127 1253 161
rect 1219 59 1253 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 391 163 425
rect 129 323 163 357
rect 223 443 257 477
rect 223 375 257 409
rect 317 375 351 409
rect 411 443 445 477
rect 411 375 445 409
rect 512 451 546 485
rect 580 451 614 485
rect 683 443 717 477
rect 683 375 717 409
rect 777 451 811 485
rect 845 451 879 485
rect 939 443 973 477
rect 939 375 973 409
rect 1041 451 1075 485
rect 1119 451 1153 485
rect 1219 443 1253 477
rect 1219 375 1253 409
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 635 497 671 523
rect 729 497 765 523
rect 891 497 927 523
rect 987 497 1023 523
rect 1171 497 1207 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 635 282 671 297
rect 729 282 765 297
rect 891 282 927 297
rect 987 282 1023 297
rect 1171 282 1207 297
rect 79 265 119 282
rect 173 265 213 282
rect 31 249 213 265
rect 31 215 47 249
rect 81 215 125 249
rect 159 215 213 249
rect 31 199 213 215
rect 89 177 119 199
rect 183 177 213 199
rect 267 259 307 282
rect 361 259 401 282
rect 267 249 401 259
rect 267 215 296 249
rect 330 215 401 249
rect 267 195 401 215
rect 455 259 495 282
rect 633 259 673 282
rect 455 249 673 259
rect 455 215 491 249
rect 525 215 583 249
rect 617 215 673 249
rect 455 205 673 215
rect 267 177 297 195
rect 371 177 401 195
rect 559 177 589 205
rect 643 177 673 205
rect 727 259 767 282
rect 889 259 929 282
rect 727 249 929 259
rect 727 215 760 249
rect 794 215 838 249
rect 872 215 929 249
rect 727 205 929 215
rect 985 259 1025 282
rect 1169 261 1209 282
rect 1169 259 1264 261
rect 985 249 1264 259
rect 985 215 1058 249
rect 1092 215 1136 249
rect 1170 215 1214 249
rect 1248 215 1264 249
rect 985 205 1264 215
rect 727 177 757 205
rect 821 177 851 205
rect 1065 177 1095 205
rect 1179 203 1264 205
rect 1179 177 1209 203
rect 89 21 119 47
rect 183 21 213 47
rect 267 21 297 47
rect 371 21 401 47
rect 559 21 589 47
rect 643 21 673 47
rect 727 21 757 47
rect 821 21 851 47
rect 1065 21 1095 47
rect 1179 21 1209 47
<< polycont >>
rect 47 215 81 249
rect 125 215 159 249
rect 296 215 330 249
rect 491 215 525 249
rect 583 215 617 249
rect 760 215 794 249
rect 838 215 872 249
rect 1058 215 1092 249
rect 1136 215 1170 249
rect 1214 215 1248 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 35 477 445 493
rect 69 459 223 477
rect 35 409 69 443
rect 257 459 411 477
rect 35 359 69 375
rect 113 391 129 425
rect 163 391 179 425
rect 113 357 179 391
rect 223 409 257 443
rect 489 485 633 527
rect 489 451 512 485
rect 546 451 580 485
rect 614 451 633 485
rect 683 477 717 493
rect 223 359 257 375
rect 317 409 351 425
rect 29 257 65 325
rect 113 323 129 357
rect 163 325 179 357
rect 317 325 351 375
rect 411 409 445 443
rect 754 485 905 527
rect 754 451 777 485
rect 811 451 845 485
rect 879 451 905 485
rect 939 477 973 493
rect 683 409 717 443
rect 445 375 683 393
rect 1025 485 1169 527
rect 1025 451 1041 485
rect 1075 451 1119 485
rect 1153 451 1169 485
rect 1219 477 1253 493
rect 939 409 973 443
rect 717 375 939 393
rect 1219 409 1253 443
rect 973 375 1219 393
rect 411 359 1253 375
rect 163 323 439 325
rect 113 291 439 323
rect 29 249 175 257
rect 29 215 47 249
rect 81 215 125 249
rect 159 215 175 249
rect 213 249 359 257
rect 213 215 296 249
rect 330 215 359 249
rect 19 161 257 177
rect 393 165 439 291
rect 475 249 651 325
rect 475 215 491 249
rect 525 215 583 249
rect 617 215 651 249
rect 744 249 915 325
rect 744 215 760 249
rect 794 215 838 249
rect 872 215 915 249
rect 1005 249 1264 325
rect 1005 215 1058 249
rect 1092 215 1136 249
rect 1170 215 1214 249
rect 1248 215 1264 249
rect 19 127 35 161
rect 69 143 223 161
rect 69 127 85 143
rect 19 93 85 127
rect 207 127 223 143
rect 291 131 317 165
rect 351 131 599 165
rect 633 131 649 165
rect 1219 161 1253 177
rect 751 127 767 161
rect 801 127 1110 161
rect 1144 127 1160 161
rect 19 59 35 93
rect 69 59 85 93
rect 129 93 163 109
rect 207 93 257 127
rect 207 59 223 93
rect 257 59 411 93
rect 445 59 461 93
rect 499 59 515 93
rect 549 59 683 93
rect 717 59 861 93
rect 895 59 921 93
rect 973 59 990 93
rect 1024 59 1050 93
rect 129 17 163 59
rect 973 17 1050 59
rect 1084 89 1160 127
rect 1084 55 1110 89
rect 1144 55 1160 89
rect 1219 93 1253 127
rect 1219 17 1253 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 855 289 889 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 855 221 889 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 125 221 159 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 1044 221 1078 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1044 289 1078 323 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1134 289 1168 323 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 765 221 799 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 765 289 799 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 580 289 614 323 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 489 289 523 323 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 401 289 435 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 580 221 614 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 220 221 254 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 401 153 435 187 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 401 221 435 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 1221 289 1255 323 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1222 221 1256 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a32oi_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 315800
string GDS_START 304374
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
