magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
<< pwell >>
rect 383 243 951 259
rect 383 224 1744 243
rect 1 187 1744 224
rect 1923 187 2111 271
rect 1 49 2111 187
rect 0 0 2112 49
<< scnmos >>
rect 80 114 110 198
rect 220 114 250 198
rect 462 149 492 233
rect 534 149 564 233
rect 620 149 650 233
rect 773 149 803 233
rect 845 149 875 233
rect 953 107 983 191
rect 1085 63 1115 191
rect 1217 89 1247 217
rect 1387 133 1417 217
rect 1477 133 1507 217
rect 1563 133 1593 217
rect 1635 133 1665 217
rect 1900 77 1930 161
rect 2002 77 2032 245
<< scpmoshvt >>
rect 80 462 110 590
rect 166 462 196 590
rect 357 533 387 617
rect 443 533 473 617
rect 529 533 559 617
rect 623 533 653 617
rect 695 533 725 617
rect 802 533 832 617
rect 1135 451 1165 619
rect 1244 449 1274 617
rect 1349 517 1379 601
rect 1467 517 1497 601
rect 1607 517 1637 601
rect 1693 517 1723 601
rect 1885 367 1915 495
rect 1987 367 2017 619
<< ndiff >>
rect 27 174 80 198
rect 27 140 35 174
rect 69 140 80 174
rect 27 114 80 140
rect 110 170 220 198
rect 110 136 121 170
rect 155 136 220 170
rect 110 114 220 136
rect 250 174 303 198
rect 250 140 261 174
rect 295 140 303 174
rect 250 114 303 140
rect 409 199 462 233
rect 409 165 417 199
rect 451 165 462 199
rect 409 149 462 165
rect 492 149 534 233
rect 564 212 620 233
rect 564 178 575 212
rect 609 178 620 212
rect 564 149 620 178
rect 650 212 773 233
rect 650 178 719 212
rect 753 178 773 212
rect 650 149 773 178
rect 803 149 845 233
rect 875 191 925 233
rect 1949 228 2002 245
rect 1137 209 1217 217
rect 1137 191 1149 209
rect 875 149 953 191
rect 903 107 953 149
rect 983 107 1085 191
rect 1005 69 1085 107
rect 1005 35 1017 69
rect 1051 63 1085 69
rect 1115 175 1149 191
rect 1183 175 1217 209
rect 1115 89 1217 175
rect 1247 189 1387 217
rect 1247 155 1305 189
rect 1339 155 1387 189
rect 1247 133 1387 155
rect 1417 133 1477 217
rect 1507 189 1563 217
rect 1507 155 1518 189
rect 1552 155 1563 189
rect 1507 133 1563 155
rect 1593 133 1635 217
rect 1665 189 1718 217
rect 1665 155 1676 189
rect 1710 155 1718 189
rect 1949 194 1957 228
rect 1991 194 2002 228
rect 1949 161 2002 194
rect 1665 133 1718 155
rect 1847 136 1900 161
rect 1247 89 1347 133
rect 1115 63 1195 89
rect 1051 35 1063 63
rect 1847 102 1855 136
rect 1889 102 1900 136
rect 1847 77 1900 102
rect 1930 119 2002 161
rect 1930 85 1955 119
rect 1989 85 2002 119
rect 1930 77 2002 85
rect 2032 233 2085 245
rect 2032 199 2043 233
rect 2077 199 2085 233
rect 2032 123 2085 199
rect 2032 89 2043 123
rect 2077 89 2085 123
rect 2032 77 2085 89
rect 1005 27 1063 35
<< pdiff >>
rect 1055 631 1113 639
rect 304 591 357 617
rect 27 578 80 590
rect 27 544 35 578
rect 69 544 80 578
rect 27 510 80 544
rect 27 476 35 510
rect 69 476 80 510
rect 27 462 80 476
rect 110 569 166 590
rect 110 535 121 569
rect 155 535 166 569
rect 110 462 166 535
rect 196 576 249 590
rect 196 542 207 576
rect 241 542 249 576
rect 196 508 249 542
rect 304 557 312 591
rect 346 557 357 591
rect 304 533 357 557
rect 387 609 443 617
rect 387 575 398 609
rect 432 575 443 609
rect 387 533 443 575
rect 473 591 529 617
rect 473 557 484 591
rect 518 557 529 591
rect 473 533 529 557
rect 559 607 623 617
rect 559 573 578 607
rect 612 573 623 607
rect 559 533 623 573
rect 653 533 695 617
rect 725 609 802 617
rect 725 575 752 609
rect 786 575 802 609
rect 725 533 802 575
rect 832 591 885 617
rect 832 557 843 591
rect 877 557 885 591
rect 832 533 885 557
rect 196 474 207 508
rect 241 474 249 508
rect 196 462 249 474
rect 1055 597 1067 631
rect 1101 619 1113 631
rect 1101 597 1135 619
rect 1055 451 1135 597
rect 1165 617 1215 619
rect 1165 493 1244 617
rect 1165 459 1190 493
rect 1224 459 1244 493
rect 1165 451 1244 459
rect 1187 449 1244 451
rect 1274 601 1327 617
rect 1930 611 1987 619
rect 1274 531 1349 601
rect 1274 497 1285 531
rect 1319 517 1349 531
rect 1379 517 1467 601
rect 1497 576 1607 601
rect 1497 542 1531 576
rect 1565 542 1607 576
rect 1497 517 1607 542
rect 1637 576 1693 601
rect 1637 542 1648 576
rect 1682 542 1693 576
rect 1637 517 1693 542
rect 1723 576 1776 601
rect 1723 542 1734 576
rect 1768 542 1776 576
rect 1723 517 1776 542
rect 1930 577 1942 611
rect 1976 577 1987 611
rect 1319 497 1327 517
rect 1274 449 1327 497
rect 1930 515 1987 577
rect 1930 495 1942 515
rect 1832 482 1885 495
rect 1832 448 1840 482
rect 1874 448 1885 482
rect 1832 414 1885 448
rect 1832 380 1840 414
rect 1874 380 1885 414
rect 1832 367 1885 380
rect 1915 481 1942 495
rect 1976 481 1987 515
rect 1915 419 1987 481
rect 1915 385 1933 419
rect 1967 385 1987 419
rect 1915 367 1987 385
rect 2017 599 2070 619
rect 2017 565 2028 599
rect 2062 565 2070 599
rect 2017 509 2070 565
rect 2017 475 2028 509
rect 2062 475 2070 509
rect 2017 419 2070 475
rect 2017 385 2028 419
rect 2062 385 2070 419
rect 2017 367 2070 385
<< ndiffc >>
rect 35 140 69 174
rect 121 136 155 170
rect 261 140 295 174
rect 417 165 451 199
rect 575 178 609 212
rect 719 178 753 212
rect 1017 35 1051 69
rect 1149 175 1183 209
rect 1305 155 1339 189
rect 1518 155 1552 189
rect 1676 155 1710 189
rect 1957 194 1991 228
rect 1855 102 1889 136
rect 1955 85 1989 119
rect 2043 199 2077 233
rect 2043 89 2077 123
<< pdiffc >>
rect 35 544 69 578
rect 35 476 69 510
rect 121 535 155 569
rect 207 542 241 576
rect 312 557 346 591
rect 398 575 432 609
rect 484 557 518 591
rect 578 573 612 607
rect 752 575 786 609
rect 843 557 877 591
rect 207 474 241 508
rect 1067 597 1101 631
rect 1190 459 1224 493
rect 1285 497 1319 531
rect 1531 542 1565 576
rect 1648 542 1682 576
rect 1734 542 1768 576
rect 1942 577 1976 611
rect 1840 448 1874 482
rect 1840 380 1874 414
rect 1942 481 1976 515
rect 1933 385 1967 419
rect 2028 565 2062 599
rect 2028 475 2062 509
rect 2028 385 2062 419
<< poly >>
rect 357 617 387 643
rect 443 617 473 643
rect 529 617 559 643
rect 623 617 653 643
rect 695 617 725 643
rect 802 617 832 643
rect 80 590 110 616
rect 166 590 196 616
rect 917 597 983 613
rect 917 563 933 597
rect 967 563 983 597
rect 80 424 110 462
rect 44 408 110 424
rect 44 374 60 408
rect 94 374 110 408
rect 44 340 110 374
rect 44 306 60 340
rect 94 306 110 340
rect 44 290 110 306
rect 80 198 110 290
rect 166 354 196 462
rect 166 338 250 354
rect 166 304 182 338
rect 216 304 250 338
rect 166 270 250 304
rect 166 236 182 270
rect 216 236 250 270
rect 166 220 250 236
rect 220 198 250 220
rect 80 88 110 114
rect 220 88 250 114
rect 357 75 387 533
rect 443 367 473 533
rect 529 481 559 533
rect 515 465 581 481
rect 515 431 531 465
rect 565 431 581 465
rect 515 415 581 431
rect 443 351 509 367
rect 443 317 459 351
rect 493 331 509 351
rect 493 317 564 331
rect 623 321 653 533
rect 695 405 725 533
rect 802 509 832 533
rect 917 529 983 563
rect 917 509 933 529
rect 802 495 933 509
rect 967 495 983 529
rect 802 479 983 495
rect 695 389 911 405
rect 695 375 861 389
rect 845 355 861 375
rect 895 355 911 389
rect 443 301 564 317
rect 462 233 492 259
rect 534 233 564 301
rect 620 305 695 321
rect 620 271 645 305
rect 679 271 695 305
rect 620 255 695 271
rect 737 311 803 327
rect 737 277 753 311
rect 787 277 803 311
rect 737 261 803 277
rect 620 233 650 255
rect 773 233 803 261
rect 845 321 911 355
rect 845 287 861 321
rect 895 287 911 321
rect 845 271 911 287
rect 845 233 875 271
rect 953 191 983 479
rect 1135 619 1165 645
rect 1244 617 1274 643
rect 1135 419 1165 451
rect 1349 601 1379 627
rect 1467 601 1497 627
rect 1607 601 1637 627
rect 1693 601 1723 627
rect 1987 619 2017 645
rect 1031 403 1165 419
rect 1244 417 1274 449
rect 1031 369 1047 403
rect 1081 389 1165 403
rect 1207 401 1274 417
rect 1081 369 1097 389
rect 1031 353 1097 369
rect 1207 367 1223 401
rect 1257 387 1274 401
rect 1349 443 1379 517
rect 1467 485 1497 517
rect 1467 469 1565 485
rect 1349 427 1425 443
rect 1349 393 1375 427
rect 1409 393 1425 427
rect 1467 435 1515 469
rect 1549 435 1565 469
rect 1467 419 1565 435
rect 1257 367 1273 387
rect 1031 279 1061 353
rect 1207 351 1273 367
rect 1349 359 1425 393
rect 1349 339 1375 359
rect 1315 325 1375 339
rect 1409 325 1425 359
rect 1315 309 1425 325
rect 1315 303 1345 309
rect 1031 263 1115 279
rect 1031 229 1047 263
rect 1081 229 1115 263
rect 1031 213 1115 229
rect 1217 273 1345 303
rect 1217 217 1247 273
rect 1387 217 1417 243
rect 1477 217 1507 419
rect 1607 377 1637 517
rect 1563 361 1637 377
rect 1693 373 1723 517
rect 1885 495 1915 521
rect 1563 327 1579 361
rect 1613 327 1637 361
rect 1563 311 1637 327
rect 1679 357 1745 373
rect 1679 323 1695 357
rect 1729 323 1745 357
rect 1563 217 1593 311
rect 1679 289 1745 323
rect 1679 269 1695 289
rect 1635 255 1695 269
rect 1729 269 1745 289
rect 1885 269 1915 367
rect 1987 333 2017 367
rect 1729 255 1915 269
rect 1957 317 2032 333
rect 1957 283 1973 317
rect 2007 283 2032 317
rect 1957 267 2032 283
rect 1635 239 1915 255
rect 2002 245 2032 267
rect 1635 217 1665 239
rect 1885 219 1915 239
rect 1085 191 1115 213
rect 462 75 492 149
rect 534 123 564 149
rect 620 123 650 149
rect 773 123 803 149
rect 845 123 875 149
rect 953 75 983 107
rect 357 45 983 75
rect 1885 189 1930 219
rect 1900 161 1930 189
rect 1387 111 1417 133
rect 1369 95 1435 111
rect 1477 107 1507 133
rect 1563 107 1593 133
rect 1635 107 1665 133
rect 1217 63 1247 89
rect 1085 37 1115 63
rect 1369 61 1385 95
rect 1419 61 1435 95
rect 1369 45 1435 61
rect 1900 51 1930 77
rect 2002 51 2032 77
<< polycont >>
rect 933 563 967 597
rect 60 374 94 408
rect 60 306 94 340
rect 182 304 216 338
rect 182 236 216 270
rect 531 431 565 465
rect 459 317 493 351
rect 933 495 967 529
rect 861 355 895 389
rect 645 271 679 305
rect 753 277 787 311
rect 861 287 895 321
rect 1047 369 1081 403
rect 1223 367 1257 401
rect 1375 393 1409 427
rect 1515 435 1549 469
rect 1375 325 1409 359
rect 1047 229 1081 263
rect 1579 327 1613 361
rect 1695 323 1729 357
rect 1695 255 1729 289
rect 1973 283 2007 317
rect 1385 61 1419 95
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 19 578 71 594
rect 19 544 35 578
rect 69 544 71 578
rect 19 510 71 544
rect 105 569 171 649
rect 382 609 448 649
rect 105 535 121 569
rect 155 535 171 569
rect 105 528 171 535
rect 205 576 257 592
rect 205 542 207 576
rect 241 542 257 576
rect 19 476 35 510
rect 69 494 71 510
rect 205 508 257 542
rect 69 476 167 494
rect 19 460 167 476
rect 19 408 94 426
rect 19 374 60 408
rect 19 340 94 374
rect 19 306 60 340
rect 19 290 94 306
rect 133 354 167 460
rect 205 474 207 508
rect 241 474 257 508
rect 296 591 348 607
rect 296 557 312 591
rect 346 557 348 591
rect 382 575 398 609
rect 432 575 448 609
rect 562 607 717 615
rect 382 569 448 575
rect 482 591 528 607
rect 296 535 348 557
rect 482 557 484 591
rect 518 557 528 591
rect 562 573 578 607
rect 612 573 717 607
rect 562 569 717 573
rect 482 535 528 557
rect 296 501 649 535
rect 205 467 257 474
rect 205 465 581 467
rect 205 431 531 465
rect 565 431 581 465
rect 205 427 581 431
rect 205 424 297 427
rect 205 390 223 424
rect 257 390 297 424
rect 615 391 649 501
rect 683 523 717 569
rect 751 609 795 649
rect 751 575 752 609
rect 786 575 795 609
rect 1051 631 1117 649
rect 751 559 795 575
rect 829 591 883 607
rect 1051 597 1067 631
rect 1101 597 1117 631
rect 829 557 843 591
rect 877 557 883 591
rect 829 523 883 557
rect 683 489 883 523
rect 917 563 933 597
rect 967 563 983 597
rect 1051 595 1117 597
rect 917 561 983 563
rect 1153 581 1479 615
rect 1153 561 1187 581
rect 917 529 1187 561
rect 917 495 933 529
rect 967 527 1187 529
rect 1274 531 1339 547
rect 967 495 983 527
rect 1274 497 1285 531
rect 1319 497 1339 531
rect 839 459 883 489
rect 1153 459 1190 493
rect 1224 459 1240 493
rect 205 388 297 390
rect 133 338 225 354
rect 133 304 182 338
rect 216 304 225 338
rect 133 270 225 304
rect 133 256 182 270
rect 19 236 182 256
rect 216 236 225 270
rect 19 220 225 236
rect 19 174 85 220
rect 19 140 35 174
rect 69 140 85 174
rect 19 124 85 140
rect 119 170 157 186
rect 119 136 121 170
rect 155 136 157 170
rect 119 17 157 136
rect 191 90 225 220
rect 259 174 297 388
rect 394 351 509 368
rect 394 317 459 351
rect 493 317 509 351
rect 394 303 509 317
rect 571 357 649 391
rect 691 424 803 436
rect 839 425 1097 459
rect 691 390 703 424
rect 737 390 803 424
rect 1031 403 1097 425
rect 691 375 803 390
rect 259 140 261 174
rect 295 140 297 174
rect 259 124 297 140
rect 331 235 537 269
rect 331 90 365 235
rect 191 56 365 90
rect 401 199 467 201
rect 401 165 417 199
rect 451 165 467 199
rect 401 17 467 165
rect 503 128 537 235
rect 571 212 611 357
rect 571 178 575 212
rect 609 178 611 212
rect 571 162 611 178
rect 645 305 679 321
rect 645 128 679 271
rect 737 311 803 375
rect 737 277 753 311
rect 787 277 803 311
rect 737 262 803 277
rect 845 389 911 391
rect 845 355 861 389
rect 895 355 911 389
rect 1031 369 1047 403
rect 1081 369 1097 403
rect 1153 453 1240 459
rect 1274 453 1339 497
rect 845 333 911 355
rect 1153 333 1187 453
rect 1221 401 1269 417
rect 1221 367 1223 401
rect 1257 367 1269 401
rect 1221 351 1269 367
rect 845 321 1187 333
rect 845 287 861 321
rect 895 299 1187 321
rect 895 287 911 299
rect 845 271 911 287
rect 1031 229 1047 263
rect 1081 229 1097 263
rect 1031 228 1097 229
rect 713 212 1097 228
rect 713 178 719 212
rect 753 186 1097 212
rect 1133 213 1187 299
rect 1133 209 1199 213
rect 753 178 829 186
rect 713 162 829 178
rect 1133 175 1149 209
rect 1183 175 1199 209
rect 1235 141 1269 351
rect 894 128 1269 141
rect 1303 273 1339 453
rect 1373 427 1411 443
rect 1373 390 1375 427
rect 1409 390 1411 427
rect 1373 359 1411 390
rect 1373 325 1375 359
rect 1409 325 1411 359
rect 1373 309 1411 325
rect 1445 377 1479 581
rect 1513 576 1581 649
rect 1513 542 1531 576
rect 1565 542 1581 576
rect 1513 526 1581 542
rect 1632 576 1693 592
rect 1632 542 1648 576
rect 1682 542 1693 576
rect 1632 485 1693 542
rect 1727 576 1784 649
rect 1727 542 1734 576
rect 1768 542 1784 576
rect 1727 526 1784 542
rect 1917 611 1992 649
rect 1917 577 1942 611
rect 1976 577 1992 611
rect 1917 515 1992 577
rect 1513 469 1693 485
rect 1513 435 1515 469
rect 1549 453 1693 469
rect 1833 482 1878 498
rect 1549 435 1799 453
rect 1513 419 1799 435
rect 1445 361 1629 377
rect 1445 327 1579 361
rect 1613 327 1629 361
rect 1445 311 1629 327
rect 1679 357 1731 373
rect 1679 323 1695 357
rect 1729 323 1731 357
rect 1679 289 1731 323
rect 1679 273 1695 289
rect 1303 255 1695 273
rect 1729 255 1731 289
rect 1303 239 1731 255
rect 1303 189 1355 239
rect 1765 205 1799 419
rect 1303 155 1305 189
rect 1339 155 1355 189
rect 1303 139 1355 155
rect 1502 189 1568 205
rect 1502 155 1518 189
rect 1552 155 1568 189
rect 503 105 1269 128
rect 503 94 967 105
rect 1101 95 1435 105
rect 1001 69 1067 71
rect 1001 35 1017 69
rect 1051 35 1067 69
rect 1101 61 1385 95
rect 1419 61 1435 95
rect 1101 51 1435 61
rect 1001 17 1067 35
rect 1502 17 1568 155
rect 1660 189 1799 205
rect 1660 155 1676 189
rect 1710 155 1799 189
rect 1660 139 1799 155
rect 1833 448 1840 482
rect 1874 448 1878 482
rect 1833 414 1878 448
rect 1833 380 1840 414
rect 1874 380 1878 414
rect 1833 333 1878 380
rect 1917 481 1942 515
rect 1976 481 1992 515
rect 1917 419 1992 481
rect 1917 385 1933 419
rect 1967 385 1992 419
rect 1917 369 1992 385
rect 2026 599 2095 615
rect 2026 565 2028 599
rect 2062 565 2095 599
rect 2026 509 2095 565
rect 2026 475 2028 509
rect 2062 475 2095 509
rect 2026 419 2095 475
rect 2026 385 2028 419
rect 2062 385 2095 419
rect 2026 369 2095 385
rect 1833 317 2007 333
rect 1833 283 1973 317
rect 1833 267 2007 283
rect 1833 136 1905 267
rect 2041 233 2095 369
rect 1833 102 1855 136
rect 1889 102 1905 136
rect 1833 86 1905 102
rect 1939 228 2007 233
rect 1939 194 1957 228
rect 1991 194 2007 228
rect 1939 119 2007 194
rect 1939 85 1955 119
rect 1989 85 2007 119
rect 1939 17 2007 85
rect 2041 199 2043 233
rect 2077 199 2095 233
rect 2041 123 2095 199
rect 2041 89 2043 123
rect 2077 89 2095 123
rect 2041 73 2095 89
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 223 390 257 424
rect 703 390 737 424
rect 1375 393 1409 424
rect 1375 390 1409 393
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 691 424 749 430
rect 691 421 703 424
rect 257 393 703 421
rect 257 390 269 393
rect 211 384 269 390
rect 691 390 703 393
rect 737 421 749 424
rect 1363 424 1421 430
rect 1363 421 1375 424
rect 737 393 1375 421
rect 737 390 749 393
rect 691 384 749 390
rect 1363 390 1375 393
rect 1409 390 1421 424
rect 1363 384 1421 390
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfrtp_1
flabel comment s 1045 321 1045 321 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2047 94 2081 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 168 2081 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 570756
string GDS_START 555284
<< end >>
