magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 337 998 704
rect -38 331 311 337
rect 656 331 998 337
<< pwell >>
rect 353 211 615 295
rect 353 157 959 211
rect 1 49 959 157
rect 0 0 960 49
<< scnmos >>
rect 436 185 466 269
rect 508 185 538 269
rect 84 47 114 131
rect 156 47 186 131
rect 242 47 272 131
rect 320 47 350 131
rect 610 101 640 185
rect 688 101 718 185
rect 774 101 804 185
rect 846 101 876 185
<< scpmoshvt >>
rect 84 409 134 609
rect 320 373 370 573
rect 578 419 628 619
rect 676 419 726 619
rect 804 419 854 619
<< ndiff >>
rect 379 229 436 269
rect 379 195 391 229
rect 425 195 436 229
rect 379 185 436 195
rect 466 185 508 269
rect 538 185 589 269
rect 553 151 610 185
rect 27 111 84 131
rect 27 77 39 111
rect 73 77 84 111
rect 27 47 84 77
rect 114 47 156 131
rect 186 103 242 131
rect 186 69 197 103
rect 231 69 242 103
rect 186 47 242 69
rect 272 47 320 131
rect 350 111 407 131
rect 350 77 361 111
rect 395 77 407 111
rect 553 117 565 151
rect 599 117 610 151
rect 553 101 610 117
rect 640 101 688 185
rect 718 151 774 185
rect 718 117 729 151
rect 763 117 774 151
rect 718 101 774 117
rect 804 101 846 185
rect 876 160 933 185
rect 876 126 887 160
rect 921 126 933 160
rect 876 101 933 126
rect 350 47 407 77
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 191 609
rect 134 563 145 597
rect 179 563 191 597
rect 521 591 578 619
rect 134 526 191 563
rect 134 492 145 526
rect 179 492 191 526
rect 134 455 191 492
rect 134 421 145 455
rect 179 421 191 455
rect 134 409 191 421
rect 263 561 320 573
rect 263 527 275 561
rect 309 527 320 561
rect 263 490 320 527
rect 263 456 275 490
rect 309 456 320 490
rect 263 419 320 456
rect 263 385 275 419
rect 309 385 320 419
rect 263 373 320 385
rect 370 527 427 573
rect 370 493 381 527
rect 415 493 427 527
rect 370 419 427 493
rect 521 557 533 591
rect 567 557 578 591
rect 521 419 578 557
rect 628 419 676 619
rect 726 596 804 619
rect 726 562 737 596
rect 771 562 804 596
rect 726 419 804 562
rect 854 597 911 619
rect 854 563 865 597
rect 899 563 911 597
rect 854 465 911 563
rect 854 431 865 465
rect 899 431 911 465
rect 854 419 911 431
rect 370 385 381 419
rect 415 385 427 419
rect 370 373 427 385
<< ndiffc >>
rect 391 195 425 229
rect 39 77 73 111
rect 197 69 231 103
rect 361 77 395 111
rect 565 117 599 151
rect 729 117 763 151
rect 887 126 921 160
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 492 179 526
rect 145 421 179 455
rect 275 527 309 561
rect 275 456 309 490
rect 275 385 309 419
rect 381 493 415 527
rect 533 557 567 591
rect 737 562 771 596
rect 865 563 899 597
rect 865 431 899 465
rect 381 385 415 419
<< poly >>
rect 84 609 134 635
rect 578 619 628 645
rect 676 619 726 645
rect 804 619 854 645
rect 320 573 370 599
rect 84 369 134 409
rect 578 387 628 419
rect 84 353 155 369
rect 84 319 105 353
rect 139 319 155 353
rect 84 285 155 319
rect 84 251 105 285
rect 139 251 155 285
rect 84 235 155 251
rect 203 274 272 290
rect 203 240 219 274
rect 253 254 272 274
rect 320 284 370 373
rect 508 371 628 387
rect 508 351 578 371
rect 436 337 578 351
rect 612 337 628 371
rect 436 321 628 337
rect 320 254 350 284
rect 436 269 466 321
rect 508 269 538 321
rect 676 273 726 419
rect 804 379 854 419
rect 774 363 854 379
rect 774 329 795 363
rect 829 329 854 363
rect 774 295 854 329
rect 253 240 350 254
rect 84 176 114 235
rect 203 224 350 240
rect 84 146 186 176
rect 84 131 114 146
rect 156 131 186 146
rect 242 131 272 224
rect 320 131 350 224
rect 610 257 718 273
rect 610 223 649 257
rect 683 223 718 257
rect 610 207 718 223
rect 610 185 640 207
rect 688 185 718 207
rect 774 261 795 295
rect 829 275 854 295
rect 829 261 876 275
rect 774 245 876 261
rect 774 185 804 245
rect 846 185 876 245
rect 436 159 466 185
rect 508 159 538 185
rect 610 75 640 101
rect 688 75 718 101
rect 774 75 804 101
rect 846 75 876 101
rect 84 21 114 47
rect 156 21 186 47
rect 242 21 272 47
rect 320 21 350 47
<< polycont >>
rect 105 319 139 353
rect 105 251 139 285
rect 219 240 253 274
rect 578 337 612 371
rect 795 329 829 363
rect 649 223 683 257
rect 795 261 829 295
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 19 597 89 613
rect 19 563 39 597
rect 73 563 89 597
rect 19 526 89 563
rect 19 492 39 526
rect 73 492 89 526
rect 19 455 89 492
rect 19 421 39 455
rect 73 421 89 455
rect 19 405 89 421
rect 129 597 195 649
rect 129 563 145 597
rect 179 563 195 597
rect 129 526 195 563
rect 129 492 145 526
rect 179 492 195 526
rect 129 455 195 492
rect 129 421 145 455
rect 179 421 195 455
rect 129 405 195 421
rect 259 591 583 613
rect 259 579 533 591
rect 259 561 325 579
rect 259 527 275 561
rect 309 527 325 561
rect 517 557 533 579
rect 567 557 583 591
rect 259 490 325 527
rect 259 456 275 490
rect 309 456 325 490
rect 259 419 325 456
rect 19 199 53 405
rect 259 385 275 419
rect 309 385 325 419
rect 259 369 325 385
rect 365 527 431 543
rect 517 536 583 557
rect 721 596 787 649
rect 721 562 737 596
rect 771 562 787 596
rect 721 536 787 562
rect 849 597 915 613
rect 849 563 865 597
rect 899 578 915 597
rect 899 563 937 578
rect 365 493 381 527
rect 415 493 431 527
rect 365 419 431 493
rect 365 385 381 419
rect 415 385 431 419
rect 89 353 167 369
rect 89 319 105 353
rect 139 319 167 353
rect 89 285 167 319
rect 365 299 431 385
rect 492 466 813 500
rect 492 299 526 466
rect 562 371 743 430
rect 562 337 578 371
rect 612 337 743 371
rect 562 335 743 337
rect 779 379 813 466
rect 849 465 937 563
rect 849 431 865 465
rect 899 431 937 465
rect 849 415 937 431
rect 779 363 845 379
rect 779 329 795 363
rect 829 329 845 363
rect 89 251 105 285
rect 139 251 167 285
rect 89 235 167 251
rect 203 274 269 290
rect 203 240 219 274
rect 253 240 269 274
rect 203 199 269 240
rect 19 165 269 199
rect 305 265 565 299
rect 779 295 845 329
rect 19 111 89 165
rect 305 135 339 265
rect 375 195 391 229
rect 425 195 481 229
rect 375 179 481 195
rect 19 77 39 111
rect 73 77 89 111
rect 19 53 89 77
rect 181 103 247 129
rect 181 69 197 103
rect 231 69 247 103
rect 181 17 247 69
rect 305 111 411 135
rect 305 77 361 111
rect 395 77 411 111
rect 305 53 411 77
rect 447 17 481 179
rect 531 171 565 265
rect 601 257 743 282
rect 601 223 649 257
rect 683 223 743 257
rect 779 261 795 295
rect 829 261 845 295
rect 779 245 845 261
rect 601 207 743 223
rect 889 189 937 415
rect 531 151 615 171
rect 531 117 565 151
rect 599 117 615 151
rect 531 97 615 117
rect 713 151 779 171
rect 713 117 729 151
rect 763 117 779 151
rect 713 17 779 117
rect 871 160 937 189
rect 871 126 887 160
rect 921 126 937 160
rect 871 88 937 126
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or3b_lp
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 94 929 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 895 464 929 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 895 538 929 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1640676
string GDS_START 1632156
<< end >>
