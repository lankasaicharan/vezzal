magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3506 1975
<< nwell >>
rect -38 331 2246 704
<< pwell >>
rect 479 217 959 229
rect 1271 217 1744 235
rect 479 211 1744 217
rect 1 157 1744 211
rect 1928 157 2202 241
rect 1 49 2202 157
rect 0 0 2208 49
<< scnmos >>
rect 80 101 110 185
rect 201 101 231 185
rect 453 78 483 162
rect 555 119 585 203
rect 641 119 671 203
rect 781 119 811 203
rect 853 119 883 203
rect 961 107 991 191
rect 1124 63 1154 191
rect 1245 63 1275 191
rect 1369 125 1399 209
rect 1477 125 1507 209
rect 1563 125 1593 209
rect 1635 125 1665 209
rect 1889 47 1919 131
rect 2007 47 2037 215
rect 2093 47 2123 215
<< scpmoshvt >>
rect 80 464 110 592
rect 166 464 196 592
rect 371 535 401 619
rect 457 535 487 619
rect 543 535 573 619
rect 637 535 667 619
rect 709 535 739 619
rect 800 535 830 619
rect 1136 451 1166 619
rect 1222 451 1252 619
rect 1327 535 1357 619
rect 1399 535 1429 619
rect 1629 535 1659 619
rect 1715 535 1745 619
rect 1905 491 1935 619
rect 2007 367 2037 619
rect 2093 367 2123 619
<< ndiff >>
rect 27 160 80 185
rect 27 126 35 160
rect 69 126 80 160
rect 27 101 80 126
rect 110 160 201 185
rect 110 126 121 160
rect 155 126 201 160
rect 110 101 201 126
rect 231 169 303 185
rect 231 135 261 169
rect 295 135 303 169
rect 231 101 303 135
rect 505 162 555 203
rect 396 124 453 162
rect 396 90 408 124
rect 442 90 453 124
rect 396 78 453 90
rect 483 119 555 162
rect 585 178 641 203
rect 585 144 596 178
rect 630 144 641 178
rect 585 119 641 144
rect 671 178 781 203
rect 671 144 736 178
rect 770 144 781 178
rect 671 119 781 144
rect 811 119 853 203
rect 883 191 933 203
rect 1297 191 1369 209
rect 883 119 961 191
rect 483 78 533 119
rect 911 107 961 119
rect 991 111 1124 191
rect 991 107 1025 111
rect 1013 77 1025 107
rect 1059 77 1124 111
rect 1013 63 1124 77
rect 1154 169 1245 191
rect 1154 135 1165 169
rect 1199 135 1245 169
rect 1154 63 1245 135
rect 1275 171 1369 191
rect 1275 137 1305 171
rect 1339 137 1369 171
rect 1275 125 1369 137
rect 1399 125 1477 209
rect 1507 174 1563 209
rect 1507 140 1518 174
rect 1552 140 1563 174
rect 1507 125 1563 140
rect 1593 125 1635 209
rect 1665 184 1718 209
rect 1665 150 1676 184
rect 1710 150 1718 184
rect 1665 125 1718 150
rect 1954 198 2007 215
rect 1954 164 1962 198
rect 1996 164 2007 198
rect 1954 131 2007 164
rect 1275 63 1347 125
rect 1836 106 1889 131
rect 1836 72 1844 106
rect 1878 72 1889 106
rect 1836 47 1889 72
rect 1919 89 2007 131
rect 1919 55 1930 89
rect 1964 55 2007 89
rect 1919 47 2007 55
rect 2037 203 2093 215
rect 2037 169 2048 203
rect 2082 169 2093 203
rect 2037 101 2093 169
rect 2037 67 2048 101
rect 2082 67 2093 101
rect 2037 47 2093 67
rect 2123 203 2176 215
rect 2123 169 2134 203
rect 2168 169 2176 203
rect 2123 93 2176 169
rect 2123 59 2134 93
rect 2168 59 2176 93
rect 2123 47 2176 59
<< pdiff >>
rect 318 594 371 619
rect 27 578 80 592
rect 27 544 35 578
rect 69 544 80 578
rect 27 510 80 544
rect 27 476 35 510
rect 69 476 80 510
rect 27 464 80 476
rect 110 570 166 592
rect 110 536 121 570
rect 155 536 166 570
rect 110 464 166 536
rect 196 578 249 592
rect 196 544 207 578
rect 241 544 249 578
rect 196 510 249 544
rect 318 560 326 594
rect 360 560 371 594
rect 318 535 371 560
rect 401 594 457 619
rect 401 560 412 594
rect 446 560 457 594
rect 401 535 457 560
rect 487 594 543 619
rect 487 560 498 594
rect 532 560 543 594
rect 487 535 543 560
rect 573 594 637 619
rect 573 560 592 594
rect 626 560 637 594
rect 573 535 637 560
rect 667 535 709 619
rect 739 594 800 619
rect 739 560 755 594
rect 789 560 800 594
rect 739 535 800 560
rect 830 594 883 619
rect 830 560 841 594
rect 875 560 883 594
rect 830 535 883 560
rect 1017 597 1136 619
rect 1017 563 1029 597
rect 1063 563 1136 597
rect 196 476 207 510
rect 241 476 249 510
rect 196 464 249 476
rect 1017 451 1136 563
rect 1166 531 1222 619
rect 1166 497 1177 531
rect 1211 497 1222 531
rect 1166 451 1222 497
rect 1252 535 1327 619
rect 1357 535 1399 619
rect 1429 594 1629 619
rect 1429 560 1457 594
rect 1491 560 1582 594
rect 1616 560 1629 594
rect 1429 535 1629 560
rect 1659 594 1715 619
rect 1659 560 1670 594
rect 1704 560 1715 594
rect 1659 535 1715 560
rect 1745 594 1798 619
rect 1745 560 1756 594
rect 1790 560 1798 594
rect 1745 535 1798 560
rect 1852 607 1905 619
rect 1852 573 1860 607
rect 1894 573 1905 607
rect 1852 539 1905 573
rect 1252 531 1305 535
rect 1252 497 1263 531
rect 1297 497 1305 531
rect 1252 451 1305 497
rect 1852 505 1860 539
rect 1894 505 1905 539
rect 1852 491 1905 505
rect 1935 607 2007 619
rect 1935 573 1946 607
rect 1980 573 2007 607
rect 1935 513 2007 573
rect 1935 491 1962 513
rect 1954 479 1962 491
rect 1996 479 2007 513
rect 1954 413 2007 479
rect 1954 379 1962 413
rect 1996 379 2007 413
rect 1954 367 2007 379
rect 2037 599 2093 619
rect 2037 565 2048 599
rect 2082 565 2093 599
rect 2037 508 2093 565
rect 2037 474 2048 508
rect 2082 474 2093 508
rect 2037 420 2093 474
rect 2037 386 2048 420
rect 2082 386 2093 420
rect 2037 367 2093 386
rect 2123 607 2176 619
rect 2123 573 2134 607
rect 2168 573 2176 607
rect 2123 513 2176 573
rect 2123 479 2134 513
rect 2168 479 2176 513
rect 2123 413 2176 479
rect 2123 379 2134 413
rect 2168 379 2176 413
rect 2123 367 2176 379
<< ndiffc >>
rect 35 126 69 160
rect 121 126 155 160
rect 261 135 295 169
rect 408 90 442 124
rect 596 144 630 178
rect 736 144 770 178
rect 1025 77 1059 111
rect 1165 135 1199 169
rect 1305 137 1339 171
rect 1518 140 1552 174
rect 1676 150 1710 184
rect 1962 164 1996 198
rect 1844 72 1878 106
rect 1930 55 1964 89
rect 2048 169 2082 203
rect 2048 67 2082 101
rect 2134 169 2168 203
rect 2134 59 2168 93
<< pdiffc >>
rect 35 544 69 578
rect 35 476 69 510
rect 121 536 155 570
rect 207 544 241 578
rect 326 560 360 594
rect 412 560 446 594
rect 498 560 532 594
rect 592 560 626 594
rect 755 560 789 594
rect 841 560 875 594
rect 1029 563 1063 597
rect 207 476 241 510
rect 1177 497 1211 531
rect 1457 560 1491 594
rect 1582 560 1616 594
rect 1670 560 1704 594
rect 1756 560 1790 594
rect 1860 573 1894 607
rect 1263 497 1297 531
rect 1860 505 1894 539
rect 1946 573 1980 607
rect 1962 479 1996 513
rect 1962 379 1996 413
rect 2048 565 2082 599
rect 2048 474 2082 508
rect 2048 386 2082 420
rect 2134 573 2168 607
rect 2134 479 2168 513
rect 2134 379 2168 413
<< poly >>
rect 371 619 401 645
rect 457 619 487 645
rect 543 619 573 645
rect 637 619 667 645
rect 709 619 739 645
rect 800 619 830 645
rect 1136 619 1166 645
rect 1222 619 1252 645
rect 1327 619 1357 645
rect 1399 619 1429 645
rect 1629 619 1659 645
rect 1715 619 1745 645
rect 1905 619 1935 645
rect 2007 619 2037 645
rect 2093 619 2123 645
rect 80 592 110 618
rect 166 592 196 618
rect 80 424 110 464
rect 44 408 110 424
rect 44 374 60 408
rect 94 374 110 408
rect 44 340 110 374
rect 166 341 196 464
rect 371 454 401 535
rect 321 424 401 454
rect 44 306 60 340
rect 94 306 110 340
rect 44 290 110 306
rect 80 185 110 290
rect 158 325 231 341
rect 158 291 174 325
rect 208 291 231 325
rect 158 257 231 291
rect 158 223 174 257
rect 208 223 231 257
rect 158 207 231 223
rect 201 185 231 207
rect 80 75 110 101
rect 201 75 231 101
rect 321 51 351 424
rect 457 376 487 535
rect 543 451 573 535
rect 529 435 595 451
rect 529 401 545 435
rect 579 401 595 435
rect 529 385 595 401
rect 399 360 487 376
rect 399 326 415 360
rect 449 346 487 360
rect 449 326 479 346
rect 399 292 479 326
rect 637 293 667 535
rect 709 441 739 535
rect 800 513 830 535
rect 800 497 997 513
rect 800 483 935 497
rect 919 463 935 483
rect 969 463 997 497
rect 919 447 997 463
rect 709 411 873 441
rect 735 347 801 363
rect 735 313 751 347
rect 785 313 801 347
rect 843 349 873 411
rect 843 333 919 349
rect 843 319 869 333
rect 735 297 801 313
rect 399 258 415 292
rect 449 272 479 292
rect 627 277 693 293
rect 449 258 585 272
rect 399 242 585 258
rect 555 203 585 242
rect 627 243 643 277
rect 677 243 693 277
rect 627 227 693 243
rect 771 271 801 297
rect 853 299 869 319
rect 903 299 919 333
rect 853 283 919 299
rect 771 241 811 271
rect 641 203 671 227
rect 781 203 811 241
rect 853 203 883 283
rect 967 243 997 447
rect 1136 419 1166 451
rect 961 213 997 243
rect 1063 403 1166 419
rect 1222 415 1252 451
rect 1327 425 1357 535
rect 1399 503 1429 535
rect 1399 487 1565 503
rect 1399 473 1515 487
rect 1477 453 1515 473
rect 1549 453 1565 487
rect 1629 467 1659 535
rect 1477 437 1565 453
rect 1607 451 1673 467
rect 1063 369 1079 403
rect 1113 389 1166 403
rect 1219 399 1285 415
rect 1113 369 1129 389
rect 1063 353 1129 369
rect 1219 365 1235 399
rect 1269 365 1285 399
rect 1063 279 1093 353
rect 1219 349 1285 365
rect 1327 409 1425 425
rect 1327 375 1375 409
rect 1409 375 1425 409
rect 1327 341 1425 375
rect 1327 307 1375 341
rect 1409 307 1425 341
rect 1245 291 1425 307
rect 1063 263 1154 279
rect 1063 229 1079 263
rect 1113 229 1154 263
rect 1063 213 1154 229
rect 453 162 483 188
rect 961 191 991 213
rect 1124 191 1154 213
rect 1245 277 1357 291
rect 1245 191 1275 277
rect 1369 209 1399 235
rect 1477 209 1507 437
rect 1607 417 1623 451
rect 1657 417 1673 451
rect 1607 383 1673 417
rect 1607 363 1623 383
rect 1563 349 1623 363
rect 1657 349 1673 383
rect 1715 399 1745 535
rect 1715 383 1787 399
rect 1715 369 1737 383
rect 1563 333 1673 349
rect 1721 349 1737 369
rect 1771 349 1787 383
rect 1905 381 1935 491
rect 1563 209 1593 333
rect 1721 315 1787 349
rect 1721 285 1737 315
rect 1635 281 1737 285
rect 1771 285 1787 315
rect 1889 351 1935 381
rect 1889 285 1919 351
rect 2007 303 2037 367
rect 1771 281 1919 285
rect 1635 255 1919 281
rect 1635 209 1665 255
rect 555 93 585 119
rect 641 93 671 119
rect 781 93 811 119
rect 853 93 883 119
rect 453 51 483 78
rect 961 51 991 107
rect 1889 131 1919 255
rect 1961 287 2037 303
rect 1961 253 1977 287
rect 2011 267 2037 287
rect 2093 267 2123 367
rect 2011 253 2123 267
rect 1961 237 2123 253
rect 2007 215 2037 237
rect 2093 215 2123 237
rect 1369 103 1399 125
rect 1369 87 1435 103
rect 1477 99 1507 125
rect 1563 99 1593 125
rect 1635 99 1665 125
rect 321 21 991 51
rect 1124 37 1154 63
rect 1245 37 1275 63
rect 1369 53 1385 87
rect 1419 53 1435 87
rect 1369 37 1435 53
rect 1889 21 1919 47
rect 2007 21 2037 47
rect 2093 21 2123 47
<< polycont >>
rect 60 374 94 408
rect 60 306 94 340
rect 174 291 208 325
rect 174 223 208 257
rect 545 401 579 435
rect 415 326 449 360
rect 935 463 969 497
rect 751 313 785 347
rect 415 258 449 292
rect 643 243 677 277
rect 869 299 903 333
rect 1515 453 1549 487
rect 1079 369 1113 403
rect 1235 365 1269 399
rect 1375 375 1409 409
rect 1375 307 1409 341
rect 1079 229 1113 263
rect 1623 417 1657 451
rect 1623 349 1657 383
rect 1737 349 1771 383
rect 1737 281 1771 315
rect 1977 253 2011 287
rect 1385 53 1419 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 19 578 71 594
rect 19 544 35 578
rect 69 544 71 578
rect 19 510 71 544
rect 105 570 171 649
rect 310 594 362 610
rect 105 536 121 570
rect 155 536 171 570
rect 105 528 171 536
rect 205 578 257 594
rect 205 544 207 578
rect 241 544 257 578
rect 19 476 35 510
rect 69 494 71 510
rect 205 510 257 544
rect 69 476 167 494
rect 19 460 167 476
rect 31 408 94 424
rect 31 374 60 408
rect 31 340 94 374
rect 31 306 60 340
rect 31 290 94 306
rect 133 341 167 460
rect 205 476 207 510
rect 241 476 257 510
rect 310 560 326 594
rect 360 560 362 594
rect 310 519 362 560
rect 396 594 462 649
rect 396 560 412 594
rect 446 560 462 594
rect 396 553 462 560
rect 496 594 540 610
rect 496 560 498 594
rect 532 560 540 594
rect 496 519 540 560
rect 574 594 717 610
rect 574 560 592 594
rect 626 560 717 594
rect 574 553 717 560
rect 310 485 649 519
rect 205 451 257 476
rect 205 435 581 451
rect 205 417 545 435
rect 259 366 295 417
rect 529 401 545 417
rect 579 401 581 435
rect 529 385 581 401
rect 259 350 365 366
rect 133 325 225 341
rect 133 291 174 325
rect 208 291 225 325
rect 133 257 225 291
rect 133 254 174 257
rect 19 223 174 254
rect 208 223 225 257
rect 19 220 225 223
rect 19 160 78 220
rect 19 126 35 160
rect 69 126 78 160
rect 19 109 78 126
rect 112 160 157 176
rect 112 126 121 160
rect 155 126 157 160
rect 112 17 157 126
rect 191 85 225 220
rect 259 316 319 350
rect 353 316 365 350
rect 259 300 365 316
rect 399 360 465 376
rect 399 326 415 360
rect 449 326 465 360
rect 615 347 649 485
rect 683 444 717 553
rect 751 594 799 649
rect 751 560 755 594
rect 789 560 799 594
rect 751 544 799 560
rect 833 594 891 610
rect 833 560 841 594
rect 875 560 891 594
rect 833 444 891 560
rect 1013 597 1065 649
rect 1013 563 1029 597
rect 1063 563 1065 597
rect 1013 547 1065 563
rect 1099 581 1407 615
rect 1099 513 1133 581
rect 925 497 1133 513
rect 925 463 935 497
rect 969 463 1133 497
rect 925 447 1133 463
rect 1167 531 1219 547
rect 1167 497 1177 531
rect 1211 497 1219 531
rect 1167 481 1219 497
rect 1253 531 1339 547
rect 1253 497 1263 531
rect 1297 497 1339 531
rect 1253 481 1339 497
rect 683 413 891 444
rect 683 403 1129 413
rect 683 384 1079 403
rect 837 369 1079 384
rect 1113 369 1129 403
rect 259 169 297 300
rect 399 292 465 326
rect 399 258 415 292
rect 449 258 465 292
rect 399 242 465 258
rect 557 313 649 347
rect 683 316 703 350
rect 737 347 801 350
rect 737 316 751 347
rect 683 313 751 316
rect 785 313 801 347
rect 1167 335 1201 481
rect 259 135 261 169
rect 295 135 297 169
rect 259 119 297 135
rect 331 174 516 208
rect 331 85 365 174
rect 191 51 365 85
rect 399 124 448 140
rect 399 90 408 124
rect 442 90 448 124
rect 399 17 448 90
rect 482 94 516 174
rect 557 194 591 313
rect 683 311 801 313
rect 853 333 1201 335
rect 853 299 869 333
rect 903 299 1201 333
rect 627 243 643 277
rect 677 243 700 277
rect 627 228 700 243
rect 557 178 632 194
rect 557 144 596 178
rect 630 144 632 178
rect 557 128 632 144
rect 666 94 700 228
rect 734 263 1129 265
rect 734 229 1079 263
rect 1113 229 1129 263
rect 734 178 776 229
rect 734 144 736 178
rect 770 144 776 178
rect 734 128 776 144
rect 810 161 1131 195
rect 810 94 844 161
rect 482 51 844 94
rect 1009 111 1063 127
rect 1009 77 1025 111
rect 1059 77 1063 111
rect 1009 17 1063 77
rect 1097 85 1131 161
rect 1165 169 1201 299
rect 1199 135 1201 169
rect 1165 119 1201 135
rect 1235 399 1271 415
rect 1269 365 1271 399
rect 1235 87 1271 365
rect 1305 245 1339 481
rect 1373 521 1407 581
rect 1441 594 1632 649
rect 1441 560 1457 594
rect 1491 560 1582 594
rect 1616 560 1632 594
rect 1441 555 1632 560
rect 1666 594 1706 610
rect 1666 560 1670 594
rect 1704 560 1706 594
rect 1666 521 1706 560
rect 1740 594 1806 649
rect 1740 560 1756 594
rect 1790 560 1806 594
rect 1740 555 1806 560
rect 1844 607 1911 615
rect 1844 573 1860 607
rect 1894 573 1911 607
rect 1844 539 1911 573
rect 1373 459 1477 521
rect 1373 409 1409 425
rect 1373 375 1375 409
rect 1373 350 1409 375
rect 1373 307 1375 350
rect 1443 403 1477 459
rect 1515 487 1767 521
rect 1844 505 1860 539
rect 1894 505 1911 539
rect 1844 503 1911 505
rect 1549 453 1565 487
rect 1515 437 1565 453
rect 1733 469 1767 487
rect 1607 417 1623 451
rect 1657 417 1699 451
rect 1733 435 1839 469
rect 1607 403 1699 417
rect 1443 383 1699 403
rect 1443 349 1623 383
rect 1657 349 1699 383
rect 1737 383 1771 399
rect 1373 291 1409 307
rect 1737 315 1771 349
rect 1445 281 1737 299
rect 1445 265 1771 281
rect 1445 245 1479 265
rect 1305 211 1479 245
rect 1805 231 1839 435
rect 1305 171 1355 211
rect 1660 197 1839 231
rect 1873 303 1911 503
rect 1945 607 2012 649
rect 1945 573 1946 607
rect 1980 573 2012 607
rect 1945 513 2012 573
rect 1945 479 1962 513
rect 1996 479 2012 513
rect 1945 413 2012 479
rect 1945 379 1962 413
rect 1996 379 2012 413
rect 1945 363 2012 379
rect 2046 599 2091 615
rect 2046 565 2048 599
rect 2082 565 2091 599
rect 2046 508 2091 565
rect 2046 474 2048 508
rect 2082 474 2091 508
rect 2046 420 2091 474
rect 2046 386 2048 420
rect 2082 386 2091 420
rect 1873 287 2012 303
rect 1873 253 1977 287
rect 2011 253 2012 287
rect 1873 237 2012 253
rect 1660 184 1726 197
rect 1339 137 1355 171
rect 1305 121 1355 137
rect 1502 174 1568 177
rect 1502 140 1518 174
rect 1552 140 1568 174
rect 1235 85 1385 87
rect 1097 53 1385 85
rect 1419 53 1435 87
rect 1097 51 1435 53
rect 1502 17 1568 140
rect 1660 150 1676 184
rect 1710 150 1726 184
rect 1873 163 1907 237
rect 2046 203 2091 386
rect 2125 607 2184 649
rect 2125 573 2134 607
rect 2168 573 2184 607
rect 2125 513 2184 573
rect 2125 479 2134 513
rect 2168 479 2184 513
rect 2125 413 2184 479
rect 2125 379 2134 413
rect 2168 379 2184 413
rect 2125 363 2184 379
rect 1660 134 1726 150
rect 1828 129 1907 163
rect 1941 198 2012 203
rect 1941 164 1962 198
rect 1996 164 2012 198
rect 1828 106 1880 129
rect 1828 72 1844 106
rect 1878 72 1880 106
rect 1941 95 2012 164
rect 1828 51 1880 72
rect 1914 89 2012 95
rect 1914 55 1930 89
rect 1964 55 2012 89
rect 1914 17 2012 55
rect 2046 169 2048 203
rect 2082 169 2091 203
rect 2046 101 2091 169
rect 2046 67 2048 101
rect 2082 67 2091 101
rect 2046 51 2091 67
rect 2125 203 2184 219
rect 2125 169 2134 203
rect 2168 169 2184 203
rect 2125 93 2184 169
rect 2125 59 2134 93
rect 2168 59 2184 93
rect 2125 17 2184 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 319 316 353 350
rect 703 316 737 350
rect 1375 341 1409 350
rect 1375 316 1409 341
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 307 350 365 356
rect 307 316 319 350
rect 353 347 365 350
rect 691 350 749 356
rect 691 347 703 350
rect 353 319 703 347
rect 353 316 365 319
rect 307 310 365 316
rect 691 316 703 319
rect 737 347 749 350
rect 1363 350 1421 356
rect 1363 347 1375 350
rect 737 319 1375 347
rect 737 316 749 319
rect 691 310 749 316
rect 1363 316 1375 319
rect 1409 316 1421 350
rect 1363 310 1421 316
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfrtp_2
flabel comment s 1075 320 1075 320 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1663 390 1697 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2047 94 2081 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 168 2081 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 464 2081 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 538 2081 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 587510
string GDS_START 570812
<< end >>
