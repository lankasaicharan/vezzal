magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 1 49 1055 167
rect 0 0 1056 49
<< scnmos >>
rect 82 57 112 141
rect 154 57 184 141
rect 240 57 270 141
rect 312 57 342 141
rect 398 57 428 141
rect 470 57 500 141
rect 556 57 586 141
rect 628 57 658 141
rect 714 57 744 141
rect 786 57 816 141
rect 872 57 902 141
rect 944 57 974 141
<< scpmoshvt >>
rect 84 409 134 609
rect 372 417 422 617
rect 470 417 520 617
rect 584 417 634 617
rect 706 417 756 617
rect 830 417 880 617
<< ndiff >>
rect 27 116 82 141
rect 27 82 37 116
rect 71 82 82 116
rect 27 57 82 82
rect 112 57 154 141
rect 184 108 240 141
rect 184 74 195 108
rect 229 74 240 108
rect 184 57 240 74
rect 270 57 312 141
rect 342 116 398 141
rect 342 82 353 116
rect 387 82 398 116
rect 342 57 398 82
rect 428 57 470 141
rect 500 116 556 141
rect 500 82 511 116
rect 545 82 556 116
rect 500 57 556 82
rect 586 57 628 141
rect 658 116 714 141
rect 658 82 669 116
rect 703 82 714 116
rect 658 57 714 82
rect 744 57 786 141
rect 816 116 872 141
rect 816 82 827 116
rect 861 82 872 116
rect 816 57 872 82
rect 902 57 944 141
rect 974 116 1029 141
rect 974 82 985 116
rect 1019 82 1029 116
rect 974 57 1029 82
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 191 609
rect 134 563 145 597
rect 179 563 191 597
rect 134 526 191 563
rect 134 492 145 526
rect 179 492 191 526
rect 134 455 191 492
rect 134 421 145 455
rect 179 421 191 455
rect 134 409 191 421
rect 311 597 372 617
rect 311 563 323 597
rect 357 563 372 597
rect 311 463 372 563
rect 311 429 323 463
rect 357 429 372 463
rect 311 417 372 429
rect 422 417 470 617
rect 520 417 584 617
rect 634 417 706 617
rect 756 605 830 617
rect 756 571 767 605
rect 801 571 830 605
rect 756 471 830 571
rect 756 437 767 471
rect 801 437 830 471
rect 756 417 830 437
rect 880 597 937 617
rect 880 563 891 597
rect 925 563 937 597
rect 880 463 937 563
rect 880 429 891 463
rect 925 429 937 463
rect 880 417 937 429
<< ndiffc >>
rect 37 82 71 116
rect 195 74 229 108
rect 353 82 387 116
rect 511 82 545 116
rect 669 82 703 116
rect 827 82 861 116
rect 985 82 1019 116
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 492 179 526
rect 145 421 179 455
rect 323 563 357 597
rect 323 429 357 463
rect 767 571 801 605
rect 767 437 801 471
rect 891 563 925 597
rect 891 429 925 463
<< poly >>
rect 84 609 134 635
rect 372 617 422 643
rect 470 617 520 643
rect 584 617 634 643
rect 706 617 756 643
rect 830 617 880 643
rect 84 369 134 409
rect 82 353 157 369
rect 82 319 107 353
rect 141 319 157 353
rect 82 285 157 319
rect 372 299 422 417
rect 82 251 107 285
rect 141 265 157 285
rect 235 283 422 299
rect 141 251 184 265
rect 82 235 184 251
rect 82 141 112 235
rect 154 141 184 235
rect 235 249 251 283
rect 285 269 422 283
rect 470 385 520 417
rect 584 385 634 417
rect 706 385 756 417
rect 470 369 536 385
rect 470 335 486 369
rect 520 335 536 369
rect 470 301 536 335
rect 285 249 342 269
rect 235 215 342 249
rect 235 181 251 215
rect 285 181 342 215
rect 470 267 486 301
rect 520 267 536 301
rect 470 251 536 267
rect 584 369 653 385
rect 584 335 603 369
rect 637 335 653 369
rect 584 301 653 335
rect 584 267 603 301
rect 637 267 653 301
rect 584 251 653 267
rect 706 369 772 385
rect 706 335 722 369
rect 756 335 772 369
rect 830 368 880 417
rect 706 301 772 335
rect 706 267 722 301
rect 756 267 772 301
rect 706 251 772 267
rect 850 352 941 368
rect 850 318 891 352
rect 925 318 941 352
rect 850 284 941 318
rect 470 186 500 251
rect 584 186 614 251
rect 714 186 744 251
rect 850 250 891 284
rect 925 264 941 284
rect 925 250 974 264
rect 850 234 974 250
rect 235 165 342 181
rect 240 141 270 165
rect 312 141 342 165
rect 398 156 500 186
rect 398 141 428 156
rect 470 141 500 156
rect 556 156 658 186
rect 556 141 586 156
rect 628 141 658 156
rect 714 156 816 186
rect 714 141 744 156
rect 786 141 816 156
rect 872 141 902 234
rect 944 141 974 234
rect 82 31 112 57
rect 154 31 184 57
rect 240 31 270 57
rect 312 31 342 57
rect 398 31 428 57
rect 470 31 500 57
rect 556 31 586 57
rect 628 31 658 57
rect 714 31 744 57
rect 786 31 816 57
rect 872 31 902 57
rect 944 31 974 57
<< polycont >>
rect 107 319 141 353
rect 107 251 141 285
rect 251 249 285 283
rect 486 335 520 369
rect 251 181 285 215
rect 486 267 520 301
rect 603 335 637 369
rect 603 267 637 301
rect 722 335 756 369
rect 722 267 756 301
rect 891 318 925 352
rect 891 250 925 284
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 21 597 89 613
rect 21 563 39 597
rect 73 563 89 597
rect 21 526 89 563
rect 21 492 39 526
rect 73 492 89 526
rect 21 455 89 492
rect 21 421 39 455
rect 73 421 89 455
rect 21 405 89 421
rect 129 597 195 649
rect 129 563 145 597
rect 179 563 195 597
rect 129 526 195 563
rect 129 492 145 526
rect 179 492 195 526
rect 129 455 195 492
rect 129 421 145 455
rect 179 421 195 455
rect 129 405 195 421
rect 307 597 373 613
rect 307 563 323 597
rect 357 563 373 597
rect 751 605 817 649
rect 307 463 373 563
rect 307 429 323 463
rect 357 429 373 463
rect 307 413 373 429
rect 21 199 55 405
rect 91 353 167 369
rect 91 319 107 353
rect 141 319 167 353
rect 91 285 167 319
rect 91 251 107 285
rect 141 251 167 285
rect 91 235 167 251
rect 235 283 301 299
rect 235 249 251 283
rect 285 249 301 283
rect 235 215 301 249
rect 235 199 251 215
rect 21 181 251 199
rect 285 181 301 215
rect 21 165 301 181
rect 337 215 373 413
rect 409 369 551 578
rect 409 335 486 369
rect 520 335 551 369
rect 409 301 551 335
rect 409 267 486 301
rect 520 267 551 301
rect 409 251 551 267
rect 587 369 653 578
rect 751 571 767 605
rect 801 571 817 605
rect 751 471 817 571
rect 751 437 767 471
rect 801 437 817 471
rect 751 421 817 437
rect 875 597 1035 613
rect 875 563 891 597
rect 925 563 1035 597
rect 875 463 1035 563
rect 875 429 891 463
rect 925 429 1035 463
rect 875 413 1035 429
rect 587 335 603 369
rect 637 335 653 369
rect 587 301 653 335
rect 587 267 603 301
rect 637 267 653 301
rect 587 251 653 267
rect 697 369 839 385
rect 697 335 722 369
rect 756 335 839 369
rect 697 301 839 335
rect 697 267 722 301
rect 756 267 839 301
rect 697 251 839 267
rect 875 352 941 368
rect 875 318 891 352
rect 925 318 941 352
rect 875 284 941 318
rect 875 250 891 284
rect 925 250 941 284
rect 875 215 941 250
rect 337 181 941 215
rect 21 116 87 165
rect 21 82 37 116
rect 71 82 87 116
rect 21 53 87 82
rect 179 108 245 129
rect 179 74 195 108
rect 229 74 245 108
rect 179 17 245 74
rect 337 116 403 181
rect 337 82 353 116
rect 387 82 403 116
rect 337 53 403 82
rect 495 116 561 145
rect 495 82 511 116
rect 545 82 561 116
rect 495 17 561 82
rect 653 116 719 181
rect 985 145 1035 413
rect 653 82 669 116
rect 703 82 719 116
rect 653 53 719 82
rect 811 116 877 145
rect 811 82 827 116
rect 861 82 877 116
rect 811 17 877 82
rect 969 116 1035 145
rect 969 82 985 116
rect 1019 82 1035 116
rect 969 53 1035 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or4b_lp
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 991 94 1025 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 991 168 1025 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 991 464 1025 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 991 538 1025 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2909472
string GDS_START 2899692
<< end >>
