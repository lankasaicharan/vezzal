magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 3026 1975
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 4 49 1727 248
rect 0 0 1728 49
<< scnmos >>
rect 87 74 117 222
rect 173 74 203 222
rect 259 74 289 222
rect 359 74 389 222
rect 445 74 475 222
rect 533 74 563 222
rect 619 74 649 222
rect 733 74 763 222
rect 933 74 963 222
rect 1077 74 1107 222
rect 1177 74 1207 222
rect 1263 74 1293 222
rect 1363 74 1393 222
rect 1614 74 1644 222
<< scpmoshvt >>
rect 86 368 116 592
rect 176 368 206 592
rect 266 368 296 592
rect 356 368 386 592
rect 446 368 476 592
rect 546 368 576 592
rect 636 368 666 592
rect 736 368 766 592
rect 836 368 866 592
rect 936 368 966 592
rect 1132 368 1162 592
rect 1242 368 1272 592
rect 1338 368 1368 592
rect 1432 368 1462 592
rect 1522 368 1552 592
rect 1612 368 1642 592
<< ndiff >>
rect 30 210 87 222
rect 30 176 42 210
rect 76 176 87 210
rect 30 120 87 176
rect 30 86 42 120
rect 76 86 87 120
rect 30 74 87 86
rect 117 152 173 222
rect 117 118 128 152
rect 162 118 173 152
rect 117 74 173 118
rect 203 210 259 222
rect 203 176 214 210
rect 248 176 259 210
rect 203 120 259 176
rect 203 86 214 120
rect 248 86 259 120
rect 203 74 259 86
rect 289 152 359 222
rect 289 118 300 152
rect 334 118 359 152
rect 289 74 359 118
rect 389 214 445 222
rect 389 180 400 214
rect 434 180 445 214
rect 389 116 445 180
rect 389 82 400 116
rect 434 82 445 116
rect 389 74 445 82
rect 475 152 533 222
rect 475 118 487 152
rect 521 118 533 152
rect 475 74 533 118
rect 563 169 619 222
rect 563 135 574 169
rect 608 135 619 169
rect 563 74 619 135
rect 649 152 733 222
rect 649 118 674 152
rect 708 118 733 152
rect 649 74 733 118
rect 763 169 820 222
rect 763 135 774 169
rect 808 135 820 169
rect 874 210 933 222
rect 874 176 887 210
rect 921 176 933 210
rect 874 164 933 176
rect 763 123 820 135
rect 763 74 813 123
rect 883 74 933 164
rect 963 143 1077 222
rect 963 109 1003 143
rect 1037 109 1077 143
rect 963 74 1077 109
rect 1107 169 1177 222
rect 1107 135 1118 169
rect 1152 135 1177 169
rect 1107 74 1177 135
rect 1207 152 1263 222
rect 1207 118 1218 152
rect 1252 118 1263 152
rect 1207 74 1263 118
rect 1293 210 1363 222
rect 1293 176 1318 210
rect 1352 176 1363 210
rect 1293 120 1363 176
rect 1293 86 1318 120
rect 1352 86 1363 120
rect 1293 74 1363 86
rect 1393 152 1614 222
rect 1393 118 1404 152
rect 1438 118 1486 152
rect 1520 118 1569 152
rect 1603 118 1614 152
rect 1393 74 1614 118
rect 1644 210 1701 222
rect 1644 176 1655 210
rect 1689 176 1701 210
rect 1644 120 1701 176
rect 1644 86 1655 120
rect 1689 86 1701 120
rect 1644 74 1701 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 504 86 546
rect 27 470 39 504
rect 73 470 86 504
rect 27 424 86 470
rect 27 390 39 424
rect 73 390 86 424
rect 27 368 86 390
rect 116 584 176 592
rect 116 550 129 584
rect 163 550 176 584
rect 116 492 176 550
rect 116 458 129 492
rect 163 458 176 492
rect 116 368 176 458
rect 206 571 266 592
rect 206 537 219 571
rect 253 537 266 571
rect 206 497 266 537
rect 206 463 219 497
rect 253 463 266 497
rect 206 424 266 463
rect 206 390 219 424
rect 253 390 266 424
rect 206 368 266 390
rect 296 584 356 592
rect 296 550 309 584
rect 343 550 356 584
rect 296 492 356 550
rect 296 458 309 492
rect 343 458 356 492
rect 296 368 356 458
rect 386 574 446 592
rect 386 540 399 574
rect 433 540 446 574
rect 386 490 446 540
rect 386 456 399 490
rect 433 456 446 490
rect 386 410 446 456
rect 386 376 399 410
rect 433 376 446 410
rect 386 368 446 376
rect 476 584 546 592
rect 476 550 489 584
rect 523 550 546 584
rect 476 498 546 550
rect 476 464 489 498
rect 523 464 546 498
rect 476 368 546 464
rect 576 580 636 592
rect 576 546 589 580
rect 623 546 636 580
rect 576 505 636 546
rect 576 471 589 505
rect 623 471 636 505
rect 576 424 636 471
rect 576 390 589 424
rect 623 390 636 424
rect 576 368 636 390
rect 666 584 736 592
rect 666 550 689 584
rect 723 550 736 584
rect 666 492 736 550
rect 666 458 689 492
rect 723 458 736 492
rect 666 368 736 458
rect 766 580 836 592
rect 766 546 789 580
rect 823 546 836 580
rect 766 505 836 546
rect 766 471 789 505
rect 823 471 836 505
rect 766 424 836 471
rect 766 390 789 424
rect 823 390 836 424
rect 766 368 836 390
rect 866 570 936 592
rect 866 536 889 570
rect 923 536 936 570
rect 866 368 936 536
rect 966 570 1132 592
rect 966 536 980 570
rect 1014 536 1085 570
rect 1119 536 1132 570
rect 966 492 1132 536
rect 966 458 980 492
rect 1014 458 1085 492
rect 1119 458 1132 492
rect 966 368 1132 458
rect 1162 570 1242 592
rect 1162 536 1185 570
rect 1219 536 1242 570
rect 1162 368 1242 536
rect 1272 584 1338 592
rect 1272 550 1285 584
rect 1319 550 1338 584
rect 1272 492 1338 550
rect 1272 458 1285 492
rect 1319 458 1338 492
rect 1272 368 1338 458
rect 1368 542 1432 592
rect 1368 508 1385 542
rect 1419 508 1432 542
rect 1368 430 1432 508
rect 1368 396 1385 430
rect 1419 396 1432 430
rect 1368 368 1432 396
rect 1462 580 1522 592
rect 1462 546 1475 580
rect 1509 546 1522 580
rect 1462 508 1522 546
rect 1462 474 1475 508
rect 1509 474 1522 508
rect 1462 368 1522 474
rect 1552 542 1612 592
rect 1552 508 1565 542
rect 1599 508 1612 542
rect 1552 430 1612 508
rect 1552 396 1565 430
rect 1599 396 1612 430
rect 1552 368 1612 396
rect 1642 580 1701 592
rect 1642 546 1655 580
rect 1689 546 1701 580
rect 1642 512 1701 546
rect 1642 478 1655 512
rect 1689 478 1701 512
rect 1642 440 1701 478
rect 1642 406 1655 440
rect 1689 406 1701 440
rect 1642 368 1701 406
<< ndiffc >>
rect 42 176 76 210
rect 42 86 76 120
rect 128 118 162 152
rect 214 176 248 210
rect 214 86 248 120
rect 300 118 334 152
rect 400 180 434 214
rect 400 82 434 116
rect 487 118 521 152
rect 574 135 608 169
rect 674 118 708 152
rect 774 135 808 169
rect 887 176 921 210
rect 1003 109 1037 143
rect 1118 135 1152 169
rect 1218 118 1252 152
rect 1318 176 1352 210
rect 1318 86 1352 120
rect 1404 118 1438 152
rect 1486 118 1520 152
rect 1569 118 1603 152
rect 1655 176 1689 210
rect 1655 86 1689 120
<< pdiffc >>
rect 39 546 73 580
rect 39 470 73 504
rect 39 390 73 424
rect 129 550 163 584
rect 129 458 163 492
rect 219 537 253 571
rect 219 463 253 497
rect 219 390 253 424
rect 309 550 343 584
rect 309 458 343 492
rect 399 540 433 574
rect 399 456 433 490
rect 399 376 433 410
rect 489 550 523 584
rect 489 464 523 498
rect 589 546 623 580
rect 589 471 623 505
rect 589 390 623 424
rect 689 550 723 584
rect 689 458 723 492
rect 789 546 823 580
rect 789 471 823 505
rect 789 390 823 424
rect 889 536 923 570
rect 980 536 1014 570
rect 1085 536 1119 570
rect 980 458 1014 492
rect 1085 458 1119 492
rect 1185 536 1219 570
rect 1285 550 1319 584
rect 1285 458 1319 492
rect 1385 508 1419 542
rect 1385 396 1419 430
rect 1475 546 1509 580
rect 1475 474 1509 508
rect 1565 508 1599 542
rect 1565 396 1599 430
rect 1655 546 1689 580
rect 1655 478 1689 512
rect 1655 406 1689 440
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 266 592 296 618
rect 356 592 386 618
rect 446 592 476 618
rect 546 592 576 618
rect 636 592 666 618
rect 736 592 766 618
rect 836 592 866 618
rect 936 592 966 618
rect 1132 592 1162 618
rect 1242 592 1272 618
rect 1338 592 1368 618
rect 1432 592 1462 618
rect 1522 592 1552 618
rect 1612 592 1642 618
rect 86 353 116 368
rect 176 353 206 368
rect 266 353 296 368
rect 356 353 386 368
rect 446 353 476 368
rect 546 353 576 368
rect 636 353 666 368
rect 736 353 766 368
rect 836 353 866 368
rect 936 353 966 368
rect 1132 353 1162 368
rect 1242 353 1272 368
rect 1338 353 1368 368
rect 1432 353 1462 368
rect 1522 353 1552 368
rect 1612 353 1642 368
rect 83 336 119 353
rect 173 336 209 353
rect 263 336 299 353
rect 353 336 389 353
rect 83 320 389 336
rect 83 286 103 320
rect 137 286 171 320
rect 205 286 239 320
rect 273 286 307 320
rect 341 286 389 320
rect 443 337 479 353
rect 543 337 579 353
rect 443 336 579 337
rect 633 336 669 353
rect 733 336 769 353
rect 443 320 769 336
rect 833 336 969 353
rect 1129 336 1165 353
rect 1239 336 1275 353
rect 833 323 1275 336
rect 443 300 491 320
rect 83 270 389 286
rect 87 222 117 270
rect 173 222 203 270
rect 259 222 289 270
rect 359 222 389 270
rect 445 286 491 300
rect 525 286 559 320
rect 593 286 627 320
rect 661 286 695 320
rect 729 300 769 320
rect 933 320 1275 323
rect 729 286 763 300
rect 445 270 763 286
rect 445 222 475 270
rect 533 222 563 270
rect 619 222 649 270
rect 733 222 763 270
rect 933 286 1021 320
rect 1055 286 1089 320
rect 1123 286 1157 320
rect 1191 294 1275 320
rect 1335 336 1371 353
rect 1429 336 1465 353
rect 1519 336 1555 353
rect 1609 336 1645 353
rect 1335 320 1645 336
rect 1191 286 1293 294
rect 933 264 1293 286
rect 1335 286 1351 320
rect 1385 286 1419 320
rect 1453 286 1487 320
rect 1521 306 1645 320
rect 1521 286 1644 306
rect 1335 270 1644 286
rect 933 222 963 264
rect 1077 222 1107 264
rect 1177 222 1207 264
rect 1263 222 1293 264
rect 1363 222 1393 270
rect 1614 222 1644 270
rect 87 48 117 74
rect 173 48 203 74
rect 259 48 289 74
rect 359 48 389 74
rect 445 48 475 74
rect 533 48 563 74
rect 619 48 649 74
rect 733 48 763 74
rect 933 48 963 74
rect 1077 48 1107 74
rect 1177 48 1207 74
rect 1263 48 1293 74
rect 1363 48 1393 74
rect 1614 48 1644 74
<< polycont >>
rect 103 286 137 320
rect 171 286 205 320
rect 239 286 273 320
rect 307 286 341 320
rect 491 286 525 320
rect 559 286 593 320
rect 627 286 661 320
rect 695 286 729 320
rect 1021 286 1055 320
rect 1089 286 1123 320
rect 1157 286 1191 320
rect 1351 286 1385 320
rect 1419 286 1453 320
rect 1487 286 1521 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 580 79 596
rect 23 546 39 580
rect 73 546 79 580
rect 23 504 79 546
rect 23 470 39 504
rect 73 470 79 504
rect 23 424 79 470
rect 113 584 179 649
rect 113 550 129 584
rect 163 550 179 584
rect 113 492 179 550
rect 113 458 129 492
rect 163 458 179 492
rect 213 571 259 587
rect 213 537 219 571
rect 253 537 259 571
rect 213 497 259 537
rect 213 463 219 497
rect 253 463 259 497
rect 213 424 259 463
rect 293 584 359 649
rect 293 550 309 584
rect 343 550 359 584
rect 293 492 359 550
rect 293 458 309 492
rect 343 458 359 492
rect 393 574 439 590
rect 393 540 399 574
rect 433 540 439 574
rect 393 490 439 540
rect 393 456 399 490
rect 433 456 439 490
rect 473 584 539 649
rect 473 550 489 584
rect 523 550 539 584
rect 473 498 539 550
rect 473 464 489 498
rect 523 464 539 498
rect 573 580 639 596
rect 573 546 589 580
rect 623 546 639 580
rect 573 505 639 546
rect 573 471 589 505
rect 623 471 639 505
rect 393 430 439 456
rect 573 430 639 471
rect 673 584 739 649
rect 673 550 689 584
rect 723 550 739 584
rect 673 492 739 550
rect 673 458 689 492
rect 723 458 739 492
rect 773 580 839 596
rect 773 546 789 580
rect 823 546 839 580
rect 773 505 839 546
rect 873 570 939 649
rect 873 536 889 570
rect 923 536 939 570
rect 873 526 939 536
rect 973 570 1135 586
rect 973 536 980 570
rect 1014 536 1085 570
rect 1119 536 1135 570
rect 773 471 789 505
rect 823 492 839 505
rect 973 492 1135 536
rect 1169 570 1235 649
rect 1169 536 1185 570
rect 1219 536 1235 570
rect 1169 526 1235 536
rect 1269 584 1705 615
rect 1269 550 1285 584
rect 1319 581 1705 584
rect 1319 550 1335 581
rect 1269 492 1335 550
rect 1475 580 1515 581
rect 823 471 980 492
rect 773 458 980 471
rect 1014 458 1085 492
rect 1119 458 1285 492
rect 1319 458 1335 492
rect 1369 542 1435 547
rect 1369 508 1385 542
rect 1419 508 1435 542
rect 393 424 639 430
rect 773 424 839 458
rect 1369 430 1435 508
rect 1509 546 1515 580
rect 1651 580 1705 581
rect 1475 508 1515 546
rect 1509 474 1515 508
rect 1475 458 1515 474
rect 1549 542 1615 547
rect 1549 508 1565 542
rect 1599 508 1615 542
rect 1369 424 1385 430
rect 23 390 39 424
rect 73 390 219 424
rect 253 410 589 424
rect 253 390 399 410
rect 383 376 399 390
rect 433 390 589 410
rect 623 390 789 424
rect 823 390 839 424
rect 889 396 1385 424
rect 1419 424 1435 430
rect 1549 430 1615 508
rect 1549 424 1565 430
rect 1419 396 1565 424
rect 1599 396 1615 430
rect 889 390 1615 396
rect 1651 546 1655 580
rect 1689 546 1705 580
rect 1651 512 1705 546
rect 1651 478 1655 512
rect 1689 478 1705 512
rect 1651 440 1705 478
rect 1651 406 1655 440
rect 1689 406 1705 440
rect 1651 390 1705 406
rect 433 376 449 390
rect 383 364 449 376
rect 25 320 349 356
rect 25 286 103 320
rect 137 286 171 320
rect 205 286 239 320
rect 273 286 307 320
rect 341 286 349 320
rect 25 270 349 286
rect 483 320 839 356
rect 483 286 491 320
rect 525 286 559 320
rect 593 286 627 320
rect 661 286 695 320
rect 729 286 839 320
rect 483 270 839 286
rect 889 236 938 390
rect 985 320 1223 356
rect 985 286 1021 320
rect 1055 286 1089 320
rect 1123 286 1157 320
rect 1191 286 1223 320
rect 985 270 1223 286
rect 1273 320 1703 356
rect 1273 286 1351 320
rect 1385 286 1419 320
rect 1453 286 1487 320
rect 1521 286 1703 320
rect 1273 270 1703 286
rect 26 214 824 236
rect 889 226 1705 236
rect 26 210 400 214
rect 26 176 42 210
rect 76 202 214 210
rect 26 120 76 176
rect 248 202 400 210
rect 26 86 42 120
rect 26 70 76 86
rect 112 152 178 168
rect 112 118 128 152
rect 162 118 178 152
rect 112 17 178 118
rect 214 120 248 176
rect 384 180 400 202
rect 434 202 824 214
rect 214 70 248 86
rect 284 152 350 168
rect 284 118 300 152
rect 334 118 350 152
rect 284 17 350 118
rect 384 116 434 180
rect 565 169 624 202
rect 384 82 400 116
rect 384 66 434 82
rect 470 152 531 168
rect 470 118 487 152
rect 521 118 531 152
rect 565 135 574 169
rect 608 135 624 169
rect 758 169 824 202
rect 565 119 624 135
rect 658 152 724 168
rect 470 85 531 118
rect 658 118 674 152
rect 708 118 724 152
rect 758 135 774 169
rect 808 135 824 169
rect 870 210 1705 226
rect 870 176 887 210
rect 921 202 1318 210
rect 921 193 1168 202
rect 921 176 937 193
rect 870 154 937 176
rect 1102 169 1168 193
rect 758 119 824 135
rect 987 143 1053 159
rect 658 85 724 118
rect 987 109 1003 143
rect 1037 109 1053 143
rect 1102 135 1118 169
rect 1152 135 1168 169
rect 1302 176 1318 202
rect 1352 202 1655 210
rect 1352 176 1368 202
rect 1102 119 1168 135
rect 1202 152 1268 168
rect 987 85 1053 109
rect 1202 118 1218 152
rect 1252 118 1268 152
rect 1202 85 1268 118
rect 470 51 1268 85
rect 1302 120 1368 176
rect 1639 176 1655 202
rect 1689 176 1705 210
rect 1302 86 1318 120
rect 1352 86 1368 120
rect 1302 70 1368 86
rect 1402 152 1605 168
rect 1402 118 1404 152
rect 1438 118 1486 152
rect 1520 118 1569 152
rect 1603 118 1605 152
rect 1402 17 1605 118
rect 1639 120 1705 176
rect 1639 86 1655 120
rect 1689 86 1705 120
rect 1639 70 1705 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a31oi_4
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 1782000
string GDS_START 1767940
<< end >>
