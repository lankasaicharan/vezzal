magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 66 49 1085 241
rect 0 0 1152 49
<< scnmos >>
rect 145 47 175 215
rect 257 47 287 215
rect 329 47 359 215
rect 478 47 508 215
rect 550 47 580 215
rect 718 47 748 215
rect 804 47 834 215
rect 890 47 920 215
rect 976 47 1006 215
<< scpmoshvt >>
rect 94 367 124 619
rect 180 367 210 619
rect 370 367 400 619
rect 456 367 486 619
rect 646 367 676 619
rect 732 367 762 619
rect 818 367 848 619
rect 904 367 934 619
rect 990 367 1020 619
<< ndiff >>
rect 92 203 145 215
rect 92 169 100 203
rect 134 169 145 203
rect 92 101 145 169
rect 92 67 100 101
rect 134 67 145 101
rect 92 47 145 67
rect 175 163 257 215
rect 175 129 199 163
rect 233 129 257 163
rect 175 89 257 129
rect 175 55 199 89
rect 233 55 257 89
rect 175 47 257 55
rect 287 47 329 215
rect 359 198 478 215
rect 359 164 433 198
rect 467 164 478 198
rect 359 89 478 164
rect 359 55 433 89
rect 467 55 478 89
rect 359 47 478 55
rect 508 47 550 215
rect 580 122 718 215
rect 580 88 591 122
rect 625 88 673 122
rect 707 88 718 122
rect 580 47 718 88
rect 748 203 804 215
rect 748 169 759 203
rect 793 169 804 203
rect 748 101 804 169
rect 748 67 759 101
rect 793 67 804 101
rect 748 47 804 67
rect 834 179 890 215
rect 834 145 845 179
rect 879 145 890 179
rect 834 93 890 145
rect 834 59 845 93
rect 879 59 890 93
rect 834 47 890 59
rect 920 203 976 215
rect 920 169 931 203
rect 965 169 976 203
rect 920 101 976 169
rect 920 67 931 101
rect 965 67 976 101
rect 920 47 976 67
rect 1006 163 1059 215
rect 1006 129 1017 163
rect 1051 129 1059 163
rect 1006 93 1059 129
rect 1006 59 1017 93
rect 1051 59 1059 93
rect 1006 47 1059 59
<< pdiff >>
rect 41 599 94 619
rect 41 565 49 599
rect 83 565 94 599
rect 41 527 94 565
rect 41 493 49 527
rect 83 493 94 527
rect 41 457 94 493
rect 41 423 49 457
rect 83 423 94 457
rect 41 367 94 423
rect 124 607 180 619
rect 124 573 135 607
rect 169 573 180 607
rect 124 526 180 573
rect 124 492 135 526
rect 169 492 180 526
rect 124 441 180 492
rect 124 407 135 441
rect 169 407 180 441
rect 124 367 180 407
rect 210 597 263 619
rect 210 563 221 597
rect 255 563 263 597
rect 210 529 263 563
rect 210 495 221 529
rect 255 495 263 529
rect 210 461 263 495
rect 210 427 221 461
rect 255 427 263 461
rect 210 367 263 427
rect 317 531 370 619
rect 317 497 325 531
rect 359 497 370 531
rect 317 457 370 497
rect 317 423 325 457
rect 359 423 370 457
rect 317 367 370 423
rect 400 451 456 619
rect 400 417 411 451
rect 445 417 456 451
rect 400 367 456 417
rect 486 607 539 619
rect 486 573 497 607
rect 531 573 539 607
rect 486 367 539 573
rect 593 599 646 619
rect 593 565 601 599
rect 635 565 646 599
rect 593 527 646 565
rect 593 493 601 527
rect 635 493 646 527
rect 593 367 646 493
rect 676 607 732 619
rect 676 573 687 607
rect 721 573 732 607
rect 676 523 732 573
rect 676 489 687 523
rect 721 489 732 523
rect 676 367 732 489
rect 762 599 818 619
rect 762 565 773 599
rect 807 565 818 599
rect 762 504 818 565
rect 762 470 773 504
rect 807 470 818 504
rect 762 413 818 470
rect 762 379 773 413
rect 807 379 818 413
rect 762 367 818 379
rect 848 611 904 619
rect 848 577 859 611
rect 893 577 904 611
rect 848 532 904 577
rect 848 498 859 532
rect 893 498 904 532
rect 848 453 904 498
rect 848 419 859 453
rect 893 419 904 453
rect 848 367 904 419
rect 934 599 990 619
rect 934 565 945 599
rect 979 565 990 599
rect 934 504 990 565
rect 934 470 945 504
rect 979 470 990 504
rect 934 413 990 470
rect 934 379 945 413
rect 979 379 990 413
rect 934 367 990 379
rect 1020 607 1073 619
rect 1020 573 1031 607
rect 1065 573 1073 607
rect 1020 533 1073 573
rect 1020 499 1031 533
rect 1065 499 1073 533
rect 1020 453 1073 499
rect 1020 419 1031 453
rect 1065 419 1073 453
rect 1020 367 1073 419
<< ndiffc >>
rect 100 169 134 203
rect 100 67 134 101
rect 199 129 233 163
rect 199 55 233 89
rect 433 164 467 198
rect 433 55 467 89
rect 591 88 625 122
rect 673 88 707 122
rect 759 169 793 203
rect 759 67 793 101
rect 845 145 879 179
rect 845 59 879 93
rect 931 169 965 203
rect 931 67 965 101
rect 1017 129 1051 163
rect 1017 59 1051 93
<< pdiffc >>
rect 49 565 83 599
rect 49 493 83 527
rect 49 423 83 457
rect 135 573 169 607
rect 135 492 169 526
rect 135 407 169 441
rect 221 563 255 597
rect 221 495 255 529
rect 221 427 255 461
rect 325 497 359 531
rect 325 423 359 457
rect 411 417 445 451
rect 497 573 531 607
rect 601 565 635 599
rect 601 493 635 527
rect 687 573 721 607
rect 687 489 721 523
rect 773 565 807 599
rect 773 470 807 504
rect 773 379 807 413
rect 859 577 893 611
rect 859 498 893 532
rect 859 419 893 453
rect 945 565 979 599
rect 945 470 979 504
rect 945 379 979 413
rect 1031 573 1065 607
rect 1031 499 1065 533
rect 1031 419 1065 453
<< poly >>
rect 94 619 124 645
rect 180 619 210 645
rect 370 619 400 645
rect 456 619 486 645
rect 646 619 676 645
rect 732 619 762 645
rect 818 619 848 645
rect 904 619 934 645
rect 990 619 1020 645
rect 94 333 124 367
rect 180 345 210 367
rect 72 317 138 333
rect 72 283 88 317
rect 122 283 138 317
rect 180 315 287 345
rect 72 267 138 283
rect 217 303 287 315
rect 370 303 400 367
rect 456 303 486 367
rect 646 303 676 367
rect 732 333 762 367
rect 818 333 848 367
rect 904 333 934 367
rect 990 333 1020 367
rect 217 269 233 303
rect 267 269 287 303
rect 72 237 175 267
rect 217 253 287 269
rect 145 215 175 237
rect 257 215 287 253
rect 329 287 400 303
rect 329 253 345 287
rect 379 253 400 287
rect 329 237 400 253
rect 442 287 508 303
rect 442 253 458 287
rect 492 253 508 287
rect 442 237 508 253
rect 329 215 359 237
rect 478 215 508 237
rect 550 287 676 303
rect 550 253 597 287
rect 631 273 676 287
rect 718 317 1056 333
rect 718 283 734 317
rect 768 283 802 317
rect 836 283 870 317
rect 904 283 938 317
rect 972 283 1006 317
rect 1040 283 1056 317
rect 631 253 647 273
rect 550 237 647 253
rect 718 267 1056 283
rect 550 215 580 237
rect 718 215 748 267
rect 804 215 834 267
rect 890 215 920 267
rect 976 215 1006 267
rect 145 21 175 47
rect 257 21 287 47
rect 329 21 359 47
rect 478 21 508 47
rect 550 21 580 47
rect 718 21 748 47
rect 804 21 834 47
rect 890 21 920 47
rect 976 21 1006 47
<< polycont >>
rect 88 283 122 317
rect 233 269 267 303
rect 345 253 379 287
rect 458 253 492 287
rect 597 253 631 287
rect 734 283 768 317
rect 802 283 836 317
rect 870 283 904 317
rect 938 283 972 317
rect 1006 283 1040 317
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 18 599 85 615
rect 18 565 49 599
rect 83 565 85 599
rect 18 527 85 565
rect 18 493 49 527
rect 83 493 85 527
rect 18 457 85 493
rect 18 423 49 457
rect 83 423 85 457
rect 18 407 85 423
rect 119 607 185 649
rect 119 573 135 607
rect 169 573 185 607
rect 119 526 185 573
rect 119 492 135 526
rect 169 492 185 526
rect 119 441 185 492
rect 119 407 135 441
rect 169 407 185 441
rect 219 607 547 615
rect 219 597 497 607
rect 219 563 221 597
rect 255 581 497 597
rect 255 563 271 581
rect 481 573 497 581
rect 531 573 547 607
rect 481 569 547 573
rect 585 599 637 615
rect 219 529 271 563
rect 585 565 601 599
rect 635 565 637 599
rect 219 495 221 529
rect 255 495 271 529
rect 219 461 271 495
rect 219 427 221 461
rect 255 427 271 461
rect 219 407 271 427
rect 309 535 359 547
rect 585 535 637 565
rect 309 531 637 535
rect 309 497 325 531
rect 359 527 637 531
rect 359 501 601 527
rect 359 497 361 501
rect 309 457 361 497
rect 585 493 601 501
rect 635 493 637 527
rect 585 477 637 493
rect 671 607 737 649
rect 671 573 687 607
rect 721 573 737 607
rect 671 523 737 573
rect 671 489 687 523
rect 721 489 737 523
rect 771 599 809 615
rect 771 565 773 599
rect 807 565 809 599
rect 771 504 809 565
rect 771 470 773 504
rect 807 470 809 504
rect 309 423 325 457
rect 359 423 361 457
rect 309 407 361 423
rect 395 451 461 467
rect 395 417 411 451
rect 445 443 461 451
rect 445 417 730 443
rect 395 407 730 417
rect 18 231 52 407
rect 86 339 651 373
rect 86 317 138 339
rect 86 283 88 317
rect 122 283 138 317
rect 86 267 138 283
rect 217 303 283 305
rect 217 269 233 303
rect 267 269 283 303
rect 217 231 283 269
rect 18 203 283 231
rect 18 169 100 203
rect 134 197 283 203
rect 317 287 381 305
rect 317 253 345 287
rect 379 253 381 287
rect 134 169 140 197
rect 18 101 140 169
rect 18 67 100 101
rect 134 67 140 101
rect 18 51 140 67
rect 174 129 199 163
rect 233 129 266 163
rect 174 89 266 129
rect 174 55 199 89
rect 233 55 266 89
rect 317 69 381 253
rect 415 287 545 305
rect 415 253 458 287
rect 492 253 545 287
rect 415 240 545 253
rect 581 287 651 339
rect 581 253 597 287
rect 631 253 651 287
rect 581 240 651 253
rect 685 317 730 407
rect 771 413 809 470
rect 843 611 909 649
rect 843 577 859 611
rect 893 577 909 611
rect 843 532 909 577
rect 843 498 859 532
rect 893 498 909 532
rect 843 453 909 498
rect 843 419 859 453
rect 893 419 909 453
rect 943 599 979 615
rect 943 565 945 599
rect 943 504 979 565
rect 943 470 945 504
rect 771 379 773 413
rect 807 385 809 413
rect 943 413 979 470
rect 1015 607 1081 649
rect 1015 573 1031 607
rect 1065 573 1081 607
rect 1015 533 1081 573
rect 1015 499 1031 533
rect 1065 499 1081 533
rect 1015 453 1081 499
rect 1015 419 1031 453
rect 1065 419 1081 453
rect 943 385 945 413
rect 807 379 945 385
rect 979 379 1132 385
rect 771 351 1132 379
rect 685 283 734 317
rect 768 283 802 317
rect 836 283 870 317
rect 904 283 938 317
rect 972 283 1006 317
rect 1040 283 1056 317
rect 685 281 1056 283
rect 685 206 719 281
rect 1092 247 1132 351
rect 417 198 719 206
rect 417 164 433 198
rect 467 172 719 198
rect 753 213 1132 247
rect 753 203 795 213
rect 467 164 506 172
rect 417 89 506 164
rect 753 169 759 203
rect 793 169 795 203
rect 929 203 974 213
rect 174 17 266 55
rect 417 55 433 89
rect 467 55 506 89
rect 417 51 506 55
rect 575 122 719 138
rect 575 88 591 122
rect 625 88 673 122
rect 707 88 719 122
rect 575 17 719 88
rect 753 101 795 169
rect 753 67 759 101
rect 793 67 795 101
rect 753 51 795 67
rect 829 145 845 179
rect 879 145 895 179
rect 829 93 895 145
rect 829 59 845 93
rect 879 59 895 93
rect 829 17 895 59
rect 929 169 931 203
rect 965 169 974 203
rect 929 101 974 169
rect 929 67 931 101
rect 965 67 974 101
rect 929 51 974 67
rect 1008 163 1053 179
rect 1008 129 1017 163
rect 1051 129 1053 163
rect 1008 93 1053 129
rect 1008 59 1017 93
rect 1051 59 1053 93
rect 1087 78 1132 213
rect 1008 17 1053 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 1087 94 1121 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1718698
string GDS_START 1708816
<< end >>
