magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 44 49 616 211
rect 0 0 672 49
<< scnmos >>
rect 143 101 173 185
rect 229 101 259 185
rect 331 101 361 185
rect 503 101 533 185
<< scpmoshvt >>
rect 119 419 169 619
rect 217 419 267 619
rect 331 419 381 619
rect 503 419 553 619
<< ndiff >>
rect 70 157 143 185
rect 70 123 82 157
rect 116 123 143 157
rect 70 101 143 123
rect 173 173 229 185
rect 173 139 184 173
rect 218 139 229 173
rect 173 101 229 139
rect 259 160 331 185
rect 259 126 286 160
rect 320 126 331 160
rect 259 101 331 126
rect 361 151 503 185
rect 361 117 405 151
rect 439 117 503 151
rect 361 101 503 117
rect 533 151 590 185
rect 533 117 544 151
rect 578 117 590 151
rect 533 101 590 117
<< pdiff >>
rect 62 607 119 619
rect 62 573 74 607
rect 108 573 119 607
rect 62 512 119 573
rect 62 478 74 512
rect 108 478 119 512
rect 62 419 119 478
rect 169 419 217 619
rect 267 597 331 619
rect 267 563 278 597
rect 312 563 331 597
rect 267 497 331 563
rect 267 463 278 497
rect 312 463 331 497
rect 267 419 331 463
rect 381 419 503 619
rect 553 607 610 619
rect 553 573 564 607
rect 598 573 610 607
rect 553 497 610 573
rect 553 463 564 497
rect 598 463 610 497
rect 553 419 610 463
<< ndiffc >>
rect 82 123 116 157
rect 184 139 218 173
rect 286 126 320 160
rect 405 117 439 151
rect 544 117 578 151
<< pdiffc >>
rect 74 573 108 607
rect 74 478 108 512
rect 278 563 312 597
rect 278 463 312 497
rect 564 573 598 607
rect 564 463 598 497
<< poly >>
rect 119 619 169 645
rect 217 619 267 645
rect 331 619 381 645
rect 503 619 553 645
rect 119 356 169 419
rect 103 340 169 356
rect 103 306 119 340
rect 153 306 169 340
rect 103 290 169 306
rect 217 356 267 419
rect 217 340 283 356
rect 217 306 233 340
rect 267 306 283 340
rect 217 290 283 306
rect 331 341 381 419
rect 503 341 553 419
rect 331 325 455 341
rect 331 291 405 325
rect 439 291 455 325
rect 139 230 169 290
rect 139 200 173 230
rect 143 185 173 200
rect 229 185 259 290
rect 331 257 455 291
rect 331 223 405 257
rect 439 223 455 257
rect 331 207 455 223
rect 503 325 569 341
rect 503 291 519 325
rect 553 291 569 325
rect 503 257 569 291
rect 503 223 519 257
rect 553 223 569 257
rect 503 207 569 223
rect 331 185 361 207
rect 503 185 533 207
rect 143 75 173 101
rect 229 75 259 101
rect 331 75 361 101
rect 503 75 533 101
<< polycont >>
rect 119 306 153 340
rect 233 306 267 340
rect 405 291 439 325
rect 405 223 439 257
rect 519 291 553 325
rect 519 223 553 257
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 58 607 124 649
rect 58 573 74 607
rect 108 573 124 607
rect 58 512 124 573
rect 58 478 74 512
rect 108 478 124 512
rect 58 462 124 478
rect 217 597 328 613
rect 217 563 278 597
rect 312 563 328 597
rect 217 497 328 563
rect 217 463 278 497
rect 312 463 328 497
rect 217 447 328 463
rect 548 607 614 649
rect 548 573 564 607
rect 598 573 614 607
rect 548 497 614 573
rect 548 463 564 497
rect 598 463 614 497
rect 548 447 614 463
rect 217 426 263 447
rect 33 392 263 426
rect 33 254 67 392
rect 319 377 639 411
rect 103 340 169 356
rect 103 306 119 340
rect 153 306 169 340
rect 103 290 169 306
rect 217 340 283 356
rect 217 306 233 340
rect 267 306 283 340
rect 217 290 283 306
rect 33 220 234 254
rect 66 157 132 184
rect 66 123 82 157
rect 116 123 132 157
rect 168 173 234 220
rect 319 189 353 377
rect 389 325 455 341
rect 389 291 405 325
rect 439 291 455 325
rect 389 257 455 291
rect 389 223 405 257
rect 439 223 455 257
rect 389 207 455 223
rect 503 325 569 341
rect 503 291 519 325
rect 553 291 569 325
rect 503 257 569 291
rect 503 223 519 257
rect 553 223 569 257
rect 503 207 569 223
rect 168 139 184 173
rect 218 139 234 173
rect 168 123 234 139
rect 270 160 353 189
rect 605 171 639 377
rect 270 126 286 160
rect 320 126 353 160
rect 66 87 132 123
rect 270 87 353 126
rect 66 53 353 87
rect 389 151 455 171
rect 389 117 405 151
rect 439 117 455 151
rect 389 17 455 117
rect 528 151 639 171
rect 528 117 544 151
rect 578 117 639 151
rect 528 97 639 117
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o22ai_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1316630
string GDS_START 1311188
<< end >>
