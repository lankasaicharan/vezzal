magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
<< pwell >>
rect 771 229 975 273
rect 1487 229 2102 247
rect 225 180 2102 229
rect 1 49 2102 180
rect 0 0 2112 49
<< scnmos >>
rect 80 70 110 154
rect 304 119 334 203
rect 399 119 429 203
rect 507 119 537 203
rect 598 119 628 203
rect 670 119 700 203
rect 866 119 896 247
rect 971 119 1001 203
rect 1095 119 1125 203
rect 1169 119 1199 203
rect 1307 75 1337 203
rect 1570 137 1600 221
rect 1703 53 1733 221
rect 1789 53 1819 221
rect 1907 53 1937 221
rect 1993 53 2023 221
<< scpmoshvt >>
rect 80 458 110 586
rect 289 463 319 591
rect 429 463 459 547
rect 515 463 545 547
rect 639 499 669 583
rect 741 463 771 547
rect 866 369 896 537
rect 952 369 982 537
rect 1127 453 1157 537
rect 1229 451 1259 535
rect 1343 451 1373 619
rect 1570 367 1600 495
rect 1703 367 1733 619
rect 1789 367 1819 619
rect 1906 367 1936 619
rect 1992 367 2022 619
<< ndiff >>
rect 797 203 866 247
rect 251 178 304 203
rect 27 128 80 154
rect 27 94 35 128
rect 69 94 80 128
rect 27 70 80 94
rect 110 128 163 154
rect 110 94 121 128
rect 155 94 163 128
rect 251 144 259 178
rect 293 144 304 178
rect 251 119 304 144
rect 334 178 399 203
rect 334 144 345 178
rect 379 144 399 178
rect 334 119 399 144
rect 429 178 507 203
rect 429 144 452 178
rect 486 144 507 178
rect 429 119 507 144
rect 537 178 598 203
rect 537 144 553 178
rect 587 144 598 178
rect 537 119 598 144
rect 628 119 670 203
rect 700 165 866 203
rect 700 131 711 165
rect 745 131 821 165
rect 855 131 866 165
rect 700 119 866 131
rect 896 235 949 247
rect 896 201 907 235
rect 941 203 949 235
rect 1513 213 1570 221
rect 941 201 971 203
rect 896 167 971 201
rect 896 133 907 167
rect 941 133 971 167
rect 896 119 971 133
rect 1001 178 1095 203
rect 1001 144 1031 178
rect 1065 144 1095 178
rect 1001 119 1095 144
rect 1125 119 1169 203
rect 1199 189 1307 203
rect 1199 155 1210 189
rect 1244 155 1307 189
rect 1199 121 1307 155
rect 1199 119 1262 121
rect 110 70 163 94
rect 1238 87 1262 119
rect 1296 87 1307 121
rect 1238 75 1307 87
rect 1337 189 1390 203
rect 1337 155 1348 189
rect 1382 155 1390 189
rect 1337 121 1390 155
rect 1513 179 1525 213
rect 1559 179 1570 213
rect 1513 137 1570 179
rect 1600 137 1703 221
rect 1337 87 1348 121
rect 1382 87 1390 121
rect 1337 75 1390 87
rect 1623 73 1703 137
rect 1623 39 1635 73
rect 1669 53 1703 73
rect 1733 213 1789 221
rect 1733 179 1744 213
rect 1778 179 1789 213
rect 1733 53 1789 179
rect 1819 73 1907 221
rect 1819 53 1846 73
rect 1669 39 1681 53
rect 1623 31 1681 39
rect 1834 39 1846 53
rect 1880 53 1907 73
rect 1937 212 1993 221
rect 1937 178 1948 212
rect 1982 178 1993 212
rect 1937 101 1993 178
rect 1937 67 1948 101
rect 1982 67 1993 101
rect 1937 53 1993 67
rect 2023 209 2076 221
rect 2023 175 2034 209
rect 2068 175 2076 209
rect 2023 99 2076 175
rect 2023 65 2034 99
rect 2068 65 2076 99
rect 2023 53 2076 65
rect 1880 39 1892 53
rect 1834 31 1892 39
<< pdiff >>
rect 27 574 80 586
rect 27 540 35 574
rect 69 540 80 574
rect 27 506 80 540
rect 27 472 35 506
rect 69 472 80 506
rect 27 458 80 472
rect 110 574 163 586
rect 110 540 121 574
rect 155 540 163 574
rect 110 506 163 540
rect 110 472 121 506
rect 155 472 163 506
rect 110 458 163 472
rect 236 577 289 591
rect 236 543 244 577
rect 278 543 289 577
rect 236 509 289 543
rect 236 475 244 509
rect 278 475 289 509
rect 236 463 289 475
rect 319 578 376 591
rect 319 544 330 578
rect 364 547 376 578
rect 567 547 639 583
rect 364 544 429 547
rect 319 463 429 544
rect 459 510 515 547
rect 459 476 470 510
rect 504 476 515 510
rect 459 463 515 476
rect 545 531 639 547
rect 545 497 575 531
rect 609 499 639 531
rect 669 547 719 583
rect 793 551 851 559
rect 793 547 805 551
rect 669 499 741 547
rect 609 497 617 499
rect 545 463 617 497
rect 691 463 741 499
rect 771 517 805 547
rect 839 537 851 551
rect 1290 607 1343 619
rect 1290 573 1298 607
rect 1332 573 1343 607
rect 839 517 866 537
rect 771 463 866 517
rect 793 369 866 463
rect 896 411 952 537
rect 896 377 907 411
rect 941 377 952 411
rect 896 369 952 377
rect 982 525 1127 537
rect 982 491 1063 525
rect 1097 491 1127 525
rect 982 453 1127 491
rect 1157 535 1207 537
rect 1290 535 1343 573
rect 1157 453 1229 535
rect 982 415 1105 453
rect 982 381 1063 415
rect 1097 381 1105 415
rect 982 369 1105 381
rect 1179 451 1229 453
rect 1259 508 1343 535
rect 1259 474 1270 508
rect 1304 474 1343 508
rect 1259 451 1343 474
rect 1373 599 1426 619
rect 1373 565 1384 599
rect 1418 565 1426 599
rect 1373 497 1426 565
rect 1642 611 1703 619
rect 1642 577 1654 611
rect 1688 577 1703 611
rect 1373 463 1384 497
rect 1418 463 1426 497
rect 1642 496 1703 577
rect 1642 495 1658 496
rect 1373 451 1426 463
rect 1517 481 1570 495
rect 1517 447 1525 481
rect 1559 447 1570 481
rect 1517 413 1570 447
rect 1517 379 1525 413
rect 1559 379 1570 413
rect 1517 367 1570 379
rect 1600 462 1658 495
rect 1692 462 1703 496
rect 1600 413 1703 462
rect 1600 379 1611 413
rect 1645 379 1703 413
rect 1600 367 1703 379
rect 1733 599 1789 619
rect 1733 565 1744 599
rect 1778 565 1789 599
rect 1733 494 1789 565
rect 1733 460 1744 494
rect 1778 460 1789 494
rect 1733 409 1789 460
rect 1733 375 1744 409
rect 1778 375 1789 409
rect 1733 367 1789 375
rect 1819 611 1906 619
rect 1819 577 1846 611
rect 1880 577 1906 611
rect 1819 511 1906 577
rect 1819 477 1846 511
rect 1880 477 1906 511
rect 1819 414 1906 477
rect 1819 380 1846 414
rect 1880 380 1906 414
rect 1819 367 1906 380
rect 1936 599 1992 619
rect 1936 565 1947 599
rect 1981 565 1992 599
rect 1936 497 1992 565
rect 1936 463 1947 497
rect 1981 463 1992 497
rect 1936 409 1992 463
rect 1936 375 1947 409
rect 1981 375 1992 409
rect 1936 367 1992 375
rect 2022 607 2075 619
rect 2022 573 2033 607
rect 2067 573 2075 607
rect 2022 508 2075 573
rect 2022 474 2033 508
rect 2067 474 2075 508
rect 2022 413 2075 474
rect 2022 379 2033 413
rect 2067 379 2075 413
rect 2022 367 2075 379
<< ndiffc >>
rect 35 94 69 128
rect 121 94 155 128
rect 259 144 293 178
rect 345 144 379 178
rect 452 144 486 178
rect 553 144 587 178
rect 711 131 745 165
rect 821 131 855 165
rect 907 201 941 235
rect 907 133 941 167
rect 1031 144 1065 178
rect 1210 155 1244 189
rect 1262 87 1296 121
rect 1348 155 1382 189
rect 1525 179 1559 213
rect 1348 87 1382 121
rect 1635 39 1669 73
rect 1744 179 1778 213
rect 1846 39 1880 73
rect 1948 178 1982 212
rect 1948 67 1982 101
rect 2034 175 2068 209
rect 2034 65 2068 99
<< pdiffc >>
rect 35 540 69 574
rect 35 472 69 506
rect 121 540 155 574
rect 121 472 155 506
rect 244 543 278 577
rect 244 475 278 509
rect 330 544 364 578
rect 470 476 504 510
rect 575 497 609 531
rect 805 517 839 551
rect 1298 573 1332 607
rect 907 377 941 411
rect 1063 491 1097 525
rect 1063 381 1097 415
rect 1270 474 1304 508
rect 1384 565 1418 599
rect 1654 577 1688 611
rect 1384 463 1418 497
rect 1525 447 1559 481
rect 1525 379 1559 413
rect 1658 462 1692 496
rect 1611 379 1645 413
rect 1744 565 1778 599
rect 1744 460 1778 494
rect 1744 375 1778 409
rect 1846 577 1880 611
rect 1846 477 1880 511
rect 1846 380 1880 414
rect 1947 565 1981 599
rect 1947 463 1981 497
rect 1947 375 1981 409
rect 2033 573 2067 607
rect 2033 474 2067 508
rect 2033 379 2067 413
<< poly >>
rect 289 615 982 645
rect 1343 619 1373 645
rect 1703 619 1733 645
rect 1789 619 1819 645
rect 1906 619 1936 645
rect 1992 619 2022 645
rect 80 586 110 612
rect 289 591 319 615
rect 639 583 669 615
rect 429 547 459 573
rect 515 547 545 573
rect 741 547 771 573
rect 639 473 669 499
rect 866 537 896 563
rect 952 537 982 615
rect 1127 537 1157 563
rect 80 310 110 458
rect 44 294 110 310
rect 44 260 60 294
rect 94 260 110 294
rect 158 404 224 420
rect 158 370 174 404
rect 208 370 224 404
rect 158 336 224 370
rect 158 302 174 336
rect 208 316 224 336
rect 289 316 319 463
rect 429 359 459 463
rect 515 431 545 463
rect 515 415 691 431
rect 741 415 771 463
rect 515 401 641 415
rect 598 381 641 401
rect 675 381 691 415
rect 598 365 691 381
rect 733 385 771 415
rect 399 343 465 359
rect 208 302 334 316
rect 158 286 334 302
rect 44 226 110 260
rect 44 192 60 226
rect 94 192 110 226
rect 304 203 334 286
rect 399 309 415 343
rect 449 309 465 343
rect 399 275 465 309
rect 399 241 415 275
rect 449 241 465 275
rect 399 225 465 241
rect 399 203 429 225
rect 507 203 537 229
rect 598 203 628 365
rect 733 291 763 385
rect 1229 535 1259 561
rect 866 337 896 369
rect 952 343 982 369
rect 670 275 763 291
rect 670 241 713 275
rect 747 241 763 275
rect 805 321 896 337
rect 1127 333 1157 453
rect 1570 495 1600 521
rect 1229 419 1259 451
rect 805 287 821 321
rect 855 287 896 321
rect 1097 303 1157 333
rect 1199 403 1265 419
rect 1199 369 1215 403
rect 1249 369 1265 403
rect 1199 335 1265 369
rect 1343 363 1373 451
rect 1097 301 1127 303
rect 805 271 896 287
rect 866 247 896 271
rect 971 285 1127 301
rect 971 251 993 285
rect 1027 271 1127 285
rect 1199 301 1215 335
rect 1249 301 1265 335
rect 1199 285 1265 301
rect 1307 347 1373 363
rect 1307 313 1323 347
rect 1357 313 1373 347
rect 1027 251 1043 271
rect 1199 255 1229 285
rect 670 225 763 241
rect 670 203 700 225
rect 44 176 110 192
rect 80 154 110 176
rect 971 235 1043 251
rect 971 203 1001 235
rect 1095 203 1125 229
rect 1169 225 1229 255
rect 1307 279 1373 313
rect 1570 303 1600 367
rect 1703 309 1733 367
rect 1789 309 1819 367
rect 1906 330 1936 367
rect 1992 330 2022 367
rect 1307 245 1323 279
rect 1357 245 1373 279
rect 1307 229 1373 245
rect 1421 287 1600 303
rect 1421 253 1437 287
rect 1471 273 1600 287
rect 1471 253 1487 273
rect 1421 237 1487 253
rect 1169 203 1199 225
rect 1307 203 1337 229
rect 1570 221 1600 273
rect 1642 293 1819 309
rect 1642 259 1658 293
rect 1692 259 1819 293
rect 1861 314 2023 330
rect 1861 280 1877 314
rect 1911 280 2023 314
rect 1861 264 2023 280
rect 1642 243 1819 259
rect 1703 221 1733 243
rect 1789 221 1819 243
rect 1907 221 1937 264
rect 1993 221 2023 264
rect 80 44 110 70
rect 304 51 334 119
rect 399 93 429 119
rect 507 51 537 119
rect 598 93 628 119
rect 670 93 700 119
rect 866 93 896 119
rect 971 93 1001 119
rect 1095 51 1125 119
rect 1169 93 1199 119
rect 1570 111 1600 137
rect 304 21 1125 51
rect 1307 49 1337 75
rect 1703 27 1733 53
rect 1789 27 1819 53
rect 1907 27 1937 53
rect 1993 27 2023 53
<< polycont >>
rect 60 260 94 294
rect 174 370 208 404
rect 174 302 208 336
rect 641 381 675 415
rect 60 192 94 226
rect 415 309 449 343
rect 415 241 449 275
rect 713 241 747 275
rect 821 287 855 321
rect 1215 369 1249 403
rect 993 251 1027 285
rect 1215 301 1249 335
rect 1323 313 1357 347
rect 1323 245 1357 279
rect 1437 253 1471 287
rect 1658 259 1692 293
rect 1877 280 1911 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 19 574 81 649
rect 19 540 35 574
rect 69 540 81 574
rect 19 506 81 540
rect 19 472 35 506
rect 69 472 81 506
rect 19 456 81 472
rect 115 574 171 590
rect 115 540 121 574
rect 155 540 171 574
rect 115 506 171 540
rect 115 472 121 506
rect 155 472 171 506
rect 115 420 171 472
rect 228 577 282 593
rect 228 543 244 577
rect 278 543 282 577
rect 228 509 282 543
rect 316 578 366 649
rect 316 544 330 578
rect 364 544 366 578
rect 316 528 366 544
rect 400 581 695 615
rect 228 475 244 509
rect 278 494 282 509
rect 400 494 434 581
rect 553 531 625 547
rect 278 475 434 494
rect 228 460 434 475
rect 470 510 519 526
rect 504 476 519 510
rect 470 460 519 476
rect 228 459 295 460
rect 115 404 208 420
rect 115 386 174 404
rect 158 370 174 386
rect 18 294 94 359
rect 18 260 60 294
rect 18 226 94 260
rect 18 192 60 226
rect 18 168 94 192
rect 158 336 208 370
rect 158 302 174 336
rect 158 144 208 302
rect 19 128 85 134
rect 19 94 35 128
rect 69 94 85 128
rect 19 17 85 94
rect 119 128 208 144
rect 243 178 295 459
rect 399 343 451 424
rect 399 309 415 343
rect 449 309 451 343
rect 399 275 451 309
rect 399 241 415 275
rect 449 241 451 275
rect 399 225 451 241
rect 485 191 519 460
rect 243 144 259 178
rect 293 144 295 178
rect 243 128 295 144
rect 329 178 395 191
rect 329 144 345 178
rect 379 144 395 178
rect 119 94 121 128
rect 155 94 208 128
rect 119 66 208 94
rect 329 17 395 144
rect 436 178 519 191
rect 436 144 452 178
rect 486 144 519 178
rect 436 125 519 144
rect 553 497 575 531
rect 609 497 625 531
rect 553 481 625 497
rect 661 481 695 581
rect 789 551 855 649
rect 789 517 805 551
rect 839 517 855 551
rect 1254 607 1346 649
rect 1254 573 1298 607
rect 1332 573 1346 607
rect 789 515 855 517
rect 1063 525 1113 541
rect 1097 491 1113 525
rect 553 345 589 481
rect 661 447 1029 481
rect 661 431 695 447
rect 625 415 695 431
rect 625 381 641 415
rect 675 381 695 415
rect 625 379 695 381
rect 891 411 957 413
rect 891 377 907 411
rect 941 377 957 411
rect 553 321 857 345
rect 553 311 821 321
rect 553 178 603 311
rect 805 287 821 311
rect 855 287 857 321
rect 697 275 763 277
rect 697 241 713 275
rect 747 241 763 275
rect 805 271 857 287
rect 697 235 763 241
rect 891 235 957 377
rect 991 285 1029 447
rect 991 251 993 285
rect 1027 251 1029 285
rect 991 235 1029 251
rect 1063 415 1113 491
rect 1254 508 1346 573
rect 1254 474 1270 508
rect 1304 474 1346 508
rect 1254 467 1346 474
rect 1380 599 1434 615
rect 1380 565 1384 599
rect 1418 565 1434 599
rect 1380 497 1434 565
rect 1609 611 1694 649
rect 1609 577 1654 611
rect 1688 577 1694 611
rect 1380 463 1384 497
rect 1418 463 1434 497
rect 1380 433 1434 463
rect 1097 381 1113 415
rect 1063 263 1113 381
rect 1199 403 1434 433
rect 1199 369 1215 403
rect 1249 397 1434 403
rect 1249 369 1265 397
rect 1199 335 1265 369
rect 1199 301 1215 335
rect 1249 301 1265 335
rect 1307 347 1359 363
rect 1307 313 1323 347
rect 1357 313 1359 347
rect 1307 279 1359 313
rect 1307 263 1323 279
rect 1063 245 1323 263
rect 1357 245 1359 279
rect 697 201 907 235
rect 941 201 957 235
rect 587 144 603 178
rect 905 167 957 201
rect 1063 229 1359 245
rect 1393 303 1434 397
rect 1509 481 1575 497
rect 1509 447 1525 481
rect 1559 447 1575 481
rect 1509 413 1575 447
rect 1509 379 1525 413
rect 1559 379 1575 413
rect 1509 366 1575 379
rect 1609 496 1694 577
rect 1609 462 1658 496
rect 1692 462 1694 496
rect 1609 413 1694 462
rect 1609 379 1611 413
rect 1645 379 1694 413
rect 1509 363 1563 366
rect 1609 363 1694 379
rect 1728 599 1794 615
rect 1728 565 1744 599
rect 1778 565 1794 599
rect 1728 494 1794 565
rect 1728 460 1744 494
rect 1778 460 1794 494
rect 1728 409 1794 460
rect 1728 375 1744 409
rect 1778 375 1794 409
rect 1521 325 1563 363
rect 1393 287 1487 303
rect 1393 253 1437 287
rect 1471 253 1487 287
rect 1393 251 1487 253
rect 1521 293 1694 325
rect 1521 259 1658 293
rect 1692 259 1694 293
rect 1063 195 1113 229
rect 1393 195 1427 251
rect 1521 217 1694 259
rect 553 128 603 144
rect 695 165 871 167
rect 695 131 711 165
rect 745 131 821 165
rect 855 131 871 165
rect 695 17 871 131
rect 905 133 907 167
rect 941 133 957 167
rect 905 117 957 133
rect 1015 178 1113 195
rect 1015 144 1031 178
rect 1065 144 1113 178
rect 1015 128 1113 144
rect 1194 189 1298 195
rect 1194 155 1210 189
rect 1244 155 1298 189
rect 1194 121 1298 155
rect 1194 87 1262 121
rect 1296 87 1298 121
rect 1194 17 1298 87
rect 1332 189 1427 195
rect 1332 155 1348 189
rect 1382 155 1427 189
rect 1509 213 1694 217
rect 1509 179 1525 213
rect 1559 179 1694 213
rect 1728 213 1794 375
rect 1830 611 1896 649
rect 1830 577 1846 611
rect 1880 577 1896 611
rect 1830 511 1896 577
rect 1830 477 1846 511
rect 1880 477 1896 511
rect 1830 414 1896 477
rect 1830 380 1846 414
rect 1880 380 1896 414
rect 1830 364 1896 380
rect 1947 599 1991 615
rect 1981 565 1991 599
rect 1947 497 1991 565
rect 1981 463 1991 497
rect 1947 409 1991 463
rect 1981 375 1991 409
rect 1728 179 1744 213
rect 1778 179 1794 213
rect 1728 177 1794 179
rect 1874 314 1911 330
rect 1874 280 1877 314
rect 1874 264 1911 280
rect 1332 143 1427 155
rect 1874 143 1908 264
rect 1947 228 1991 375
rect 2025 607 2083 649
rect 2025 573 2033 607
rect 2067 573 2083 607
rect 2025 508 2083 573
rect 2025 474 2033 508
rect 2067 474 2083 508
rect 2025 413 2083 474
rect 2025 379 2033 413
rect 2067 379 2083 413
rect 2025 363 2083 379
rect 1332 121 1908 143
rect 1332 87 1348 121
rect 1382 109 1908 121
rect 1944 212 1991 228
rect 1944 178 1948 212
rect 1982 178 1991 212
rect 1382 87 1427 109
rect 1332 71 1427 87
rect 1944 101 1991 178
rect 1619 73 1685 75
rect 1619 39 1635 73
rect 1669 39 1685 73
rect 1619 17 1685 39
rect 1830 73 1896 75
rect 1830 39 1846 73
rect 1880 39 1896 73
rect 1944 67 1948 101
rect 1982 67 1991 101
rect 1944 51 1991 67
rect 2025 209 2084 225
rect 2025 175 2034 209
rect 2068 175 2084 209
rect 2025 99 2084 175
rect 2025 65 2034 99
rect 2068 65 2084 99
rect 1830 17 1896 39
rect 2025 17 2084 65
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfxbp_2
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1759 316 1793 350 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1759 390 1793 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1759 464 1793 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1759 538 1793 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 94 1985 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1951 168 1985 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1951 390 1985 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1951 464 1985 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1951 538 1985 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2394996
string GDS_START 2378954
<< end >>
