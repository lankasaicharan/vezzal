magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
rect 780 319 1060 331
<< pwell >>
rect 1347 257 1535 273
rect 1052 241 1535 257
rect 20 157 294 172
rect 822 157 1535 241
rect 20 49 1535 157
rect 0 0 1536 49
<< scnmos >>
rect 99 62 129 146
rect 185 62 215 146
rect 434 47 464 131
rect 538 47 568 131
rect 610 47 640 131
rect 718 47 748 131
rect 790 47 820 131
rect 901 47 931 215
rect 1131 63 1161 231
rect 1236 147 1266 231
rect 1426 79 1456 247
<< scpmoshvt >>
rect 113 419 143 547
rect 199 419 229 547
rect 420 491 450 619
rect 506 491 536 619
rect 578 491 608 619
rect 683 491 713 575
rect 758 491 788 575
rect 941 355 971 607
rect 1131 367 1161 619
rect 1236 367 1266 495
rect 1426 367 1456 619
<< ndiff >>
rect 46 118 99 146
rect 46 84 54 118
rect 88 84 99 118
rect 46 62 99 84
rect 129 118 185 146
rect 129 84 140 118
rect 174 84 185 118
rect 129 62 185 84
rect 215 123 268 146
rect 215 89 226 123
rect 260 89 268 123
rect 215 62 268 89
rect 1373 235 1426 247
rect 848 161 901 215
rect 848 131 856 161
rect 381 106 434 131
rect 381 72 389 106
rect 423 72 434 106
rect 381 47 434 72
rect 464 99 538 131
rect 464 65 484 99
rect 518 65 538 99
rect 464 47 538 65
rect 568 47 610 131
rect 640 99 718 131
rect 640 65 661 99
rect 695 65 718 99
rect 640 47 718 65
rect 748 47 790 131
rect 820 127 856 131
rect 890 127 901 161
rect 820 93 901 127
rect 820 59 831 93
rect 865 59 901 93
rect 820 47 901 59
rect 931 185 988 215
rect 931 151 946 185
rect 980 151 988 185
rect 931 101 988 151
rect 931 67 946 101
rect 980 67 988 101
rect 931 47 988 67
rect 1078 203 1131 231
rect 1078 169 1086 203
rect 1120 169 1131 203
rect 1078 118 1131 169
rect 1078 84 1086 118
rect 1120 84 1131 118
rect 1078 63 1131 84
rect 1161 218 1236 231
rect 1161 184 1180 218
rect 1214 184 1236 218
rect 1161 147 1236 184
rect 1266 208 1319 231
rect 1266 174 1277 208
rect 1311 174 1319 208
rect 1266 147 1319 174
rect 1373 201 1381 235
rect 1415 201 1426 235
rect 1161 109 1214 147
rect 1373 125 1426 201
rect 1161 75 1172 109
rect 1206 75 1214 109
rect 1373 91 1381 125
rect 1415 91 1426 125
rect 1373 79 1426 91
rect 1456 235 1509 247
rect 1456 201 1467 235
rect 1501 201 1509 235
rect 1456 125 1509 201
rect 1456 91 1467 125
rect 1501 91 1509 125
rect 1456 79 1509 91
rect 1161 63 1214 75
<< pdiff >>
rect 367 605 420 619
rect 367 571 375 605
rect 409 571 420 605
rect 60 535 113 547
rect 60 501 68 535
rect 102 501 113 535
rect 60 465 113 501
rect 60 431 68 465
rect 102 431 113 465
rect 60 419 113 431
rect 143 535 199 547
rect 143 501 154 535
rect 188 501 199 535
rect 143 465 199 501
rect 143 431 154 465
rect 188 431 199 465
rect 143 419 199 431
rect 229 535 282 547
rect 229 501 240 535
rect 274 501 282 535
rect 229 465 282 501
rect 367 537 420 571
rect 367 503 375 537
rect 409 503 420 537
rect 367 491 420 503
rect 450 603 506 619
rect 450 569 461 603
rect 495 569 506 603
rect 450 491 506 569
rect 536 491 578 619
rect 608 595 661 619
rect 608 561 619 595
rect 653 575 661 595
rect 888 595 941 607
rect 888 575 896 595
rect 653 561 683 575
rect 608 491 683 561
rect 713 491 758 575
rect 788 561 896 575
rect 930 561 941 595
rect 788 548 941 561
rect 788 514 805 548
rect 839 527 941 548
rect 839 514 896 527
rect 788 493 896 514
rect 930 493 941 527
rect 788 491 941 493
rect 229 431 240 465
rect 274 431 282 465
rect 229 419 282 431
rect 888 459 941 491
rect 888 425 896 459
rect 930 425 941 459
rect 888 355 941 425
rect 971 595 1024 607
rect 971 561 982 595
rect 1016 561 1024 595
rect 971 503 1024 561
rect 971 469 982 503
rect 1016 469 1024 503
rect 971 405 1024 469
rect 971 371 982 405
rect 1016 371 1024 405
rect 971 355 1024 371
rect 1078 599 1131 619
rect 1078 565 1086 599
rect 1120 565 1131 599
rect 1078 503 1131 565
rect 1078 469 1086 503
rect 1120 469 1131 503
rect 1078 413 1131 469
rect 1078 379 1086 413
rect 1120 379 1131 413
rect 1078 367 1131 379
rect 1161 607 1214 619
rect 1161 573 1172 607
rect 1206 573 1214 607
rect 1161 507 1214 573
rect 1373 607 1426 619
rect 1373 573 1381 607
rect 1415 573 1426 607
rect 1161 473 1172 507
rect 1206 495 1214 507
rect 1373 508 1426 573
rect 1206 473 1236 495
rect 1161 413 1236 473
rect 1161 379 1182 413
rect 1216 379 1236 413
rect 1161 367 1236 379
rect 1266 483 1319 495
rect 1266 449 1277 483
rect 1311 449 1319 483
rect 1266 413 1319 449
rect 1266 379 1277 413
rect 1311 379 1319 413
rect 1266 367 1319 379
rect 1373 474 1381 508
rect 1415 474 1426 508
rect 1373 413 1426 474
rect 1373 379 1381 413
rect 1415 379 1426 413
rect 1373 367 1426 379
rect 1456 599 1509 619
rect 1456 565 1467 599
rect 1501 565 1509 599
rect 1456 502 1509 565
rect 1456 468 1467 502
rect 1501 468 1509 502
rect 1456 413 1509 468
rect 1456 379 1467 413
rect 1501 379 1509 413
rect 1456 367 1509 379
<< ndiffc >>
rect 54 84 88 118
rect 140 84 174 118
rect 226 89 260 123
rect 389 72 423 106
rect 484 65 518 99
rect 661 65 695 99
rect 856 127 890 161
rect 831 59 865 93
rect 946 151 980 185
rect 946 67 980 101
rect 1086 169 1120 203
rect 1086 84 1120 118
rect 1180 184 1214 218
rect 1277 174 1311 208
rect 1381 201 1415 235
rect 1172 75 1206 109
rect 1381 91 1415 125
rect 1467 201 1501 235
rect 1467 91 1501 125
<< pdiffc >>
rect 375 571 409 605
rect 68 501 102 535
rect 68 431 102 465
rect 154 501 188 535
rect 154 431 188 465
rect 240 501 274 535
rect 375 503 409 537
rect 461 569 495 603
rect 619 561 653 595
rect 896 561 930 595
rect 805 514 839 548
rect 896 493 930 527
rect 240 431 274 465
rect 896 425 930 459
rect 982 561 1016 595
rect 982 469 1016 503
rect 982 371 1016 405
rect 1086 565 1120 599
rect 1086 469 1120 503
rect 1086 379 1120 413
rect 1172 573 1206 607
rect 1381 573 1415 607
rect 1172 473 1206 507
rect 1182 379 1216 413
rect 1277 449 1311 483
rect 1277 379 1311 413
rect 1381 474 1415 508
rect 1381 379 1415 413
rect 1467 565 1501 599
rect 1467 468 1501 502
rect 1467 379 1501 413
<< poly >>
rect 420 619 450 645
rect 506 619 536 645
rect 578 619 608 645
rect 113 547 143 573
rect 199 547 229 573
rect 941 607 971 633
rect 1131 619 1161 645
rect 1426 619 1456 645
rect 683 575 713 601
rect 758 575 788 601
rect 420 469 450 491
rect 398 439 450 469
rect 113 302 143 419
rect 77 286 143 302
rect 77 252 93 286
rect 127 252 143 286
rect 77 218 143 252
rect 77 184 93 218
rect 127 184 143 218
rect 199 202 229 419
rect 398 283 428 439
rect 506 397 536 491
rect 470 381 536 397
rect 470 347 486 381
rect 520 347 536 381
rect 470 331 536 347
rect 398 267 464 283
rect 398 233 414 267
rect 448 233 464 267
rect 398 217 464 233
rect 77 168 143 184
rect 185 186 356 202
rect 185 172 306 186
rect 99 146 129 168
rect 185 146 215 172
rect 290 152 306 172
rect 340 152 356 186
rect 290 118 356 152
rect 434 131 464 217
rect 506 225 536 331
rect 578 339 608 491
rect 683 459 713 491
rect 650 443 716 459
rect 650 409 666 443
rect 700 409 716 443
rect 650 393 716 409
rect 758 397 788 491
rect 758 381 856 397
rect 758 359 806 381
rect 790 347 806 359
rect 840 347 856 381
rect 1236 495 1266 521
rect 578 323 644 339
rect 578 289 594 323
rect 628 303 644 323
rect 790 313 856 347
rect 628 289 748 303
rect 578 273 748 289
rect 506 195 568 225
rect 538 131 568 195
rect 610 203 676 219
rect 610 169 626 203
rect 660 169 676 203
rect 610 153 676 169
rect 610 131 640 153
rect 718 131 748 273
rect 790 279 806 313
rect 840 279 856 313
rect 941 303 971 355
rect 790 255 856 279
rect 901 287 971 303
rect 790 131 820 255
rect 901 253 917 287
rect 951 253 971 287
rect 1013 303 1079 319
rect 1013 269 1029 303
rect 1063 283 1079 303
rect 1131 283 1161 367
rect 1236 283 1266 367
rect 1426 335 1456 367
rect 1063 269 1266 283
rect 1381 319 1456 335
rect 1381 285 1397 319
rect 1431 285 1456 319
rect 1381 269 1456 285
rect 1013 253 1266 269
rect 901 237 971 253
rect 901 215 931 237
rect 1131 231 1161 253
rect 1236 231 1266 253
rect 1426 247 1456 269
rect 290 84 306 118
rect 340 84 356 118
rect 290 68 356 84
rect 99 36 129 62
rect 185 36 215 62
rect 1236 121 1266 147
rect 434 21 464 47
rect 538 21 568 47
rect 610 21 640 47
rect 718 21 748 47
rect 790 21 820 47
rect 901 21 931 47
rect 1131 37 1161 63
rect 1426 53 1456 79
<< polycont >>
rect 93 252 127 286
rect 93 184 127 218
rect 486 347 520 381
rect 414 233 448 267
rect 306 152 340 186
rect 666 409 700 443
rect 806 347 840 381
rect 594 289 628 323
rect 626 169 660 203
rect 806 279 840 313
rect 917 253 951 287
rect 1029 269 1063 303
rect 1397 285 1431 319
rect 306 84 340 118
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 52 535 111 551
rect 52 501 68 535
rect 102 501 111 535
rect 52 465 111 501
rect 52 431 68 465
rect 102 431 111 465
rect 52 381 111 431
rect 145 535 197 649
rect 359 605 425 615
rect 359 571 375 605
rect 409 571 425 605
rect 145 501 154 535
rect 188 501 197 535
rect 145 465 197 501
rect 145 431 154 465
rect 188 431 197 465
rect 145 415 197 431
rect 231 535 290 551
rect 231 501 240 535
rect 274 501 290 535
rect 231 465 290 501
rect 359 537 425 571
rect 459 603 511 649
rect 459 569 461 603
rect 495 569 511 603
rect 459 553 511 569
rect 603 595 770 615
rect 603 561 619 595
rect 653 561 770 595
rect 603 553 770 561
rect 359 503 375 537
rect 409 519 425 537
rect 409 503 702 519
rect 359 485 702 503
rect 231 431 240 465
rect 274 451 290 465
rect 274 431 628 451
rect 231 415 628 431
rect 17 347 486 381
rect 520 347 536 381
rect 17 341 536 347
rect 17 134 57 341
rect 578 323 628 415
rect 578 307 594 323
rect 91 286 183 302
rect 91 252 93 286
rect 127 252 183 286
rect 91 218 183 252
rect 91 184 93 218
rect 127 184 183 218
rect 91 168 183 184
rect 217 289 594 307
rect 217 273 628 289
rect 662 443 702 485
rect 662 409 666 443
rect 700 409 702 443
rect 217 267 464 273
rect 217 257 414 267
rect 17 118 98 134
rect 17 84 54 118
rect 88 84 98 118
rect 17 68 98 84
rect 132 118 183 134
rect 132 84 140 118
rect 174 84 183 118
rect 132 17 183 84
rect 217 123 272 257
rect 398 233 414 257
rect 448 233 464 267
rect 662 237 702 409
rect 217 89 226 123
rect 260 89 272 123
rect 217 73 272 89
rect 306 186 355 223
rect 398 217 464 233
rect 340 152 355 186
rect 610 203 702 237
rect 736 229 770 553
rect 804 595 946 649
rect 804 561 896 595
rect 930 561 946 595
rect 804 548 946 561
rect 804 514 805 548
rect 839 527 946 548
rect 839 514 896 527
rect 804 493 896 514
rect 930 493 946 527
rect 804 471 946 493
rect 880 459 946 471
rect 880 425 896 459
rect 930 425 946 459
rect 880 423 946 425
rect 980 595 1032 611
rect 980 561 982 595
rect 1016 561 1032 595
rect 980 503 1032 561
rect 980 469 982 503
rect 1016 469 1032 503
rect 980 405 1032 469
rect 804 389 842 397
rect 980 389 982 405
rect 804 381 982 389
rect 804 347 806 381
rect 840 371 982 381
rect 1016 371 1032 405
rect 840 355 1032 371
rect 1070 599 1133 615
rect 1070 565 1086 599
rect 1120 565 1133 599
rect 1070 503 1133 565
rect 1070 469 1086 503
rect 1120 469 1133 503
rect 1070 413 1133 469
rect 1070 379 1086 413
rect 1120 379 1133 413
rect 1070 363 1133 379
rect 1167 607 1227 649
rect 1167 573 1172 607
rect 1206 573 1227 607
rect 1167 507 1227 573
rect 1167 473 1172 507
rect 1206 473 1227 507
rect 1365 607 1431 649
rect 1365 573 1381 607
rect 1415 573 1431 607
rect 1365 508 1431 573
rect 1167 413 1227 473
rect 1167 379 1182 413
rect 1216 379 1227 413
rect 1167 363 1227 379
rect 1261 483 1327 499
rect 1261 449 1277 483
rect 1311 449 1327 483
rect 1261 413 1327 449
rect 1261 379 1277 413
rect 1311 379 1327 413
rect 840 347 842 355
rect 804 313 842 347
rect 804 279 806 313
rect 840 279 842 313
rect 987 319 1032 355
rect 987 303 1063 319
rect 804 263 842 279
rect 876 287 951 303
rect 876 253 917 287
rect 876 237 951 253
rect 987 269 1029 303
rect 987 253 1063 269
rect 876 229 910 237
rect 610 183 626 203
rect 306 118 355 152
rect 340 84 355 118
rect 306 51 355 84
rect 389 169 626 183
rect 660 169 662 203
rect 389 149 662 169
rect 736 195 910 229
rect 987 201 1021 253
rect 1099 219 1133 363
rect 1261 335 1327 379
rect 1365 474 1381 508
rect 1415 474 1431 508
rect 1365 413 1431 474
rect 1365 379 1381 413
rect 1415 379 1431 413
rect 1365 369 1431 379
rect 1465 599 1519 615
rect 1465 565 1467 599
rect 1501 565 1519 599
rect 1465 502 1519 565
rect 1465 468 1467 502
rect 1501 468 1519 502
rect 1465 413 1519 468
rect 1465 379 1467 413
rect 1501 379 1519 413
rect 1261 319 1431 335
rect 1261 285 1397 319
rect 1261 269 1431 285
rect 736 167 770 195
rect 389 106 427 149
rect 696 133 770 167
rect 944 185 1021 201
rect 696 115 730 133
rect 423 72 427 106
rect 389 56 427 72
rect 468 99 534 115
rect 468 65 484 99
rect 518 65 534 99
rect 468 17 534 65
rect 645 99 730 115
rect 645 65 661 99
rect 695 65 730 99
rect 645 55 730 65
rect 815 127 856 161
rect 890 127 906 161
rect 815 93 906 127
rect 815 59 831 93
rect 865 59 906 93
rect 815 17 906 59
rect 944 151 946 185
rect 980 151 1021 185
rect 944 101 1021 151
rect 944 67 946 101
rect 980 67 1021 101
rect 944 51 1021 67
rect 1070 203 1133 219
rect 1070 169 1086 203
rect 1120 169 1133 203
rect 1070 118 1133 169
rect 1070 84 1086 118
rect 1120 84 1133 118
rect 1070 51 1133 84
rect 1167 218 1227 234
rect 1167 184 1180 218
rect 1214 184 1227 218
rect 1167 109 1227 184
rect 1261 208 1327 269
rect 1465 235 1519 379
rect 1261 174 1277 208
rect 1311 174 1327 208
rect 1261 158 1327 174
rect 1365 201 1381 235
rect 1415 201 1431 235
rect 1167 75 1172 109
rect 1206 75 1227 109
rect 1167 17 1227 75
rect 1365 125 1431 201
rect 1365 91 1381 125
rect 1415 91 1431 125
rect 1365 17 1431 91
rect 1465 201 1467 235
rect 1501 201 1519 235
rect 1465 125 1519 201
rect 1465 91 1467 125
rect 1501 91 1519 125
rect 1465 75 1519 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlxbp_1
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1471 94 1505 128 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1471 168 1505 202 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1471 390 1505 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1471 464 1505 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1471 538 1505 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1087 94 1121 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2293442
string GDS_START 2280380
<< end >>
