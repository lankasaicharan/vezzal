magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 20 49 606 243
rect 0 0 672 49
<< scnmos >>
rect 103 133 133 217
rect 221 49 251 217
rect 307 49 337 217
rect 425 133 455 217
rect 497 133 527 217
<< scpmoshvt >>
rect 81 367 111 451
rect 186 367 216 619
rect 272 367 302 619
rect 411 367 441 451
rect 497 367 527 451
<< ndiff >>
rect 46 192 103 217
rect 46 158 54 192
rect 88 158 103 192
rect 46 133 103 158
rect 133 133 221 217
rect 148 69 221 133
rect 148 35 160 69
rect 194 49 221 69
rect 251 209 307 217
rect 251 175 262 209
rect 296 175 307 209
rect 251 49 307 175
rect 337 133 425 217
rect 455 133 497 217
rect 527 195 580 217
rect 527 161 538 195
rect 572 161 580 195
rect 527 133 580 161
rect 337 69 410 133
rect 337 49 364 69
rect 194 35 206 49
rect 148 27 206 35
rect 352 35 364 49
rect 398 35 410 69
rect 352 27 410 35
<< pdiff >>
rect 133 607 186 619
rect 133 573 141 607
rect 175 573 186 607
rect 133 516 186 573
rect 133 482 141 516
rect 175 482 186 516
rect 133 451 186 482
rect 28 426 81 451
rect 28 392 36 426
rect 70 392 81 426
rect 28 367 81 392
rect 111 434 186 451
rect 111 400 122 434
rect 156 400 186 434
rect 111 367 186 400
rect 216 599 272 619
rect 216 565 227 599
rect 261 565 272 599
rect 216 502 272 565
rect 216 468 227 502
rect 261 468 272 502
rect 216 413 272 468
rect 216 379 227 413
rect 261 379 272 413
rect 216 367 272 379
rect 302 607 355 619
rect 302 573 313 607
rect 347 573 355 607
rect 302 507 355 573
rect 302 473 313 507
rect 347 473 355 507
rect 302 451 355 473
rect 302 427 411 451
rect 302 393 366 427
rect 400 393 411 427
rect 302 367 411 393
rect 441 426 497 451
rect 441 392 452 426
rect 486 392 497 426
rect 441 367 497 392
rect 527 432 580 451
rect 527 398 538 432
rect 572 398 580 432
rect 527 367 580 398
<< ndiffc >>
rect 54 158 88 192
rect 160 35 194 69
rect 262 175 296 209
rect 538 161 572 195
rect 364 35 398 69
<< pdiffc >>
rect 141 573 175 607
rect 141 482 175 516
rect 36 392 70 426
rect 122 400 156 434
rect 227 565 261 599
rect 227 468 261 502
rect 227 379 261 413
rect 313 573 347 607
rect 313 473 347 507
rect 366 393 400 427
rect 452 392 486 426
rect 538 398 572 432
<< poly >>
rect 186 619 216 645
rect 272 619 302 645
rect 81 451 111 477
rect 411 451 441 477
rect 497 451 527 477
rect 81 308 111 367
rect 72 292 138 308
rect 72 258 88 292
rect 122 258 138 292
rect 72 242 138 258
rect 186 299 216 367
rect 272 335 302 367
rect 272 319 347 335
rect 272 299 297 319
rect 186 285 297 299
rect 331 285 347 319
rect 411 305 441 367
rect 186 269 347 285
rect 389 289 455 305
rect 103 217 133 242
rect 186 239 251 269
rect 221 217 251 239
rect 307 217 337 269
rect 389 255 405 289
rect 439 255 455 289
rect 389 239 455 255
rect 425 217 455 239
rect 497 269 527 367
rect 497 239 533 269
rect 497 217 527 239
rect 103 107 133 133
rect 425 107 455 133
rect 497 111 527 133
rect 221 23 251 49
rect 307 23 337 49
rect 497 95 563 111
rect 497 61 513 95
rect 547 61 563 95
rect 497 45 563 61
<< polycont >>
rect 88 258 122 292
rect 297 285 331 319
rect 405 255 439 289
rect 513 61 547 95
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 120 607 184 649
rect 120 573 141 607
rect 175 573 184 607
rect 120 516 184 573
rect 120 482 141 516
rect 175 482 184 516
rect 18 426 86 442
rect 18 392 36 426
rect 70 392 86 426
rect 18 384 86 392
rect 120 434 184 482
rect 120 400 122 434
rect 156 400 184 434
rect 120 384 184 400
rect 218 599 263 615
rect 218 565 227 599
rect 261 565 263 599
rect 218 502 263 565
rect 218 468 227 502
rect 261 468 263 502
rect 218 413 263 468
rect 18 203 52 384
rect 218 379 227 413
rect 261 379 263 413
rect 297 607 416 649
rect 297 573 313 607
rect 347 573 416 607
rect 297 507 416 573
rect 297 473 313 507
rect 347 473 416 507
rect 297 427 416 473
rect 297 393 366 427
rect 400 393 416 427
rect 450 426 488 442
rect 88 292 184 350
rect 122 258 184 292
rect 88 237 184 258
rect 218 225 263 379
rect 450 392 452 426
rect 486 392 488 426
rect 522 432 588 649
rect 522 398 538 432
rect 572 398 588 432
rect 522 393 588 398
rect 450 359 488 392
rect 297 325 632 359
rect 297 319 347 325
rect 331 285 347 319
rect 297 269 347 285
rect 389 289 547 291
rect 389 255 405 289
rect 439 255 547 289
rect 389 240 547 255
rect 218 209 312 225
rect 18 192 104 203
rect 18 158 54 192
rect 88 158 104 192
rect 218 175 262 209
rect 296 175 312 209
rect 581 206 632 325
rect 522 195 632 206
rect 18 141 104 158
rect 522 161 538 195
rect 572 161 632 195
rect 522 145 632 161
rect 18 111 486 141
rect 18 107 563 111
rect 452 95 563 107
rect 144 69 210 73
rect 144 35 160 69
rect 194 35 210 69
rect 144 17 210 35
rect 348 69 414 73
rect 348 35 364 69
rect 398 35 414 69
rect 452 61 513 95
rect 547 61 563 95
rect 452 51 563 61
rect 348 17 414 35
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and2b_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5126662
string GDS_START 5120406
<< end >>
