magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1288 -1260 2888 1289
use sky130_fd_pr__dfl1sd__example_5595914180868  sky130_fd_pr__dfl1sd__example_5595914180868_0
timestamp 1627201311
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180868  sky130_fd_pr__dfl1sd__example_5595914180868_1
timestamp 1627201311
transform 1 0 1600 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 1628 29 1628 29 0 FreeSans 300 0 0 0 D
flabel comment s -28 29 -28 29 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 38324904
string GDS_START 38323982
<< end >>
