magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3890 1975
<< nwell >>
rect -38 394 2630 704
rect -38 331 1677 394
rect 1931 331 2630 394
rect 1931 307 2299 331
<< pwell >>
rect 1780 241 1889 313
rect 1780 208 2589 241
rect 1206 201 2589 208
rect 1 157 197 167
rect 788 157 2589 201
rect 1 49 2589 157
rect 0 0 2592 49
<< scnmos >>
rect 84 57 114 141
rect 282 47 312 131
rect 501 47 531 131
rect 587 47 617 131
rect 689 47 719 131
rect 767 47 797 131
rect 887 47 917 175
rect 973 47 1003 175
rect 1091 47 1121 175
rect 1289 54 1319 182
rect 1367 54 1397 182
rect 1469 98 1499 182
rect 1547 98 1577 182
rect 1675 54 1705 182
rect 1761 54 1791 182
rect 1878 54 1908 182
rect 2075 131 2105 215
rect 2177 47 2207 215
rect 2374 131 2404 215
rect 2476 47 2506 215
<< scpmoshvt >>
rect 114 481 144 609
rect 312 463 342 591
rect 537 463 567 547
rect 623 463 653 547
rect 725 463 755 547
rect 803 463 833 547
rect 930 379 960 547
rect 1016 379 1046 547
rect 1094 379 1124 547
rect 1182 379 1212 547
rect 1277 428 1307 596
rect 1389 512 1419 596
rect 1547 512 1577 596
rect 1689 430 1719 598
rect 1793 430 1823 598
rect 1875 430 1905 598
rect 2074 343 2104 471
rect 2176 343 2206 595
rect 2374 367 2404 495
rect 2476 367 2506 619
<< ndiff >>
rect 27 116 84 141
rect 27 82 39 116
rect 73 82 84 116
rect 27 57 84 82
rect 114 116 171 141
rect 1806 275 1863 287
rect 1806 241 1818 275
rect 1852 241 1863 275
rect 1806 182 1863 241
rect 814 131 887 175
rect 114 82 125 116
rect 159 82 171 116
rect 114 57 171 82
rect 225 111 282 131
rect 225 77 237 111
rect 271 77 282 111
rect 225 47 282 77
rect 312 97 501 131
rect 312 63 369 97
rect 403 63 501 97
rect 312 47 501 63
rect 531 111 587 131
rect 531 77 542 111
rect 576 77 587 111
rect 531 47 587 77
rect 617 108 689 131
rect 617 74 644 108
rect 678 74 689 108
rect 617 47 689 74
rect 719 47 767 131
rect 797 126 887 131
rect 797 92 826 126
rect 860 92 887 126
rect 797 47 887 92
rect 917 131 973 175
rect 917 97 928 131
rect 962 97 973 131
rect 917 47 973 97
rect 1003 160 1091 175
rect 1003 126 1030 160
rect 1064 126 1091 160
rect 1003 47 1091 126
rect 1121 99 1178 175
rect 1121 65 1132 99
rect 1166 65 1178 99
rect 1121 47 1178 65
rect 1232 100 1289 182
rect 1232 66 1244 100
rect 1278 66 1289 100
rect 1232 54 1289 66
rect 1319 54 1367 182
rect 1397 163 1469 182
rect 1397 129 1408 163
rect 1442 129 1469 163
rect 1397 98 1469 129
rect 1499 98 1547 182
rect 1577 118 1675 182
rect 1577 98 1614 118
rect 1397 54 1454 98
rect 1602 84 1614 98
rect 1648 84 1675 118
rect 1602 54 1675 84
rect 1705 103 1761 182
rect 1705 69 1716 103
rect 1750 69 1761 103
rect 1705 54 1761 69
rect 1791 54 1878 182
rect 1908 103 1964 182
rect 2018 180 2075 215
rect 2018 146 2030 180
rect 2064 146 2075 180
rect 2018 131 2075 146
rect 2105 184 2177 215
rect 2105 150 2132 184
rect 2166 150 2177 184
rect 2105 131 2177 150
rect 1908 69 1919 103
rect 1953 69 1964 103
rect 1908 54 1964 69
rect 2120 93 2177 131
rect 2120 59 2132 93
rect 2166 59 2177 93
rect 2120 47 2177 59
rect 2207 185 2264 215
rect 2207 151 2218 185
rect 2252 151 2264 185
rect 2207 103 2264 151
rect 2318 190 2374 215
rect 2318 156 2329 190
rect 2363 156 2374 190
rect 2318 131 2374 156
rect 2404 171 2476 215
rect 2404 137 2431 171
rect 2465 137 2476 171
rect 2404 131 2476 137
rect 2207 69 2218 103
rect 2252 69 2264 103
rect 2207 47 2264 69
rect 2419 93 2476 131
rect 2419 59 2431 93
rect 2465 59 2476 93
rect 2419 47 2476 59
rect 2506 203 2563 215
rect 2506 169 2517 203
rect 2551 169 2563 203
rect 2506 103 2563 169
rect 2506 69 2517 103
rect 2551 69 2563 103
rect 2506 47 2563 69
<< pdiff >>
rect 41 597 114 609
rect 41 563 53 597
rect 87 563 114 597
rect 41 527 114 563
rect 41 493 53 527
rect 87 493 114 527
rect 41 481 114 493
rect 144 597 201 609
rect 144 563 155 597
rect 189 563 201 597
rect 144 527 201 563
rect 144 493 155 527
rect 189 493 201 527
rect 144 481 201 493
rect 255 579 312 591
rect 255 545 267 579
rect 301 545 312 579
rect 255 509 312 545
rect 255 475 267 509
rect 301 475 312 509
rect 255 463 312 475
rect 342 573 415 591
rect 342 539 369 573
rect 403 547 415 573
rect 857 586 915 598
rect 1632 596 1689 598
rect 857 552 869 586
rect 903 552 915 586
rect 857 547 915 552
rect 1227 547 1277 596
rect 403 539 537 547
rect 342 463 537 539
rect 567 522 623 547
rect 567 488 578 522
rect 612 488 623 522
rect 567 463 623 488
rect 653 533 725 547
rect 653 499 680 533
rect 714 499 725 533
rect 653 463 725 499
rect 755 463 803 547
rect 833 463 930 547
rect 857 379 930 463
rect 960 535 1016 547
rect 960 501 971 535
rect 1005 501 1016 535
rect 960 442 1016 501
rect 960 408 971 442
rect 1005 408 1016 442
rect 960 379 1016 408
rect 1046 379 1094 547
rect 1124 523 1182 547
rect 1124 489 1135 523
rect 1169 489 1182 523
rect 1124 379 1182 489
rect 1212 428 1277 547
rect 1307 575 1389 596
rect 1307 541 1344 575
rect 1378 541 1389 575
rect 1307 512 1389 541
rect 1419 512 1547 596
rect 1577 586 1689 596
rect 1577 552 1644 586
rect 1678 552 1689 586
rect 1577 512 1689 552
rect 1307 428 1357 512
rect 1212 379 1262 428
rect 1632 430 1689 512
rect 1719 586 1793 598
rect 1719 552 1748 586
rect 1782 552 1793 586
rect 1719 479 1793 552
rect 1719 445 1748 479
rect 1782 445 1793 479
rect 1719 430 1793 445
rect 1823 430 1875 598
rect 1905 573 1962 598
rect 2419 607 2476 619
rect 1905 539 1916 573
rect 1950 539 1962 573
rect 1905 430 1962 539
rect 2119 572 2176 595
rect 2119 538 2131 572
rect 2165 538 2176 572
rect 2119 471 2176 538
rect 2017 389 2074 471
rect 2017 355 2029 389
rect 2063 355 2074 389
rect 2017 343 2074 355
rect 2104 343 2176 471
rect 2206 583 2263 595
rect 2206 549 2217 583
rect 2251 549 2263 583
rect 2206 486 2263 549
rect 2419 573 2431 607
rect 2465 573 2476 607
rect 2419 510 2476 573
rect 2419 495 2431 510
rect 2206 452 2217 486
rect 2251 452 2263 486
rect 2206 389 2263 452
rect 2206 355 2217 389
rect 2251 355 2263 389
rect 2317 483 2374 495
rect 2317 449 2329 483
rect 2363 449 2374 483
rect 2317 413 2374 449
rect 2317 379 2329 413
rect 2363 379 2374 413
rect 2317 367 2374 379
rect 2404 476 2431 495
rect 2465 476 2476 510
rect 2404 413 2476 476
rect 2404 379 2431 413
rect 2465 379 2476 413
rect 2404 367 2476 379
rect 2506 597 2563 619
rect 2506 563 2517 597
rect 2551 563 2563 597
rect 2506 505 2563 563
rect 2506 471 2517 505
rect 2551 471 2563 505
rect 2506 413 2563 471
rect 2506 379 2517 413
rect 2551 379 2563 413
rect 2506 367 2563 379
rect 2206 343 2263 355
<< ndiffc >>
rect 39 82 73 116
rect 1818 241 1852 275
rect 125 82 159 116
rect 237 77 271 111
rect 369 63 403 97
rect 542 77 576 111
rect 644 74 678 108
rect 826 92 860 126
rect 928 97 962 131
rect 1030 126 1064 160
rect 1132 65 1166 99
rect 1244 66 1278 100
rect 1408 129 1442 163
rect 1614 84 1648 118
rect 1716 69 1750 103
rect 2030 146 2064 180
rect 2132 150 2166 184
rect 1919 69 1953 103
rect 2132 59 2166 93
rect 2218 151 2252 185
rect 2329 156 2363 190
rect 2431 137 2465 171
rect 2218 69 2252 103
rect 2431 59 2465 93
rect 2517 169 2551 203
rect 2517 69 2551 103
<< pdiffc >>
rect 53 563 87 597
rect 53 493 87 527
rect 155 563 189 597
rect 155 493 189 527
rect 267 545 301 579
rect 267 475 301 509
rect 369 539 403 573
rect 869 552 903 586
rect 578 488 612 522
rect 680 499 714 533
rect 971 501 1005 535
rect 971 408 1005 442
rect 1135 489 1169 523
rect 1344 541 1378 575
rect 1644 552 1678 586
rect 1748 552 1782 586
rect 1748 445 1782 479
rect 1916 539 1950 573
rect 2131 538 2165 572
rect 2029 355 2063 389
rect 2217 549 2251 583
rect 2431 573 2465 607
rect 2217 452 2251 486
rect 2217 355 2251 389
rect 2329 449 2363 483
rect 2329 379 2363 413
rect 2431 476 2465 510
rect 2431 379 2465 413
rect 2517 563 2551 597
rect 2517 471 2551 505
rect 2517 379 2551 413
<< poly >>
rect 114 609 144 635
rect 312 615 1307 645
rect 312 591 342 615
rect 114 466 144 481
rect 61 436 144 466
rect 537 547 567 573
rect 623 547 653 573
rect 725 547 755 615
rect 1277 596 1307 615
rect 1389 596 1419 622
rect 1547 596 1577 622
rect 1689 598 1719 624
rect 1793 598 1823 624
rect 1875 598 1905 624
rect 803 547 833 573
rect 930 547 960 573
rect 1016 547 1046 573
rect 1094 547 1124 573
rect 1182 547 1212 573
rect 61 315 91 436
rect 25 299 91 315
rect 25 265 41 299
rect 75 265 91 299
rect 25 231 91 265
rect 139 372 205 388
rect 139 338 155 372
rect 189 338 205 372
rect 139 304 205 338
rect 139 270 155 304
rect 189 297 205 304
rect 312 297 342 463
rect 537 448 567 463
rect 426 418 567 448
rect 426 411 456 418
rect 390 395 456 411
rect 390 361 406 395
rect 440 361 456 395
rect 623 376 653 463
rect 725 437 755 463
rect 390 345 456 361
rect 534 360 719 376
rect 534 326 550 360
rect 584 326 719 360
rect 803 347 833 463
rect 1389 480 1419 512
rect 1389 464 1455 480
rect 1389 430 1405 464
rect 1439 430 1455 464
rect 1277 413 1307 428
rect 1389 414 1455 430
rect 1277 383 1347 413
rect 1547 398 1577 512
rect 2176 595 2206 621
rect 2476 619 2506 645
rect 2074 471 2104 497
rect 1689 398 1719 430
rect 930 355 960 379
rect 534 310 719 326
rect 189 270 492 297
rect 139 267 492 270
rect 139 254 205 267
rect 25 197 41 231
rect 75 206 91 231
rect 75 197 114 206
rect 25 176 114 197
rect 84 141 114 176
rect 282 131 312 267
rect 462 261 492 267
rect 462 231 617 261
rect 354 203 420 219
rect 354 169 370 203
rect 404 183 420 203
rect 404 169 531 183
rect 354 153 531 169
rect 501 131 531 153
rect 587 131 617 231
rect 689 131 719 310
rect 767 331 833 347
rect 767 297 783 331
rect 817 297 833 331
rect 767 281 833 297
rect 875 331 960 355
rect 875 297 891 331
rect 925 325 960 331
rect 925 297 941 325
rect 875 281 941 297
rect 767 131 797 281
rect 887 175 917 281
rect 1016 277 1046 379
rect 983 261 1049 277
rect 1094 263 1124 379
rect 1182 335 1212 379
rect 1317 366 1347 383
rect 1545 382 1611 398
rect 1317 336 1499 366
rect 1182 305 1275 335
rect 1245 288 1275 305
rect 1245 272 1319 288
rect 983 233 999 261
rect 973 227 999 233
rect 1033 227 1049 261
rect 973 203 1049 227
rect 1091 247 1203 263
rect 1091 213 1153 247
rect 1187 213 1203 247
rect 1245 238 1261 272
rect 1295 238 1319 272
rect 1245 222 1319 238
rect 1361 272 1427 288
rect 1361 238 1377 272
rect 1411 238 1427 272
rect 1361 222 1427 238
rect 973 175 1003 203
rect 1091 197 1203 213
rect 1091 175 1121 197
rect 1289 182 1319 222
rect 1367 182 1397 222
rect 1469 182 1499 336
rect 1545 348 1561 382
rect 1595 348 1611 382
rect 1545 332 1611 348
rect 1653 382 1719 398
rect 1793 393 1823 430
rect 1653 348 1669 382
rect 1703 348 1719 382
rect 1653 332 1719 348
rect 1761 377 1827 393
rect 1761 343 1777 377
rect 1811 343 1827 377
rect 1547 182 1577 332
rect 1675 182 1705 332
rect 1761 327 1827 343
rect 1875 332 1905 430
rect 2374 495 2404 521
rect 1761 182 1791 327
rect 1875 302 2002 332
rect 2074 303 2104 343
rect 2176 303 2206 343
rect 1878 295 2002 302
rect 1878 261 1952 295
rect 1986 261 2002 295
rect 1878 245 2002 261
rect 2044 287 2110 303
rect 2044 253 2060 287
rect 2094 253 2110 287
rect 1878 182 1908 245
rect 2044 237 2110 253
rect 2153 287 2219 303
rect 2153 253 2169 287
rect 2203 267 2219 287
rect 2374 267 2404 367
rect 2476 327 2506 367
rect 2203 253 2404 267
rect 2446 311 2512 327
rect 2446 277 2462 311
rect 2496 277 2512 311
rect 2446 261 2512 277
rect 2153 237 2404 253
rect 2075 215 2105 237
rect 2177 215 2207 237
rect 2374 215 2404 237
rect 2476 215 2506 261
rect 84 31 114 57
rect 1469 72 1499 98
rect 1547 72 1577 98
rect 2075 105 2105 131
rect 282 21 312 47
rect 501 21 531 47
rect 587 21 617 47
rect 689 21 719 47
rect 767 21 797 47
rect 887 21 917 47
rect 973 21 1003 47
rect 1091 21 1121 47
rect 1289 28 1319 54
rect 1367 28 1397 54
rect 1675 28 1705 54
rect 1761 28 1791 54
rect 1878 28 1908 54
rect 2374 105 2404 131
rect 2177 21 2207 47
rect 2476 21 2506 47
<< polycont >>
rect 41 265 75 299
rect 155 338 189 372
rect 155 270 189 304
rect 406 361 440 395
rect 550 326 584 360
rect 1405 430 1439 464
rect 41 197 75 231
rect 370 169 404 203
rect 783 297 817 331
rect 891 297 925 331
rect 999 227 1033 261
rect 1153 213 1187 247
rect 1261 238 1295 272
rect 1377 238 1411 272
rect 1561 348 1595 382
rect 1669 348 1703 382
rect 1777 343 1811 377
rect 1952 261 1986 295
rect 2060 253 2094 287
rect 2169 253 2203 287
rect 2462 277 2496 311
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 37 597 103 649
rect 37 563 53 597
rect 87 563 103 597
rect 37 527 103 563
rect 37 493 53 527
rect 87 493 103 527
rect 37 477 103 493
rect 139 597 205 613
rect 139 563 155 597
rect 189 563 205 597
rect 139 527 205 563
rect 139 493 155 527
rect 189 493 205 527
rect 25 299 91 430
rect 25 265 41 299
rect 75 265 91 299
rect 25 231 91 265
rect 25 197 41 231
rect 75 197 91 231
rect 25 181 91 197
rect 139 372 205 493
rect 139 338 155 372
rect 189 338 205 372
rect 139 304 205 338
rect 139 270 155 304
rect 189 270 205 304
rect 139 254 205 270
rect 251 579 317 595
rect 251 545 267 579
rect 301 545 317 579
rect 251 509 317 545
rect 353 573 419 649
rect 353 539 369 573
rect 403 539 419 573
rect 853 586 919 649
rect 853 552 869 586
rect 903 552 919 586
rect 353 517 419 539
rect 562 522 628 551
rect 251 475 267 509
rect 301 481 317 509
rect 562 488 578 522
rect 612 488 628 522
rect 301 475 526 481
rect 251 447 526 475
rect 139 145 175 254
rect 23 116 73 145
rect 23 82 39 116
rect 23 17 73 82
rect 109 116 175 145
rect 251 135 317 447
rect 354 395 456 411
rect 354 361 406 395
rect 440 361 456 395
rect 354 203 456 361
rect 492 376 526 447
rect 562 446 628 488
rect 664 533 740 551
rect 853 536 919 552
rect 664 499 680 533
rect 714 499 740 533
rect 971 535 1021 551
rect 1005 501 1021 535
rect 971 500 1021 501
rect 664 482 740 499
rect 562 412 670 446
rect 492 360 600 376
rect 492 326 550 360
rect 584 326 600 360
rect 492 312 600 326
rect 492 276 551 312
rect 492 242 511 276
rect 545 242 551 276
rect 492 236 551 242
rect 354 169 370 203
rect 404 169 456 203
rect 636 200 670 412
rect 354 153 456 169
rect 526 166 670 200
rect 706 245 740 482
rect 776 466 1021 500
rect 776 331 833 466
rect 971 442 1021 466
rect 1119 523 1185 649
rect 1119 489 1135 523
rect 1169 489 1185 523
rect 1328 575 1394 600
rect 1328 541 1344 575
rect 1378 550 1394 575
rect 1628 586 1694 649
rect 1628 552 1644 586
rect 1678 552 1694 586
rect 1378 541 1517 550
rect 1328 516 1517 541
rect 1628 536 1694 552
rect 1748 586 1798 602
rect 1782 552 1798 586
rect 1119 462 1185 489
rect 1361 464 1447 480
rect 776 297 783 331
rect 817 297 833 331
rect 776 281 833 297
rect 875 424 935 430
rect 875 390 895 424
rect 929 390 935 424
rect 1005 426 1021 442
rect 1361 430 1405 464
rect 1439 430 1447 464
rect 1005 408 1311 426
rect 971 392 1311 408
rect 875 356 935 390
rect 875 331 941 356
rect 875 297 891 331
rect 925 297 941 331
rect 875 281 941 297
rect 983 261 1040 277
rect 983 245 999 261
rect 706 227 999 245
rect 1033 227 1040 261
rect 706 211 1040 227
rect 109 82 125 116
rect 159 82 175 116
rect 109 53 175 82
rect 221 111 317 135
rect 221 77 237 111
rect 271 77 317 111
rect 221 53 317 77
rect 353 97 419 117
rect 353 63 369 97
rect 403 63 419 97
rect 353 17 419 63
rect 526 111 592 166
rect 706 130 740 211
rect 1076 175 1110 392
rect 1245 272 1311 392
rect 526 77 542 111
rect 576 77 592 111
rect 526 53 592 77
rect 628 108 740 130
rect 628 74 644 108
rect 678 96 740 108
rect 810 126 876 175
rect 678 74 694 96
rect 628 53 694 74
rect 810 92 826 126
rect 860 92 876 126
rect 810 17 876 92
rect 912 131 978 175
rect 912 97 928 131
rect 962 97 978 131
rect 1014 160 1110 175
rect 1014 126 1030 160
rect 1064 141 1110 160
rect 1146 247 1203 263
rect 1146 213 1153 247
rect 1187 213 1203 247
rect 1245 238 1261 272
rect 1295 238 1311 272
rect 1245 222 1311 238
rect 1361 414 1447 430
rect 1361 276 1427 414
rect 1483 296 1517 516
rect 1748 500 1798 552
rect 1900 573 1966 649
rect 1900 539 1916 573
rect 1950 539 1966 573
rect 1900 511 1966 539
rect 2115 572 2181 649
rect 2415 607 2465 649
rect 2115 538 2131 572
rect 2165 538 2181 572
rect 2115 511 2181 538
rect 2217 583 2289 599
rect 2251 549 2289 583
rect 1553 479 1798 500
rect 1553 466 1748 479
rect 1553 382 1611 466
rect 1782 475 1798 479
rect 2217 486 2289 549
rect 2415 573 2431 607
rect 2415 510 2465 573
rect 1782 445 2181 475
rect 1748 441 2181 445
rect 1553 348 1561 382
rect 1595 348 1611 382
rect 1553 332 1611 348
rect 1653 424 1712 430
rect 1748 429 1897 441
rect 1653 390 1663 424
rect 1697 390 1712 424
rect 1653 382 1712 390
rect 1653 348 1669 382
rect 1703 348 1712 382
rect 1653 332 1712 348
rect 1748 377 1827 393
rect 1748 343 1777 377
rect 1811 343 1827 377
rect 1748 327 1827 343
rect 1748 296 1782 327
rect 1361 242 1375 276
rect 1409 272 1427 276
rect 1361 238 1377 242
rect 1411 238 1427 272
rect 1361 222 1427 238
rect 1463 262 1782 296
rect 1863 291 1897 429
rect 1818 275 1897 291
rect 1146 186 1203 213
rect 1463 186 1497 262
rect 1852 241 1897 275
rect 1818 225 1897 241
rect 1936 389 2079 405
rect 1936 355 2029 389
rect 2063 355 2079 389
rect 1936 339 2079 355
rect 1936 295 2002 339
rect 2147 303 2181 441
rect 2251 452 2289 486
rect 2217 389 2289 452
rect 2251 355 2289 389
rect 2217 339 2289 355
rect 1936 261 1952 295
rect 1986 261 2002 295
rect 1146 152 1348 186
rect 1064 126 1080 141
rect 1014 123 1080 126
rect 912 87 978 97
rect 1116 99 1182 105
rect 1116 87 1132 99
rect 912 65 1132 87
rect 1166 65 1182 99
rect 912 53 1182 65
rect 1228 100 1278 116
rect 1228 66 1244 100
rect 1228 17 1278 66
rect 1314 87 1348 152
rect 1392 163 1497 186
rect 1392 129 1408 163
rect 1442 129 1497 163
rect 1392 123 1497 129
rect 1533 189 1782 223
rect 1936 200 2002 261
rect 2041 287 2110 303
rect 2041 253 2060 287
rect 2094 253 2110 287
rect 2041 236 2110 253
rect 2147 287 2219 303
rect 2147 253 2169 287
rect 2203 253 2219 287
rect 2147 237 2219 253
rect 2255 201 2289 339
rect 2329 483 2379 499
rect 2363 449 2379 483
rect 2329 413 2379 449
rect 2363 379 2379 413
rect 2329 327 2379 379
rect 2415 476 2431 510
rect 2415 413 2465 476
rect 2415 379 2431 413
rect 2415 363 2465 379
rect 2501 597 2574 613
rect 2501 563 2517 597
rect 2551 563 2574 597
rect 2501 505 2574 563
rect 2501 471 2517 505
rect 2551 471 2574 505
rect 2501 413 2574 471
rect 2501 379 2517 413
rect 2551 379 2574 413
rect 2501 363 2574 379
rect 2329 311 2504 327
rect 2329 293 2462 311
rect 2431 277 2462 293
rect 2496 277 2504 311
rect 2431 261 2504 277
rect 2431 257 2465 261
rect 1936 189 2080 200
rect 1533 87 1567 189
rect 1748 180 2080 189
rect 1748 155 2030 180
rect 1314 53 1567 87
rect 1614 118 1664 153
rect 2014 146 2030 155
rect 2064 146 2080 180
rect 2014 127 2080 146
rect 2116 184 2166 200
rect 2116 150 2132 184
rect 1648 84 1664 118
rect 1614 17 1664 84
rect 1700 103 1969 119
rect 1700 69 1716 103
rect 1750 69 1919 103
rect 1953 69 1969 103
rect 1700 53 1969 69
rect 2116 93 2166 150
rect 2116 59 2132 93
rect 2116 17 2166 59
rect 2202 185 2289 201
rect 2202 151 2218 185
rect 2252 151 2289 185
rect 2202 103 2289 151
rect 2329 223 2465 257
rect 2329 190 2379 223
rect 2540 219 2574 363
rect 2363 156 2379 190
rect 2501 203 2574 219
rect 2329 127 2379 156
rect 2415 171 2465 187
rect 2415 137 2431 171
rect 2202 69 2218 103
rect 2252 69 2289 103
rect 2202 53 2289 69
rect 2415 93 2465 137
rect 2415 59 2431 93
rect 2415 17 2465 59
rect 2501 169 2517 203
rect 2551 169 2574 203
rect 2501 103 2574 169
rect 2501 69 2517 103
rect 2551 69 2574 103
rect 2501 53 2574 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 511 242 545 276
rect 895 390 929 424
rect 1663 390 1697 424
rect 1375 272 1409 276
rect 1375 242 1377 272
rect 1377 242 1409 272
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 883 424 941 430
rect 883 390 895 424
rect 929 421 941 424
rect 1651 424 1709 430
rect 1651 421 1663 424
rect 929 393 1663 421
rect 929 390 941 393
rect 883 384 941 390
rect 1651 390 1663 393
rect 1697 390 1709 424
rect 1651 384 1709 390
rect 499 276 557 282
rect 499 242 511 276
rect 545 273 557 276
rect 1363 276 1421 282
rect 1363 273 1375 276
rect 545 245 1375 273
rect 545 242 557 245
rect 499 236 557 242
rect 1363 242 1375 245
rect 1409 242 1421 276
rect 1363 236 1421 242
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
flabel pwell s 0 0 2592 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2592 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfbbp_1
flabel metal1 s 0 617 2592 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2592 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 2239 390 2273 424 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2239 464 2273 498 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2239 538 2273 572 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2527 94 2561 128 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2527 168 2561 202 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 SET_B
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2592 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 7023142
string GDS_START 7004108
<< end >>
