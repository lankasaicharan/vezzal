magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3026 1975
<< nwell >>
rect -38 344 1766 704
rect -38 331 1079 344
rect 1595 331 1766 344
rect 388 319 1079 331
<< pwell >>
rect 1 157 607 211
rect 1121 158 1553 302
rect 1121 157 1703 158
rect 1 49 1703 157
rect 0 0 1728 49
<< scnmos >>
rect 84 101 114 185
rect 162 101 192 185
rect 248 101 278 185
rect 320 101 350 185
rect 406 101 436 185
rect 478 101 508 185
rect 1204 192 1234 276
rect 1276 192 1306 276
rect 1362 192 1392 276
rect 1440 192 1470 276
rect 696 47 726 131
rect 782 47 812 131
rect 860 47 890 131
rect 986 47 1016 131
rect 1064 47 1094 131
rect 1518 48 1548 132
rect 1590 48 1620 132
<< scpmoshvt >>
rect 150 376 200 576
rect 248 376 298 576
rect 397 376 447 576
rect 648 405 698 605
rect 754 405 804 605
rect 860 405 910 605
rect 973 405 1023 605
rect 1228 416 1278 616
rect 1334 416 1384 616
rect 1440 416 1490 616
rect 1578 416 1628 616
<< ndiff >>
rect 27 151 84 185
rect 27 117 39 151
rect 73 117 84 151
rect 27 101 84 117
rect 114 101 162 185
rect 192 160 248 185
rect 192 126 203 160
rect 237 126 248 160
rect 192 101 248 126
rect 278 101 320 185
rect 350 151 406 185
rect 350 117 361 151
rect 395 117 406 151
rect 350 101 406 117
rect 436 101 478 185
rect 508 173 581 185
rect 508 139 535 173
rect 569 139 581 173
rect 508 101 581 139
rect 1147 251 1204 276
rect 1147 217 1159 251
rect 1193 217 1204 251
rect 1147 192 1204 217
rect 1234 192 1276 276
rect 1306 251 1362 276
rect 1306 217 1317 251
rect 1351 217 1362 251
rect 1306 192 1362 217
rect 1392 192 1440 276
rect 1470 251 1527 276
rect 1470 217 1481 251
rect 1515 217 1527 251
rect 1470 192 1527 217
rect 639 111 696 131
rect 639 77 651 111
rect 685 77 696 111
rect 639 47 696 77
rect 726 111 782 131
rect 726 77 737 111
rect 771 77 782 111
rect 726 47 782 77
rect 812 47 860 131
rect 890 106 986 131
rect 890 72 901 106
rect 935 72 986 106
rect 890 47 986 72
rect 1016 47 1064 131
rect 1094 111 1151 131
rect 1094 77 1105 111
rect 1139 77 1151 111
rect 1094 47 1151 77
rect 1457 107 1518 132
rect 1457 73 1469 107
rect 1503 73 1518 107
rect 1457 48 1518 73
rect 1548 48 1590 132
rect 1620 103 1677 132
rect 1620 69 1631 103
rect 1665 69 1677 103
rect 1620 48 1677 69
<< pdiff >>
rect 313 627 371 639
rect 313 593 325 627
rect 359 593 371 627
rect 1505 618 1563 630
rect 1505 616 1517 618
rect 313 576 371 593
rect 591 592 648 605
rect 93 564 150 576
rect 93 530 105 564
rect 139 530 150 564
rect 93 495 150 530
rect 93 461 105 495
rect 139 461 150 495
rect 93 427 150 461
rect 93 393 105 427
rect 139 393 150 427
rect 93 376 150 393
rect 200 376 248 576
rect 298 376 397 576
rect 447 401 520 576
rect 591 558 603 592
rect 637 558 648 592
rect 591 405 648 558
rect 698 451 754 605
rect 698 417 709 451
rect 743 417 754 451
rect 698 405 754 417
rect 804 405 860 605
rect 910 589 973 605
rect 910 555 921 589
rect 955 555 973 589
rect 910 405 973 555
rect 1023 593 1080 605
rect 1023 559 1034 593
rect 1068 559 1080 593
rect 1023 516 1080 559
rect 1023 482 1034 516
rect 1068 482 1080 516
rect 1023 405 1080 482
rect 1171 462 1228 616
rect 1171 428 1183 462
rect 1217 428 1228 462
rect 1171 416 1228 428
rect 1278 603 1334 616
rect 1278 569 1289 603
rect 1323 569 1334 603
rect 1278 416 1334 569
rect 1384 462 1440 616
rect 1384 428 1395 462
rect 1429 428 1440 462
rect 1384 416 1440 428
rect 1490 584 1517 616
rect 1551 616 1563 618
rect 1551 584 1578 616
rect 1490 416 1578 584
rect 1628 597 1685 616
rect 1628 563 1639 597
rect 1673 563 1685 597
rect 1628 462 1685 563
rect 1628 428 1639 462
rect 1673 428 1685 462
rect 1628 416 1685 428
rect 447 376 474 401
rect 462 367 474 376
rect 508 367 520 401
rect 462 355 520 367
<< ndiffc >>
rect 39 117 73 151
rect 203 126 237 160
rect 361 117 395 151
rect 535 139 569 173
rect 1159 217 1193 251
rect 1317 217 1351 251
rect 1481 217 1515 251
rect 651 77 685 111
rect 737 77 771 111
rect 901 72 935 106
rect 1105 77 1139 111
rect 1469 73 1503 107
rect 1631 69 1665 103
<< pdiffc >>
rect 325 593 359 627
rect 105 530 139 564
rect 105 461 139 495
rect 105 393 139 427
rect 603 558 637 592
rect 709 417 743 451
rect 921 555 955 589
rect 1034 559 1068 593
rect 1034 482 1068 516
rect 1183 428 1217 462
rect 1289 569 1323 603
rect 1395 428 1429 462
rect 1517 584 1551 618
rect 1639 563 1673 597
rect 1639 428 1673 462
rect 474 367 508 401
<< poly >>
rect 150 576 200 602
rect 248 576 298 602
rect 648 605 698 631
rect 754 605 804 631
rect 860 605 910 631
rect 973 605 1023 631
rect 1228 616 1278 642
rect 1334 616 1384 642
rect 1440 616 1490 642
rect 397 576 447 602
rect 1578 616 1628 642
rect 150 341 200 376
rect 45 325 200 341
rect 45 291 61 325
rect 95 291 200 325
rect 45 257 200 291
rect 45 223 61 257
rect 95 237 200 257
rect 248 344 298 376
rect 397 344 447 376
rect 648 344 698 405
rect 754 365 804 405
rect 860 373 910 405
rect 248 328 314 344
rect 248 294 264 328
rect 298 294 314 328
rect 248 278 314 294
rect 356 328 447 344
rect 356 294 372 328
rect 406 294 447 328
rect 356 278 447 294
rect 574 328 698 344
rect 574 294 590 328
rect 624 294 698 328
rect 746 349 812 365
rect 746 315 762 349
rect 796 315 812 349
rect 746 299 812 315
rect 860 357 931 373
rect 860 323 881 357
rect 915 323 931 357
rect 860 307 931 323
rect 574 278 698 294
rect 95 223 192 237
rect 45 207 192 223
rect 84 185 114 207
rect 162 185 192 207
rect 248 230 278 278
rect 406 230 436 278
rect 668 251 698 278
rect 248 200 350 230
rect 248 185 278 200
rect 320 185 350 200
rect 406 200 626 230
rect 668 221 812 251
rect 406 185 436 200
rect 478 185 508 200
rect 596 179 626 200
rect 596 149 726 179
rect 696 131 726 149
rect 782 131 812 221
rect 860 131 890 307
rect 973 219 1023 405
rect 1065 357 1131 373
rect 1065 323 1081 357
rect 1115 337 1131 357
rect 1228 337 1278 416
rect 1115 323 1278 337
rect 1065 321 1278 323
rect 1334 321 1384 416
rect 1440 321 1490 416
rect 1578 401 1628 416
rect 1578 371 1695 401
rect 1551 321 1617 329
rect 1065 307 1392 321
rect 1204 291 1392 307
rect 1204 276 1234 291
rect 1276 276 1306 291
rect 1362 276 1392 291
rect 1440 313 1617 321
rect 1440 291 1567 313
rect 1440 276 1470 291
rect 1551 279 1567 291
rect 1601 279 1617 313
rect 986 203 1053 219
rect 986 169 1003 203
rect 1037 177 1053 203
rect 1551 263 1617 279
rect 1665 221 1695 371
rect 1555 205 1695 221
rect 1037 169 1094 177
rect 986 147 1094 169
rect 1204 166 1234 192
rect 1276 166 1306 192
rect 1362 166 1392 192
rect 1440 166 1470 192
rect 1555 177 1571 205
rect 1518 171 1571 177
rect 1605 171 1695 205
rect 986 131 1016 147
rect 1064 131 1094 147
rect 1518 147 1695 171
rect 1518 132 1548 147
rect 1590 132 1620 147
rect 84 75 114 101
rect 162 75 192 101
rect 248 75 278 101
rect 320 75 350 101
rect 406 75 436 101
rect 478 75 508 101
rect 696 21 726 47
rect 782 21 812 47
rect 860 21 890 47
rect 986 21 1016 47
rect 1064 21 1094 47
rect 1518 22 1548 48
rect 1590 22 1620 48
<< polycont >>
rect 61 291 95 325
rect 61 223 95 257
rect 264 294 298 328
rect 372 294 406 328
rect 590 294 624 328
rect 762 315 796 349
rect 881 323 915 357
rect 1081 323 1115 357
rect 1567 279 1601 313
rect 1003 169 1037 203
rect 1571 171 1605 205
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 309 627 375 649
rect 309 593 325 627
rect 359 593 375 627
rect 411 592 653 609
rect 89 564 155 580
rect 89 530 105 564
rect 139 557 155 564
rect 411 558 603 592
rect 637 558 653 592
rect 411 557 653 558
rect 905 589 971 649
rect 139 530 445 557
rect 905 555 921 589
rect 955 555 971 589
rect 905 536 971 555
rect 1018 593 1084 609
rect 1018 559 1034 593
rect 1068 559 1084 593
rect 1273 603 1339 649
rect 1273 569 1289 603
rect 1323 569 1339 603
rect 1273 568 1339 569
rect 1501 618 1567 649
rect 1501 584 1517 618
rect 1551 584 1567 618
rect 1501 568 1567 584
rect 1623 597 1703 613
rect 89 523 445 530
rect 1018 532 1084 559
rect 1623 563 1639 597
rect 1673 563 1703 597
rect 89 495 181 523
rect 89 461 105 495
rect 139 461 181 495
rect 481 487 829 521
rect 1018 516 1585 532
rect 1018 500 1034 516
rect 89 427 181 461
rect 356 453 515 487
rect 89 393 105 427
rect 139 393 181 427
rect 89 377 181 393
rect 25 325 111 341
rect 25 291 61 325
rect 95 291 111 325
rect 25 257 111 291
rect 25 223 61 257
rect 95 223 111 257
rect 25 207 111 223
rect 147 242 181 377
rect 217 328 314 430
rect 217 294 264 328
rect 298 294 314 328
rect 217 278 314 294
rect 356 328 422 453
rect 676 417 709 451
rect 743 417 759 451
rect 356 294 372 328
rect 406 294 422 328
rect 356 278 422 294
rect 458 401 524 417
rect 458 367 474 401
rect 508 367 524 401
rect 458 344 524 367
rect 676 401 759 417
rect 458 328 640 344
rect 458 294 590 328
rect 624 294 640 328
rect 458 278 640 294
rect 147 208 481 242
rect 23 151 89 171
rect 23 117 39 151
rect 73 117 89 151
rect 23 17 89 117
rect 147 160 253 208
rect 147 126 203 160
rect 237 126 253 160
rect 147 97 253 126
rect 345 151 411 172
rect 345 117 361 151
rect 395 117 411 151
rect 345 17 411 117
rect 447 87 481 208
rect 560 189 594 278
rect 519 173 594 189
rect 676 210 710 401
rect 795 365 829 487
rect 746 349 829 365
rect 746 315 762 349
rect 796 315 829 349
rect 865 482 1034 500
rect 1068 498 1585 516
rect 1068 482 1084 498
rect 865 466 1084 482
rect 865 357 931 466
rect 865 323 881 357
rect 915 323 931 357
rect 865 316 931 323
rect 985 357 1131 430
rect 985 323 1081 357
rect 1115 323 1131 357
rect 985 316 1131 323
rect 1167 428 1183 462
rect 1217 428 1233 462
rect 1167 412 1233 428
rect 746 299 829 315
rect 795 280 829 299
rect 1167 280 1209 412
rect 1269 350 1303 498
rect 1379 428 1395 462
rect 1429 446 1445 462
rect 1429 428 1515 446
rect 1379 412 1515 428
rect 795 251 1209 280
rect 795 246 1159 251
rect 1143 217 1159 246
rect 1193 217 1209 251
rect 676 203 1053 210
rect 676 176 1003 203
rect 519 139 535 173
rect 569 139 594 173
rect 519 123 594 139
rect 635 111 701 135
rect 635 87 651 111
rect 447 77 651 87
rect 685 77 701 111
rect 447 53 701 77
rect 737 111 787 176
rect 987 169 1003 176
rect 1037 169 1053 203
rect 1143 188 1209 217
rect 1245 316 1303 350
rect 987 153 1053 169
rect 1245 135 1279 316
rect 771 77 787 111
rect 737 53 787 77
rect 885 106 951 135
rect 885 72 901 106
rect 935 72 951 106
rect 885 17 951 72
rect 1089 111 1279 135
rect 1089 77 1105 111
rect 1139 101 1279 111
rect 1317 251 1367 280
rect 1351 217 1367 251
rect 1139 77 1155 101
rect 1089 53 1155 77
rect 1317 17 1367 217
rect 1465 251 1515 412
rect 1551 329 1585 498
rect 1623 462 1703 563
rect 1623 428 1639 462
rect 1673 428 1703 462
rect 1623 412 1703 428
rect 1551 313 1617 329
rect 1551 279 1567 313
rect 1601 279 1617 313
rect 1551 263 1617 279
rect 1465 217 1481 251
rect 1515 217 1621 221
rect 1465 205 1621 217
rect 1465 187 1571 205
rect 1555 171 1571 187
rect 1605 171 1621 205
rect 1555 155 1621 171
rect 1453 107 1519 136
rect 1657 119 1703 412
rect 1453 73 1469 107
rect 1503 73 1519 107
rect 1453 17 1519 73
rect 1615 103 1703 119
rect 1615 69 1631 103
rect 1665 69 1703 103
rect 1615 53 1703 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdlclkp_lp
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1087 390 1121 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 1663 94 1697 128 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1663 168 1697 202 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1663 390 1697 424 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1663 464 1697 498 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1450618
string GDS_START 1438602
<< end >>
