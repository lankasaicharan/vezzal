magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 17 49 765 167
rect 0 0 768 49
<< scnmos >>
rect 100 57 130 141
rect 178 57 208 141
rect 264 57 294 141
rect 336 57 366 141
rect 422 57 452 141
rect 494 57 524 141
rect 580 57 610 141
rect 652 57 682 141
<< scpmoshvt >>
rect 86 409 136 609
rect 202 409 252 609
rect 308 409 358 609
rect 414 409 464 609
rect 632 409 682 609
<< ndiff >>
rect 43 116 100 141
rect 43 82 55 116
rect 89 82 100 116
rect 43 57 100 82
rect 130 57 178 141
rect 208 107 264 141
rect 208 73 219 107
rect 253 73 264 107
rect 208 57 264 73
rect 294 57 336 141
rect 366 116 422 141
rect 366 82 377 116
rect 411 82 422 116
rect 366 57 422 82
rect 452 57 494 141
rect 524 107 580 141
rect 524 73 535 107
rect 569 73 580 107
rect 524 57 580 73
rect 610 57 652 141
rect 682 116 739 141
rect 682 82 693 116
rect 727 82 739 116
rect 682 57 739 82
<< pdiff >>
rect 29 597 86 609
rect 29 563 41 597
rect 75 563 86 597
rect 29 526 86 563
rect 29 492 41 526
rect 75 492 86 526
rect 29 455 86 492
rect 29 421 41 455
rect 75 421 86 455
rect 29 409 86 421
rect 136 597 202 609
rect 136 563 147 597
rect 181 563 202 597
rect 136 524 202 563
rect 136 490 147 524
rect 181 490 202 524
rect 136 409 202 490
rect 252 597 308 609
rect 252 563 263 597
rect 297 563 308 597
rect 252 526 308 563
rect 252 492 263 526
rect 297 492 308 526
rect 252 455 308 492
rect 252 421 263 455
rect 297 421 308 455
rect 252 409 308 421
rect 358 409 414 609
rect 464 597 521 609
rect 464 563 475 597
rect 509 563 521 597
rect 464 526 521 563
rect 464 492 475 526
rect 509 492 521 526
rect 464 455 521 492
rect 464 421 475 455
rect 509 421 521 455
rect 464 409 521 421
rect 575 597 632 609
rect 575 563 587 597
rect 621 563 632 597
rect 575 524 632 563
rect 575 490 587 524
rect 621 490 632 524
rect 575 409 632 490
rect 682 597 739 609
rect 682 563 693 597
rect 727 563 739 597
rect 682 526 739 563
rect 682 492 693 526
rect 727 492 739 526
rect 682 455 739 492
rect 682 421 693 455
rect 727 421 739 455
rect 682 409 739 421
<< ndiffc >>
rect 55 82 89 116
rect 219 73 253 107
rect 377 82 411 116
rect 535 73 569 107
rect 693 82 727 116
<< pdiffc >>
rect 41 563 75 597
rect 41 492 75 526
rect 41 421 75 455
rect 147 563 181 597
rect 147 490 181 524
rect 263 563 297 597
rect 263 492 297 526
rect 263 421 297 455
rect 475 563 509 597
rect 475 492 509 526
rect 475 421 509 455
rect 587 563 621 597
rect 587 490 621 524
rect 693 563 727 597
rect 693 492 727 526
rect 693 421 727 455
<< poly >>
rect 86 609 136 635
rect 202 609 252 635
rect 308 609 358 635
rect 414 609 464 635
rect 632 609 682 635
rect 86 325 136 409
rect 202 368 252 409
rect 308 368 358 409
rect 414 368 464 409
rect 178 352 252 368
rect 31 309 130 325
rect 31 275 47 309
rect 81 275 130 309
rect 31 241 130 275
rect 31 207 47 241
rect 81 207 130 241
rect 31 191 130 207
rect 100 141 130 191
rect 178 318 202 352
rect 236 318 252 352
rect 178 284 252 318
rect 178 250 202 284
rect 236 250 252 284
rect 178 234 252 250
rect 300 352 366 368
rect 300 318 316 352
rect 350 318 366 352
rect 300 284 366 318
rect 300 250 316 284
rect 350 250 366 284
rect 178 141 208 234
rect 300 186 366 250
rect 414 352 480 368
rect 414 318 430 352
rect 464 318 480 352
rect 414 284 480 318
rect 632 298 682 409
rect 414 250 430 284
rect 464 264 480 284
rect 575 282 682 298
rect 464 250 524 264
rect 414 234 524 250
rect 264 156 366 186
rect 264 141 294 156
rect 336 141 366 156
rect 422 141 452 234
rect 494 141 524 234
rect 575 248 591 282
rect 625 248 682 282
rect 575 214 682 248
rect 575 180 591 214
rect 625 180 682 214
rect 575 164 682 180
rect 580 141 610 164
rect 652 141 682 164
rect 100 31 130 57
rect 178 31 208 57
rect 264 31 294 57
rect 336 31 366 57
rect 422 31 452 57
rect 494 31 524 57
rect 580 31 610 57
rect 652 31 682 57
<< polycont >>
rect 47 275 81 309
rect 47 207 81 241
rect 202 318 236 352
rect 202 250 236 284
rect 316 318 350 352
rect 316 250 350 284
rect 430 318 464 352
rect 430 250 464 284
rect 591 248 625 282
rect 591 180 625 214
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 25 597 91 613
rect 25 563 41 597
rect 75 563 91 597
rect 25 526 91 563
rect 25 492 41 526
rect 75 492 91 526
rect 25 455 91 492
rect 131 597 197 649
rect 131 563 147 597
rect 181 563 197 597
rect 131 524 197 563
rect 131 490 147 524
rect 181 490 197 524
rect 131 474 197 490
rect 247 597 313 613
rect 247 563 263 597
rect 297 563 313 597
rect 247 526 313 563
rect 247 492 263 526
rect 297 492 313 526
rect 25 421 41 455
rect 75 438 91 455
rect 247 455 313 492
rect 247 438 263 455
rect 75 421 263 438
rect 297 421 313 455
rect 25 404 313 421
rect 459 597 525 613
rect 459 563 475 597
rect 509 563 525 597
rect 459 526 525 563
rect 459 492 475 526
rect 509 492 525 526
rect 459 455 525 492
rect 571 597 637 649
rect 571 563 587 597
rect 621 563 637 597
rect 571 524 637 563
rect 571 490 587 524
rect 621 490 637 524
rect 571 474 637 490
rect 677 597 743 613
rect 677 563 693 597
rect 727 563 743 597
rect 677 526 743 563
rect 677 492 693 526
rect 727 492 743 526
rect 459 421 475 455
rect 509 438 525 455
rect 677 455 743 492
rect 509 421 609 438
rect 459 404 609 421
rect 25 309 97 356
rect 25 275 47 309
rect 81 275 97 309
rect 25 241 97 275
rect 25 207 47 241
rect 81 207 97 241
rect 186 352 263 368
rect 186 318 202 352
rect 236 318 263 352
rect 186 284 263 318
rect 186 250 202 284
rect 236 250 263 284
rect 186 234 263 250
rect 300 352 366 368
rect 300 318 316 352
rect 350 318 366 352
rect 300 284 366 318
rect 300 250 316 284
rect 350 250 366 284
rect 300 234 366 250
rect 409 352 480 368
rect 409 318 430 352
rect 464 318 480 352
rect 409 284 480 318
rect 409 250 430 284
rect 464 250 480 284
rect 409 234 480 250
rect 575 298 609 404
rect 677 421 693 455
rect 727 421 743 455
rect 575 282 641 298
rect 575 248 591 282
rect 625 248 641 282
rect 25 191 97 207
rect 575 214 641 248
rect 575 198 591 214
rect 133 180 591 198
rect 625 180 641 214
rect 133 164 641 180
rect 133 145 167 164
rect 39 116 167 145
rect 39 82 55 116
rect 89 111 167 116
rect 89 82 105 111
rect 39 53 105 82
rect 203 107 269 128
rect 203 73 219 107
rect 253 73 269 107
rect 203 17 269 73
rect 361 116 427 164
rect 361 82 377 116
rect 411 82 427 116
rect 361 53 427 82
rect 519 107 585 128
rect 519 73 535 107
rect 569 73 585 107
rect 519 17 585 73
rect 677 116 743 421
rect 677 82 693 116
rect 727 82 743 116
rect 677 53 743 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a211o_lp
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1976512
string GDS_START 1968624
<< end >>
