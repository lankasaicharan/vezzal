magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2034 1852
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 11 21 669 203
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 465 47 495 177
rect 559 47 589 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
<< ndiff >>
rect 37 93 89 177
rect 37 59 45 93
rect 79 59 89 93
rect 37 47 89 59
rect 119 101 183 177
rect 119 67 129 101
rect 163 67 183 101
rect 119 47 183 67
rect 213 93 277 177
rect 213 59 223 93
rect 257 59 277 93
rect 213 47 277 59
rect 307 101 371 177
rect 307 67 317 101
rect 351 67 371 101
rect 307 47 371 67
rect 401 93 465 177
rect 401 59 411 93
rect 445 59 465 93
rect 401 47 465 59
rect 495 101 559 177
rect 495 67 505 101
rect 539 67 559 101
rect 495 47 559 67
rect 589 94 643 177
rect 589 60 599 94
rect 633 60 643 94
rect 589 47 643 60
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 349 551 383
rect 493 315 505 349
rect 539 315 551 349
rect 493 297 551 315
rect 587 485 643 497
rect 587 451 599 485
rect 633 451 643 485
rect 587 297 643 451
<< ndiffc >>
rect 45 59 79 93
rect 129 67 163 101
rect 223 59 257 93
rect 317 67 351 101
rect 411 59 445 93
rect 505 67 539 101
rect 599 60 633 94
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 505 451 539 485
rect 505 383 539 417
rect 505 315 539 349
rect 599 451 633 485
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 57 249 589 265
rect 57 215 90 249
rect 124 215 192 249
rect 226 215 291 249
rect 325 215 385 249
rect 419 215 479 249
rect 513 215 589 249
rect 57 199 589 215
rect 89 177 119 199
rect 183 177 213 199
rect 277 177 307 199
rect 371 177 401 199
rect 465 177 495 199
rect 559 177 589 199
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 465 21 495 47
rect 559 21 589 47
<< polycont >>
rect 90 215 124 249
rect 192 215 226 249
rect 291 215 325 249
rect 385 215 419 249
rect 479 215 513 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 35 485 69 527
rect 35 417 69 451
rect 35 349 69 383
rect 35 299 69 315
rect 103 485 179 493
rect 103 451 129 485
rect 163 451 179 485
rect 103 417 179 451
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 223 485 257 527
rect 223 417 257 451
rect 223 367 257 383
rect 291 485 367 493
rect 291 451 317 485
rect 351 451 367 485
rect 291 417 367 451
rect 291 383 317 417
rect 351 383 367 417
rect 103 315 129 349
rect 163 333 179 349
rect 291 349 367 383
rect 411 485 445 527
rect 411 417 445 451
rect 411 367 445 383
rect 479 485 555 493
rect 479 451 505 485
rect 539 451 555 485
rect 479 417 555 451
rect 599 485 633 527
rect 599 435 633 451
rect 479 383 505 417
rect 539 383 555 417
rect 291 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 479 349 555 383
rect 479 333 505 349
rect 351 315 505 333
rect 539 337 555 349
rect 539 315 653 337
rect 103 299 653 315
rect 57 249 539 265
rect 57 215 90 249
rect 124 215 192 249
rect 226 215 291 249
rect 325 215 385 249
rect 419 215 479 249
rect 513 215 539 249
rect 573 181 653 299
rect 129 145 653 181
rect 26 93 79 109
rect 26 59 45 93
rect 26 17 79 59
rect 129 101 163 145
rect 129 51 163 67
rect 223 93 257 109
rect 223 17 257 59
rect 317 101 351 145
rect 317 51 351 67
rect 411 93 445 109
rect 411 17 445 59
rect 505 101 539 145
rect 505 51 539 67
rect 573 94 633 110
rect 573 60 599 94
rect 573 17 633 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 599 153 633 187 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 599 221 633 255 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 599 289 633 323 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 82 221 116 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 280 238 280 238 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel locali s 372 238 372 238 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel locali s 464 238 464 238 0 FreeSans 340 0 0 0 A
port 1 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional
rlabel comment s 3 0 3 0 4 inv_6
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2135642
string GDS_START 2129276
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
