magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4178 1975
<< nwell >>
rect -38 331 2918 704
<< pwell >>
rect 1624 229 1745 282
rect 2601 242 2875 250
rect 650 222 1745 229
rect 650 191 1860 222
rect 1 178 1860 191
rect 2220 178 2875 242
rect 1 49 2875 178
rect 0 0 2880 49
<< scnmos >>
rect 80 81 110 165
rect 293 81 323 165
rect 365 81 395 165
rect 456 81 486 165
rect 545 81 575 165
rect 631 81 661 165
rect 729 119 759 203
rect 815 119 845 203
rect 925 119 955 203
rect 1011 119 1041 203
rect 1233 119 1263 203
rect 1319 119 1349 203
rect 1391 119 1421 203
rect 1463 119 1493 203
rect 1605 68 1635 196
rect 1749 68 1779 196
rect 1849 68 1879 152
rect 1951 68 1981 152
rect 2037 68 2067 152
rect 2109 68 2139 152
rect 2299 48 2329 216
rect 2385 48 2415 216
rect 2490 48 2520 132
rect 2680 56 2710 224
rect 2766 56 2796 224
<< scpmoshvt >>
rect 171 489 201 617
rect 257 489 287 617
rect 329 489 359 617
rect 415 489 445 617
rect 509 489 539 617
rect 617 489 647 617
rect 818 367 848 619
rect 904 367 934 619
rect 1132 463 1162 547
rect 1218 463 1248 547
rect 1290 463 1320 547
rect 1422 463 1452 547
rect 1625 379 1655 547
rect 1740 412 1770 580
rect 1855 496 1885 580
rect 1963 496 1993 580
rect 2088 496 2118 580
rect 2174 496 2204 580
rect 2295 367 2325 619
rect 2381 367 2411 619
rect 2486 367 2516 495
rect 2680 367 2710 619
rect 2766 367 2796 619
<< ndiff >>
rect 27 143 80 165
rect 27 109 35 143
rect 69 109 80 143
rect 27 81 80 109
rect 110 137 163 165
rect 110 103 121 137
rect 155 103 163 137
rect 110 81 163 103
rect 676 165 729 203
rect 240 137 293 165
rect 240 103 248 137
rect 282 103 293 137
rect 240 81 293 103
rect 323 81 365 165
rect 395 157 456 165
rect 395 123 411 157
rect 445 123 456 157
rect 395 81 456 123
rect 486 81 545 165
rect 575 123 631 165
rect 575 89 586 123
rect 620 89 631 123
rect 575 81 631 89
rect 661 140 729 165
rect 661 106 672 140
rect 706 119 729 140
rect 759 181 815 203
rect 759 147 770 181
rect 804 147 815 181
rect 759 119 815 147
rect 845 138 925 203
rect 845 119 868 138
rect 706 106 714 119
rect 661 81 714 106
rect 860 104 868 119
rect 902 119 925 138
rect 955 174 1011 203
rect 955 140 966 174
rect 1000 140 1011 174
rect 955 119 1011 140
rect 1041 165 1094 203
rect 1041 131 1052 165
rect 1086 131 1094 165
rect 1041 119 1094 131
rect 1180 180 1233 203
rect 1180 146 1188 180
rect 1222 146 1233 180
rect 1180 119 1233 146
rect 1263 172 1319 203
rect 1263 138 1274 172
rect 1308 138 1319 172
rect 1263 119 1319 138
rect 1349 119 1391 203
rect 1421 119 1463 203
rect 1493 196 1590 203
rect 1650 246 1719 256
rect 1650 212 1662 246
rect 1696 212 1719 246
rect 1650 196 1719 212
rect 1493 119 1605 196
rect 902 104 910 119
rect 860 88 910 104
rect 1518 110 1605 119
rect 1518 76 1535 110
rect 1569 76 1605 110
rect 1518 68 1605 76
rect 1635 68 1749 196
rect 1779 152 1834 196
rect 2246 164 2299 216
rect 1779 114 1849 152
rect 1779 80 1804 114
rect 1838 80 1849 114
rect 1779 68 1849 80
rect 1879 68 1951 152
rect 1981 118 2037 152
rect 1981 84 1992 118
rect 2026 84 2037 118
rect 1981 68 2037 84
rect 2067 68 2109 152
rect 2139 127 2192 152
rect 2139 93 2150 127
rect 2184 93 2192 127
rect 2139 68 2192 93
rect 2246 130 2254 164
rect 2288 130 2299 164
rect 2246 94 2299 130
rect 2246 60 2254 94
rect 2288 60 2299 94
rect 2246 48 2299 60
rect 2329 204 2385 216
rect 2329 170 2340 204
rect 2374 170 2385 204
rect 2329 101 2385 170
rect 2329 67 2340 101
rect 2374 67 2385 101
rect 2329 48 2385 67
rect 2415 203 2468 216
rect 2415 169 2426 203
rect 2460 169 2468 203
rect 2415 132 2468 169
rect 2627 196 2680 224
rect 2627 162 2635 196
rect 2669 162 2680 196
rect 2415 94 2490 132
rect 2415 60 2445 94
rect 2479 60 2490 94
rect 2415 48 2490 60
rect 2520 107 2573 132
rect 2520 73 2531 107
rect 2565 73 2573 107
rect 2520 48 2573 73
rect 2627 102 2680 162
rect 2627 68 2635 102
rect 2669 68 2680 102
rect 2627 56 2680 68
rect 2710 212 2766 224
rect 2710 178 2721 212
rect 2755 178 2766 212
rect 2710 101 2766 178
rect 2710 67 2721 101
rect 2755 67 2766 101
rect 2710 56 2766 67
rect 2796 212 2849 224
rect 2796 178 2807 212
rect 2841 178 2849 212
rect 2796 102 2849 178
rect 2796 68 2807 102
rect 2841 68 2849 102
rect 2796 56 2849 68
<< pdiff >>
rect 118 604 171 617
rect 118 570 126 604
rect 160 570 171 604
rect 118 535 171 570
rect 118 501 126 535
rect 160 501 171 535
rect 118 489 171 501
rect 201 605 257 617
rect 201 571 212 605
rect 246 571 257 605
rect 201 537 257 571
rect 201 503 212 537
rect 246 503 257 537
rect 201 489 257 503
rect 287 489 329 617
rect 359 604 415 617
rect 359 570 370 604
rect 404 570 415 604
rect 359 535 415 570
rect 359 501 370 535
rect 404 501 415 535
rect 359 489 415 501
rect 445 489 509 617
rect 539 605 617 617
rect 539 571 550 605
rect 584 571 617 605
rect 539 489 617 571
rect 647 604 700 617
rect 647 570 658 604
rect 692 570 700 604
rect 647 535 700 570
rect 647 501 658 535
rect 692 501 700 535
rect 647 489 700 501
rect 765 447 818 619
rect 765 413 773 447
rect 807 413 818 447
rect 765 367 818 413
rect 848 603 904 619
rect 848 569 859 603
rect 893 569 904 603
rect 848 367 904 569
rect 934 447 987 619
rect 934 413 945 447
rect 979 413 987 447
rect 934 367 987 413
rect 1335 570 1407 583
rect 2234 607 2295 619
rect 2234 580 2246 607
rect 1335 547 1354 570
rect 1074 515 1132 547
rect 1074 481 1087 515
rect 1121 481 1132 515
rect 1074 463 1132 481
rect 1162 523 1218 547
rect 1162 489 1173 523
rect 1207 489 1218 523
rect 1162 463 1218 489
rect 1248 463 1290 547
rect 1320 536 1354 547
rect 1388 547 1407 570
rect 1670 547 1740 580
rect 1388 536 1422 547
rect 1320 463 1422 536
rect 1452 523 1505 547
rect 1452 489 1463 523
rect 1497 489 1505 523
rect 1452 463 1505 489
rect 1563 535 1625 547
rect 1563 501 1571 535
rect 1605 501 1625 535
rect 1563 467 1625 501
rect 1563 433 1571 467
rect 1605 433 1625 467
rect 1563 379 1625 433
rect 1655 539 1740 547
rect 1655 505 1680 539
rect 1714 505 1740 539
rect 1655 471 1740 505
rect 1655 437 1666 471
rect 1700 437 1740 471
rect 1655 412 1740 437
rect 1770 563 1855 580
rect 1770 529 1781 563
rect 1815 529 1855 563
rect 1770 496 1855 529
rect 1885 496 1963 580
rect 1993 555 2088 580
rect 1993 521 2021 555
rect 2055 521 2088 555
rect 1993 496 2088 521
rect 2118 555 2174 580
rect 2118 521 2129 555
rect 2163 521 2174 555
rect 2118 496 2174 521
rect 2204 573 2246 580
rect 2280 573 2295 607
rect 2204 496 2295 573
rect 1770 471 1823 496
rect 1770 437 1781 471
rect 1815 437 1823 471
rect 1770 412 1823 437
rect 1655 379 1705 412
rect 2234 490 2295 496
rect 2234 456 2246 490
rect 2280 456 2295 490
rect 2234 367 2295 456
rect 2325 599 2381 619
rect 2325 565 2336 599
rect 2370 565 2381 599
rect 2325 498 2381 565
rect 2325 464 2336 498
rect 2370 464 2381 498
rect 2325 409 2381 464
rect 2325 375 2336 409
rect 2370 375 2381 409
rect 2325 367 2381 375
rect 2411 607 2464 619
rect 2411 573 2422 607
rect 2456 573 2464 607
rect 2411 509 2464 573
rect 2627 607 2680 619
rect 2627 573 2635 607
rect 2669 573 2680 607
rect 2411 475 2422 509
rect 2456 495 2464 509
rect 2627 510 2680 573
rect 2456 475 2486 495
rect 2411 409 2486 475
rect 2411 375 2431 409
rect 2465 375 2486 409
rect 2411 367 2486 375
rect 2516 483 2569 495
rect 2516 449 2527 483
rect 2561 449 2569 483
rect 2516 413 2569 449
rect 2516 379 2527 413
rect 2561 379 2569 413
rect 2516 367 2569 379
rect 2627 476 2635 510
rect 2669 476 2680 510
rect 2627 413 2680 476
rect 2627 379 2635 413
rect 2669 379 2680 413
rect 2627 367 2680 379
rect 2710 599 2766 619
rect 2710 565 2721 599
rect 2755 565 2766 599
rect 2710 495 2766 565
rect 2710 461 2721 495
rect 2755 461 2766 495
rect 2710 413 2766 461
rect 2710 379 2721 413
rect 2755 379 2766 413
rect 2710 367 2766 379
rect 2796 607 2849 619
rect 2796 573 2807 607
rect 2841 573 2849 607
rect 2796 510 2849 573
rect 2796 476 2807 510
rect 2841 476 2849 510
rect 2796 413 2849 476
rect 2796 379 2807 413
rect 2841 379 2849 413
rect 2796 367 2849 379
<< ndiffc >>
rect 35 109 69 143
rect 121 103 155 137
rect 248 103 282 137
rect 411 123 445 157
rect 586 89 620 123
rect 672 106 706 140
rect 770 147 804 181
rect 868 104 902 138
rect 966 140 1000 174
rect 1052 131 1086 165
rect 1188 146 1222 180
rect 1274 138 1308 172
rect 1662 212 1696 246
rect 1535 76 1569 110
rect 1804 80 1838 114
rect 1992 84 2026 118
rect 2150 93 2184 127
rect 2254 130 2288 164
rect 2254 60 2288 94
rect 2340 170 2374 204
rect 2340 67 2374 101
rect 2426 169 2460 203
rect 2635 162 2669 196
rect 2445 60 2479 94
rect 2531 73 2565 107
rect 2635 68 2669 102
rect 2721 178 2755 212
rect 2721 67 2755 101
rect 2807 178 2841 212
rect 2807 68 2841 102
<< pdiffc >>
rect 126 570 160 604
rect 126 501 160 535
rect 212 571 246 605
rect 212 503 246 537
rect 370 570 404 604
rect 370 501 404 535
rect 550 571 584 605
rect 658 570 692 604
rect 658 501 692 535
rect 773 413 807 447
rect 859 569 893 603
rect 945 413 979 447
rect 1087 481 1121 515
rect 1173 489 1207 523
rect 1354 536 1388 570
rect 1463 489 1497 523
rect 1571 501 1605 535
rect 1571 433 1605 467
rect 1680 505 1714 539
rect 1666 437 1700 471
rect 1781 529 1815 563
rect 2021 521 2055 555
rect 2129 521 2163 555
rect 2246 573 2280 607
rect 1781 437 1815 471
rect 2246 456 2280 490
rect 2336 565 2370 599
rect 2336 464 2370 498
rect 2336 375 2370 409
rect 2422 573 2456 607
rect 2635 573 2669 607
rect 2422 475 2456 509
rect 2431 375 2465 409
rect 2527 449 2561 483
rect 2527 379 2561 413
rect 2635 476 2669 510
rect 2635 379 2669 413
rect 2721 565 2755 599
rect 2721 461 2755 495
rect 2721 379 2755 413
rect 2807 573 2841 607
rect 2807 476 2841 510
rect 2807 379 2841 413
<< poly >>
rect 171 617 201 643
rect 257 617 287 643
rect 329 617 359 643
rect 415 617 445 643
rect 509 617 539 643
rect 617 617 647 643
rect 818 619 848 645
rect 904 619 934 645
rect 171 467 201 489
rect 257 467 287 489
rect 171 437 287 467
rect 171 369 201 437
rect 80 353 261 369
rect 80 319 143 353
rect 177 319 211 353
rect 245 319 261 353
rect 80 303 261 319
rect 80 165 110 303
rect 329 299 359 489
rect 415 455 445 489
rect 509 455 539 489
rect 401 439 467 455
rect 401 405 417 439
rect 451 405 467 439
rect 401 389 467 405
rect 509 439 575 455
rect 509 405 525 439
rect 559 405 575 439
rect 509 371 575 405
rect 617 440 647 489
rect 617 424 731 440
rect 617 390 681 424
rect 715 390 731 424
rect 617 374 731 390
rect 509 337 525 371
rect 559 337 575 371
rect 509 321 575 337
rect 309 283 375 299
rect 178 237 251 253
rect 178 203 201 237
rect 235 203 251 237
rect 309 249 325 283
rect 359 263 375 283
rect 437 263 503 279
rect 359 249 395 263
rect 309 233 395 249
rect 178 187 251 203
rect 80 55 110 81
rect 178 59 225 187
rect 293 165 323 191
rect 365 165 395 233
rect 437 229 453 263
rect 487 229 503 263
rect 437 213 503 229
rect 456 165 486 213
rect 545 165 575 321
rect 631 165 661 374
rect 1002 615 1770 645
rect 2295 619 2325 645
rect 2381 619 2411 645
rect 2680 619 2710 645
rect 2766 619 2796 645
rect 818 322 848 367
rect 729 306 848 322
rect 729 272 783 306
rect 817 272 848 306
rect 729 218 848 272
rect 904 322 934 367
rect 1002 322 1032 615
rect 1132 547 1162 573
rect 1218 547 1248 615
rect 1290 547 1320 573
rect 1740 580 1770 615
rect 1855 580 1885 606
rect 1963 580 1993 606
rect 2088 580 2118 606
rect 2174 580 2204 606
rect 1422 547 1452 573
rect 1625 547 1655 573
rect 1132 356 1162 463
rect 1218 437 1248 463
rect 1290 431 1320 463
rect 1422 448 1452 463
rect 1290 415 1380 431
rect 1422 429 1533 448
rect 1426 426 1533 429
rect 1431 422 1533 426
rect 1437 418 1533 422
rect 1290 381 1324 415
rect 1358 398 1380 415
rect 1463 415 1533 418
rect 1358 392 1388 398
rect 1358 383 1400 392
rect 1358 381 1411 383
rect 1290 379 1411 381
rect 1463 381 1481 415
rect 1515 381 1533 415
rect 1290 365 1421 379
rect 1362 360 1421 365
rect 904 306 1032 322
rect 904 272 920 306
rect 954 272 1032 306
rect 1074 340 1162 356
rect 1370 353 1421 360
rect 1074 306 1090 340
rect 1124 320 1162 340
rect 1384 336 1421 353
rect 1124 318 1311 320
rect 1124 311 1319 318
rect 1124 306 1349 311
rect 1074 290 1349 306
rect 1284 287 1349 290
rect 1293 279 1349 287
rect 904 256 1032 272
rect 925 248 1032 256
rect 925 218 1263 248
rect 729 203 759 218
rect 815 203 845 218
rect 925 203 955 218
rect 1011 203 1041 218
rect 1233 203 1263 218
rect 1319 203 1349 279
rect 1391 203 1421 336
rect 1463 364 1533 381
rect 1855 464 1885 496
rect 1855 448 1921 464
rect 1855 414 1871 448
rect 1905 414 1921 448
rect 1463 203 1493 364
rect 1625 347 1655 379
rect 1577 331 1655 347
rect 1577 297 1593 331
rect 1627 297 1655 331
rect 1740 356 1770 412
rect 1855 398 1921 414
rect 1740 326 1879 356
rect 1577 281 1655 297
rect 729 93 759 119
rect 815 93 845 119
rect 1605 196 1635 281
rect 1741 268 1807 284
rect 1741 234 1757 268
rect 1791 234 1807 268
rect 1741 218 1807 234
rect 1749 196 1779 218
rect 925 93 955 119
rect 1011 93 1041 119
rect 1233 93 1263 119
rect 1319 93 1349 119
rect 1391 93 1421 119
rect 293 59 323 81
rect 178 29 323 59
rect 365 55 395 81
rect 456 55 486 81
rect 545 55 575 81
rect 631 51 661 81
rect 1463 51 1493 119
rect 1849 152 1879 326
rect 1963 240 1993 496
rect 2088 464 2118 496
rect 2035 448 2118 464
rect 2035 414 2051 448
rect 2085 414 2118 448
rect 2035 398 2118 414
rect 1923 224 1993 240
rect 1923 190 1939 224
rect 1973 190 1993 224
rect 1923 174 1993 190
rect 1951 152 1981 174
rect 2037 152 2067 398
rect 2174 356 2204 496
rect 2486 495 2516 521
rect 2109 336 2204 356
rect 2109 302 2125 336
rect 2159 306 2204 336
rect 2295 306 2325 367
rect 2381 306 2411 367
rect 2486 306 2516 367
rect 2680 312 2710 367
rect 2766 312 2796 367
rect 2159 302 2520 306
rect 2109 276 2520 302
rect 2109 152 2139 276
rect 2299 216 2329 276
rect 2385 216 2415 276
rect 631 21 1493 51
rect 1605 42 1635 68
rect 1749 42 1779 68
rect 1849 42 1879 68
rect 1951 42 1981 68
rect 2037 42 2067 68
rect 2109 42 2139 68
rect 2490 132 2520 276
rect 2631 296 2796 312
rect 2631 262 2647 296
rect 2681 262 2796 296
rect 2631 246 2796 262
rect 2680 224 2710 246
rect 2766 224 2796 246
rect 2299 22 2329 48
rect 2385 22 2415 48
rect 2490 22 2520 48
rect 2680 30 2710 56
rect 2766 30 2796 56
<< polycont >>
rect 143 319 177 353
rect 211 319 245 353
rect 417 405 451 439
rect 525 405 559 439
rect 681 390 715 424
rect 525 337 559 371
rect 201 203 235 237
rect 325 249 359 283
rect 453 229 487 263
rect 783 272 817 306
rect 1324 381 1358 415
rect 1481 381 1515 415
rect 920 272 954 306
rect 1090 306 1124 340
rect 1871 414 1905 448
rect 1593 297 1627 331
rect 1757 234 1791 268
rect 2051 414 2085 448
rect 1939 190 1973 224
rect 2125 302 2159 336
rect 2647 262 2681 296
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 106 604 176 615
rect 106 570 126 604
rect 160 570 176 604
rect 106 535 176 570
rect 106 501 126 535
rect 160 501 176 535
rect 106 453 176 501
rect 210 605 262 649
rect 210 571 212 605
rect 246 571 262 605
rect 210 537 262 571
rect 210 503 212 537
rect 246 503 262 537
rect 210 487 262 503
rect 354 604 420 615
rect 354 570 370 604
rect 404 570 420 604
rect 354 535 420 570
rect 534 605 600 649
rect 534 571 550 605
rect 584 571 600 605
rect 534 567 600 571
rect 642 604 708 615
rect 642 570 658 604
rect 692 570 708 604
rect 354 501 370 535
rect 404 531 420 535
rect 642 535 708 570
rect 843 603 909 649
rect 843 569 859 603
rect 893 569 909 603
rect 843 565 909 569
rect 1338 570 1404 649
rect 642 531 658 535
rect 404 501 658 531
rect 692 531 708 535
rect 692 515 1125 531
rect 692 501 1087 515
rect 354 497 1087 501
rect 354 489 629 497
rect 106 439 467 453
rect 19 405 417 439
rect 451 405 467 439
rect 19 403 467 405
rect 505 439 561 455
rect 505 405 525 439
rect 559 405 561 439
rect 19 253 73 403
rect 505 371 561 405
rect 107 353 471 369
rect 107 319 143 353
rect 177 319 211 353
rect 245 335 471 353
rect 245 319 269 335
rect 107 303 269 319
rect 314 283 361 299
rect 19 237 251 253
rect 19 203 201 237
rect 235 203 251 237
rect 19 187 251 203
rect 314 249 325 283
rect 359 249 361 283
rect 19 143 71 187
rect 314 168 361 249
rect 437 279 471 335
rect 505 337 525 371
rect 559 337 561 371
rect 505 313 561 337
rect 437 263 503 279
rect 437 229 453 263
rect 487 229 503 263
rect 437 227 503 229
rect 595 193 629 489
rect 1071 481 1087 497
rect 1121 481 1125 515
rect 1071 465 1125 481
rect 773 447 823 463
rect 665 424 739 440
rect 665 390 681 424
rect 737 390 739 424
rect 665 384 739 390
rect 807 420 823 447
rect 937 447 1017 463
rect 807 413 903 420
rect 773 386 903 413
rect 663 306 835 350
rect 663 272 783 306
rect 817 272 835 306
rect 663 242 835 272
rect 869 322 903 386
rect 937 413 945 447
rect 979 429 1017 447
rect 979 413 1024 429
rect 937 363 1024 413
rect 1078 424 1125 465
rect 1159 523 1304 539
rect 1338 536 1354 570
rect 1388 536 1404 570
rect 1338 535 1404 536
rect 1159 489 1173 523
rect 1207 501 1304 523
rect 1438 523 1513 539
rect 1438 501 1463 523
rect 1207 489 1463 501
rect 1497 489 1513 523
rect 1159 467 1513 489
rect 1555 535 1605 649
rect 1555 501 1571 535
rect 1555 467 1605 501
rect 1159 458 1290 467
rect 1078 390 1222 424
rect 990 356 1024 363
rect 990 340 1154 356
rect 869 306 956 322
rect 869 272 920 306
rect 954 272 956 306
rect 869 256 956 272
rect 990 306 1090 340
rect 1124 306 1154 340
rect 869 208 903 256
rect 990 231 1154 306
rect 981 222 1154 231
rect 395 159 629 193
rect 760 181 903 208
rect 395 157 461 159
rect 19 109 35 143
rect 69 109 71 143
rect 19 93 71 109
rect 105 137 171 153
rect 105 103 121 137
rect 155 103 171 137
rect 105 17 171 103
rect 223 137 283 153
rect 223 103 248 137
rect 282 103 298 137
rect 395 123 411 157
rect 445 123 461 157
rect 670 140 722 156
rect 395 121 461 123
rect 570 123 636 125
rect 223 87 298 103
rect 570 89 586 123
rect 620 89 636 123
rect 570 87 636 89
rect 223 53 636 87
rect 670 106 672 140
rect 706 106 722 140
rect 760 147 770 181
rect 804 172 903 181
rect 954 215 1154 222
rect 954 210 1024 215
rect 954 174 1018 210
rect 804 147 812 172
rect 760 119 812 147
rect 954 140 966 174
rect 1000 140 1018 174
rect 670 17 722 106
rect 852 104 868 138
rect 902 104 918 138
rect 954 119 1018 140
rect 1052 165 1086 181
rect 852 17 918 104
rect 1052 17 1086 131
rect 1120 96 1154 215
rect 1188 180 1222 390
rect 1188 130 1222 146
rect 1256 178 1290 458
rect 1324 415 1358 431
rect 1324 247 1358 381
rect 1392 329 1426 467
rect 1555 433 1571 467
rect 1460 424 1521 431
rect 1460 390 1471 424
rect 1505 415 1521 424
rect 1555 417 1605 433
rect 1662 539 1726 582
rect 1662 505 1680 539
rect 1714 505 1726 539
rect 1662 471 1726 505
rect 1662 437 1666 471
rect 1700 437 1726 471
rect 1460 381 1481 390
rect 1515 381 1521 415
rect 1460 365 1521 381
rect 1662 416 1726 437
rect 1765 563 1831 582
rect 1942 570 2091 649
rect 2230 607 2296 649
rect 2230 573 2246 607
rect 2280 573 2296 607
rect 1765 529 1781 563
rect 1815 534 1831 563
rect 2021 555 2091 570
rect 1815 529 1987 534
rect 1765 498 1987 529
rect 2055 521 2091 555
rect 2021 505 2091 521
rect 2125 555 2179 571
rect 2125 521 2129 555
rect 2163 521 2179 555
rect 1765 471 1821 498
rect 1765 437 1781 471
rect 1815 437 1821 471
rect 1765 416 1821 437
rect 1855 448 1919 464
rect 1593 331 1628 347
rect 1392 297 1593 329
rect 1627 297 1628 331
rect 1392 281 1628 297
rect 1662 247 1712 416
rect 1855 414 1871 448
rect 1905 414 1919 448
rect 1855 398 1919 414
rect 1855 380 1903 398
rect 1324 246 1712 247
rect 1324 212 1662 246
rect 1696 212 1712 246
rect 1746 340 1903 380
rect 1953 352 1987 498
rect 2125 494 2179 521
rect 2025 448 2101 460
rect 2025 424 2051 448
rect 2025 390 2041 424
rect 2085 414 2101 448
rect 2075 390 2101 414
rect 2025 388 2101 390
rect 2135 422 2179 494
rect 2230 490 2296 573
rect 2230 456 2246 490
rect 2280 456 2296 490
rect 2330 599 2383 615
rect 2330 565 2336 599
rect 2370 565 2383 599
rect 2330 498 2383 565
rect 2330 464 2336 498
rect 2370 464 2383 498
rect 2135 388 2247 422
rect 1746 268 1814 340
rect 1953 336 2175 352
rect 1953 306 2125 336
rect 1746 234 1757 268
rect 1791 234 1814 268
rect 1746 193 1814 234
rect 1741 186 1814 193
rect 1734 178 1814 186
rect 1256 172 1324 178
rect 1256 138 1274 172
rect 1308 138 1324 172
rect 1256 130 1324 138
rect 1449 164 1814 178
rect 1848 302 2125 306
rect 2159 302 2175 336
rect 1848 286 2175 302
rect 1848 272 1991 286
rect 1449 155 1780 164
rect 1449 144 1770 155
rect 1449 96 1485 144
rect 1848 130 1889 272
rect 2213 252 2247 388
rect 2025 238 2247 252
rect 1923 224 2247 238
rect 1923 190 1939 224
rect 1973 214 2247 224
rect 2330 409 2383 464
rect 2330 375 2336 409
rect 2370 375 2383 409
rect 1973 190 2200 214
rect 1923 172 2200 190
rect 2330 204 2383 375
rect 2417 607 2481 649
rect 2417 573 2422 607
rect 2456 573 2481 607
rect 2417 509 2481 573
rect 2417 475 2422 509
rect 2456 475 2481 509
rect 2619 607 2681 649
rect 2619 573 2635 607
rect 2669 573 2681 607
rect 2619 510 2681 573
rect 2417 409 2481 475
rect 2417 375 2431 409
rect 2465 375 2481 409
rect 2417 359 2481 375
rect 2515 483 2577 499
rect 2515 449 2527 483
rect 2561 449 2577 483
rect 2515 413 2577 449
rect 2515 379 2527 413
rect 2561 379 2577 413
rect 2515 312 2577 379
rect 2619 476 2635 510
rect 2669 476 2681 510
rect 2619 413 2681 476
rect 2619 379 2635 413
rect 2669 379 2681 413
rect 2619 363 2681 379
rect 2715 599 2762 615
rect 2715 565 2721 599
rect 2755 565 2762 599
rect 2715 495 2762 565
rect 2715 461 2721 495
rect 2755 461 2762 495
rect 2715 413 2762 461
rect 2715 379 2721 413
rect 2755 379 2762 413
rect 2515 296 2681 312
rect 2515 262 2647 296
rect 2515 246 2681 262
rect 1804 114 1889 130
rect 1120 62 1485 96
rect 1519 76 1535 110
rect 1569 76 1585 110
rect 1519 17 1585 76
rect 1838 80 1889 114
rect 1804 51 1889 80
rect 1976 118 2042 134
rect 1976 84 1992 118
rect 2026 84 2042 118
rect 1976 17 2042 84
rect 2134 127 2200 172
rect 2134 93 2150 127
rect 2184 93 2200 127
rect 2134 66 2200 93
rect 2238 164 2296 180
rect 2238 130 2254 164
rect 2288 130 2296 164
rect 2238 94 2296 130
rect 2238 60 2254 94
rect 2288 60 2296 94
rect 2238 17 2296 60
rect 2330 170 2340 204
rect 2374 170 2383 204
rect 2330 101 2383 170
rect 2330 67 2340 101
rect 2374 67 2383 101
rect 2330 51 2383 67
rect 2417 203 2481 219
rect 2417 169 2426 203
rect 2460 169 2481 203
rect 2417 94 2481 169
rect 2417 60 2445 94
rect 2479 60 2481 94
rect 2417 17 2481 60
rect 2515 107 2581 246
rect 2715 212 2762 379
rect 2796 607 2857 649
rect 2796 573 2807 607
rect 2841 573 2857 607
rect 2796 510 2857 573
rect 2796 476 2807 510
rect 2841 476 2857 510
rect 2796 413 2857 476
rect 2796 379 2807 413
rect 2841 379 2857 413
rect 2796 363 2857 379
rect 2515 73 2531 107
rect 2565 73 2581 107
rect 2515 57 2581 73
rect 2619 196 2681 212
rect 2619 162 2635 196
rect 2669 162 2681 196
rect 2619 102 2681 162
rect 2619 68 2635 102
rect 2669 68 2681 102
rect 2619 17 2681 68
rect 2715 178 2721 212
rect 2755 178 2762 212
rect 2715 101 2762 178
rect 2715 67 2721 101
rect 2755 67 2762 101
rect 2715 51 2762 67
rect 2796 212 2857 228
rect 2796 178 2807 212
rect 2841 178 2857 212
rect 2796 102 2857 178
rect 2796 68 2807 102
rect 2841 68 2857 102
rect 2796 17 2857 68
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 703 390 715 424
rect 715 390 737 424
rect 1471 415 1505 424
rect 1471 390 1481 415
rect 1481 390 1505 415
rect 2041 414 2051 424
rect 2051 414 2075 424
rect 2041 390 2075 414
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 691 424 749 430
rect 691 390 703 424
rect 737 421 749 424
rect 1459 424 1517 430
rect 1459 421 1471 424
rect 737 393 1471 421
rect 737 390 749 393
rect 691 384 749 390
rect 1459 390 1471 393
rect 1505 421 1517 424
rect 2029 424 2087 430
rect 2029 421 2041 424
rect 1505 393 2041 421
rect 1505 390 1517 393
rect 1459 384 1517 390
rect 2029 390 2041 393
rect 2075 390 2087 424
rect 2029 384 2087 390
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel comment s 1368 630 1368 630 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 sdfrbp_2
flabel comment s 1061 36 1061 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel metal1 s 2047 390 2081 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2719 242 2753 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2719 316 2753 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2719 390 2753 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2719 464 2753 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2719 538 2753 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 2335 94 2369 128 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2335 168 2369 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2335 242 2369 276 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2335 316 2369 350 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2335 390 2369 424 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2335 464 2369 498 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2335 538 2369 572 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2880 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry R90
string GDS_END 6195420
string GDS_START 6171652
<< end >>
