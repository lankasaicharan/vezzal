magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1490 1975
<< nwell >>
rect -38 331 230 704
<< pwell >>
rect 1 49 191 289
rect 0 0 192 49
<< ndiff >>
rect 27 251 165 263
rect 27 217 39 251
rect 73 217 119 251
rect 153 217 165 251
rect 27 172 165 217
rect 27 138 39 172
rect 73 138 119 172
rect 153 138 165 172
rect 27 93 165 138
rect 27 59 39 93
rect 73 59 119 93
rect 153 59 165 93
rect 27 47 165 59
<< ndiffc >>
rect 39 217 73 251
rect 119 217 153 251
rect 39 138 73 172
rect 119 138 153 172
rect 39 59 73 93
rect 119 59 153 93
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 18 251 174 615
rect 18 217 39 251
rect 73 217 119 251
rect 153 217 174 251
rect 18 172 174 217
rect 18 138 39 172
rect 73 138 119 172
rect 153 138 174 172
rect 18 93 174 138
rect 18 59 39 93
rect 73 59 119 93
rect 153 59 174 93
rect 18 51 174 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 31 -17 65 17
rect 127 -17 161 17
<< metal1 >>
rect 0 683 192 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 192 683
rect 0 617 192 649
rect 0 17 192 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 192 17
rect 0 -49 192 -17
<< labels >>
flabel pwell s 0 0 192 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 192 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 127 538 161 572 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 31 168 65 202 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 127 168 161 202 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 31 94 65 128 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 127 464 161 498 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 127 242 161 276 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 127 390 161 424 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 31 390 65 424 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 31 464 65 498 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 31 538 65 572 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 127 94 161 128 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 31 316 65 350 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 127 316 161 350 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
flabel locali s 31 242 65 276 0 FreeSans 200 0 0 0 DIODE
port 1 nsew default bidirectional
rlabel comment s 0 0 0 0 4 diode_1
flabel metal1 s 0 617 192 666 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 192 49 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE ANTENNACELL
string FIXED_BBOX 0 0 192 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4378192
string GDS_START 4374374
<< end >>
