magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 671 259 1135 263
rect 191 161 1135 259
rect 1 49 1135 161
rect 0 0 1152 49
<< scnmos >>
rect 80 51 110 135
rect 270 65 300 233
rect 356 65 386 233
rect 456 65 486 233
rect 556 65 586 233
rect 766 69 796 237
rect 852 69 882 237
rect 938 69 968 237
rect 1026 69 1056 237
<< scpmoshvt >>
rect 145 367 175 451
rect 270 367 300 619
rect 356 367 386 619
rect 456 367 486 619
rect 544 367 574 619
rect 766 367 796 619
rect 852 367 882 619
rect 938 367 968 619
rect 1024 367 1054 619
<< ndiff >>
rect 217 221 270 233
rect 217 187 225 221
rect 259 187 270 221
rect 27 110 80 135
rect 27 76 35 110
rect 69 76 80 110
rect 27 51 80 76
rect 110 101 163 135
rect 110 67 121 101
rect 155 67 163 101
rect 110 51 163 67
rect 217 111 270 187
rect 217 77 225 111
rect 259 77 270 111
rect 217 65 270 77
rect 300 225 356 233
rect 300 191 311 225
rect 345 191 356 225
rect 300 153 356 191
rect 300 119 311 153
rect 345 119 356 153
rect 300 65 356 119
rect 386 181 456 233
rect 386 147 411 181
rect 445 147 456 181
rect 386 107 456 147
rect 386 73 411 107
rect 445 73 456 107
rect 386 65 456 73
rect 486 111 556 233
rect 486 77 511 111
rect 545 77 556 111
rect 486 65 556 77
rect 586 179 639 233
rect 586 145 597 179
rect 631 145 639 179
rect 586 65 639 145
rect 697 225 766 237
rect 697 191 705 225
rect 739 191 766 225
rect 697 153 766 191
rect 697 119 705 153
rect 739 119 766 153
rect 697 69 766 119
rect 796 183 852 237
rect 796 149 807 183
rect 841 149 852 183
rect 796 111 852 149
rect 796 77 807 111
rect 841 77 852 111
rect 796 69 852 77
rect 882 225 938 237
rect 882 191 893 225
rect 927 191 938 225
rect 882 115 938 191
rect 882 81 893 115
rect 927 81 938 115
rect 882 69 938 81
rect 968 183 1026 237
rect 968 149 981 183
rect 1015 149 1026 183
rect 968 111 1026 149
rect 968 77 981 111
rect 1015 77 1026 111
rect 968 69 1026 77
rect 1056 225 1109 237
rect 1056 191 1067 225
rect 1101 191 1109 225
rect 1056 115 1109 191
rect 1056 81 1067 115
rect 1101 81 1109 115
rect 1056 69 1109 81
<< pdiff >>
rect 213 611 270 619
rect 213 577 225 611
rect 259 577 270 611
rect 213 511 270 577
rect 213 477 225 511
rect 259 477 270 511
rect 213 451 270 477
rect 92 429 145 451
rect 92 395 100 429
rect 134 395 145 429
rect 92 367 145 395
rect 175 413 270 451
rect 175 379 191 413
rect 225 379 270 413
rect 175 367 270 379
rect 300 599 356 619
rect 300 565 311 599
rect 345 565 356 599
rect 300 515 356 565
rect 300 481 311 515
rect 345 481 356 515
rect 300 434 356 481
rect 300 400 311 434
rect 345 400 356 434
rect 300 367 356 400
rect 386 607 456 619
rect 386 573 404 607
rect 438 573 456 607
rect 386 494 456 573
rect 386 460 404 494
rect 438 460 456 494
rect 386 367 456 460
rect 486 599 544 619
rect 486 565 499 599
rect 533 565 544 599
rect 486 508 544 565
rect 486 474 499 508
rect 533 474 544 508
rect 486 418 544 474
rect 486 384 499 418
rect 533 384 544 418
rect 486 367 544 384
rect 574 607 766 619
rect 574 573 585 607
rect 619 573 653 607
rect 687 573 721 607
rect 755 573 766 607
rect 574 492 766 573
rect 574 458 585 492
rect 619 458 653 492
rect 687 458 721 492
rect 755 458 766 492
rect 574 367 766 458
rect 796 599 852 619
rect 796 565 807 599
rect 841 565 852 599
rect 796 508 852 565
rect 796 474 807 508
rect 841 474 852 508
rect 796 424 852 474
rect 796 390 807 424
rect 841 390 852 424
rect 796 367 852 390
rect 882 607 938 619
rect 882 573 893 607
rect 927 573 938 607
rect 882 495 938 573
rect 882 461 893 495
rect 927 461 938 495
rect 882 367 938 461
rect 968 599 1024 619
rect 968 565 979 599
rect 1013 565 1024 599
rect 968 516 1024 565
rect 968 482 979 516
rect 1013 482 1024 516
rect 968 434 1024 482
rect 968 400 979 434
rect 1013 400 1024 434
rect 968 367 1024 400
rect 1054 607 1107 619
rect 1054 573 1065 607
rect 1099 573 1107 607
rect 1054 508 1107 573
rect 1054 474 1065 508
rect 1099 474 1107 508
rect 1054 418 1107 474
rect 1054 384 1065 418
rect 1099 384 1107 418
rect 1054 367 1107 384
<< ndiffc >>
rect 225 187 259 221
rect 35 76 69 110
rect 121 67 155 101
rect 225 77 259 111
rect 311 191 345 225
rect 311 119 345 153
rect 411 147 445 181
rect 411 73 445 107
rect 511 77 545 111
rect 597 145 631 179
rect 705 191 739 225
rect 705 119 739 153
rect 807 149 841 183
rect 807 77 841 111
rect 893 191 927 225
rect 893 81 927 115
rect 981 149 1015 183
rect 981 77 1015 111
rect 1067 191 1101 225
rect 1067 81 1101 115
<< pdiffc >>
rect 225 577 259 611
rect 225 477 259 511
rect 100 395 134 429
rect 191 379 225 413
rect 311 565 345 599
rect 311 481 345 515
rect 311 400 345 434
rect 404 573 438 607
rect 404 460 438 494
rect 499 565 533 599
rect 499 474 533 508
rect 499 384 533 418
rect 585 573 619 607
rect 653 573 687 607
rect 721 573 755 607
rect 585 458 619 492
rect 653 458 687 492
rect 721 458 755 492
rect 807 565 841 599
rect 807 474 841 508
rect 807 390 841 424
rect 893 573 927 607
rect 893 461 927 495
rect 979 565 1013 599
rect 979 482 1013 516
rect 979 400 1013 434
rect 1065 573 1099 607
rect 1065 474 1099 508
rect 1065 384 1099 418
<< poly >>
rect 270 619 300 645
rect 356 619 386 645
rect 456 619 486 645
rect 544 619 574 645
rect 766 619 796 645
rect 852 619 882 645
rect 938 619 968 645
rect 1024 619 1054 645
rect 145 451 175 477
rect 145 325 175 367
rect 270 335 300 367
rect 356 335 386 367
rect 21 309 175 325
rect 21 275 37 309
rect 71 295 175 309
rect 217 319 386 335
rect 71 275 110 295
rect 21 241 110 275
rect 217 285 233 319
rect 267 285 301 319
rect 335 285 386 319
rect 217 269 386 285
rect 21 207 37 241
rect 71 207 110 241
rect 270 233 300 269
rect 356 233 386 269
rect 456 335 486 367
rect 544 335 574 367
rect 766 335 796 367
rect 852 335 882 367
rect 456 319 574 335
rect 456 285 474 319
rect 508 299 574 319
rect 748 319 882 335
rect 508 285 586 299
rect 456 269 586 285
rect 748 285 764 319
rect 798 285 832 319
rect 866 285 882 319
rect 748 269 882 285
rect 456 233 486 269
rect 556 233 586 269
rect 766 237 796 269
rect 852 237 882 269
rect 938 335 968 367
rect 1024 335 1054 367
rect 938 319 1056 335
rect 938 285 1003 319
rect 1037 285 1056 319
rect 938 269 1056 285
rect 938 237 968 269
rect 1026 237 1056 269
rect 21 191 110 207
rect 80 135 110 191
rect 80 25 110 51
rect 270 39 300 65
rect 356 39 386 65
rect 456 39 486 65
rect 556 39 586 65
rect 766 43 796 69
rect 852 43 882 69
rect 938 43 968 69
rect 1026 43 1056 69
<< polycont >>
rect 37 275 71 309
rect 233 285 267 319
rect 301 285 335 319
rect 37 207 71 241
rect 474 285 508 319
rect 764 285 798 319
rect 832 285 866 319
rect 1003 285 1037 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 191 611 267 649
rect 191 577 225 611
rect 259 577 267 611
rect 191 511 267 577
rect 191 477 225 511
rect 259 477 267 511
rect 84 429 157 445
rect 84 395 100 429
rect 134 395 157 429
rect 84 379 157 395
rect 121 329 157 379
rect 191 413 267 477
rect 225 379 267 413
rect 301 599 354 615
rect 301 565 311 599
rect 345 565 354 599
rect 301 515 354 565
rect 301 481 311 515
rect 345 481 354 515
rect 301 434 354 481
rect 388 607 454 649
rect 388 573 404 607
rect 438 573 454 607
rect 388 494 454 573
rect 388 460 404 494
rect 438 460 454 494
rect 388 452 454 460
rect 488 599 535 615
rect 488 565 499 599
rect 533 565 535 599
rect 488 508 535 565
rect 488 474 499 508
rect 533 474 535 508
rect 301 400 311 434
rect 345 418 354 434
rect 488 424 535 474
rect 569 607 771 649
rect 569 573 585 607
rect 619 573 653 607
rect 687 573 721 607
rect 755 573 771 607
rect 569 492 771 573
rect 569 458 585 492
rect 619 458 653 492
rect 687 458 721 492
rect 755 458 771 492
rect 805 599 843 615
rect 805 565 807 599
rect 841 565 843 599
rect 805 508 843 565
rect 805 474 807 508
rect 841 474 843 508
rect 805 424 843 474
rect 877 607 943 649
rect 877 573 893 607
rect 927 573 943 607
rect 877 495 943 573
rect 877 461 893 495
rect 927 461 943 495
rect 877 452 943 461
rect 977 599 1015 615
rect 977 565 979 599
rect 1013 565 1015 599
rect 977 516 1015 565
rect 977 482 979 516
rect 1013 482 1015 516
rect 488 418 807 424
rect 345 400 499 418
rect 301 384 499 400
rect 533 390 807 418
rect 841 418 843 424
rect 977 434 1015 482
rect 977 418 979 434
rect 841 400 979 418
rect 1013 400 1015 434
rect 841 390 1015 400
rect 533 384 1015 390
rect 1049 607 1115 649
rect 1049 573 1065 607
rect 1099 573 1115 607
rect 1049 508 1115 573
rect 1049 474 1065 508
rect 1099 474 1115 508
rect 1049 418 1115 474
rect 1049 384 1065 418
rect 1099 384 1115 418
rect 191 363 267 379
rect 21 309 87 325
rect 21 275 37 309
rect 71 275 87 309
rect 21 241 87 275
rect 21 207 37 241
rect 71 207 87 241
rect 121 319 351 329
rect 121 285 233 319
rect 267 285 301 319
rect 335 285 351 319
rect 121 283 351 285
rect 385 319 547 350
rect 385 285 474 319
rect 508 285 547 319
rect 385 283 547 285
rect 121 173 157 283
rect 581 249 643 384
rect 677 319 943 350
rect 677 285 764 319
rect 798 285 832 319
rect 866 285 943 319
rect 977 319 1121 350
rect 977 285 1003 319
rect 1037 285 1121 319
rect 31 139 157 173
rect 209 221 261 237
rect 209 187 225 221
rect 259 187 261 221
rect 31 110 69 139
rect 31 76 35 110
rect 209 111 261 187
rect 295 225 643 249
rect 295 191 311 225
rect 345 215 643 225
rect 689 225 1121 251
rect 345 191 361 215
rect 295 153 361 191
rect 689 191 705 225
rect 739 217 893 225
rect 739 191 755 217
rect 295 119 311 153
rect 345 119 361 153
rect 395 147 411 181
rect 445 179 647 181
rect 445 147 597 179
rect 395 145 597 147
rect 631 145 647 179
rect 31 60 69 76
rect 105 101 171 105
rect 105 67 121 101
rect 155 67 171 101
rect 105 17 171 67
rect 209 77 225 111
rect 259 85 261 111
rect 395 107 461 145
rect 595 129 647 145
rect 689 153 755 191
rect 891 191 893 217
rect 927 217 1067 225
rect 927 191 931 217
rect 689 119 705 153
rect 739 119 755 153
rect 791 149 807 183
rect 841 149 857 183
rect 791 111 857 149
rect 395 85 411 107
rect 259 77 411 85
rect 209 73 411 77
rect 445 73 461 107
rect 209 51 461 73
rect 495 77 511 111
rect 545 85 561 111
rect 791 85 807 111
rect 545 77 807 85
rect 841 77 857 111
rect 495 51 857 77
rect 891 115 931 191
rect 1065 191 1067 217
rect 1101 191 1121 225
rect 891 81 893 115
rect 927 81 931 115
rect 891 65 931 81
rect 965 149 981 183
rect 1015 149 1031 183
rect 965 111 1031 149
rect 965 77 981 111
rect 1015 77 1031 111
rect 965 17 1031 77
rect 1065 115 1121 191
rect 1065 81 1067 115
rect 1101 81 1121 115
rect 1065 65 1121 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4b_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 648716
string GDS_START 638372
<< end >>
