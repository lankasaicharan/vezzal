magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2954 1852
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 1 21 1631 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 173 47 203 177
rect 267 47 297 177
rect 361 47 391 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 747 47 777 177
rect 831 47 861 177
rect 925 47 955 177
rect 1019 47 1049 177
rect 1113 47 1143 177
rect 1207 47 1237 177
rect 1301 47 1331 177
rect 1395 47 1425 177
rect 1499 47 1529 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
rect 1209 297 1245 497
rect 1303 297 1339 497
rect 1397 297 1433 497
rect 1491 297 1527 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 97 173 177
rect 109 63 129 97
rect 163 63 173 97
rect 109 47 173 63
rect 203 165 267 177
rect 203 131 223 165
rect 257 131 267 165
rect 203 97 267 131
rect 203 63 223 97
rect 257 63 267 97
rect 203 47 267 63
rect 297 97 361 177
rect 297 63 317 97
rect 351 63 361 97
rect 297 47 361 63
rect 391 165 455 177
rect 391 131 411 165
rect 445 131 455 165
rect 391 97 455 131
rect 391 63 411 97
rect 445 63 455 97
rect 391 47 455 63
rect 485 97 549 177
rect 485 63 505 97
rect 539 63 549 97
rect 485 47 549 63
rect 579 165 643 177
rect 579 131 599 165
rect 633 131 643 165
rect 579 97 643 131
rect 579 63 599 97
rect 633 63 643 97
rect 579 47 643 63
rect 673 97 747 177
rect 673 63 693 97
rect 727 63 747 97
rect 673 47 747 63
rect 777 165 831 177
rect 777 131 787 165
rect 821 131 831 165
rect 777 97 831 131
rect 777 63 787 97
rect 821 63 831 97
rect 777 47 831 63
rect 861 165 925 177
rect 861 131 881 165
rect 915 131 925 165
rect 861 47 925 131
rect 955 97 1019 177
rect 955 63 975 97
rect 1009 63 1019 97
rect 955 47 1019 63
rect 1049 165 1113 177
rect 1049 131 1069 165
rect 1103 131 1113 165
rect 1049 47 1113 131
rect 1143 97 1207 177
rect 1143 63 1163 97
rect 1197 63 1207 97
rect 1143 47 1207 63
rect 1237 165 1301 177
rect 1237 131 1257 165
rect 1291 131 1301 165
rect 1237 47 1301 131
rect 1331 97 1395 177
rect 1331 63 1351 97
rect 1385 63 1395 97
rect 1331 47 1395 63
rect 1425 165 1499 177
rect 1425 131 1445 165
rect 1479 131 1499 165
rect 1425 47 1499 131
rect 1529 165 1605 177
rect 1529 131 1559 165
rect 1593 131 1605 165
rect 1529 97 1605 131
rect 1529 63 1559 97
rect 1593 63 1605 97
rect 1529 47 1605 63
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 349 551 383
rect 493 315 505 349
rect 539 315 551 349
rect 493 297 551 315
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 417 645 451
rect 587 383 599 417
rect 633 383 645 417
rect 587 297 645 383
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 349 739 383
rect 681 315 693 349
rect 727 315 739 349
rect 681 297 739 315
rect 775 485 833 497
rect 775 451 787 485
rect 821 451 833 485
rect 775 417 833 451
rect 775 383 787 417
rect 821 383 833 417
rect 775 297 833 383
rect 869 485 927 497
rect 869 451 881 485
rect 915 451 927 485
rect 869 417 927 451
rect 869 383 881 417
rect 915 383 927 417
rect 869 349 927 383
rect 869 315 881 349
rect 915 315 927 349
rect 869 297 927 315
rect 963 485 1021 497
rect 963 451 975 485
rect 1009 451 1021 485
rect 963 417 1021 451
rect 963 383 975 417
rect 1009 383 1021 417
rect 963 297 1021 383
rect 1057 485 1115 497
rect 1057 451 1069 485
rect 1103 451 1115 485
rect 1057 417 1115 451
rect 1057 383 1069 417
rect 1103 383 1115 417
rect 1057 349 1115 383
rect 1057 315 1069 349
rect 1103 315 1115 349
rect 1057 297 1115 315
rect 1151 485 1209 497
rect 1151 451 1163 485
rect 1197 451 1209 485
rect 1151 417 1209 451
rect 1151 383 1163 417
rect 1197 383 1209 417
rect 1151 297 1209 383
rect 1245 485 1303 497
rect 1245 451 1257 485
rect 1291 451 1303 485
rect 1245 417 1303 451
rect 1245 383 1257 417
rect 1291 383 1303 417
rect 1245 349 1303 383
rect 1245 315 1257 349
rect 1291 315 1303 349
rect 1245 297 1303 315
rect 1339 485 1397 497
rect 1339 451 1351 485
rect 1385 451 1397 485
rect 1339 417 1397 451
rect 1339 383 1351 417
rect 1385 383 1397 417
rect 1339 297 1397 383
rect 1433 485 1491 497
rect 1433 451 1445 485
rect 1479 451 1491 485
rect 1433 417 1491 451
rect 1433 383 1445 417
rect 1479 383 1491 417
rect 1433 349 1491 383
rect 1433 315 1445 349
rect 1479 315 1491 349
rect 1433 297 1491 315
rect 1527 485 1605 497
rect 1527 451 1559 485
rect 1593 451 1605 485
rect 1527 417 1605 451
rect 1527 383 1559 417
rect 1593 383 1605 417
rect 1527 349 1605 383
rect 1527 315 1559 349
rect 1593 315 1605 349
rect 1527 297 1605 315
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 129 63 163 97
rect 223 131 257 165
rect 223 63 257 97
rect 317 63 351 97
rect 411 131 445 165
rect 411 63 445 97
rect 505 63 539 97
rect 599 131 633 165
rect 599 63 633 97
rect 693 63 727 97
rect 787 131 821 165
rect 787 63 821 97
rect 881 131 915 165
rect 975 63 1009 97
rect 1069 131 1103 165
rect 1163 63 1197 97
rect 1257 131 1291 165
rect 1351 63 1385 97
rect 1445 131 1479 165
rect 1559 131 1593 165
rect 1559 63 1593 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 505 451 539 485
rect 505 383 539 417
rect 505 315 539 349
rect 599 451 633 485
rect 599 383 633 417
rect 693 451 727 485
rect 693 383 727 417
rect 693 315 727 349
rect 787 451 821 485
rect 787 383 821 417
rect 881 451 915 485
rect 881 383 915 417
rect 881 315 915 349
rect 975 451 1009 485
rect 975 383 1009 417
rect 1069 451 1103 485
rect 1069 383 1103 417
rect 1069 315 1103 349
rect 1163 451 1197 485
rect 1163 383 1197 417
rect 1257 451 1291 485
rect 1257 383 1291 417
rect 1257 315 1291 349
rect 1351 451 1385 485
rect 1351 383 1385 417
rect 1445 451 1479 485
rect 1445 383 1479 417
rect 1445 315 1479 349
rect 1559 451 1593 485
rect 1559 383 1593 417
rect 1559 315 1593 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 1209 497 1245 523
rect 1303 497 1339 523
rect 1397 497 1433 523
rect 1491 497 1527 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 1209 282 1245 297
rect 1303 282 1339 297
rect 1397 282 1433 297
rect 1491 282 1527 297
rect 79 259 119 282
rect 173 259 213 282
rect 267 259 307 282
rect 361 259 401 282
rect 455 259 495 282
rect 549 259 589 282
rect 643 259 683 282
rect 737 259 777 282
rect 79 249 777 259
rect 79 215 128 249
rect 162 215 223 249
rect 257 215 317 249
rect 351 215 411 249
rect 445 215 505 249
rect 539 215 599 249
rect 633 215 693 249
rect 727 215 777 249
rect 79 205 777 215
rect 79 177 109 205
rect 173 177 203 205
rect 267 177 297 205
rect 361 177 391 205
rect 455 177 485 205
rect 549 177 579 205
rect 643 177 673 205
rect 747 177 777 205
rect 831 259 871 282
rect 925 259 965 282
rect 1019 259 1059 282
rect 1113 259 1153 282
rect 1207 259 1247 282
rect 1301 259 1341 282
rect 1395 259 1435 282
rect 1489 259 1529 282
rect 831 249 1529 259
rect 831 215 975 249
rect 1009 215 1069 249
rect 1103 215 1163 249
rect 1197 215 1257 249
rect 1291 215 1351 249
rect 1385 215 1529 249
rect 831 205 1529 215
rect 831 177 861 205
rect 925 177 955 205
rect 1019 177 1049 205
rect 1113 177 1143 205
rect 1207 177 1237 205
rect 1301 177 1331 205
rect 1395 177 1425 205
rect 1499 177 1529 205
rect 79 21 109 47
rect 173 21 203 47
rect 267 21 297 47
rect 361 21 391 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 747 21 777 47
rect 831 21 861 47
rect 925 21 955 47
rect 1019 21 1049 47
rect 1113 21 1143 47
rect 1207 21 1237 47
rect 1301 21 1331 47
rect 1395 21 1425 47
rect 1499 21 1529 47
<< polycont >>
rect 128 215 162 249
rect 223 215 257 249
rect 317 215 351 249
rect 411 215 445 249
rect 505 215 539 249
rect 599 215 633 249
rect 693 215 727 249
rect 975 215 1009 249
rect 1069 215 1103 249
rect 1163 215 1197 249
rect 1257 215 1291 249
rect 1351 215 1385 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 485 179 493
rect 103 451 129 485
rect 163 451 179 485
rect 103 417 179 451
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 223 485 257 527
rect 223 417 257 451
rect 223 367 257 383
rect 291 485 367 493
rect 291 451 317 485
rect 351 451 367 485
rect 291 417 367 451
rect 291 383 317 417
rect 351 383 367 417
rect 103 315 129 349
rect 163 333 179 349
rect 291 349 367 383
rect 411 485 445 527
rect 411 417 445 451
rect 411 367 445 383
rect 479 485 555 493
rect 479 451 505 485
rect 539 451 555 485
rect 479 417 555 451
rect 479 383 505 417
rect 539 383 555 417
rect 291 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 479 349 555 383
rect 599 485 633 527
rect 599 417 633 451
rect 599 367 633 383
rect 667 485 743 493
rect 667 451 693 485
rect 727 451 743 485
rect 667 417 743 451
rect 667 383 693 417
rect 727 383 743 417
rect 479 333 505 349
rect 351 315 505 333
rect 539 333 555 349
rect 667 349 743 383
rect 787 485 821 527
rect 787 417 821 451
rect 787 367 821 383
rect 855 485 931 493
rect 855 451 881 485
rect 915 451 931 485
rect 855 417 931 451
rect 855 383 881 417
rect 915 383 931 417
rect 667 333 693 349
rect 539 315 693 333
rect 727 333 743 349
rect 855 349 931 383
rect 975 485 1009 527
rect 975 417 1009 451
rect 975 367 1009 383
rect 1043 485 1119 493
rect 1043 451 1069 485
rect 1103 451 1119 485
rect 1043 417 1119 451
rect 1043 383 1069 417
rect 1103 383 1119 417
rect 855 333 881 349
rect 727 315 881 333
rect 915 333 931 349
rect 1043 349 1119 383
rect 1163 485 1197 527
rect 1163 417 1197 451
rect 1163 367 1197 383
rect 1231 485 1307 493
rect 1231 451 1257 485
rect 1291 451 1307 485
rect 1231 417 1307 451
rect 1231 383 1257 417
rect 1291 383 1307 417
rect 1043 333 1069 349
rect 915 315 1069 333
rect 1103 333 1119 349
rect 1231 349 1307 383
rect 1351 485 1385 527
rect 1351 417 1385 451
rect 1351 367 1385 383
rect 1419 485 1495 493
rect 1419 451 1445 485
rect 1479 451 1495 485
rect 1419 417 1495 451
rect 1419 383 1445 417
rect 1479 383 1495 417
rect 1231 333 1257 349
rect 1103 315 1257 333
rect 1291 333 1307 349
rect 1419 349 1495 383
rect 1419 333 1445 349
rect 1291 315 1445 333
rect 1479 315 1495 349
rect 103 293 1495 315
rect 1543 485 1614 527
rect 1543 451 1559 485
rect 1593 451 1614 485
rect 1543 417 1614 451
rect 1543 383 1559 417
rect 1593 383 1614 417
rect 1543 349 1614 383
rect 1543 315 1559 349
rect 1593 315 1614 349
rect 1543 299 1614 315
rect 102 249 743 259
rect 102 215 128 249
rect 162 215 223 249
rect 257 215 317 249
rect 351 215 411 249
rect 445 215 505 249
rect 539 215 599 249
rect 633 215 693 249
rect 727 215 743 249
rect 808 215 914 293
rect 948 249 1401 255
rect 948 215 975 249
rect 1009 215 1069 249
rect 1103 215 1163 249
rect 1197 215 1257 249
rect 1291 215 1351 249
rect 1385 215 1401 249
rect 855 181 914 215
rect 1445 181 1495 293
rect 18 165 821 181
rect 18 131 35 165
rect 69 147 223 165
rect 69 131 85 147
rect 18 97 85 131
rect 197 131 223 147
rect 257 147 411 165
rect 257 131 273 147
rect 18 63 35 97
rect 69 63 85 97
rect 18 51 85 63
rect 129 97 163 113
rect 129 17 163 63
rect 197 97 273 131
rect 385 131 411 147
rect 445 147 599 165
rect 445 131 461 147
rect 197 63 223 97
rect 257 63 273 97
rect 197 51 273 63
rect 317 97 351 113
rect 317 17 351 63
rect 385 97 461 131
rect 573 131 599 147
rect 633 147 787 165
rect 633 131 649 147
rect 385 63 411 97
rect 445 63 461 97
rect 385 51 461 63
rect 505 97 539 113
rect 505 17 539 63
rect 573 97 649 131
rect 761 131 787 147
rect 855 165 1495 181
rect 855 131 881 165
rect 915 131 1069 165
rect 1103 131 1257 165
rect 1291 131 1445 165
rect 1479 131 1495 165
rect 1539 165 1614 181
rect 1539 131 1559 165
rect 1593 131 1614 165
rect 573 63 599 97
rect 633 63 649 97
rect 573 51 649 63
rect 693 97 727 113
rect 693 17 727 63
rect 761 97 821 131
rect 1539 97 1614 131
rect 761 63 787 97
rect 821 63 975 97
rect 1009 63 1163 97
rect 1197 63 1351 97
rect 1385 63 1559 97
rect 1593 63 1614 97
rect 761 51 1614 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel locali s 1041 221 1075 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 1317 221 1351 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 857 289 891 323 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 857 221 891 255 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 1225 221 1259 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 1133 221 1167 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2_8
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1656 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2202794
string GDS_START 2189702
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
