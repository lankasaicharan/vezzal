magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 1 49 1053 241
rect 0 0 1056 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 252 47 282 215
rect 338 47 368 215
rect 424 47 454 215
rect 510 47 540 215
rect 596 47 626 215
rect 682 47 712 215
rect 768 47 798 215
rect 854 47 884 215
rect 940 47 970 215
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 252 367 282 619
rect 338 367 368 619
rect 424 367 454 619
rect 510 367 540 619
rect 596 367 626 619
rect 682 367 712 619
rect 768 367 798 619
rect 854 367 884 619
rect 940 367 970 619
<< ndiff >>
rect 27 185 80 215
rect 27 151 35 185
rect 69 151 80 185
rect 27 111 80 151
rect 27 77 35 111
rect 69 77 80 111
rect 27 47 80 77
rect 110 118 166 215
rect 110 84 121 118
rect 155 84 166 118
rect 110 47 166 84
rect 196 185 252 215
rect 196 151 207 185
rect 241 151 252 185
rect 196 111 252 151
rect 196 77 207 111
rect 241 77 252 111
rect 196 47 252 77
rect 282 159 338 215
rect 282 125 293 159
rect 327 125 338 159
rect 282 91 338 125
rect 282 57 293 91
rect 327 57 338 91
rect 282 47 338 57
rect 368 185 424 215
rect 368 151 379 185
rect 413 151 424 185
rect 368 111 424 151
rect 368 77 379 111
rect 413 77 424 111
rect 368 47 424 77
rect 454 159 510 215
rect 454 125 465 159
rect 499 125 510 159
rect 454 91 510 125
rect 454 57 465 91
rect 499 57 510 91
rect 454 47 510 57
rect 540 185 596 215
rect 540 151 551 185
rect 585 151 596 185
rect 540 111 596 151
rect 540 77 551 111
rect 585 77 596 111
rect 540 47 596 77
rect 626 159 682 215
rect 626 125 637 159
rect 671 125 682 159
rect 626 91 682 125
rect 626 57 637 91
rect 671 57 682 91
rect 626 47 682 57
rect 712 185 768 215
rect 712 151 723 185
rect 757 151 768 185
rect 712 111 768 151
rect 712 77 723 111
rect 757 77 768 111
rect 712 47 768 77
rect 798 159 854 215
rect 798 125 809 159
rect 843 125 854 159
rect 798 91 854 125
rect 798 57 809 91
rect 843 57 854 91
rect 798 47 854 57
rect 884 185 940 215
rect 884 151 895 185
rect 929 151 940 185
rect 884 111 940 151
rect 884 77 895 111
rect 929 77 940 111
rect 884 47 940 77
rect 970 159 1027 215
rect 970 125 981 159
rect 1015 125 1027 159
rect 970 91 1027 125
rect 970 57 981 91
rect 1015 57 1027 91
rect 970 47 1027 57
<< pdiff >>
rect 27 580 80 619
rect 27 546 35 580
rect 69 546 80 580
rect 27 506 80 546
rect 27 472 35 506
rect 69 472 80 506
rect 27 432 80 472
rect 27 398 35 432
rect 69 398 80 432
rect 27 367 80 398
rect 110 605 166 619
rect 110 571 121 605
rect 155 571 166 605
rect 110 537 166 571
rect 110 503 121 537
rect 155 503 166 537
rect 110 469 166 503
rect 110 435 121 469
rect 155 435 166 469
rect 110 367 166 435
rect 196 580 252 619
rect 196 546 207 580
rect 241 546 252 580
rect 196 506 252 546
rect 196 472 207 506
rect 241 472 252 506
rect 196 432 252 472
rect 196 398 207 432
rect 241 398 252 432
rect 196 367 252 398
rect 282 605 338 619
rect 282 571 293 605
rect 327 571 338 605
rect 282 537 338 571
rect 282 503 293 537
rect 327 503 338 537
rect 282 469 338 503
rect 282 435 293 469
rect 327 435 338 469
rect 282 367 338 435
rect 368 580 424 619
rect 368 546 379 580
rect 413 546 424 580
rect 368 506 424 546
rect 368 472 379 506
rect 413 472 424 506
rect 368 432 424 472
rect 368 398 379 432
rect 413 398 424 432
rect 368 367 424 398
rect 454 605 510 619
rect 454 571 465 605
rect 499 571 510 605
rect 454 537 510 571
rect 454 503 465 537
rect 499 503 510 537
rect 454 469 510 503
rect 454 435 465 469
rect 499 435 510 469
rect 454 367 510 435
rect 540 580 596 619
rect 540 546 551 580
rect 585 546 596 580
rect 540 506 596 546
rect 540 472 551 506
rect 585 472 596 506
rect 540 432 596 472
rect 540 398 551 432
rect 585 398 596 432
rect 540 367 596 398
rect 626 605 682 619
rect 626 571 637 605
rect 671 571 682 605
rect 626 537 682 571
rect 626 503 637 537
rect 671 503 682 537
rect 626 469 682 503
rect 626 435 637 469
rect 671 435 682 469
rect 626 367 682 435
rect 712 580 768 619
rect 712 546 723 580
rect 757 546 768 580
rect 712 506 768 546
rect 712 472 723 506
rect 757 472 768 506
rect 712 432 768 472
rect 712 398 723 432
rect 757 398 768 432
rect 712 367 768 398
rect 798 605 854 619
rect 798 571 809 605
rect 843 571 854 605
rect 798 537 854 571
rect 798 503 809 537
rect 843 503 854 537
rect 798 469 854 503
rect 798 435 809 469
rect 843 435 854 469
rect 798 367 854 435
rect 884 580 940 619
rect 884 546 895 580
rect 929 546 940 580
rect 884 506 940 546
rect 884 472 895 506
rect 929 472 940 506
rect 884 432 940 472
rect 884 398 895 432
rect 929 398 940 432
rect 884 367 940 398
rect 970 605 1027 619
rect 970 571 981 605
rect 1015 571 1027 605
rect 970 537 1027 571
rect 970 503 981 537
rect 1015 503 1027 537
rect 970 469 1027 503
rect 970 435 981 469
rect 1015 435 1027 469
rect 970 367 1027 435
<< ndiffc >>
rect 35 151 69 185
rect 35 77 69 111
rect 121 84 155 118
rect 207 151 241 185
rect 207 77 241 111
rect 293 125 327 159
rect 293 57 327 91
rect 379 151 413 185
rect 379 77 413 111
rect 465 125 499 159
rect 465 57 499 91
rect 551 151 585 185
rect 551 77 585 111
rect 637 125 671 159
rect 637 57 671 91
rect 723 151 757 185
rect 723 77 757 111
rect 809 125 843 159
rect 809 57 843 91
rect 895 151 929 185
rect 895 77 929 111
rect 981 125 1015 159
rect 981 57 1015 91
<< pdiffc >>
rect 35 546 69 580
rect 35 472 69 506
rect 35 398 69 432
rect 121 571 155 605
rect 121 503 155 537
rect 121 435 155 469
rect 207 546 241 580
rect 207 472 241 506
rect 207 398 241 432
rect 293 571 327 605
rect 293 503 327 537
rect 293 435 327 469
rect 379 546 413 580
rect 379 472 413 506
rect 379 398 413 432
rect 465 571 499 605
rect 465 503 499 537
rect 465 435 499 469
rect 551 546 585 580
rect 551 472 585 506
rect 551 398 585 432
rect 637 571 671 605
rect 637 503 671 537
rect 637 435 671 469
rect 723 546 757 580
rect 723 472 757 506
rect 723 398 757 432
rect 809 571 843 605
rect 809 503 843 537
rect 809 435 843 469
rect 895 546 929 580
rect 895 472 929 506
rect 895 398 929 432
rect 981 571 1015 605
rect 981 503 1015 537
rect 981 435 1015 469
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 252 619 282 645
rect 338 619 368 645
rect 424 619 454 645
rect 510 619 540 645
rect 596 619 626 645
rect 682 619 712 645
rect 768 619 798 645
rect 854 619 884 645
rect 940 619 970 645
rect 80 329 110 367
rect 166 329 196 367
rect 252 329 282 367
rect 67 313 282 329
rect 67 279 83 313
rect 117 279 151 313
rect 185 279 219 313
rect 253 279 282 313
rect 67 263 282 279
rect 80 215 110 263
rect 166 215 196 263
rect 252 215 282 263
rect 338 329 368 367
rect 424 329 454 367
rect 510 329 540 367
rect 596 329 626 367
rect 682 329 712 367
rect 768 329 798 367
rect 854 329 884 367
rect 940 329 970 367
rect 338 313 970 329
rect 338 279 354 313
rect 388 279 422 313
rect 456 279 490 313
rect 524 279 558 313
rect 592 279 626 313
rect 660 279 694 313
rect 728 279 762 313
rect 796 279 830 313
rect 864 279 898 313
rect 932 279 970 313
rect 338 263 970 279
rect 338 215 368 263
rect 424 215 454 263
rect 510 215 540 263
rect 596 215 626 263
rect 682 215 712 263
rect 768 215 798 263
rect 854 215 884 263
rect 940 215 970 263
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 424 21 454 47
rect 510 21 540 47
rect 596 21 626 47
rect 682 21 712 47
rect 768 21 798 47
rect 854 21 884 47
rect 940 21 970 47
<< polycont >>
rect 83 279 117 313
rect 151 279 185 313
rect 219 279 253 313
rect 354 279 388 313
rect 422 279 456 313
rect 490 279 524 313
rect 558 279 592 313
rect 626 279 660 313
rect 694 279 728 313
rect 762 279 796 313
rect 830 279 864 313
rect 898 279 932 313
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 112 605 164 649
rect 19 580 78 596
rect 19 546 35 580
rect 69 546 78 580
rect 19 506 78 546
rect 19 472 35 506
rect 69 472 78 506
rect 19 432 78 472
rect 19 398 35 432
rect 69 398 78 432
rect 112 571 121 605
rect 155 571 164 605
rect 284 605 339 649
rect 112 537 164 571
rect 112 503 121 537
rect 155 503 164 537
rect 112 469 164 503
rect 112 435 121 469
rect 155 435 164 469
rect 112 419 164 435
rect 198 580 250 596
rect 198 546 207 580
rect 241 546 250 580
rect 198 506 250 546
rect 198 472 207 506
rect 241 472 250 506
rect 198 432 250 472
rect 19 385 78 398
rect 198 398 207 432
rect 241 398 250 432
rect 284 571 293 605
rect 327 571 339 605
rect 455 605 507 649
rect 284 537 339 571
rect 284 503 293 537
rect 327 503 339 537
rect 284 469 339 503
rect 284 435 293 469
rect 327 435 339 469
rect 284 419 339 435
rect 373 580 421 596
rect 373 546 379 580
rect 413 546 421 580
rect 373 506 421 546
rect 373 472 379 506
rect 413 472 421 506
rect 373 432 421 472
rect 198 385 250 398
rect 373 398 379 432
rect 413 398 421 432
rect 455 571 465 605
rect 499 571 507 605
rect 629 605 680 649
rect 455 537 507 571
rect 455 503 465 537
rect 499 503 507 537
rect 455 469 507 503
rect 455 435 465 469
rect 499 435 507 469
rect 455 419 507 435
rect 541 580 595 596
rect 541 546 551 580
rect 585 546 595 580
rect 541 506 595 546
rect 541 472 551 506
rect 585 472 595 506
rect 541 432 595 472
rect 373 385 421 398
rect 541 398 551 432
rect 585 398 595 432
rect 629 571 637 605
rect 671 571 680 605
rect 800 605 852 649
rect 629 537 680 571
rect 629 503 637 537
rect 671 503 680 537
rect 629 469 680 503
rect 629 435 637 469
rect 671 435 680 469
rect 629 419 680 435
rect 714 580 766 596
rect 714 546 723 580
rect 757 546 766 580
rect 714 506 766 546
rect 714 472 723 506
rect 757 472 766 506
rect 714 432 766 472
rect 541 385 595 398
rect 714 398 723 432
rect 757 398 766 432
rect 800 571 809 605
rect 843 571 852 605
rect 972 605 1019 649
rect 800 537 852 571
rect 800 503 809 537
rect 843 503 852 537
rect 800 469 852 503
rect 800 435 809 469
rect 843 435 852 469
rect 800 419 852 435
rect 886 580 938 596
rect 886 546 895 580
rect 929 546 938 580
rect 886 506 938 546
rect 886 472 895 506
rect 929 472 938 506
rect 886 432 938 472
rect 714 385 766 398
rect 886 398 895 432
rect 929 398 938 432
rect 972 571 981 605
rect 1015 571 1019 605
rect 972 537 1019 571
rect 972 503 981 537
rect 1015 503 1019 537
rect 972 469 1019 503
rect 972 435 981 469
rect 1015 435 1019 469
rect 972 419 1019 435
rect 886 385 938 398
rect 19 349 339 385
rect 373 349 1038 385
rect 305 315 339 349
rect 19 313 269 315
rect 19 279 83 313
rect 117 279 151 313
rect 185 279 219 313
rect 253 279 269 313
rect 19 277 269 279
rect 305 313 948 315
rect 305 279 354 313
rect 388 279 422 313
rect 456 279 490 313
rect 524 279 558 313
rect 592 279 626 313
rect 660 279 694 313
rect 728 279 762 313
rect 796 279 830 313
rect 864 279 898 313
rect 932 279 948 313
rect 19 236 176 277
rect 305 243 339 279
rect 982 245 1038 349
rect 210 209 339 243
rect 373 209 1038 245
rect 210 202 250 209
rect 19 185 250 202
rect 19 151 35 185
rect 69 168 207 185
rect 69 151 78 168
rect 19 111 78 151
rect 198 151 207 168
rect 241 151 250 185
rect 373 185 422 209
rect 19 77 35 111
rect 69 77 78 111
rect 19 61 78 77
rect 112 118 164 134
rect 112 84 121 118
rect 155 84 164 118
rect 112 17 164 84
rect 198 111 250 151
rect 198 77 207 111
rect 241 77 250 111
rect 198 61 250 77
rect 284 159 339 175
rect 284 125 293 159
rect 327 125 339 159
rect 284 91 339 125
rect 284 57 293 91
rect 327 57 339 91
rect 373 151 379 185
rect 413 151 422 185
rect 542 185 593 209
rect 373 111 422 151
rect 373 77 379 111
rect 413 77 422 111
rect 373 61 422 77
rect 456 159 508 175
rect 456 125 465 159
rect 499 125 508 159
rect 456 91 508 125
rect 284 17 339 57
rect 456 57 465 91
rect 499 57 508 91
rect 542 151 551 185
rect 585 151 593 185
rect 714 185 766 209
rect 542 111 593 151
rect 542 77 551 111
rect 585 77 593 111
rect 542 61 593 77
rect 627 159 680 175
rect 627 125 637 159
rect 671 125 680 159
rect 627 91 680 125
rect 456 17 508 57
rect 627 57 637 91
rect 671 57 680 91
rect 714 151 723 185
rect 757 151 766 185
rect 886 185 937 209
rect 714 111 766 151
rect 714 77 723 111
rect 757 77 766 111
rect 714 61 766 77
rect 800 159 852 175
rect 800 125 809 159
rect 843 125 852 159
rect 800 91 852 125
rect 627 17 680 57
rect 800 57 809 91
rect 843 57 852 91
rect 886 151 895 185
rect 929 151 937 185
rect 886 111 937 151
rect 886 77 895 111
rect 929 77 937 111
rect 886 61 937 77
rect 971 159 1031 175
rect 971 125 981 159
rect 1015 125 1031 159
rect 971 91 1031 125
rect 800 17 852 57
rect 971 57 981 91
rect 1015 57 1031 91
rect 971 17 1031 57
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 buf_8
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6027014
string GDS_START 6017362
<< end >>
