magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 1 157 490 241
rect 1 49 671 157
rect 0 0 672 49
<< scnmos >>
rect 98 47 128 215
rect 184 47 214 215
rect 284 47 314 215
rect 384 47 414 215
rect 486 47 516 131
rect 558 47 588 131
<< scpmoshvt >>
rect 98 367 128 619
rect 184 367 214 619
rect 270 367 300 619
rect 356 367 386 619
rect 479 377 509 505
rect 557 377 587 505
<< ndiff >>
rect 27 203 98 215
rect 27 169 39 203
rect 73 169 98 203
rect 27 93 98 169
rect 27 59 39 93
rect 73 59 98 93
rect 27 47 98 59
rect 128 203 184 215
rect 128 169 139 203
rect 173 169 184 203
rect 128 101 184 169
rect 128 67 139 101
rect 173 67 184 101
rect 128 47 184 67
rect 214 186 284 215
rect 214 152 239 186
rect 273 152 284 186
rect 214 47 284 152
rect 314 203 384 215
rect 314 169 339 203
rect 373 169 384 203
rect 314 101 384 169
rect 314 67 339 101
rect 373 67 384 101
rect 314 47 384 67
rect 414 131 464 215
rect 414 93 486 131
rect 414 59 439 93
rect 473 59 486 93
rect 414 47 486 59
rect 516 47 558 131
rect 588 110 645 131
rect 588 76 599 110
rect 633 76 645 110
rect 588 47 645 76
<< pdiff >>
rect 27 607 98 619
rect 27 573 39 607
rect 73 573 98 607
rect 27 510 98 573
rect 27 476 39 510
rect 73 476 98 510
rect 27 413 98 476
rect 27 379 39 413
rect 73 379 98 413
rect 27 367 98 379
rect 128 599 184 619
rect 128 565 139 599
rect 173 565 184 599
rect 128 506 184 565
rect 128 472 139 506
rect 173 472 184 506
rect 128 413 184 472
rect 128 379 139 413
rect 173 379 184 413
rect 128 367 184 379
rect 214 531 270 619
rect 214 497 225 531
rect 259 497 270 531
rect 214 413 270 497
rect 214 379 225 413
rect 259 379 270 413
rect 214 367 270 379
rect 300 599 356 619
rect 300 565 311 599
rect 345 565 356 599
rect 300 506 356 565
rect 300 472 311 506
rect 345 472 356 506
rect 300 413 356 472
rect 300 379 311 413
rect 345 379 356 413
rect 300 367 356 379
rect 386 607 457 619
rect 386 573 411 607
rect 445 573 457 607
rect 386 510 457 573
rect 386 476 411 510
rect 445 505 457 510
rect 445 476 479 505
rect 386 413 479 476
rect 386 379 411 413
rect 445 379 479 413
rect 386 377 479 379
rect 509 377 557 505
rect 587 493 644 505
rect 587 459 598 493
rect 632 459 644 493
rect 587 423 644 459
rect 587 389 598 423
rect 632 389 644 423
rect 587 377 644 389
rect 386 367 457 377
<< ndiffc >>
rect 39 169 73 203
rect 39 59 73 93
rect 139 169 173 203
rect 139 67 173 101
rect 239 152 273 186
rect 339 169 373 203
rect 339 67 373 101
rect 439 59 473 93
rect 599 76 633 110
<< pdiffc >>
rect 39 573 73 607
rect 39 476 73 510
rect 39 379 73 413
rect 139 565 173 599
rect 139 472 173 506
rect 139 379 173 413
rect 225 497 259 531
rect 225 379 259 413
rect 311 565 345 599
rect 311 472 345 506
rect 311 379 345 413
rect 411 573 445 607
rect 411 476 445 510
rect 411 379 445 413
rect 598 459 632 493
rect 598 389 632 423
<< poly >>
rect 98 619 128 645
rect 184 619 214 645
rect 270 619 300 645
rect 356 619 386 645
rect 479 505 509 531
rect 557 505 587 531
rect 98 283 128 367
rect 184 283 214 367
rect 270 283 300 367
rect 356 319 386 367
rect 356 303 431 319
rect 356 283 381 303
rect 98 269 381 283
rect 415 269 431 303
rect 98 253 431 269
rect 479 277 509 377
rect 557 355 587 377
rect 557 325 588 355
rect 558 277 588 325
rect 479 261 588 277
rect 98 215 128 253
rect 184 215 214 253
rect 284 215 314 253
rect 384 215 414 253
rect 479 227 511 261
rect 545 227 588 261
rect 479 211 588 227
rect 486 131 516 211
rect 558 131 588 211
rect 98 21 128 47
rect 184 21 214 47
rect 284 21 314 47
rect 384 21 414 47
rect 486 21 516 47
rect 558 21 588 47
<< polycont >>
rect 381 269 415 303
rect 511 227 545 261
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 607 89 649
rect 23 573 39 607
rect 73 573 89 607
rect 23 510 89 573
rect 23 476 39 510
rect 73 476 89 510
rect 23 413 89 476
rect 23 379 39 413
rect 73 379 89 413
rect 23 363 89 379
rect 123 599 361 615
rect 123 565 139 599
rect 173 581 311 599
rect 123 506 173 565
rect 345 565 361 599
rect 123 472 139 506
rect 123 413 173 472
rect 123 379 139 413
rect 123 363 173 379
rect 209 531 275 547
rect 209 497 225 531
rect 259 497 275 531
rect 209 413 275 497
rect 209 379 225 413
rect 259 379 275 413
rect 209 310 275 379
rect 311 506 361 565
rect 345 472 361 506
rect 311 413 361 472
rect 345 379 361 413
rect 311 363 361 379
rect 395 607 461 649
rect 395 573 411 607
rect 445 573 461 607
rect 395 510 461 573
rect 395 476 411 510
rect 445 476 461 510
rect 395 413 461 476
rect 395 379 411 413
rect 445 379 461 413
rect 395 363 461 379
rect 223 219 275 310
rect 365 303 457 319
rect 365 269 381 303
rect 415 269 457 303
rect 365 253 457 269
rect 23 203 89 219
rect 23 169 39 203
rect 73 169 89 203
rect 23 93 89 169
rect 23 59 39 93
rect 73 59 89 93
rect 23 17 89 59
rect 123 203 189 219
rect 123 169 139 203
rect 173 169 189 203
rect 123 101 189 169
rect 223 186 289 219
rect 223 152 239 186
rect 273 152 289 186
rect 223 119 289 152
rect 323 203 389 219
rect 323 169 339 203
rect 373 169 389 203
rect 123 67 139 101
rect 173 85 189 101
rect 323 101 389 169
rect 423 177 457 253
rect 495 261 561 578
rect 495 227 511 261
rect 545 227 561 261
rect 495 211 561 227
rect 598 493 649 509
rect 632 459 649 493
rect 598 423 649 459
rect 632 389 649 423
rect 598 177 649 389
rect 423 143 649 177
rect 583 110 649 143
rect 323 85 339 101
rect 173 67 339 85
rect 373 67 389 101
rect 123 51 389 67
rect 423 93 489 109
rect 423 59 439 93
rect 473 59 489 93
rect 423 17 489 59
rect 583 76 599 110
rect 633 76 649 110
rect 583 51 649 76
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 buflp_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6968572
string GDS_START 6962350
<< end >>
