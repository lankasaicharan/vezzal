magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
rect 167 327 1396 331
rect 167 309 335 327
<< pwell >>
rect 24 157 298 245
rect 1043 241 1441 271
rect 838 157 1631 241
rect 24 49 1631 157
rect 0 0 1632 49
<< scnmos >>
rect 103 135 133 219
rect 189 135 219 219
rect 438 47 468 131
rect 524 47 554 131
rect 596 47 626 131
rect 704 47 734 131
rect 812 47 842 131
rect 917 47 947 215
rect 1122 161 1152 245
rect 1332 77 1362 245
rect 1522 47 1552 215
<< scpmoshvt >>
rect 87 407 117 535
rect 189 407 219 535
rect 416 483 446 611
rect 554 483 584 611
rect 626 483 656 611
rect 734 483 764 567
rect 806 483 836 567
rect 960 363 990 615
rect 1179 365 1209 493
rect 1277 365 1307 617
rect 1522 367 1552 619
<< ndiff >>
rect 50 191 103 219
rect 50 157 58 191
rect 92 157 103 191
rect 50 135 103 157
rect 133 191 189 219
rect 133 157 144 191
rect 178 157 189 191
rect 133 135 189 157
rect 219 207 272 219
rect 219 173 230 207
rect 264 173 272 207
rect 219 135 272 173
rect 1069 221 1122 245
rect 864 203 917 215
rect 864 169 872 203
rect 906 169 917 203
rect 864 131 917 169
rect 385 107 438 131
rect 385 73 393 107
rect 427 73 438 107
rect 385 47 438 73
rect 468 97 524 131
rect 468 63 479 97
rect 513 63 524 97
rect 468 47 524 63
rect 554 47 596 131
rect 626 93 704 131
rect 626 59 649 93
rect 683 59 704 93
rect 626 47 704 59
rect 734 47 812 131
rect 842 93 917 131
rect 842 59 864 93
rect 898 59 917 93
rect 842 47 917 59
rect 947 203 1000 215
rect 947 169 958 203
rect 992 169 1000 203
rect 947 101 1000 169
rect 1069 187 1077 221
rect 1111 187 1122 221
rect 1069 161 1122 187
rect 1152 165 1332 245
rect 1152 161 1217 165
rect 947 67 958 101
rect 992 67 1000 101
rect 1209 131 1217 161
rect 1251 131 1332 165
rect 1209 77 1332 131
rect 1362 233 1415 245
rect 1362 199 1373 233
rect 1407 199 1415 233
rect 1362 77 1415 199
rect 1469 93 1522 215
rect 947 47 1000 67
rect 1469 59 1477 93
rect 1511 59 1522 93
rect 1469 47 1522 59
rect 1552 203 1605 215
rect 1552 169 1563 203
rect 1597 169 1605 203
rect 1552 101 1605 169
rect 1552 67 1563 101
rect 1597 67 1605 101
rect 1552 47 1605 67
<< pdiff >>
rect 363 599 416 611
rect 363 565 371 599
rect 405 565 416 599
rect 34 523 87 535
rect 34 489 42 523
rect 76 489 87 523
rect 34 453 87 489
rect 34 419 42 453
rect 76 419 87 453
rect 34 407 87 419
rect 117 527 189 535
rect 117 493 144 527
rect 178 493 189 527
rect 117 407 189 493
rect 219 407 299 535
rect 363 531 416 565
rect 363 497 371 531
rect 405 497 416 531
rect 363 483 416 497
rect 446 603 554 611
rect 446 569 486 603
rect 520 569 554 603
rect 446 483 554 569
rect 584 483 626 611
rect 656 597 709 611
rect 656 563 667 597
rect 701 567 709 597
rect 904 603 960 615
rect 904 569 912 603
rect 946 569 960 603
rect 904 567 960 569
rect 701 563 734 567
rect 656 529 734 563
rect 656 495 689 529
rect 723 495 734 529
rect 656 483 734 495
rect 764 483 806 567
rect 836 541 960 567
rect 836 507 847 541
rect 881 535 960 541
rect 881 507 915 535
rect 836 501 915 507
rect 949 501 960 535
rect 836 483 960 501
rect 241 387 299 407
rect 241 353 253 387
rect 287 353 299 387
rect 241 345 299 353
rect 904 363 960 483
rect 990 599 1043 615
rect 990 565 1001 599
rect 1035 565 1043 599
rect 990 512 1043 565
rect 1224 605 1277 617
rect 1224 571 1232 605
rect 1266 571 1277 605
rect 990 478 1001 512
rect 1035 478 1043 512
rect 1224 505 1277 571
rect 1224 493 1232 505
rect 990 423 1043 478
rect 990 389 1001 423
rect 1035 389 1043 423
rect 990 363 1043 389
rect 1126 481 1179 493
rect 1126 447 1134 481
rect 1168 447 1179 481
rect 1126 411 1179 447
rect 1126 377 1134 411
rect 1168 377 1179 411
rect 1126 365 1179 377
rect 1209 471 1232 493
rect 1266 471 1277 505
rect 1209 411 1277 471
rect 1209 377 1225 411
rect 1259 377 1277 411
rect 1209 365 1277 377
rect 1307 599 1360 617
rect 1307 565 1318 599
rect 1352 565 1360 599
rect 1307 503 1360 565
rect 1307 469 1318 503
rect 1352 469 1360 503
rect 1307 411 1360 469
rect 1307 377 1318 411
rect 1352 377 1360 411
rect 1307 365 1360 377
rect 1469 607 1522 619
rect 1469 573 1477 607
rect 1511 573 1522 607
rect 1469 539 1522 573
rect 1469 505 1477 539
rect 1511 505 1522 539
rect 1469 413 1522 505
rect 1469 379 1477 413
rect 1511 379 1522 413
rect 1469 367 1522 379
rect 1552 599 1605 619
rect 1552 565 1563 599
rect 1597 565 1605 599
rect 1552 503 1605 565
rect 1552 469 1563 503
rect 1597 469 1605 503
rect 1552 413 1605 469
rect 1552 379 1563 413
rect 1597 379 1605 413
rect 1552 367 1605 379
<< ndiffc >>
rect 58 157 92 191
rect 144 157 178 191
rect 230 173 264 207
rect 872 169 906 203
rect 393 73 427 107
rect 479 63 513 97
rect 649 59 683 93
rect 864 59 898 93
rect 958 169 992 203
rect 1077 187 1111 221
rect 958 67 992 101
rect 1217 131 1251 165
rect 1373 199 1407 233
rect 1477 59 1511 93
rect 1563 169 1597 203
rect 1563 67 1597 101
<< pdiffc >>
rect 371 565 405 599
rect 42 489 76 523
rect 42 419 76 453
rect 144 493 178 527
rect 371 497 405 531
rect 486 569 520 603
rect 667 563 701 597
rect 912 569 946 603
rect 689 495 723 529
rect 847 507 881 541
rect 915 501 949 535
rect 253 353 287 387
rect 1001 565 1035 599
rect 1232 571 1266 605
rect 1001 478 1035 512
rect 1001 389 1035 423
rect 1134 447 1168 481
rect 1134 377 1168 411
rect 1232 471 1266 505
rect 1225 377 1259 411
rect 1318 565 1352 599
rect 1318 469 1352 503
rect 1318 377 1352 411
rect 1477 573 1511 607
rect 1477 505 1511 539
rect 1477 379 1511 413
rect 1563 565 1597 599
rect 1563 469 1597 503
rect 1563 379 1597 413
<< poly >>
rect 416 611 446 637
rect 554 611 584 637
rect 626 611 656 637
rect 960 615 990 641
rect 1277 617 1307 643
rect 1522 619 1552 645
rect 87 535 117 561
rect 189 535 219 561
rect 734 567 764 593
rect 806 567 836 593
rect 87 375 117 407
rect 75 359 141 375
rect 75 325 91 359
rect 125 325 141 359
rect 75 291 141 325
rect 75 257 91 291
rect 125 257 141 291
rect 75 241 141 257
rect 189 271 219 407
rect 416 373 446 483
rect 554 451 584 483
rect 374 357 446 373
rect 374 323 390 357
rect 424 343 446 357
rect 488 435 584 451
rect 488 401 504 435
rect 538 421 584 435
rect 626 451 656 483
rect 626 435 692 451
rect 538 401 554 421
rect 488 367 554 401
rect 626 401 642 435
rect 676 401 692 435
rect 626 385 692 401
rect 424 323 440 343
rect 374 289 440 323
rect 488 333 504 367
rect 538 333 554 367
rect 734 337 764 483
rect 806 451 836 483
rect 806 435 872 451
rect 806 401 822 435
rect 856 401 872 435
rect 806 385 872 401
rect 488 317 554 333
rect 518 307 554 317
rect 189 241 317 271
rect 103 219 133 241
rect 189 219 219 241
rect 103 109 133 135
rect 189 109 219 135
rect 287 113 317 241
rect 374 255 390 289
rect 424 269 440 289
rect 424 255 468 269
rect 374 239 468 255
rect 438 131 468 239
rect 524 131 554 307
rect 596 321 764 337
rect 596 287 612 321
rect 646 307 764 321
rect 646 287 662 307
rect 596 253 662 287
rect 596 219 612 253
rect 646 219 662 253
rect 596 203 662 219
rect 704 203 770 219
rect 596 131 626 203
rect 704 169 720 203
rect 754 169 770 203
rect 704 153 770 169
rect 704 131 734 153
rect 812 131 842 385
rect 1179 493 1209 519
rect 960 321 990 363
rect 917 305 990 321
rect 917 271 933 305
rect 967 271 990 305
rect 1179 297 1209 365
rect 1277 333 1307 365
rect 917 255 990 271
rect 1122 267 1209 297
rect 1257 317 1362 333
rect 1257 283 1273 317
rect 1307 283 1362 317
rect 1522 303 1552 367
rect 1257 267 1362 283
rect 917 215 947 255
rect 1122 245 1152 267
rect 1332 245 1362 267
rect 1459 287 1552 303
rect 1459 253 1475 287
rect 1509 253 1552 287
rect 287 97 353 113
rect 287 63 303 97
rect 337 63 353 97
rect 287 47 353 63
rect 1122 135 1152 161
rect 1115 119 1181 135
rect 1115 85 1131 119
rect 1165 85 1181 119
rect 1115 69 1181 85
rect 1459 237 1552 253
rect 1522 215 1552 237
rect 1332 51 1362 77
rect 438 21 468 47
rect 524 21 554 47
rect 596 21 626 47
rect 704 21 734 47
rect 812 21 842 47
rect 917 21 947 47
rect 1522 21 1552 47
<< polycont >>
rect 91 325 125 359
rect 91 257 125 291
rect 390 323 424 357
rect 504 401 538 435
rect 642 401 676 435
rect 504 333 538 367
rect 822 401 856 435
rect 390 255 424 289
rect 612 287 646 321
rect 612 219 646 253
rect 720 169 754 203
rect 933 271 967 305
rect 1273 283 1307 317
rect 1475 253 1509 287
rect 303 63 337 97
rect 1131 85 1165 119
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 21 523 92 539
rect 21 489 42 523
rect 76 489 92 523
rect 128 527 194 649
rect 128 493 144 527
rect 178 493 194 527
rect 128 491 194 493
rect 355 599 421 615
rect 355 565 371 599
rect 405 565 421 599
rect 470 603 536 649
rect 470 569 486 603
rect 520 569 536 603
rect 470 565 536 569
rect 663 597 746 613
rect 355 531 421 565
rect 355 497 371 531
rect 405 527 421 531
rect 663 563 667 597
rect 701 563 746 597
rect 663 529 746 563
rect 405 497 629 527
rect 355 491 629 497
rect 21 457 92 489
rect 21 453 554 457
rect 21 419 42 453
rect 76 435 554 453
rect 76 423 504 435
rect 76 419 92 423
rect 21 409 92 419
rect 21 207 55 409
rect 488 401 504 423
rect 538 401 554 435
rect 214 387 440 389
rect 91 359 180 375
rect 125 325 180 359
rect 91 291 180 325
rect 125 257 180 291
rect 91 241 180 257
rect 214 353 253 387
rect 287 357 440 387
rect 287 353 390 357
rect 214 323 390 353
rect 424 323 440 357
rect 214 289 440 323
rect 488 367 554 401
rect 595 445 629 491
rect 663 495 689 529
rect 723 513 746 529
rect 831 603 951 649
rect 831 569 912 603
rect 946 569 951 603
rect 831 541 951 569
rect 723 495 786 513
rect 663 479 786 495
rect 831 507 847 541
rect 881 535 951 541
rect 881 507 915 535
rect 831 501 915 507
rect 949 501 951 535
rect 831 485 951 501
rect 985 599 1048 615
rect 985 565 1001 599
rect 1035 565 1048 599
rect 985 512 1048 565
rect 595 435 716 445
rect 595 401 642 435
rect 676 401 716 435
rect 595 385 716 401
rect 488 333 504 367
rect 538 333 554 367
rect 488 317 554 333
rect 596 321 648 337
rect 214 255 390 289
rect 424 273 440 289
rect 596 287 612 321
rect 646 287 648 321
rect 596 273 648 287
rect 424 255 648 273
rect 214 253 648 255
rect 214 239 612 253
rect 214 207 303 239
rect 21 191 101 207
rect 21 157 58 191
rect 92 157 101 191
rect 21 139 101 157
rect 135 191 178 207
rect 135 157 144 191
rect 214 173 230 207
rect 264 173 303 207
rect 596 219 612 239
rect 646 219 648 253
rect 596 203 648 219
rect 682 219 716 385
rect 752 349 786 479
rect 985 478 1001 512
rect 1035 478 1048 512
rect 1218 605 1270 649
rect 1218 571 1232 605
rect 1266 571 1270 605
rect 1218 505 1270 571
rect 985 451 1048 478
rect 820 435 1048 451
rect 820 401 822 435
rect 856 423 1048 435
rect 856 401 1001 423
rect 820 389 1001 401
rect 1035 389 1048 423
rect 820 385 1048 389
rect 1118 481 1184 497
rect 1118 447 1134 481
rect 1168 447 1184 481
rect 1118 411 1184 447
rect 752 315 824 349
rect 790 289 824 315
rect 917 305 969 321
rect 917 289 933 305
rect 790 271 933 289
rect 967 271 969 305
rect 790 255 969 271
rect 682 203 756 219
rect 214 169 303 173
rect 682 169 720 203
rect 754 169 756 203
rect 135 17 178 157
rect 389 135 756 169
rect 212 97 355 135
rect 212 63 303 97
rect 337 63 355 97
rect 212 51 355 63
rect 389 107 427 135
rect 389 73 393 107
rect 389 57 427 73
rect 463 97 529 101
rect 790 97 824 255
rect 1003 219 1039 385
rect 1118 377 1134 411
rect 1168 377 1184 411
rect 1118 327 1184 377
rect 1218 471 1232 505
rect 1266 471 1270 505
rect 1218 411 1270 471
rect 1218 377 1225 411
rect 1259 377 1270 411
rect 1218 361 1270 377
rect 1318 599 1425 615
rect 1352 565 1425 599
rect 1318 503 1425 565
rect 1352 469 1425 503
rect 1318 411 1425 469
rect 1352 377 1425 411
rect 1318 361 1425 377
rect 1461 607 1527 649
rect 1461 573 1477 607
rect 1511 573 1527 607
rect 1461 539 1527 573
rect 1461 505 1477 539
rect 1511 505 1527 539
rect 1461 413 1527 505
rect 1461 379 1477 413
rect 1511 379 1527 413
rect 1461 363 1527 379
rect 1561 599 1613 615
rect 1561 565 1563 599
rect 1597 565 1613 599
rect 1561 503 1613 565
rect 1561 469 1563 503
rect 1597 469 1613 503
rect 1561 413 1613 469
rect 1561 379 1563 413
rect 1597 379 1613 413
rect 1118 317 1323 327
rect 463 63 479 97
rect 513 63 529 97
rect 463 17 529 63
rect 633 93 824 97
rect 633 59 649 93
rect 683 59 824 93
rect 633 55 824 59
rect 858 203 920 219
rect 858 169 872 203
rect 906 169 920 203
rect 858 93 920 169
rect 858 59 864 93
rect 898 59 920 93
rect 858 17 920 59
rect 954 203 1039 219
rect 954 169 958 203
rect 992 169 1039 203
rect 1073 283 1273 317
rect 1307 283 1323 317
rect 1073 221 1111 283
rect 1073 187 1077 221
rect 1073 171 1111 187
rect 1145 215 1323 249
rect 954 135 1039 169
rect 1145 135 1179 215
rect 954 119 1179 135
rect 954 101 1131 119
rect 954 67 958 101
rect 992 85 1131 101
rect 1165 85 1179 119
rect 992 67 1179 85
rect 954 51 1179 67
rect 1213 165 1255 181
rect 1213 131 1217 165
rect 1251 131 1255 165
rect 1289 165 1323 215
rect 1357 233 1425 361
rect 1357 199 1373 233
rect 1407 199 1425 233
rect 1459 287 1525 303
rect 1459 253 1475 287
rect 1509 253 1525 287
rect 1459 165 1525 253
rect 1289 131 1525 165
rect 1561 203 1613 379
rect 1561 169 1563 203
rect 1597 169 1613 203
rect 1213 17 1255 131
rect 1561 101 1613 169
rect 1461 93 1527 97
rect 1461 59 1477 93
rect 1511 59 1527 93
rect 1461 17 1527 59
rect 1561 67 1563 101
rect 1597 67 1613 101
rect 1561 51 1613 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlxbn_1
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1375 390 1409 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1375 464 1409 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1375 538 1409 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5939342
string GDS_START 5925726
<< end >>
