magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
<< pwell >>
rect 452 241 2055 259
rect 1 49 2055 241
rect 0 0 2112 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 252 47 282 215
rect 338 47 368 215
rect 531 65 561 233
rect 617 65 647 233
rect 703 65 733 233
rect 789 65 819 233
rect 891 65 921 233
rect 977 65 1007 233
rect 1063 65 1093 233
rect 1149 65 1179 233
rect 1344 65 1374 233
rect 1430 65 1460 233
rect 1516 65 1546 233
rect 1602 65 1632 233
rect 1688 65 1718 233
rect 1774 65 1804 233
rect 1860 65 1890 233
rect 1946 65 1976 233
<< scpmoshvt >>
rect 83 367 113 619
rect 169 367 199 619
rect 255 367 285 619
rect 341 367 371 619
rect 427 367 457 619
rect 517 367 547 619
rect 603 367 633 619
rect 775 367 805 619
rect 861 367 891 619
rect 947 367 977 619
rect 1033 367 1063 619
rect 1151 367 1181 619
rect 1237 367 1267 619
rect 1323 367 1353 619
rect 1409 367 1439 619
rect 1599 367 1629 619
rect 1685 367 1715 619
rect 1771 367 1801 619
rect 1857 367 1887 619
rect 1943 367 1973 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 93 80 169
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 192 166 215
rect 110 158 121 192
rect 155 158 166 192
rect 110 101 166 158
rect 110 67 121 101
rect 155 67 166 101
rect 110 47 166 67
rect 196 126 252 215
rect 196 92 207 126
rect 241 92 252 126
rect 196 47 252 92
rect 282 192 338 215
rect 282 158 293 192
rect 327 158 338 192
rect 282 101 338 158
rect 282 67 293 101
rect 327 67 338 101
rect 282 47 338 67
rect 368 118 421 215
rect 368 84 379 118
rect 413 84 421 118
rect 368 47 421 84
rect 478 111 531 233
rect 478 77 486 111
rect 520 77 531 111
rect 478 65 531 77
rect 561 201 617 233
rect 561 167 572 201
rect 606 167 617 201
rect 561 65 617 167
rect 647 111 703 233
rect 647 77 658 111
rect 692 77 703 111
rect 647 65 703 77
rect 733 225 789 233
rect 733 191 744 225
rect 778 191 789 225
rect 733 153 789 191
rect 733 119 744 153
rect 778 119 789 153
rect 733 65 789 119
rect 819 179 891 233
rect 819 145 846 179
rect 880 145 891 179
rect 819 107 891 145
rect 819 73 846 107
rect 880 73 891 107
rect 819 65 891 73
rect 921 169 977 233
rect 921 135 932 169
rect 966 135 977 169
rect 921 65 977 135
rect 1007 111 1063 233
rect 1007 77 1018 111
rect 1052 77 1063 111
rect 1007 65 1063 77
rect 1093 201 1149 233
rect 1093 167 1104 201
rect 1138 167 1149 201
rect 1093 65 1149 167
rect 1179 111 1232 233
rect 1179 77 1190 111
rect 1224 77 1232 111
rect 1179 65 1232 77
rect 1291 113 1344 233
rect 1291 79 1299 113
rect 1333 79 1344 113
rect 1291 65 1344 79
rect 1374 225 1430 233
rect 1374 191 1385 225
rect 1419 191 1430 225
rect 1374 157 1430 191
rect 1374 123 1385 157
rect 1419 123 1430 157
rect 1374 65 1430 123
rect 1460 113 1516 233
rect 1460 79 1471 113
rect 1505 79 1516 113
rect 1460 65 1516 79
rect 1546 225 1602 233
rect 1546 191 1557 225
rect 1591 191 1602 225
rect 1546 157 1602 191
rect 1546 123 1557 157
rect 1591 123 1602 157
rect 1546 65 1602 123
rect 1632 190 1688 233
rect 1632 156 1643 190
rect 1677 156 1688 190
rect 1632 111 1688 156
rect 1632 77 1643 111
rect 1677 77 1688 111
rect 1632 65 1688 77
rect 1718 130 1774 233
rect 1718 96 1729 130
rect 1763 96 1774 130
rect 1718 65 1774 96
rect 1804 192 1860 233
rect 1804 158 1815 192
rect 1849 158 1860 192
rect 1804 113 1860 158
rect 1804 79 1815 113
rect 1849 79 1860 113
rect 1804 65 1860 79
rect 1890 130 1946 233
rect 1890 96 1901 130
rect 1935 96 1946 130
rect 1890 65 1946 96
rect 1976 192 2029 233
rect 1976 158 1987 192
rect 2021 158 2029 192
rect 1976 113 2029 158
rect 1976 79 1987 113
rect 2021 79 2029 113
rect 1976 65 2029 79
<< pdiff >>
rect 30 599 83 619
rect 30 565 38 599
rect 72 565 83 599
rect 30 509 83 565
rect 30 475 38 509
rect 72 475 83 509
rect 30 415 83 475
rect 30 381 38 415
rect 72 381 83 415
rect 30 367 83 381
rect 113 547 169 619
rect 113 513 124 547
rect 158 513 169 547
rect 113 479 169 513
rect 113 445 124 479
rect 158 445 169 479
rect 113 411 169 445
rect 113 377 124 411
rect 158 377 169 411
rect 113 367 169 377
rect 199 599 255 619
rect 199 565 210 599
rect 244 565 255 599
rect 199 517 255 565
rect 199 483 210 517
rect 244 483 255 517
rect 199 442 255 483
rect 199 408 210 442
rect 244 408 255 442
rect 199 367 255 408
rect 285 547 341 619
rect 285 513 296 547
rect 330 513 341 547
rect 285 479 341 513
rect 285 445 296 479
rect 330 445 341 479
rect 285 411 341 445
rect 285 377 296 411
rect 330 377 341 411
rect 285 367 341 377
rect 371 599 427 619
rect 371 565 382 599
rect 416 565 427 599
rect 371 471 427 565
rect 371 437 382 471
rect 416 437 427 471
rect 371 367 427 437
rect 457 611 517 619
rect 457 577 472 611
rect 506 577 517 611
rect 457 541 517 577
rect 457 507 472 541
rect 506 507 517 541
rect 457 367 517 507
rect 547 599 603 619
rect 547 565 558 599
rect 592 565 603 599
rect 547 471 603 565
rect 547 437 558 471
rect 592 437 603 471
rect 547 367 603 437
rect 633 611 775 619
rect 633 577 648 611
rect 682 577 716 611
rect 750 577 775 611
rect 633 530 775 577
rect 633 496 648 530
rect 682 496 716 530
rect 750 496 775 530
rect 633 367 775 496
rect 805 611 861 619
rect 805 577 816 611
rect 850 577 861 611
rect 805 538 861 577
rect 805 504 816 538
rect 850 504 861 538
rect 805 461 861 504
rect 805 427 816 461
rect 850 427 861 461
rect 805 367 861 427
rect 891 611 947 619
rect 891 577 902 611
rect 936 577 947 611
rect 891 541 947 577
rect 891 507 902 541
rect 936 507 947 541
rect 891 367 947 507
rect 977 599 1033 619
rect 977 565 988 599
rect 1022 565 1033 599
rect 977 503 1033 565
rect 977 469 988 503
rect 1022 469 1033 503
rect 977 413 1033 469
rect 977 379 988 413
rect 1022 379 1033 413
rect 977 367 1033 379
rect 1063 607 1151 619
rect 1063 573 1090 607
rect 1124 573 1151 607
rect 1063 529 1151 573
rect 1063 495 1090 529
rect 1124 495 1151 529
rect 1063 455 1151 495
rect 1063 421 1090 455
rect 1124 421 1151 455
rect 1063 367 1151 421
rect 1181 599 1237 619
rect 1181 565 1192 599
rect 1226 565 1237 599
rect 1181 509 1237 565
rect 1181 475 1192 509
rect 1226 475 1237 509
rect 1181 413 1237 475
rect 1181 379 1192 413
rect 1226 379 1237 413
rect 1181 367 1237 379
rect 1267 607 1323 619
rect 1267 573 1278 607
rect 1312 573 1323 607
rect 1267 529 1323 573
rect 1267 495 1278 529
rect 1312 495 1323 529
rect 1267 455 1323 495
rect 1267 421 1278 455
rect 1312 421 1323 455
rect 1267 367 1323 421
rect 1353 599 1409 619
rect 1353 565 1364 599
rect 1398 565 1409 599
rect 1353 509 1409 565
rect 1353 475 1364 509
rect 1398 475 1409 509
rect 1353 413 1409 475
rect 1353 379 1364 413
rect 1398 379 1409 413
rect 1353 367 1409 379
rect 1439 607 1599 619
rect 1439 573 1450 607
rect 1484 573 1554 607
rect 1588 573 1599 607
rect 1439 529 1599 573
rect 1439 495 1450 529
rect 1484 495 1554 529
rect 1588 495 1599 529
rect 1439 455 1599 495
rect 1439 421 1450 455
rect 1484 421 1554 455
rect 1588 421 1599 455
rect 1439 367 1599 421
rect 1629 599 1685 619
rect 1629 565 1640 599
rect 1674 565 1685 599
rect 1629 509 1685 565
rect 1629 475 1640 509
rect 1674 475 1685 509
rect 1629 413 1685 475
rect 1629 379 1640 413
rect 1674 379 1685 413
rect 1629 367 1685 379
rect 1715 607 1771 619
rect 1715 573 1726 607
rect 1760 573 1771 607
rect 1715 529 1771 573
rect 1715 495 1726 529
rect 1760 495 1771 529
rect 1715 455 1771 495
rect 1715 421 1726 455
rect 1760 421 1771 455
rect 1715 367 1771 421
rect 1801 599 1857 619
rect 1801 565 1812 599
rect 1846 565 1857 599
rect 1801 509 1857 565
rect 1801 475 1812 509
rect 1846 475 1857 509
rect 1801 413 1857 475
rect 1801 379 1812 413
rect 1846 379 1857 413
rect 1801 367 1857 379
rect 1887 607 1943 619
rect 1887 573 1898 607
rect 1932 573 1943 607
rect 1887 529 1943 573
rect 1887 495 1898 529
rect 1932 495 1943 529
rect 1887 455 1943 495
rect 1887 421 1898 455
rect 1932 421 1943 455
rect 1887 367 1943 421
rect 1973 599 2026 619
rect 1973 565 1984 599
rect 2018 565 2026 599
rect 1973 509 2026 565
rect 1973 475 1984 509
rect 2018 475 2026 509
rect 1973 413 2026 475
rect 1973 379 1984 413
rect 2018 379 2026 413
rect 1973 367 2026 379
<< ndiffc >>
rect 35 169 69 203
rect 35 59 69 93
rect 121 158 155 192
rect 121 67 155 101
rect 207 92 241 126
rect 293 158 327 192
rect 293 67 327 101
rect 379 84 413 118
rect 486 77 520 111
rect 572 167 606 201
rect 658 77 692 111
rect 744 191 778 225
rect 744 119 778 153
rect 846 145 880 179
rect 846 73 880 107
rect 932 135 966 169
rect 1018 77 1052 111
rect 1104 167 1138 201
rect 1190 77 1224 111
rect 1299 79 1333 113
rect 1385 191 1419 225
rect 1385 123 1419 157
rect 1471 79 1505 113
rect 1557 191 1591 225
rect 1557 123 1591 157
rect 1643 156 1677 190
rect 1643 77 1677 111
rect 1729 96 1763 130
rect 1815 158 1849 192
rect 1815 79 1849 113
rect 1901 96 1935 130
rect 1987 158 2021 192
rect 1987 79 2021 113
<< pdiffc >>
rect 38 565 72 599
rect 38 475 72 509
rect 38 381 72 415
rect 124 513 158 547
rect 124 445 158 479
rect 124 377 158 411
rect 210 565 244 599
rect 210 483 244 517
rect 210 408 244 442
rect 296 513 330 547
rect 296 445 330 479
rect 296 377 330 411
rect 382 565 416 599
rect 382 437 416 471
rect 472 577 506 611
rect 472 507 506 541
rect 558 565 592 599
rect 558 437 592 471
rect 648 577 682 611
rect 716 577 750 611
rect 648 496 682 530
rect 716 496 750 530
rect 816 577 850 611
rect 816 504 850 538
rect 816 427 850 461
rect 902 577 936 611
rect 902 507 936 541
rect 988 565 1022 599
rect 988 469 1022 503
rect 988 379 1022 413
rect 1090 573 1124 607
rect 1090 495 1124 529
rect 1090 421 1124 455
rect 1192 565 1226 599
rect 1192 475 1226 509
rect 1192 379 1226 413
rect 1278 573 1312 607
rect 1278 495 1312 529
rect 1278 421 1312 455
rect 1364 565 1398 599
rect 1364 475 1398 509
rect 1364 379 1398 413
rect 1450 573 1484 607
rect 1554 573 1588 607
rect 1450 495 1484 529
rect 1554 495 1588 529
rect 1450 421 1484 455
rect 1554 421 1588 455
rect 1640 565 1674 599
rect 1640 475 1674 509
rect 1640 379 1674 413
rect 1726 573 1760 607
rect 1726 495 1760 529
rect 1726 421 1760 455
rect 1812 565 1846 599
rect 1812 475 1846 509
rect 1812 379 1846 413
rect 1898 573 1932 607
rect 1898 495 1932 529
rect 1898 421 1932 455
rect 1984 565 2018 599
rect 1984 475 2018 509
rect 1984 379 2018 413
<< poly >>
rect 83 619 113 645
rect 169 619 199 645
rect 255 619 285 645
rect 341 619 371 645
rect 427 619 457 645
rect 517 619 547 645
rect 603 619 633 645
rect 775 619 805 645
rect 861 619 891 645
rect 947 619 977 645
rect 1033 619 1063 645
rect 1151 619 1181 645
rect 1237 619 1267 645
rect 1323 619 1353 645
rect 1409 619 1439 645
rect 1599 619 1629 645
rect 1685 619 1715 645
rect 1771 619 1801 645
rect 1857 619 1887 645
rect 1943 619 1973 645
rect 83 303 113 367
rect 169 303 199 367
rect 255 303 285 367
rect 341 345 371 367
rect 335 315 371 345
rect 427 331 457 367
rect 517 331 547 367
rect 603 331 633 367
rect 775 331 805 367
rect 413 315 819 331
rect 335 303 365 315
rect 27 287 365 303
rect 27 253 43 287
rect 77 253 111 287
rect 145 253 179 287
rect 213 253 247 287
rect 281 253 315 287
rect 349 267 365 287
rect 413 281 429 315
rect 463 281 497 315
rect 531 281 565 315
rect 599 281 633 315
rect 667 281 701 315
rect 735 281 769 315
rect 803 281 819 315
rect 349 253 368 267
rect 413 265 819 281
rect 27 237 368 253
rect 80 215 110 237
rect 166 215 196 237
rect 252 215 282 237
rect 338 215 368 237
rect 531 233 561 265
rect 617 233 647 265
rect 703 233 733 265
rect 789 233 819 265
rect 861 321 891 367
rect 947 321 977 367
rect 1033 321 1063 367
rect 1151 321 1181 367
rect 1237 321 1267 367
rect 1323 321 1353 367
rect 1409 321 1439 367
rect 1599 321 1629 367
rect 1685 321 1715 367
rect 1771 321 1801 367
rect 1857 321 1887 367
rect 1943 321 1973 367
rect 861 305 1195 321
rect 861 271 941 305
rect 975 271 1009 305
rect 1043 271 1077 305
rect 1111 271 1145 305
rect 1179 271 1195 305
rect 861 255 1195 271
rect 1237 305 1643 321
rect 1237 271 1253 305
rect 1287 271 1321 305
rect 1355 271 1389 305
rect 1423 271 1457 305
rect 1491 271 1525 305
rect 1559 271 1593 305
rect 1627 271 1643 305
rect 1237 255 1643 271
rect 1685 305 2091 321
rect 1685 271 1701 305
rect 1735 271 1769 305
rect 1803 271 1837 305
rect 1871 271 1905 305
rect 1939 271 1973 305
rect 2007 271 2041 305
rect 2075 271 2091 305
rect 1685 255 2091 271
rect 891 233 921 255
rect 977 233 1007 255
rect 1063 233 1093 255
rect 1149 233 1179 255
rect 1344 233 1374 255
rect 1430 233 1460 255
rect 1516 233 1546 255
rect 1602 233 1632 255
rect 1688 233 1718 255
rect 1774 233 1804 255
rect 1860 233 1890 255
rect 1946 233 1976 255
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 531 39 561 65
rect 617 39 647 65
rect 703 39 733 65
rect 789 39 819 65
rect 891 39 921 65
rect 977 39 1007 65
rect 1063 39 1093 65
rect 1149 39 1179 65
rect 1344 39 1374 65
rect 1430 39 1460 65
rect 1516 39 1546 65
rect 1602 39 1632 65
rect 1688 39 1718 65
rect 1774 39 1804 65
rect 1860 39 1890 65
rect 1946 39 1976 65
<< polycont >>
rect 43 253 77 287
rect 111 253 145 287
rect 179 253 213 287
rect 247 253 281 287
rect 315 253 349 287
rect 429 281 463 315
rect 497 281 531 315
rect 565 281 599 315
rect 633 281 667 315
rect 701 281 735 315
rect 769 281 803 315
rect 941 271 975 305
rect 1009 271 1043 305
rect 1077 271 1111 305
rect 1145 271 1179 305
rect 1253 271 1287 305
rect 1321 271 1355 305
rect 1389 271 1423 305
rect 1457 271 1491 305
rect 1525 271 1559 305
rect 1593 271 1627 305
rect 1701 271 1735 305
rect 1769 271 1803 305
rect 1837 271 1871 305
rect 1905 271 1939 305
rect 1973 271 2007 305
rect 2041 271 2075 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 22 599 422 615
rect 22 565 38 599
rect 72 581 210 599
rect 72 565 74 581
rect 22 509 74 565
rect 208 565 210 581
rect 244 581 382 599
rect 244 565 246 581
rect 22 475 38 509
rect 72 475 74 509
rect 22 415 74 475
rect 22 381 38 415
rect 72 381 74 415
rect 22 365 74 381
rect 108 513 124 547
rect 158 513 174 547
rect 108 479 174 513
rect 108 445 124 479
rect 158 445 174 479
rect 108 411 174 445
rect 108 377 124 411
rect 158 377 174 411
rect 208 517 246 565
rect 380 565 382 581
rect 416 565 422 599
rect 208 483 210 517
rect 244 483 246 517
rect 208 442 246 483
rect 208 408 210 442
rect 244 408 246 442
rect 208 392 246 408
rect 280 513 296 547
rect 330 513 346 547
rect 280 479 346 513
rect 280 445 296 479
rect 330 445 346 479
rect 280 411 346 445
rect 380 471 422 565
rect 456 611 522 649
rect 456 577 472 611
rect 506 577 522 611
rect 456 541 522 577
rect 456 507 472 541
rect 506 507 522 541
rect 456 491 522 507
rect 556 599 598 615
rect 556 565 558 599
rect 592 565 598 599
rect 380 437 382 471
rect 416 457 422 471
rect 556 471 598 565
rect 632 611 766 649
rect 632 577 648 611
rect 682 577 716 611
rect 750 577 766 611
rect 632 530 766 577
rect 632 496 648 530
rect 682 496 716 530
rect 750 496 766 530
rect 632 493 766 496
rect 800 611 866 615
rect 800 577 816 611
rect 850 577 866 611
rect 800 538 866 577
rect 800 504 816 538
rect 850 504 866 538
rect 556 457 558 471
rect 416 437 558 457
rect 592 457 598 471
rect 800 461 866 504
rect 900 611 944 649
rect 900 577 902 611
rect 936 577 944 611
rect 900 541 944 577
rect 900 507 902 541
rect 936 507 944 541
rect 900 491 944 507
rect 978 599 1026 615
rect 978 565 988 599
rect 1022 565 1026 599
rect 978 503 1026 565
rect 800 457 816 461
rect 592 437 816 457
rect 380 427 816 437
rect 850 457 866 461
rect 978 469 988 503
rect 1022 469 1026 503
rect 978 457 1026 469
rect 850 427 1026 457
rect 380 421 1026 427
rect 1074 607 1140 649
rect 1074 573 1090 607
rect 1124 573 1140 607
rect 1074 529 1140 573
rect 1074 495 1090 529
rect 1124 495 1140 529
rect 1074 455 1140 495
rect 1074 421 1090 455
rect 1124 421 1140 455
rect 1176 599 1228 615
rect 1176 565 1192 599
rect 1226 565 1228 599
rect 1176 509 1228 565
rect 1176 475 1192 509
rect 1226 475 1228 509
rect 108 358 174 377
rect 280 377 296 411
rect 330 387 346 411
rect 972 413 1026 421
rect 330 377 891 387
rect 280 358 891 377
rect 108 349 891 358
rect 972 379 988 413
rect 1022 385 1026 413
rect 1176 413 1228 475
rect 1262 607 1328 649
rect 1262 573 1278 607
rect 1312 573 1328 607
rect 1262 529 1328 573
rect 1262 495 1278 529
rect 1312 495 1328 529
rect 1262 455 1328 495
rect 1262 421 1278 455
rect 1312 421 1328 455
rect 1362 599 1400 615
rect 1362 565 1364 599
rect 1398 565 1400 599
rect 1362 509 1400 565
rect 1362 475 1364 509
rect 1398 475 1400 509
rect 1176 385 1192 413
rect 1022 379 1192 385
rect 1226 385 1228 413
rect 1362 413 1400 475
rect 1434 607 1604 649
rect 1434 573 1450 607
rect 1484 573 1554 607
rect 1588 573 1604 607
rect 1434 529 1604 573
rect 1434 495 1450 529
rect 1484 495 1554 529
rect 1588 495 1604 529
rect 1434 455 1604 495
rect 1434 421 1450 455
rect 1484 421 1554 455
rect 1588 421 1604 455
rect 1638 599 1676 615
rect 1638 565 1640 599
rect 1674 565 1676 599
rect 1638 509 1676 565
rect 1638 475 1640 509
rect 1674 475 1676 509
rect 1362 385 1364 413
rect 1226 379 1364 385
rect 1398 385 1400 413
rect 1638 413 1676 475
rect 1710 607 1776 649
rect 1710 573 1726 607
rect 1760 573 1776 607
rect 1710 529 1776 573
rect 1710 495 1726 529
rect 1760 495 1776 529
rect 1710 455 1776 495
rect 1710 421 1726 455
rect 1760 421 1776 455
rect 1810 599 1848 615
rect 1810 565 1812 599
rect 1846 565 1848 599
rect 1810 509 1848 565
rect 1810 475 1812 509
rect 1846 475 1848 509
rect 1638 385 1640 413
rect 1398 379 1640 385
rect 1674 385 1676 413
rect 1810 413 1848 475
rect 1882 607 1948 649
rect 1882 573 1898 607
rect 1932 573 1948 607
rect 1882 529 1948 573
rect 1882 495 1898 529
rect 1932 495 1948 529
rect 1882 455 1948 495
rect 1882 421 1898 455
rect 1932 421 1948 455
rect 1982 599 2034 615
rect 1982 565 1984 599
rect 2018 565 2034 599
rect 1982 509 2034 565
rect 1982 475 1984 509
rect 2018 475 2034 509
rect 1810 385 1812 413
rect 1674 379 1812 385
rect 1846 385 1848 413
rect 1982 413 2034 475
rect 1982 385 1984 413
rect 1846 379 1984 385
rect 2018 379 2034 413
rect 972 351 2034 379
rect 108 321 363 349
rect 20 253 43 287
rect 77 253 111 287
rect 145 253 179 287
rect 213 253 247 287
rect 281 253 315 287
rect 349 253 365 287
rect 413 281 429 315
rect 463 281 497 315
rect 531 281 565 315
rect 599 281 633 315
rect 667 281 701 315
rect 735 281 769 315
rect 803 281 819 315
rect 20 242 365 253
rect 511 242 641 281
rect 853 247 891 349
rect 728 225 891 247
rect 925 305 1195 317
rect 925 271 941 305
rect 975 271 1009 305
rect 1043 271 1077 305
rect 1111 271 1145 305
rect 1179 271 1195 305
rect 925 239 1195 271
rect 1237 305 1643 317
rect 1237 271 1253 305
rect 1287 271 1321 305
rect 1355 271 1389 305
rect 1423 271 1457 305
rect 1491 271 1525 305
rect 1559 271 1593 305
rect 1627 271 1643 305
rect 1685 305 2091 317
rect 1685 271 1701 305
rect 1735 271 1769 305
rect 1803 271 1837 305
rect 1871 271 1905 305
rect 1939 271 1973 305
rect 2007 271 2041 305
rect 2075 271 2091 305
rect 1237 263 1507 271
rect 1469 231 1507 263
rect 1685 240 2091 271
rect 728 208 744 225
rect 19 203 85 208
rect 19 169 35 203
rect 69 169 85 203
rect 19 93 85 169
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 119 201 744 208
rect 119 192 572 201
rect 119 158 121 192
rect 155 171 293 192
rect 155 158 157 171
rect 119 101 157 158
rect 291 158 293 171
rect 327 167 572 192
rect 606 191 744 201
rect 778 213 891 225
rect 1369 225 1435 229
rect 778 191 794 213
rect 1369 205 1385 225
rect 606 167 794 191
rect 930 201 1385 205
rect 327 163 794 167
rect 327 158 329 163
rect 119 67 121 101
rect 155 67 157 101
rect 119 51 157 67
rect 191 126 257 137
rect 191 92 207 126
rect 241 92 257 126
rect 191 17 257 92
rect 291 101 329 158
rect 728 153 794 163
rect 291 67 293 101
rect 327 67 329 101
rect 291 51 329 67
rect 363 118 429 129
rect 363 84 379 118
rect 413 84 429 118
rect 363 17 429 84
rect 470 111 694 129
rect 728 119 744 153
rect 778 119 794 153
rect 830 145 846 179
rect 880 145 896 179
rect 470 77 486 111
rect 520 77 658 111
rect 692 85 694 111
rect 830 107 896 145
rect 930 169 1104 201
rect 930 135 932 169
rect 966 167 1104 169
rect 1138 191 1385 201
rect 1419 197 1435 225
rect 1541 225 1607 229
rect 1541 197 1557 225
rect 1419 191 1557 197
rect 1591 191 1607 225
rect 1138 167 1607 191
rect 966 163 1607 167
rect 966 135 980 163
rect 930 119 980 135
rect 1369 157 1435 163
rect 830 85 846 107
rect 692 77 846 85
rect 470 73 846 77
rect 880 85 896 107
rect 1014 111 1228 129
rect 1014 85 1018 111
rect 880 77 1018 85
rect 1052 77 1190 111
rect 1224 77 1228 111
rect 880 73 1228 77
rect 470 51 1228 73
rect 1295 113 1335 129
rect 1369 123 1385 157
rect 1419 123 1435 157
rect 1541 157 1607 163
rect 1295 79 1299 113
rect 1333 85 1335 113
rect 1469 113 1507 129
rect 1541 123 1557 157
rect 1591 123 1607 157
rect 1643 192 2037 206
rect 1643 190 1815 192
rect 1677 172 1815 190
rect 1677 156 1679 172
rect 1469 85 1471 113
rect 1333 79 1471 85
rect 1505 85 1507 113
rect 1643 111 1679 156
rect 1813 158 1815 172
rect 1849 172 1987 192
rect 1849 158 1851 172
rect 1505 79 1643 85
rect 1295 77 1643 79
rect 1677 77 1679 111
rect 1295 51 1679 77
rect 1713 130 1779 138
rect 1713 96 1729 130
rect 1763 96 1779 130
rect 1713 17 1779 96
rect 1813 113 1851 158
rect 1985 158 1987 172
rect 2021 158 2037 192
rect 1813 79 1815 113
rect 1849 79 1851 113
rect 1813 63 1851 79
rect 1885 130 1951 138
rect 1885 96 1901 130
rect 1935 96 1951 130
rect 1885 17 1951 96
rect 1985 113 2037 158
rect 1985 79 1987 113
rect 2021 79 2037 113
rect 1985 63 2037 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a41oi_4
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1373272
string GDS_START 1355166
<< end >>
