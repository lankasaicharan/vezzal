magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 1 49 627 241
rect 0 0 672 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 252 47 282 215
rect 338 47 368 215
rect 432 47 462 215
rect 518 47 548 215
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 252 367 282 619
rect 346 367 376 619
rect 432 367 462 619
rect 518 367 548 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 93 80 169
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 203 166 215
rect 110 169 121 203
rect 155 169 166 203
rect 110 103 166 169
rect 110 69 121 103
rect 155 69 166 103
rect 110 47 166 69
rect 196 169 252 215
rect 196 135 207 169
rect 241 135 252 169
rect 196 47 252 135
rect 282 123 338 215
rect 282 89 293 123
rect 327 89 338 123
rect 282 47 338 89
rect 368 127 432 215
rect 368 93 383 127
rect 417 93 432 127
rect 368 47 432 93
rect 462 203 518 215
rect 462 169 473 203
rect 507 169 518 203
rect 462 101 518 169
rect 462 67 473 101
rect 507 67 518 101
rect 462 47 518 67
rect 548 167 601 215
rect 548 133 559 167
rect 593 133 601 167
rect 548 93 601 133
rect 548 59 559 93
rect 593 59 601 93
rect 548 47 601 59
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 516 80 565
rect 27 482 35 516
rect 69 482 80 516
rect 27 425 80 482
rect 27 391 35 425
rect 69 391 80 425
rect 27 367 80 391
rect 110 607 166 619
rect 110 573 121 607
rect 155 573 166 607
rect 110 501 166 573
rect 110 467 121 501
rect 155 467 166 501
rect 110 367 166 467
rect 196 599 252 619
rect 196 565 207 599
rect 241 565 252 599
rect 196 516 252 565
rect 196 482 207 516
rect 241 482 252 516
rect 196 425 252 482
rect 196 391 207 425
rect 241 391 252 425
rect 196 367 252 391
rect 282 607 346 619
rect 282 573 297 607
rect 331 573 346 607
rect 282 501 346 573
rect 282 467 297 501
rect 331 467 346 501
rect 282 367 346 467
rect 376 599 432 619
rect 376 565 387 599
rect 421 565 432 599
rect 376 516 432 565
rect 376 482 387 516
rect 421 482 432 516
rect 376 441 432 482
rect 376 407 387 441
rect 421 407 432 441
rect 376 367 432 407
rect 462 541 518 619
rect 462 507 473 541
rect 507 507 518 541
rect 462 420 518 507
rect 462 386 473 420
rect 507 386 518 420
rect 462 367 518 386
rect 548 599 601 619
rect 548 565 559 599
rect 593 565 601 599
rect 548 504 601 565
rect 548 470 559 504
rect 593 470 601 504
rect 548 367 601 470
<< ndiffc >>
rect 35 169 69 203
rect 35 59 69 93
rect 121 169 155 203
rect 121 69 155 103
rect 207 135 241 169
rect 293 89 327 123
rect 383 93 417 127
rect 473 169 507 203
rect 473 67 507 101
rect 559 133 593 167
rect 559 59 593 93
<< pdiffc >>
rect 35 565 69 599
rect 35 482 69 516
rect 35 391 69 425
rect 121 573 155 607
rect 121 467 155 501
rect 207 565 241 599
rect 207 482 241 516
rect 207 391 241 425
rect 297 573 331 607
rect 297 467 331 501
rect 387 565 421 599
rect 387 482 421 516
rect 387 407 421 441
rect 473 507 507 541
rect 473 386 507 420
rect 559 565 593 599
rect 559 470 593 504
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 252 619 282 645
rect 346 619 376 645
rect 432 619 462 645
rect 518 619 548 645
rect 80 325 110 367
rect 25 309 110 325
rect 25 275 41 309
rect 75 275 110 309
rect 25 259 110 275
rect 80 215 110 259
rect 166 303 196 367
rect 252 303 282 367
rect 346 335 376 367
rect 432 335 462 367
rect 518 335 548 367
rect 166 287 282 303
rect 166 253 182 287
rect 216 253 282 287
rect 324 319 390 335
rect 324 285 340 319
rect 374 285 390 319
rect 324 269 390 285
rect 432 319 548 335
rect 432 285 448 319
rect 482 285 548 319
rect 432 269 548 285
rect 166 237 282 253
rect 166 215 196 237
rect 252 215 282 237
rect 338 215 368 269
rect 432 215 462 269
rect 518 215 548 269
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 432 21 462 47
rect 518 21 548 47
<< polycont >>
rect 41 275 75 309
rect 182 253 216 287
rect 340 285 374 319
rect 448 285 482 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 19 599 71 615
rect 19 565 35 599
rect 69 565 71 599
rect 19 516 71 565
rect 19 482 35 516
rect 69 482 71 516
rect 19 425 71 482
rect 105 607 171 649
rect 105 573 121 607
rect 155 573 171 607
rect 105 501 171 573
rect 105 467 121 501
rect 155 467 171 501
rect 105 459 171 467
rect 205 599 247 615
rect 205 565 207 599
rect 241 565 247 599
rect 205 516 247 565
rect 205 482 207 516
rect 241 482 247 516
rect 205 425 247 482
rect 281 607 347 649
rect 281 573 297 607
rect 331 573 347 607
rect 281 501 347 573
rect 281 467 297 501
rect 331 467 347 501
rect 281 459 347 467
rect 381 599 609 615
rect 381 565 387 599
rect 421 581 559 599
rect 421 565 423 581
rect 381 516 423 565
rect 557 565 559 581
rect 593 565 609 599
rect 381 482 387 516
rect 421 482 423 516
rect 381 441 423 482
rect 381 425 387 441
rect 19 391 35 425
rect 69 391 207 425
rect 241 407 387 425
rect 421 407 423 441
rect 241 391 423 407
rect 457 541 523 547
rect 457 507 473 541
rect 507 507 523 541
rect 457 420 523 507
rect 557 504 609 565
rect 557 470 559 504
rect 593 470 609 504
rect 557 454 609 470
rect 457 386 473 420
rect 507 386 655 420
rect 25 335 353 357
rect 25 321 374 335
rect 25 309 91 321
rect 25 275 41 309
rect 75 275 91 309
rect 305 319 374 321
rect 25 259 91 275
rect 125 253 182 287
rect 216 253 271 287
rect 305 285 340 319
rect 408 319 560 352
rect 408 285 448 319
rect 482 285 560 319
rect 305 269 374 285
rect 125 241 271 253
rect 594 235 655 386
rect 19 203 71 219
rect 469 207 655 235
rect 19 169 35 203
rect 69 169 71 203
rect 19 93 71 169
rect 19 59 35 93
rect 69 59 71 93
rect 19 17 71 59
rect 105 203 171 207
rect 105 169 121 203
rect 155 169 171 203
rect 105 103 171 169
rect 205 203 655 207
rect 205 173 473 203
rect 205 169 252 173
rect 205 135 207 169
rect 241 135 252 169
rect 467 169 473 173
rect 507 201 655 203
rect 507 169 509 201
rect 205 119 252 135
rect 286 123 333 139
rect 105 69 121 103
rect 155 85 171 103
rect 286 89 293 123
rect 327 89 333 123
rect 286 85 333 89
rect 155 69 333 85
rect 105 51 333 69
rect 367 127 433 139
rect 367 93 383 127
rect 417 93 433 127
rect 367 17 433 93
rect 467 101 509 169
rect 467 67 473 101
rect 507 67 509 101
rect 467 51 509 67
rect 543 133 559 167
rect 593 133 609 167
rect 543 93 609 133
rect 543 59 559 93
rect 593 59 609 93
rect 543 17 609 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21oi_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3596356
string GDS_START 3589732
<< end >>
