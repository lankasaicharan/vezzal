magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2586 1852
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 108 157 1030 203
rect 1 21 1287 157
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 131
rect 184 47 214 177
rect 278 47 308 177
rect 372 47 402 177
rect 466 47 496 177
rect 576 47 606 177
rect 689 47 719 177
rect 806 47 836 177
rect 912 47 942 177
rect 1169 47 1199 131
<< scpmoshvt >>
rect 81 413 117 497
rect 186 297 222 497
rect 280 297 316 497
rect 374 297 410 497
rect 468 297 504 497
rect 578 297 614 497
rect 691 297 727 497
rect 808 297 844 497
rect 914 297 950 497
rect 1171 413 1207 497
<< ndiff >>
rect 134 131 184 177
rect 27 101 89 131
rect 27 67 35 101
rect 69 67 89 101
rect 27 47 89 67
rect 119 93 184 131
rect 119 59 140 93
rect 174 59 184 93
rect 119 47 184 59
rect 214 101 278 177
rect 214 67 234 101
rect 268 67 278 101
rect 214 47 278 67
rect 308 94 372 177
rect 308 60 328 94
rect 362 60 372 94
rect 308 47 372 60
rect 402 101 466 177
rect 402 67 422 101
rect 456 67 466 101
rect 402 47 466 67
rect 496 89 576 177
rect 496 55 510 89
rect 544 55 576 89
rect 496 47 576 55
rect 606 47 689 177
rect 719 47 806 177
rect 836 47 912 177
rect 942 162 1004 177
rect 942 128 962 162
rect 996 128 1004 162
rect 942 94 1004 128
rect 942 60 962 94
rect 996 60 1004 94
rect 942 47 1004 60
rect 1077 93 1169 131
rect 1077 59 1093 93
rect 1127 59 1169 93
rect 1077 47 1169 59
rect 1199 101 1261 131
rect 1199 67 1219 101
rect 1253 67 1261 101
rect 1199 47 1261 67
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 413 81 443
rect 117 485 186 497
rect 117 451 129 485
rect 163 451 186 485
rect 117 413 186 451
rect 134 297 186 413
rect 222 343 280 497
rect 222 309 234 343
rect 268 309 280 343
rect 222 297 280 309
rect 316 485 374 497
rect 316 451 328 485
rect 362 451 374 485
rect 316 297 374 451
rect 410 343 468 497
rect 410 309 422 343
rect 456 309 468 343
rect 410 297 468 309
rect 504 485 578 497
rect 504 451 516 485
rect 550 451 578 485
rect 504 297 578 451
rect 614 343 691 497
rect 614 309 638 343
rect 672 309 691 343
rect 614 297 691 309
rect 727 485 808 497
rect 727 451 752 485
rect 786 451 808 485
rect 727 297 808 451
rect 844 343 914 497
rect 844 309 860 343
rect 894 309 914 343
rect 844 297 914 309
rect 950 485 1171 497
rect 950 451 978 485
rect 1012 451 1046 485
rect 1080 451 1114 485
rect 1148 451 1171 485
rect 950 413 1171 451
rect 1207 477 1261 497
rect 1207 443 1219 477
rect 1253 443 1261 477
rect 1207 413 1261 443
rect 950 297 1004 413
<< ndiffc >>
rect 35 67 69 101
rect 140 59 174 93
rect 234 67 268 101
rect 328 60 362 94
rect 422 67 456 101
rect 510 55 544 89
rect 962 128 996 162
rect 962 60 996 94
rect 1093 59 1127 93
rect 1219 67 1253 101
<< pdiffc >>
rect 35 443 69 477
rect 129 451 163 485
rect 234 309 268 343
rect 328 451 362 485
rect 422 309 456 343
rect 516 451 550 485
rect 638 309 672 343
rect 752 451 786 485
rect 860 309 894 343
rect 978 451 1012 485
rect 1046 451 1080 485
rect 1114 451 1148 485
rect 1219 443 1253 477
<< poly >>
rect 81 497 117 523
rect 186 497 222 523
rect 280 497 316 523
rect 374 497 410 523
rect 468 497 504 523
rect 578 497 614 523
rect 691 497 727 523
rect 808 497 844 523
rect 914 497 950 523
rect 1171 497 1207 523
rect 81 398 117 413
rect 79 265 119 398
rect 1171 398 1207 413
rect 186 282 222 297
rect 280 282 316 297
rect 374 282 410 297
rect 468 282 504 297
rect 578 282 614 297
rect 691 282 727 297
rect 808 282 844 297
rect 914 282 950 297
rect 184 275 224 282
rect 278 275 318 282
rect 372 275 412 282
rect 466 275 504 282
rect 76 249 140 265
rect 76 215 86 249
rect 120 215 140 249
rect 76 199 140 215
rect 184 259 504 275
rect 576 265 616 282
rect 689 265 729 282
rect 806 265 846 282
rect 912 275 952 282
rect 184 249 496 259
rect 184 215 328 249
rect 362 215 396 249
rect 430 215 496 249
rect 184 205 496 215
rect 89 131 119 199
rect 184 177 214 205
rect 278 177 308 205
rect 372 177 402 205
rect 466 177 496 205
rect 576 249 647 265
rect 576 215 586 249
rect 620 215 647 249
rect 576 199 647 215
rect 689 249 764 265
rect 689 215 710 249
rect 744 215 764 249
rect 689 199 764 215
rect 806 249 870 265
rect 806 215 816 249
rect 850 215 870 249
rect 806 199 870 215
rect 912 249 1126 275
rect 912 215 1072 249
rect 1106 215 1126 249
rect 912 205 1126 215
rect 1169 265 1209 398
rect 1169 249 1241 265
rect 1169 215 1187 249
rect 1221 215 1241 249
rect 576 177 606 199
rect 689 177 719 199
rect 806 177 836 199
rect 912 177 942 205
rect 1169 199 1241 215
rect 1169 131 1199 199
rect 89 21 119 47
rect 184 21 214 47
rect 278 21 308 47
rect 372 21 402 47
rect 466 21 496 47
rect 576 21 606 47
rect 689 21 719 47
rect 806 21 836 47
rect 912 21 942 47
rect 1169 21 1199 47
<< polycont >>
rect 86 215 120 249
rect 328 215 362 249
rect 396 215 430 249
rect 586 215 620 249
rect 710 215 744 249
rect 816 215 850 249
rect 1072 215 1106 249
rect 1187 215 1221 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 477 69 493
rect 17 443 35 477
rect 103 485 179 527
rect 103 451 129 485
rect 163 451 179 485
rect 302 485 378 527
rect 302 451 328 485
rect 362 451 378 485
rect 490 485 566 527
rect 490 451 516 485
rect 550 451 566 485
rect 736 485 802 527
rect 736 451 752 485
rect 786 451 802 485
rect 962 485 1164 527
rect 962 451 978 485
rect 1012 451 1046 485
rect 1080 451 1114 485
rect 1148 451 1164 485
rect 1219 477 1253 493
rect 17 417 69 443
rect 1219 417 1253 443
rect 17 383 988 417
rect 17 117 52 383
rect 86 249 166 327
rect 120 215 166 249
rect 86 153 166 215
rect 202 309 234 343
rect 268 309 422 343
rect 456 309 472 343
rect 506 309 638 343
rect 672 309 860 343
rect 894 309 910 343
rect 202 164 268 309
rect 506 249 540 309
rect 954 275 988 383
rect 302 215 328 249
rect 362 215 396 249
rect 430 215 540 249
rect 202 130 456 164
rect 17 101 69 117
rect 17 67 35 101
rect 234 101 268 130
rect 17 51 69 67
rect 124 93 190 94
rect 124 59 140 93
rect 174 59 190 93
rect 124 17 190 59
rect 422 101 456 130
rect 506 157 540 215
rect 581 249 639 265
rect 581 215 586 249
rect 620 215 639 249
rect 581 199 639 215
rect 673 249 768 265
rect 673 215 710 249
rect 744 215 768 249
rect 506 123 639 157
rect 673 128 768 215
rect 816 249 988 275
rect 850 241 988 249
rect 1072 383 1253 417
rect 1072 249 1106 383
rect 850 215 860 241
rect 816 199 860 215
rect 1072 165 1106 215
rect 1187 249 1269 324
rect 1221 215 1269 249
rect 1187 199 1269 215
rect 942 128 962 162
rect 996 128 1012 162
rect 1072 131 1253 165
rect 234 51 268 67
rect 302 60 328 94
rect 362 60 378 94
rect 302 17 378 60
rect 595 94 639 123
rect 942 94 1012 128
rect 422 51 456 67
rect 494 55 510 89
rect 544 55 560 89
rect 595 60 962 94
rect 996 60 1012 94
rect 1219 101 1253 131
rect 494 17 560 55
rect 1077 59 1093 93
rect 1127 59 1143 93
rect 1077 17 1143 59
rect 1219 51 1253 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 673 141 707 175 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 1187 199 1269 324 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 1196 238 1196 238 0 FreeSans 200 0 0 0 A_N
port 1 nsew
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 214 289 248 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 132 153 166 187 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel locali s 132 289 166 323 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel locali s 217 153 251 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 132 221 166 255 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4bb_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1897630
string GDS_START 1888588
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
