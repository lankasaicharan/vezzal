magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 9 157 469 241
rect 9 49 863 157
rect 0 0 864 49
<< scnmos >>
rect 92 131 122 215
rect 164 131 194 215
rect 278 47 308 215
rect 356 47 386 215
rect 678 47 708 131
rect 750 47 780 131
<< scpmoshvt >>
rect 86 483 116 611
rect 164 483 194 611
rect 485 367 515 619
rect 563 367 593 619
rect 672 401 702 529
rect 750 401 780 529
<< ndiff >>
rect 35 188 92 215
rect 35 154 47 188
rect 81 154 92 188
rect 35 131 92 154
rect 122 131 164 215
rect 194 187 278 215
rect 194 153 229 187
rect 263 153 278 187
rect 194 131 278 153
rect 217 93 278 131
rect 217 59 229 93
rect 263 59 278 93
rect 217 47 278 59
rect 308 47 356 215
rect 386 186 443 215
rect 386 152 397 186
rect 431 152 443 186
rect 386 47 443 152
rect 621 105 678 131
rect 621 71 633 105
rect 667 71 678 105
rect 621 47 678 71
rect 708 47 750 131
rect 780 110 837 131
rect 780 76 791 110
rect 825 76 837 110
rect 780 47 837 76
<< pdiff >>
rect 29 599 86 611
rect 29 565 41 599
rect 75 565 86 599
rect 29 529 86 565
rect 29 495 41 529
rect 75 495 86 529
rect 29 483 86 495
rect 116 483 164 611
rect 194 599 331 611
rect 194 565 285 599
rect 319 565 331 599
rect 194 529 331 565
rect 194 495 285 529
rect 319 495 331 529
rect 194 483 331 495
rect 428 599 485 619
rect 428 565 440 599
rect 474 565 485 599
rect 428 527 485 565
rect 428 493 440 527
rect 474 493 485 527
rect 428 455 485 493
rect 428 421 440 455
rect 474 421 485 455
rect 428 367 485 421
rect 515 367 563 619
rect 593 607 650 619
rect 593 573 604 607
rect 638 573 650 607
rect 593 529 650 573
rect 593 510 672 529
rect 593 476 604 510
rect 638 476 672 510
rect 593 413 672 476
rect 593 379 604 413
rect 638 401 672 413
rect 702 401 750 529
rect 780 517 837 529
rect 780 483 791 517
rect 825 483 837 517
rect 780 447 837 483
rect 780 413 791 447
rect 825 413 837 447
rect 780 401 837 413
rect 638 379 650 401
rect 593 367 650 379
<< ndiffc >>
rect 47 154 81 188
rect 229 153 263 187
rect 229 59 263 93
rect 397 152 431 186
rect 633 71 667 105
rect 791 76 825 110
<< pdiffc >>
rect 41 565 75 599
rect 41 495 75 529
rect 285 565 319 599
rect 285 495 319 529
rect 440 565 474 599
rect 440 493 474 527
rect 440 421 474 455
rect 604 573 638 607
rect 604 476 638 510
rect 604 379 638 413
rect 791 483 825 517
rect 791 413 825 447
<< poly >>
rect 86 611 116 637
rect 164 611 194 637
rect 485 619 515 645
rect 563 619 593 645
rect 86 383 116 483
rect 164 383 194 483
rect 86 367 194 383
rect 672 529 702 555
rect 750 529 780 555
rect 86 333 114 367
rect 148 333 194 367
rect 485 335 515 367
rect 86 299 194 333
rect 356 319 515 335
rect 86 265 114 299
rect 148 265 194 299
rect 86 249 194 265
rect 92 215 122 249
rect 164 215 194 249
rect 242 287 308 303
rect 242 253 258 287
rect 292 253 308 287
rect 242 237 308 253
rect 278 215 308 237
rect 356 285 397 319
rect 431 305 515 319
rect 431 285 447 305
rect 356 269 447 285
rect 356 215 386 269
rect 563 265 593 367
rect 672 301 702 401
rect 750 379 780 401
rect 750 349 832 379
rect 672 285 754 301
rect 672 265 704 285
rect 563 251 704 265
rect 738 265 754 285
rect 802 265 832 349
rect 738 251 832 265
rect 563 235 832 251
rect 92 105 122 131
rect 164 105 194 131
rect 678 131 708 235
rect 750 131 780 235
rect 278 21 308 47
rect 356 21 386 47
rect 678 21 708 47
rect 750 21 780 47
<< polycont >>
rect 114 333 148 367
rect 114 265 148 299
rect 258 253 292 287
rect 397 285 431 319
rect 704 251 738 285
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 25 599 91 615
rect 25 565 41 599
rect 75 565 91 599
rect 25 529 91 565
rect 25 495 41 529
rect 75 513 91 529
rect 269 599 335 649
rect 269 565 285 599
rect 319 565 335 599
rect 269 529 335 565
rect 75 495 235 513
rect 25 479 235 495
rect 269 495 285 529
rect 319 495 335 529
rect 269 479 335 495
rect 424 599 490 615
rect 424 565 440 599
rect 474 578 490 599
rect 588 607 654 649
rect 474 565 551 578
rect 424 527 551 565
rect 424 493 440 527
rect 474 493 551 527
rect 25 215 59 479
rect 98 367 167 430
rect 98 333 114 367
rect 148 333 167 367
rect 201 371 235 479
rect 424 455 551 493
rect 424 421 440 455
rect 474 421 551 455
rect 424 405 551 421
rect 201 337 447 371
rect 98 299 167 333
rect 381 319 447 337
rect 98 265 114 299
rect 148 265 167 299
rect 98 249 167 265
rect 242 287 347 303
rect 242 253 258 287
rect 292 253 347 287
rect 381 285 397 319
rect 431 285 447 319
rect 381 269 447 285
rect 242 237 347 253
rect 25 188 97 215
rect 25 154 47 188
rect 81 154 97 188
rect 25 127 97 154
rect 213 187 279 203
rect 213 153 229 187
rect 263 153 279 187
rect 213 93 279 153
rect 213 59 229 93
rect 263 59 279 93
rect 213 17 279 59
rect 313 85 347 237
rect 481 235 551 405
rect 588 573 604 607
rect 638 573 654 607
rect 588 510 654 573
rect 588 476 604 510
rect 638 476 654 510
rect 588 413 654 476
rect 588 379 604 413
rect 638 379 654 413
rect 775 517 841 533
rect 775 483 791 517
rect 825 483 841 517
rect 775 447 841 483
rect 775 413 791 447
rect 825 413 841 447
rect 775 397 841 413
rect 588 363 654 379
rect 688 285 754 356
rect 688 251 704 285
rect 738 251 754 285
rect 688 235 754 251
rect 381 201 515 235
rect 807 201 841 397
rect 381 186 481 201
rect 381 152 397 186
rect 431 152 481 186
rect 381 119 481 152
rect 549 167 841 201
rect 549 85 583 167
rect 313 51 583 85
rect 617 105 683 133
rect 617 71 633 105
rect 667 71 683 105
rect 617 17 683 71
rect 775 110 841 167
rect 775 76 791 110
rect 825 76 841 110
rect 775 51 841 76
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ebufn_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3345586
string GDS_START 3338706
<< end >>
