magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2678 1852
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 1 21 1359 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 267 47 297 177
rect 371 47 401 177
rect 465 47 495 177
rect 561 47 591 177
rect 667 47 697 177
rect 761 47 791 177
rect 969 47 999 177
rect 1063 47 1093 177
rect 1157 47 1187 177
rect 1251 47 1281 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 563 297 599 497
rect 669 297 705 497
rect 763 297 799 497
rect 961 297 997 497
rect 1055 297 1091 497
rect 1149 297 1185 497
rect 1243 297 1279 497
<< ndiff >>
rect 27 165 89 177
rect 27 131 35 165
rect 69 131 89 165
rect 27 97 89 131
rect 27 63 35 97
rect 69 63 89 97
rect 27 47 89 63
rect 119 47 183 177
rect 213 47 267 177
rect 297 113 371 177
rect 297 79 317 113
rect 351 79 371 113
rect 297 47 371 79
rect 401 47 465 177
rect 495 47 561 177
rect 591 90 667 177
rect 591 56 619 90
rect 653 56 667 90
rect 591 47 667 56
rect 697 161 761 177
rect 697 127 717 161
rect 751 127 761 161
rect 697 93 761 127
rect 697 59 717 93
rect 751 59 761 93
rect 697 47 761 59
rect 791 97 969 177
rect 791 63 827 97
rect 861 63 899 97
rect 933 63 969 97
rect 791 47 969 63
rect 999 165 1063 177
rect 999 131 1009 165
rect 1043 131 1063 165
rect 999 47 1063 131
rect 1093 97 1157 177
rect 1093 63 1103 97
rect 1137 63 1157 97
rect 1093 47 1157 63
rect 1187 165 1251 177
rect 1187 131 1197 165
rect 1231 131 1251 165
rect 1187 47 1251 131
rect 1281 97 1333 177
rect 1281 63 1291 97
rect 1325 63 1333 97
rect 1281 47 1333 63
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 407 81 443
rect 27 373 35 407
rect 69 373 81 407
rect 27 297 81 373
rect 117 459 175 497
rect 117 425 129 459
rect 163 425 175 459
rect 117 297 175 425
rect 211 477 269 497
rect 211 443 223 477
rect 257 443 269 477
rect 211 407 269 443
rect 211 373 223 407
rect 257 373 269 407
rect 211 297 269 373
rect 305 459 363 497
rect 305 425 317 459
rect 351 425 363 459
rect 305 297 363 425
rect 399 477 457 497
rect 399 443 411 477
rect 445 443 457 477
rect 399 407 457 443
rect 399 373 411 407
rect 445 373 457 407
rect 399 297 457 373
rect 493 459 563 497
rect 493 425 505 459
rect 539 425 563 459
rect 493 297 563 425
rect 599 477 669 497
rect 599 443 623 477
rect 657 443 669 477
rect 599 407 669 443
rect 599 373 623 407
rect 657 373 669 407
rect 599 297 669 373
rect 705 423 763 497
rect 705 389 717 423
rect 751 389 763 423
rect 705 343 763 389
rect 705 309 717 343
rect 751 309 763 343
rect 705 297 763 309
rect 799 477 853 497
rect 799 443 811 477
rect 845 443 853 477
rect 799 409 853 443
rect 799 375 811 409
rect 845 375 853 409
rect 799 297 853 375
rect 907 459 961 497
rect 907 425 915 459
rect 949 425 961 459
rect 907 297 961 425
rect 997 477 1055 497
rect 997 443 1009 477
rect 1043 443 1055 477
rect 997 407 1055 443
rect 997 373 1009 407
rect 1043 373 1055 407
rect 997 297 1055 373
rect 1091 459 1149 497
rect 1091 425 1103 459
rect 1137 425 1149 459
rect 1091 297 1149 425
rect 1185 477 1243 497
rect 1185 443 1197 477
rect 1231 443 1243 477
rect 1185 407 1243 443
rect 1185 373 1197 407
rect 1231 373 1243 407
rect 1185 297 1243 373
rect 1279 459 1333 497
rect 1279 425 1291 459
rect 1325 425 1333 459
rect 1279 297 1333 425
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 317 79 351 113
rect 619 56 653 90
rect 717 127 751 161
rect 717 59 751 93
rect 827 63 861 97
rect 899 63 933 97
rect 1009 131 1043 165
rect 1103 63 1137 97
rect 1197 131 1231 165
rect 1291 63 1325 97
<< pdiffc >>
rect 35 443 69 477
rect 35 373 69 407
rect 129 425 163 459
rect 223 443 257 477
rect 223 373 257 407
rect 317 425 351 459
rect 411 443 445 477
rect 411 373 445 407
rect 505 425 539 459
rect 623 443 657 477
rect 623 373 657 407
rect 717 389 751 423
rect 717 309 751 343
rect 811 443 845 477
rect 811 375 845 409
rect 915 425 949 459
rect 1009 443 1043 477
rect 1009 373 1043 407
rect 1103 425 1137 459
rect 1197 443 1231 477
rect 1197 373 1231 407
rect 1291 425 1325 459
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 563 497 599 523
rect 669 497 705 523
rect 763 497 799 523
rect 961 497 997 523
rect 1055 497 1091 523
rect 1149 497 1185 523
rect 1243 497 1279 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 563 282 599 297
rect 669 282 705 297
rect 763 282 799 297
rect 961 282 997 297
rect 1055 282 1091 297
rect 1149 282 1185 297
rect 1243 282 1279 297
rect 79 265 119 282
rect 173 265 213 282
rect 45 249 119 265
rect 45 215 55 249
rect 89 215 119 249
rect 45 199 119 215
rect 161 249 225 265
rect 161 215 171 249
rect 205 215 225 249
rect 161 199 225 215
rect 267 259 307 282
rect 361 259 401 282
rect 455 265 495 282
rect 561 265 601 282
rect 667 265 707 282
rect 761 265 801 282
rect 959 265 999 282
rect 1053 265 1093 282
rect 1147 265 1187 282
rect 1241 265 1281 282
rect 267 249 401 259
rect 267 215 316 249
rect 350 215 401 249
rect 267 205 401 215
rect 89 177 119 199
rect 183 177 213 199
rect 267 177 297 205
rect 371 177 401 205
rect 443 249 507 265
rect 443 215 453 249
rect 487 215 507 249
rect 443 199 507 215
rect 561 249 625 265
rect 561 215 571 249
rect 605 215 625 249
rect 561 199 625 215
rect 667 259 801 265
rect 667 249 861 259
rect 667 215 811 249
rect 845 215 861 249
rect 667 205 861 215
rect 951 249 1281 265
rect 951 215 961 249
rect 995 215 1039 249
rect 1073 215 1117 249
rect 1151 215 1195 249
rect 1229 215 1281 249
rect 667 199 791 205
rect 951 199 1281 215
rect 465 177 495 199
rect 561 177 591 199
rect 667 177 697 199
rect 761 177 791 199
rect 969 177 999 199
rect 1063 177 1093 199
rect 1157 177 1187 199
rect 1251 177 1281 199
rect 89 21 119 47
rect 183 21 213 47
rect 267 21 297 47
rect 371 21 401 47
rect 465 21 495 47
rect 561 21 591 47
rect 667 21 697 47
rect 761 21 791 47
rect 969 21 999 47
rect 1063 21 1093 47
rect 1157 21 1187 47
rect 1251 21 1281 47
<< polycont >>
rect 55 215 89 249
rect 171 215 205 249
rect 316 215 350 249
rect 453 215 487 249
rect 571 215 605 249
rect 811 215 845 249
rect 961 215 995 249
rect 1039 215 1073 249
rect 1117 215 1151 249
rect 1195 215 1229 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 35 477 69 493
rect 35 407 69 443
rect 103 459 179 527
rect 103 425 129 459
rect 163 425 179 459
rect 223 477 257 493
rect 223 407 257 443
rect 291 459 367 527
rect 291 425 317 459
rect 351 425 367 459
rect 411 477 445 493
rect 69 373 223 391
rect 411 407 445 443
rect 479 459 555 527
rect 479 425 505 459
rect 539 425 555 459
rect 623 477 845 493
rect 657 459 811 477
rect 257 373 411 391
rect 623 407 657 443
rect 445 373 623 391
rect 35 357 657 373
rect 691 389 717 423
rect 751 389 767 423
rect 691 343 767 389
rect 811 409 845 443
rect 899 459 965 527
rect 899 425 915 459
rect 949 425 965 459
rect 1009 477 1043 493
rect 1009 407 1043 443
rect 1077 459 1153 527
rect 1077 425 1103 459
rect 1137 425 1153 459
rect 1197 477 1231 493
rect 811 359 845 375
rect 987 373 1009 391
rect 1197 407 1231 443
rect 1265 459 1341 527
rect 1265 425 1291 459
rect 1325 425 1341 459
rect 1043 373 1197 391
rect 1231 373 1356 391
rect 987 357 1356 373
rect 29 289 631 323
rect 29 249 105 289
rect 29 215 55 249
rect 89 215 105 249
rect 155 249 251 255
rect 155 215 171 249
rect 205 215 251 249
rect 291 249 371 255
rect 291 215 316 249
rect 350 215 371 249
rect 437 249 513 255
rect 437 215 453 249
rect 487 215 513 249
rect 555 249 631 289
rect 555 215 571 249
rect 605 215 631 249
rect 691 309 717 343
rect 751 325 767 343
rect 751 309 964 325
rect 691 291 964 309
rect 155 181 251 215
rect 437 181 474 215
rect 35 165 69 181
rect 155 147 474 181
rect 691 174 739 291
rect 930 265 964 291
rect 785 249 891 257
rect 785 215 811 249
rect 845 215 891 249
rect 520 161 739 174
rect 35 97 69 131
rect 520 140 717 161
rect 520 113 554 140
rect 291 79 317 113
rect 351 79 554 113
rect 691 127 717 140
rect 751 127 767 161
rect 843 149 891 215
rect 930 249 1271 265
rect 930 215 961 249
rect 995 215 1039 249
rect 1073 215 1117 249
rect 1151 215 1195 249
rect 1229 215 1271 249
rect 930 199 1271 215
rect 1317 165 1356 357
rect 981 131 1009 165
rect 1043 131 1197 165
rect 1231 131 1356 165
rect 590 90 657 106
rect 35 17 69 63
rect 590 56 619 90
rect 653 56 657 90
rect 691 93 767 127
rect 691 59 717 93
rect 751 59 767 93
rect 827 97 933 113
rect 861 63 899 97
rect 590 17 657 56
rect 827 17 933 63
rect 1077 63 1103 97
rect 1137 63 1153 97
rect 1077 17 1153 63
rect 1265 63 1291 97
rect 1325 63 1341 97
rect 1265 17 1341 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 846 153 880 187 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 213 153 247 187 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 846 221 880 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1317 221 1351 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 1317 153 1351 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 1317 357 1351 391 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1317 289 1351 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1385746
string GDS_START 1375540
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
