magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 3026 1975
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 1 49 1727 256
rect 0 0 1728 49
<< scpmos >>
rect 87 368 117 592
rect 177 368 207 592
rect 267 368 297 592
rect 367 368 397 592
rect 457 368 487 592
rect 557 368 587 592
rect 701 368 731 592
rect 791 368 821 592
rect 1003 368 1033 592
rect 1093 368 1123 592
rect 1183 368 1213 592
rect 1273 368 1303 592
rect 1373 368 1403 592
rect 1612 368 1642 592
<< nmoslvt >>
rect 84 82 114 230
rect 184 82 214 230
rect 270 82 300 230
rect 370 82 400 230
rect 456 82 486 230
rect 604 82 634 230
rect 704 82 734 230
rect 790 82 820 230
rect 876 82 906 230
rect 1064 82 1094 230
rect 1150 82 1180 230
rect 1270 82 1300 230
rect 1356 82 1386 230
rect 1442 82 1472 230
rect 1528 82 1558 230
rect 1614 82 1644 230
<< ndiff >>
rect 27 218 84 230
rect 27 184 39 218
rect 73 184 84 218
rect 27 128 84 184
rect 27 94 39 128
rect 73 94 84 128
rect 27 82 84 94
rect 114 131 184 230
rect 114 97 139 131
rect 173 97 184 131
rect 114 82 184 97
rect 214 218 270 230
rect 214 184 225 218
rect 259 184 270 218
rect 214 82 270 184
rect 300 131 370 230
rect 300 97 311 131
rect 345 97 370 131
rect 300 82 370 97
rect 400 218 456 230
rect 400 184 411 218
rect 445 184 456 218
rect 400 128 456 184
rect 400 94 411 128
rect 445 94 456 128
rect 400 82 456 94
rect 486 151 604 230
rect 486 117 528 151
rect 562 117 604 151
rect 486 82 604 117
rect 634 218 704 230
rect 634 184 645 218
rect 679 184 704 218
rect 634 128 704 184
rect 634 94 645 128
rect 679 94 704 128
rect 634 82 704 94
rect 734 148 790 230
rect 734 114 745 148
rect 779 114 790 148
rect 734 82 790 114
rect 820 218 876 230
rect 820 184 831 218
rect 865 184 876 218
rect 820 128 876 184
rect 820 94 831 128
rect 865 94 876 128
rect 820 82 876 94
rect 906 84 1064 230
rect 906 82 933 84
rect 921 50 933 82
rect 967 50 1003 84
rect 1037 82 1064 84
rect 1094 140 1150 230
rect 1094 106 1105 140
rect 1139 106 1150 140
rect 1094 82 1150 106
rect 1180 82 1270 230
rect 1300 131 1356 230
rect 1300 97 1311 131
rect 1345 97 1356 131
rect 1300 82 1356 97
rect 1386 218 1442 230
rect 1386 184 1397 218
rect 1431 184 1442 218
rect 1386 82 1442 184
rect 1472 131 1528 230
rect 1472 97 1483 131
rect 1517 97 1528 131
rect 1472 82 1528 97
rect 1558 218 1614 230
rect 1558 184 1569 218
rect 1603 184 1614 218
rect 1558 82 1614 184
rect 1644 218 1701 230
rect 1644 184 1655 218
rect 1689 184 1701 218
rect 1644 131 1701 184
rect 1644 97 1655 131
rect 1689 97 1701 131
rect 1644 82 1701 97
rect 1037 50 1049 82
rect 921 38 1049 50
rect 1195 48 1208 82
rect 1242 48 1255 82
rect 1195 36 1255 48
<< pdiff >>
rect 28 580 87 592
rect 28 546 40 580
rect 74 546 87 580
rect 28 510 87 546
rect 28 476 40 510
rect 74 476 87 510
rect 28 440 87 476
rect 28 406 40 440
rect 74 406 87 440
rect 28 368 87 406
rect 117 580 177 592
rect 117 546 130 580
rect 164 546 177 580
rect 117 508 177 546
rect 117 474 130 508
rect 164 474 177 508
rect 117 368 177 474
rect 207 580 267 592
rect 207 546 220 580
rect 254 546 267 580
rect 207 510 267 546
rect 207 476 220 510
rect 254 476 267 510
rect 207 440 267 476
rect 207 406 220 440
rect 254 406 267 440
rect 207 368 267 406
rect 297 580 367 592
rect 297 546 310 580
rect 344 546 367 580
rect 297 508 367 546
rect 297 474 310 508
rect 344 474 367 508
rect 297 368 367 474
rect 397 580 457 592
rect 397 546 410 580
rect 444 546 457 580
rect 397 497 457 546
rect 397 463 410 497
rect 444 463 457 497
rect 397 414 457 463
rect 397 380 410 414
rect 444 380 457 414
rect 397 368 457 380
rect 487 580 557 592
rect 487 546 510 580
rect 544 546 557 580
rect 487 508 557 546
rect 487 474 510 508
rect 544 474 557 508
rect 487 368 557 474
rect 587 531 701 592
rect 587 497 610 531
rect 644 497 701 531
rect 587 440 701 497
rect 587 406 610 440
rect 644 406 701 440
rect 587 368 701 406
rect 731 578 791 592
rect 731 544 744 578
rect 778 544 791 578
rect 731 368 791 544
rect 821 527 890 592
rect 821 493 844 527
rect 878 493 890 527
rect 821 368 890 493
rect 944 531 1003 592
rect 944 497 956 531
rect 990 497 1003 531
rect 944 424 1003 497
rect 944 390 956 424
rect 990 390 1003 424
rect 944 368 1003 390
rect 1033 580 1093 592
rect 1033 546 1046 580
rect 1080 546 1093 580
rect 1033 508 1093 546
rect 1033 474 1046 508
rect 1080 474 1093 508
rect 1033 368 1093 474
rect 1123 531 1183 592
rect 1123 497 1136 531
rect 1170 497 1183 531
rect 1123 440 1183 497
rect 1123 406 1136 440
rect 1170 406 1183 440
rect 1123 368 1183 406
rect 1213 580 1273 592
rect 1213 546 1226 580
rect 1260 546 1273 580
rect 1213 508 1273 546
rect 1213 474 1226 508
rect 1260 474 1273 508
rect 1213 368 1273 474
rect 1303 580 1373 592
rect 1303 546 1326 580
rect 1360 546 1373 580
rect 1303 510 1373 546
rect 1303 476 1326 510
rect 1360 476 1373 510
rect 1303 440 1373 476
rect 1303 406 1326 440
rect 1360 406 1373 440
rect 1303 368 1373 406
rect 1403 580 1612 592
rect 1403 546 1416 580
rect 1450 546 1494 580
rect 1528 546 1565 580
rect 1599 546 1612 580
rect 1403 508 1612 546
rect 1403 474 1416 508
rect 1450 474 1494 508
rect 1528 474 1565 508
rect 1599 474 1612 508
rect 1403 368 1612 474
rect 1642 580 1701 592
rect 1642 546 1655 580
rect 1689 546 1701 580
rect 1642 497 1701 546
rect 1642 463 1655 497
rect 1689 463 1701 497
rect 1642 414 1701 463
rect 1642 380 1655 414
rect 1689 380 1701 414
rect 1642 368 1701 380
<< ndiffc >>
rect 39 184 73 218
rect 39 94 73 128
rect 139 97 173 131
rect 225 184 259 218
rect 311 97 345 131
rect 411 184 445 218
rect 411 94 445 128
rect 528 117 562 151
rect 645 184 679 218
rect 645 94 679 128
rect 745 114 779 148
rect 831 184 865 218
rect 831 94 865 128
rect 933 50 967 84
rect 1003 50 1037 84
rect 1105 106 1139 140
rect 1311 97 1345 131
rect 1397 184 1431 218
rect 1483 97 1517 131
rect 1569 184 1603 218
rect 1655 184 1689 218
rect 1655 97 1689 131
rect 1208 48 1242 82
<< pdiffc >>
rect 40 546 74 580
rect 40 476 74 510
rect 40 406 74 440
rect 130 546 164 580
rect 130 474 164 508
rect 220 546 254 580
rect 220 476 254 510
rect 220 406 254 440
rect 310 546 344 580
rect 310 474 344 508
rect 410 546 444 580
rect 410 463 444 497
rect 410 380 444 414
rect 510 546 544 580
rect 510 474 544 508
rect 610 497 644 531
rect 610 406 644 440
rect 744 544 778 578
rect 844 493 878 527
rect 956 497 990 531
rect 956 390 990 424
rect 1046 546 1080 580
rect 1046 474 1080 508
rect 1136 497 1170 531
rect 1136 406 1170 440
rect 1226 546 1260 580
rect 1226 474 1260 508
rect 1326 546 1360 580
rect 1326 476 1360 510
rect 1326 406 1360 440
rect 1416 546 1450 580
rect 1494 546 1528 580
rect 1565 546 1599 580
rect 1416 474 1450 508
rect 1494 474 1528 508
rect 1565 474 1599 508
rect 1655 546 1689 580
rect 1655 463 1689 497
rect 1655 380 1689 414
<< poly >>
rect 87 592 117 618
rect 177 592 207 618
rect 267 592 297 618
rect 367 592 397 618
rect 457 592 487 618
rect 557 592 587 618
rect 701 592 731 618
rect 791 592 821 618
rect 1003 592 1033 618
rect 1093 592 1123 618
rect 1183 592 1213 618
rect 1273 592 1303 618
rect 1373 592 1403 618
rect 1612 592 1642 618
rect 87 353 117 368
rect 177 353 207 368
rect 267 353 297 368
rect 367 353 397 368
rect 457 353 487 368
rect 557 353 587 368
rect 701 353 731 368
rect 791 353 821 368
rect 1003 353 1033 368
rect 1093 353 1123 368
rect 1183 353 1213 368
rect 1273 353 1303 368
rect 1373 353 1403 368
rect 1612 353 1642 368
rect 84 336 120 353
rect 174 336 210 353
rect 264 336 300 353
rect 84 320 300 336
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 300 300 320
rect 364 300 400 353
rect 454 300 490 353
rect 554 336 590 353
rect 698 336 734 353
rect 788 336 821 353
rect 1000 336 1036 353
rect 1090 336 1126 353
rect 1180 336 1216 353
rect 532 320 820 336
rect 532 300 548 320
rect 270 286 400 300
rect 84 270 400 286
rect 84 230 114 270
rect 184 230 214 270
rect 270 230 300 270
rect 370 230 400 270
rect 456 286 548 300
rect 582 286 616 320
rect 650 286 684 320
rect 718 306 820 320
rect 718 286 734 306
rect 456 270 734 286
rect 456 230 486 270
rect 604 230 634 270
rect 704 230 734 270
rect 790 230 820 306
rect 967 326 1216 336
rect 1270 326 1303 353
rect 1370 336 1406 353
rect 967 320 1300 326
rect 967 300 983 320
rect 876 286 983 300
rect 1017 286 1051 320
rect 1085 286 1119 320
rect 1153 296 1300 320
rect 1153 286 1180 296
rect 876 270 1180 286
rect 876 230 906 270
rect 1064 230 1094 270
rect 1150 230 1180 270
rect 1270 230 1300 296
rect 1356 320 1558 336
rect 1356 286 1372 320
rect 1406 286 1440 320
rect 1474 286 1508 320
rect 1542 300 1558 320
rect 1609 300 1645 353
rect 1542 286 1645 300
rect 1356 270 1645 286
rect 1356 230 1386 270
rect 1442 230 1472 270
rect 1528 230 1558 270
rect 1614 245 1645 270
rect 1614 230 1644 245
rect 84 56 114 82
rect 184 56 214 82
rect 270 56 300 82
rect 370 56 400 82
rect 456 56 486 82
rect 604 56 634 82
rect 704 56 734 82
rect 790 56 820 82
rect 876 56 906 82
rect 1064 56 1094 82
rect 1150 56 1180 82
rect 1270 56 1300 82
rect 1356 56 1386 82
rect 1442 56 1472 82
rect 1528 56 1558 82
rect 1614 56 1644 82
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 236 286 270 320
rect 548 286 582 320
rect 616 286 650 320
rect 684 286 718 320
rect 983 286 1017 320
rect 1051 286 1085 320
rect 1119 286 1153 320
rect 1372 286 1406 320
rect 1440 286 1474 320
rect 1508 286 1542 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 24 580 74 596
rect 24 546 40 580
rect 24 510 74 546
rect 24 476 40 510
rect 24 440 74 476
rect 114 580 180 649
rect 114 546 130 580
rect 164 546 180 580
rect 114 508 180 546
rect 114 474 130 508
rect 164 474 180 508
rect 114 458 180 474
rect 220 580 254 596
rect 220 510 254 546
rect 24 406 40 440
rect 220 440 254 476
rect 294 580 360 649
rect 294 546 310 580
rect 344 546 360 580
rect 294 508 360 546
rect 294 474 310 508
rect 344 474 360 508
rect 294 458 360 474
rect 394 580 460 596
rect 394 546 410 580
rect 444 546 460 580
rect 394 497 460 546
rect 394 463 410 497
rect 444 463 460 497
rect 74 406 220 424
rect 394 424 460 463
rect 494 581 1276 615
rect 494 580 560 581
rect 494 546 510 580
rect 544 546 560 580
rect 728 578 794 581
rect 494 508 560 546
rect 494 474 510 508
rect 544 474 560 508
rect 494 458 560 474
rect 594 531 660 547
rect 728 544 744 578
rect 778 544 794 578
rect 1030 580 1080 581
rect 728 542 794 544
rect 594 497 610 531
rect 644 508 660 531
rect 828 527 894 547
rect 828 508 844 527
rect 644 497 844 508
rect 594 493 844 497
rect 878 493 894 527
rect 594 474 894 493
rect 940 531 994 547
rect 940 497 956 531
rect 990 497 994 531
rect 594 440 660 474
rect 594 424 610 440
rect 254 414 610 424
rect 254 406 410 414
rect 24 390 410 406
rect 394 380 410 390
rect 444 406 610 414
rect 644 406 660 440
rect 940 430 994 497
rect 1030 546 1046 580
rect 1226 580 1276 581
rect 1030 508 1080 546
rect 1030 474 1046 508
rect 1030 458 1080 474
rect 1120 531 1186 547
rect 1120 497 1136 531
rect 1170 497 1186 531
rect 444 390 660 406
rect 793 424 994 430
rect 1120 440 1186 497
rect 1260 546 1276 580
rect 1226 508 1276 546
rect 1260 474 1276 508
rect 1226 458 1276 474
rect 1310 580 1376 596
rect 1310 546 1326 580
rect 1360 546 1376 580
rect 1310 510 1376 546
rect 1310 476 1326 510
rect 1360 476 1376 510
rect 1120 424 1136 440
rect 793 390 956 424
rect 990 406 1136 424
rect 1170 424 1186 440
rect 1310 440 1376 476
rect 1410 580 1605 649
rect 1410 546 1416 580
rect 1450 546 1494 580
rect 1528 546 1565 580
rect 1599 546 1605 580
rect 1410 508 1605 546
rect 1410 474 1416 508
rect 1450 474 1494 508
rect 1528 474 1565 508
rect 1599 474 1605 508
rect 1410 458 1605 474
rect 1639 580 1705 596
rect 1639 546 1655 580
rect 1689 546 1705 580
rect 1639 497 1705 546
rect 1639 463 1655 497
rect 1689 463 1705 497
rect 1310 424 1326 440
rect 1170 406 1326 424
rect 1360 424 1376 440
rect 1639 424 1705 463
rect 1360 414 1705 424
rect 1360 406 1655 414
rect 990 390 1655 406
rect 444 380 460 390
rect 394 364 460 380
rect 25 320 359 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 359 320
rect 25 270 359 286
rect 505 320 743 356
rect 505 286 548 320
rect 582 286 616 320
rect 650 286 684 320
rect 718 286 743 320
rect 793 310 933 390
rect 1639 380 1655 390
rect 1689 380 1705 414
rect 1639 364 1705 380
rect 505 270 743 286
rect 899 236 933 310
rect 967 320 1223 356
rect 967 286 983 320
rect 1017 286 1051 320
rect 1085 286 1119 320
rect 1153 286 1223 320
rect 967 270 1223 286
rect 1273 320 1558 356
rect 1273 286 1372 320
rect 1406 286 1440 320
rect 1474 286 1508 320
rect 1542 286 1558 320
rect 1273 270 1558 286
rect 23 218 865 236
rect 23 184 39 218
rect 73 184 225 218
rect 259 184 411 218
rect 445 202 645 218
rect 445 184 461 202
rect 23 128 89 184
rect 23 94 39 128
rect 73 94 89 128
rect 23 78 89 94
rect 123 131 189 150
rect 123 97 139 131
rect 173 97 189 131
rect 123 17 189 97
rect 295 131 361 150
rect 295 97 311 131
rect 345 97 361 131
rect 295 17 361 97
rect 395 128 461 184
rect 629 184 645 202
rect 679 202 831 218
rect 679 184 695 202
rect 395 94 411 128
rect 445 94 461 128
rect 395 78 461 94
rect 499 151 592 161
rect 499 117 528 151
rect 562 117 592 151
rect 499 17 592 117
rect 629 128 695 184
rect 899 218 1619 236
rect 899 202 1397 218
rect 1381 184 1397 202
rect 1431 184 1569 218
rect 1603 184 1619 218
rect 1653 218 1705 234
rect 1653 184 1655 218
rect 1689 184 1705 218
rect 831 168 865 184
rect 629 94 645 128
rect 679 94 695 128
rect 629 78 695 94
rect 729 148 795 168
rect 729 114 745 148
rect 779 114 795 148
rect 729 17 795 114
rect 831 150 1155 168
rect 831 140 1361 150
rect 831 134 1105 140
rect 831 128 865 134
rect 1089 106 1105 134
rect 1139 131 1361 140
rect 1139 116 1311 131
rect 1139 106 1155 116
rect 831 78 865 94
rect 917 84 1053 100
rect 917 50 933 84
rect 967 50 1003 84
rect 1037 50 1053 84
rect 1089 78 1155 106
rect 1295 97 1311 116
rect 1345 112 1361 131
rect 1467 131 1533 150
rect 1467 112 1483 131
rect 1345 97 1483 112
rect 1517 112 1533 131
rect 1653 131 1705 184
rect 1653 112 1655 131
rect 1517 97 1655 112
rect 1689 97 1705 131
rect 917 17 1053 50
rect 1191 48 1208 82
rect 1242 48 1259 82
rect 1295 78 1705 97
rect 1191 17 1259 48
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o31ai_4
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 295936
string GDS_START 282224
<< end >>
