magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 753 157
rect 0 0 768 49
<< scnmos >>
rect 80 47 110 131
rect 245 47 275 131
rect 333 47 363 131
rect 425 47 455 131
rect 533 47 563 131
rect 641 47 671 131
<< scpmoshvt >>
rect 153 429 183 557
rect 239 429 269 557
rect 344 429 374 557
rect 449 429 479 557
rect 539 429 569 557
rect 625 429 655 557
<< ndiff >>
rect 27 101 80 131
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 95 245 131
rect 110 61 121 95
rect 155 61 200 95
rect 234 61 245 95
rect 110 47 245 61
rect 275 47 333 131
rect 363 47 425 131
rect 455 106 533 131
rect 455 72 476 106
rect 510 72 533 106
rect 455 47 533 72
rect 563 47 641 131
rect 671 106 727 131
rect 671 72 685 106
rect 719 72 727 106
rect 671 47 727 72
<< pdiff >>
rect 100 545 153 557
rect 100 511 108 545
rect 142 511 153 545
rect 100 475 153 511
rect 100 441 108 475
rect 142 441 153 475
rect 100 429 153 441
rect 183 545 239 557
rect 183 511 194 545
rect 228 511 239 545
rect 183 475 239 511
rect 183 441 194 475
rect 228 441 239 475
rect 183 429 239 441
rect 269 545 344 557
rect 269 511 291 545
rect 325 511 344 545
rect 269 475 344 511
rect 269 441 291 475
rect 325 441 344 475
rect 269 429 344 441
rect 374 549 449 557
rect 374 515 389 549
rect 423 515 449 549
rect 374 475 449 515
rect 374 441 389 475
rect 423 441 449 475
rect 374 429 449 441
rect 479 543 539 557
rect 479 509 490 543
rect 524 509 539 543
rect 479 475 539 509
rect 479 441 490 475
rect 524 441 539 475
rect 479 429 539 441
rect 569 545 625 557
rect 569 511 580 545
rect 614 511 625 545
rect 569 471 625 511
rect 569 437 580 471
rect 614 437 625 471
rect 569 429 625 437
rect 655 545 708 557
rect 655 511 666 545
rect 700 511 708 545
rect 655 475 708 511
rect 655 441 666 475
rect 700 441 708 475
rect 655 429 708 441
<< ndiffc >>
rect 35 67 69 101
rect 121 61 155 95
rect 200 61 234 95
rect 476 72 510 106
rect 685 72 719 106
<< pdiffc >>
rect 108 511 142 545
rect 108 441 142 475
rect 194 511 228 545
rect 194 441 228 475
rect 291 511 325 545
rect 291 441 325 475
rect 389 515 423 549
rect 389 441 423 475
rect 490 509 524 543
rect 490 441 524 475
rect 580 511 614 545
rect 580 437 614 471
rect 666 511 700 545
rect 666 441 700 475
<< poly >>
rect 153 557 183 583
rect 239 557 269 583
rect 344 557 374 583
rect 449 557 479 583
rect 539 557 569 583
rect 625 557 655 583
rect 153 399 183 429
rect 80 375 183 399
rect 80 341 101 375
rect 135 369 183 375
rect 135 341 151 369
rect 80 307 151 341
rect 239 321 269 429
rect 344 337 374 429
rect 317 321 383 337
rect 80 273 101 307
rect 135 273 151 307
rect 80 257 151 273
rect 193 305 275 321
rect 193 271 209 305
rect 243 271 275 305
rect 80 131 110 257
rect 193 237 275 271
rect 193 203 209 237
rect 243 203 275 237
rect 317 287 333 321
rect 367 287 383 321
rect 449 302 479 429
rect 539 302 569 429
rect 625 380 655 429
rect 625 350 711 380
rect 681 325 711 350
rect 681 309 747 325
rect 317 253 383 287
rect 317 219 333 253
rect 367 219 383 253
rect 317 203 383 219
rect 425 286 491 302
rect 425 252 441 286
rect 475 252 491 286
rect 425 218 491 252
rect 193 187 275 203
rect 245 131 275 187
rect 333 131 363 203
rect 425 184 441 218
rect 475 184 491 218
rect 425 168 491 184
rect 533 286 599 302
rect 533 252 549 286
rect 583 252 599 286
rect 533 218 599 252
rect 681 275 697 309
rect 731 275 747 309
rect 681 241 747 275
rect 681 221 697 241
rect 533 184 549 218
rect 583 184 599 218
rect 533 168 599 184
rect 641 207 697 221
rect 731 207 747 241
rect 641 191 747 207
rect 425 131 455 168
rect 533 131 563 168
rect 641 131 671 191
rect 80 21 110 47
rect 245 21 275 47
rect 333 21 363 47
rect 425 21 455 47
rect 533 21 563 47
rect 641 21 671 47
<< polycont >>
rect 101 341 135 375
rect 101 273 135 307
rect 209 271 243 305
rect 209 203 243 237
rect 333 287 367 321
rect 333 219 367 253
rect 441 252 475 286
rect 441 184 475 218
rect 549 252 583 286
rect 697 275 731 309
rect 549 184 583 218
rect 697 207 731 241
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 545 151 587
rect 17 511 108 545
rect 142 511 151 545
rect 17 475 151 511
rect 17 441 108 475
rect 142 441 151 475
rect 17 425 151 441
rect 185 545 241 649
rect 185 511 194 545
rect 228 511 241 545
rect 185 475 241 511
rect 185 441 194 475
rect 228 441 241 475
rect 185 425 241 441
rect 275 545 339 561
rect 275 511 291 545
rect 325 511 339 545
rect 275 475 339 511
rect 275 441 291 475
rect 325 441 339 475
rect 373 549 439 649
rect 373 515 389 549
rect 423 515 439 549
rect 373 475 439 515
rect 373 441 389 475
rect 423 441 439 475
rect 473 579 720 613
rect 473 543 530 579
rect 664 545 720 579
rect 473 509 490 543
rect 524 509 530 543
rect 473 475 530 509
rect 473 441 490 475
rect 524 441 530 475
rect 17 117 67 425
rect 275 407 339 441
rect 473 407 530 441
rect 275 406 530 407
rect 101 375 151 391
rect 135 341 151 375
rect 295 373 530 406
rect 564 511 580 545
rect 614 511 630 545
rect 564 471 630 511
rect 564 437 580 471
rect 614 437 630 471
rect 564 391 630 437
rect 664 511 666 545
rect 700 511 720 545
rect 664 475 720 511
rect 664 441 666 475
rect 700 441 720 475
rect 664 425 720 441
rect 101 307 151 341
rect 135 273 151 307
rect 101 169 151 273
rect 193 349 261 372
rect 564 357 651 391
rect 193 305 270 349
rect 193 271 209 305
rect 243 271 270 305
rect 193 237 270 271
rect 193 203 209 237
rect 243 203 270 237
rect 304 321 370 337
rect 304 287 333 321
rect 367 287 370 321
rect 304 253 370 287
rect 304 219 333 253
rect 367 219 370 253
rect 304 203 370 219
rect 404 286 475 302
rect 404 252 441 286
rect 404 218 475 252
rect 404 184 441 218
rect 101 135 370 169
rect 404 156 475 184
rect 509 286 583 302
rect 509 252 549 286
rect 509 218 583 252
rect 509 184 549 218
rect 509 156 583 184
rect 319 122 370 135
rect 617 122 651 357
rect 685 309 751 370
rect 685 275 697 309
rect 731 275 751 309
rect 685 241 751 275
rect 685 207 697 241
rect 731 207 751 241
rect 685 156 751 207
rect 17 101 71 117
rect 319 106 651 122
rect 17 67 35 101
rect 69 67 71 101
rect 17 51 71 67
rect 105 95 250 101
rect 105 61 121 95
rect 155 61 200 95
rect 234 61 250 95
rect 105 17 250 61
rect 319 72 476 106
rect 510 72 651 106
rect 319 56 651 72
rect 685 106 735 122
rect 719 72 735 106
rect 685 17 735 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a32o_0
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2036860
string GDS_START 2028578
<< end >>
