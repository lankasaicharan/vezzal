magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2218 1852
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 855 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 371 47 401 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 747 47 777 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
<< ndiff >>
rect 27 161 89 177
rect 27 127 35 161
rect 69 127 89 161
rect 27 93 89 127
rect 27 59 35 93
rect 69 59 89 93
rect 27 47 89 59
rect 119 93 183 177
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 161 277 177
rect 213 127 223 161
rect 257 127 277 161
rect 213 93 277 127
rect 213 59 223 93
rect 257 59 277 93
rect 213 47 277 59
rect 307 93 371 177
rect 307 59 317 93
rect 351 59 371 93
rect 307 47 371 59
rect 401 161 455 177
rect 401 127 411 161
rect 445 127 455 161
rect 401 93 455 127
rect 401 59 411 93
rect 445 59 455 93
rect 401 47 455 59
rect 485 161 549 177
rect 485 127 505 161
rect 539 127 549 161
rect 485 47 549 127
rect 579 93 643 177
rect 579 59 599 93
rect 633 59 643 93
rect 579 47 643 59
rect 673 161 747 177
rect 673 127 693 161
rect 727 127 747 161
rect 673 47 747 127
rect 777 161 829 177
rect 777 127 787 161
rect 821 127 829 161
rect 777 93 829 127
rect 777 59 787 93
rect 821 59 829 93
rect 777 47 829 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 349 551 383
rect 493 315 505 349
rect 539 315 551 349
rect 493 297 551 315
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 417 645 451
rect 587 383 599 417
rect 633 383 645 417
rect 587 297 645 383
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 349 739 383
rect 681 315 693 349
rect 727 315 739 349
rect 681 297 739 315
rect 775 485 829 497
rect 775 451 787 485
rect 821 451 829 485
rect 775 417 829 451
rect 775 383 787 417
rect 821 383 829 417
rect 775 297 829 383
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 59 163 93
rect 223 127 257 161
rect 223 59 257 93
rect 317 59 351 93
rect 411 127 445 161
rect 411 59 445 93
rect 505 127 539 161
rect 599 59 633 93
rect 693 127 727 161
rect 787 127 821 161
rect 787 59 821 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 505 451 539 485
rect 505 383 539 417
rect 505 315 539 349
rect 599 451 633 485
rect 599 383 633 417
rect 693 451 727 485
rect 693 383 727 417
rect 693 315 727 349
rect 787 451 821 485
rect 787 383 821 417
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 22 249 401 265
rect 22 215 38 249
rect 72 215 129 249
rect 163 215 223 249
rect 257 215 317 249
rect 351 215 401 249
rect 22 199 401 215
rect 89 177 119 199
rect 183 177 213 199
rect 277 177 307 199
rect 371 177 401 199
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 455 249 777 265
rect 455 215 599 249
rect 633 215 693 249
rect 727 215 777 249
rect 455 199 777 215
rect 455 177 485 199
rect 549 177 579 199
rect 643 177 673 199
rect 747 177 777 199
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 371 21 401 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 747 21 777 47
<< polycont >>
rect 38 215 72 249
rect 129 215 163 249
rect 223 215 257 249
rect 317 215 351 249
rect 599 215 633 249
rect 693 215 727 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 485 179 493
rect 103 451 129 485
rect 163 451 179 485
rect 103 417 179 451
rect 103 383 129 417
rect 163 383 179 417
rect 103 349 179 383
rect 223 485 257 527
rect 223 417 257 451
rect 223 367 257 383
rect 291 485 367 493
rect 291 451 317 485
rect 351 451 367 485
rect 291 417 367 451
rect 291 383 317 417
rect 351 383 367 417
rect 103 315 129 349
rect 163 333 179 349
rect 291 349 367 383
rect 411 485 445 527
rect 411 417 445 451
rect 411 367 445 383
rect 479 485 555 493
rect 479 451 505 485
rect 539 451 555 485
rect 479 417 555 451
rect 479 383 505 417
rect 539 383 555 417
rect 291 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 479 349 555 383
rect 599 485 633 527
rect 599 417 633 451
rect 599 367 633 383
rect 667 485 743 493
rect 667 451 693 485
rect 727 451 743 485
rect 667 417 743 451
rect 667 383 693 417
rect 727 383 743 417
rect 479 333 505 349
rect 351 315 505 333
rect 539 333 555 349
rect 667 349 743 383
rect 787 485 837 527
rect 821 451 837 485
rect 787 417 837 451
rect 821 383 837 417
rect 787 367 837 383
rect 667 333 693 349
rect 539 315 693 333
rect 727 315 743 349
rect 103 299 743 315
rect 22 249 376 265
rect 22 215 38 249
rect 72 215 129 249
rect 163 215 223 249
rect 257 215 317 249
rect 351 215 376 249
rect 18 161 445 181
rect 18 127 35 161
rect 69 143 223 161
rect 69 127 85 143
rect 18 93 85 127
rect 197 127 223 143
rect 257 143 411 161
rect 257 127 273 143
rect 18 59 35 93
rect 69 59 85 93
rect 18 51 85 59
rect 129 93 163 109
rect 129 17 163 59
rect 197 93 273 127
rect 385 127 411 143
rect 479 161 539 299
rect 573 249 823 265
rect 573 215 599 249
rect 633 215 693 249
rect 727 215 823 249
rect 787 161 837 177
rect 479 127 505 161
rect 539 127 693 161
rect 727 127 743 161
rect 821 127 837 161
rect 197 59 223 93
rect 257 59 273 93
rect 197 51 273 59
rect 317 93 351 109
rect 317 17 351 59
rect 385 93 445 127
rect 787 93 837 127
rect 385 59 411 93
rect 445 59 599 93
rect 633 59 787 93
rect 821 59 837 93
rect 385 51 837 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 489 221 523 255 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 489 289 523 323 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 673 221 707 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2189644
string GDS_START 2181726
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
