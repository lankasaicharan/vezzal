magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2678 1852
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 873 157 1343 203
rect 11 21 1343 157
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 131
rect 173 47 203 131
rect 381 47 411 131
rect 470 47 500 131
rect 574 47 604 119
rect 678 47 708 131
rect 750 47 780 131
rect 951 47 981 177
rect 1032 47 1062 177
rect 1139 47 1169 177
rect 1223 47 1253 177
<< scpmoshvt >>
rect 81 363 117 491
rect 175 363 211 491
rect 373 369 409 497
rect 467 369 503 497
rect 572 413 608 497
rect 666 413 702 497
rect 762 413 798 497
rect 943 297 979 497
rect 1037 297 1073 497
rect 1131 297 1167 497
rect 1225 297 1261 497
<< ndiff >>
rect 37 106 89 131
rect 37 72 45 106
rect 79 72 89 106
rect 37 47 89 72
rect 119 93 173 131
rect 119 59 129 93
rect 163 59 173 93
rect 119 47 173 59
rect 203 106 255 131
rect 203 72 213 106
rect 247 72 255 106
rect 203 47 255 72
rect 329 119 381 131
rect 329 85 337 119
rect 371 85 381 119
rect 329 47 381 85
rect 411 89 470 131
rect 411 55 421 89
rect 455 55 470 89
rect 411 47 470 55
rect 500 119 550 131
rect 899 165 951 177
rect 899 131 907 165
rect 941 131 951 165
rect 628 119 678 131
rect 500 47 574 119
rect 604 106 678 119
rect 604 72 624 106
rect 658 72 678 106
rect 604 47 678 72
rect 708 47 750 131
rect 780 106 832 131
rect 780 72 790 106
rect 824 72 832 106
rect 780 47 832 72
rect 899 93 951 131
rect 899 59 907 93
rect 941 59 951 93
rect 899 47 951 59
rect 981 47 1032 177
rect 1062 165 1139 177
rect 1062 131 1079 165
rect 1113 131 1139 165
rect 1062 93 1139 131
rect 1062 59 1079 93
rect 1113 59 1139 93
rect 1062 47 1139 59
rect 1169 161 1223 177
rect 1169 127 1179 161
rect 1213 127 1223 161
rect 1169 93 1223 127
rect 1169 59 1179 93
rect 1213 59 1223 93
rect 1169 47 1223 59
rect 1253 161 1317 177
rect 1253 127 1275 161
rect 1309 127 1317 161
rect 1253 93 1317 127
rect 1253 59 1275 93
rect 1309 59 1317 93
rect 1253 47 1317 59
<< pdiff >>
rect 27 477 81 491
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 363 81 375
rect 117 461 175 491
rect 117 427 129 461
rect 163 427 175 461
rect 117 363 175 427
rect 211 477 265 491
rect 211 443 223 477
rect 257 443 265 477
rect 211 409 265 443
rect 211 375 223 409
rect 257 375 265 409
rect 211 363 265 375
rect 319 483 373 497
rect 319 449 327 483
rect 361 449 373 483
rect 319 415 373 449
rect 319 381 327 415
rect 361 381 373 415
rect 319 369 373 381
rect 409 485 467 497
rect 409 451 421 485
rect 455 451 467 485
rect 409 417 467 451
rect 409 383 421 417
rect 455 383 467 417
rect 409 369 467 383
rect 503 413 572 497
rect 608 472 666 497
rect 608 438 620 472
rect 654 438 666 472
rect 608 413 666 438
rect 702 413 762 497
rect 798 477 943 497
rect 798 443 810 477
rect 844 443 892 477
rect 926 443 943 477
rect 798 413 943 443
rect 503 369 555 413
rect 886 297 943 413
rect 979 477 1037 497
rect 979 443 991 477
rect 1025 443 1037 477
rect 979 409 1037 443
rect 979 375 991 409
rect 1025 375 1037 409
rect 979 341 1037 375
rect 979 307 991 341
rect 1025 307 1037 341
rect 979 297 1037 307
rect 1073 485 1131 497
rect 1073 451 1085 485
rect 1119 451 1131 485
rect 1073 411 1131 451
rect 1073 377 1085 411
rect 1119 377 1131 411
rect 1073 297 1131 377
rect 1167 485 1225 497
rect 1167 451 1179 485
rect 1213 451 1225 485
rect 1167 417 1225 451
rect 1167 383 1179 417
rect 1213 383 1225 417
rect 1167 349 1225 383
rect 1167 315 1179 349
rect 1213 315 1225 349
rect 1167 297 1225 315
rect 1261 485 1317 497
rect 1261 451 1275 485
rect 1309 451 1317 485
rect 1261 417 1317 451
rect 1261 383 1275 417
rect 1309 383 1317 417
rect 1261 349 1317 383
rect 1261 315 1275 349
rect 1309 315 1317 349
rect 1261 297 1317 315
<< ndiffc >>
rect 45 72 79 106
rect 129 59 163 93
rect 213 72 247 106
rect 337 85 371 119
rect 421 55 455 89
rect 907 131 941 165
rect 624 72 658 106
rect 790 72 824 106
rect 907 59 941 93
rect 1079 131 1113 165
rect 1079 59 1113 93
rect 1179 127 1213 161
rect 1179 59 1213 93
rect 1275 127 1309 161
rect 1275 59 1309 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 427 163 461
rect 223 443 257 477
rect 223 375 257 409
rect 327 449 361 483
rect 327 381 361 415
rect 421 451 455 485
rect 421 383 455 417
rect 620 438 654 472
rect 810 443 844 477
rect 892 443 926 477
rect 991 443 1025 477
rect 991 375 1025 409
rect 991 307 1025 341
rect 1085 451 1119 485
rect 1085 377 1119 411
rect 1179 451 1213 485
rect 1179 383 1213 417
rect 1179 315 1213 349
rect 1275 451 1309 485
rect 1275 383 1309 417
rect 1275 315 1309 349
<< poly >>
rect 81 491 117 517
rect 175 491 211 517
rect 373 497 409 523
rect 467 497 503 523
rect 572 497 608 523
rect 666 497 702 523
rect 762 497 798 523
rect 943 497 979 523
rect 1037 497 1073 523
rect 1131 497 1167 523
rect 1225 497 1261 523
rect 572 398 608 413
rect 666 398 702 413
rect 762 398 798 413
rect 81 348 117 363
rect 175 348 211 363
rect 373 354 409 369
rect 467 354 503 369
rect 45 318 119 348
rect 173 318 213 348
rect 45 280 87 318
rect 33 264 87 280
rect 173 274 203 318
rect 33 230 43 264
rect 77 230 87 264
rect 33 214 87 230
rect 129 264 203 274
rect 371 265 411 354
rect 129 230 145 264
rect 179 230 203 264
rect 129 220 203 230
rect 45 176 87 214
rect 45 146 119 176
rect 89 131 119 146
rect 173 131 203 220
rect 293 249 411 265
rect 293 215 303 249
rect 337 215 411 249
rect 465 219 505 354
rect 570 327 610 398
rect 664 375 704 398
rect 547 305 610 327
rect 652 365 718 375
rect 652 331 668 365
rect 702 331 718 365
rect 652 321 718 331
rect 760 373 800 398
rect 760 357 852 373
rect 760 323 804 357
rect 838 323 852 357
rect 547 271 557 305
rect 591 279 610 305
rect 760 307 852 323
rect 760 285 790 307
rect 591 271 708 279
rect 547 249 708 271
rect 293 199 411 215
rect 381 131 411 199
rect 453 203 507 219
rect 453 169 463 203
rect 497 169 507 203
rect 453 153 507 169
rect 556 197 622 207
rect 556 163 572 197
rect 606 163 622 197
rect 470 131 500 153
rect 556 147 622 163
rect 574 119 604 147
rect 678 131 708 249
rect 750 255 790 285
rect 943 282 979 297
rect 1037 282 1073 297
rect 1131 282 1167 297
rect 1225 282 1261 297
rect 941 265 981 282
rect 1035 265 1075 282
rect 1129 265 1169 282
rect 1223 265 1263 282
rect 750 131 780 255
rect 832 249 981 265
rect 832 215 842 249
rect 876 235 981 249
rect 876 215 886 235
rect 832 199 886 215
rect 951 177 981 235
rect 1023 249 1077 265
rect 1023 215 1033 249
rect 1067 215 1077 249
rect 1023 199 1077 215
rect 1119 249 1263 265
rect 1119 215 1129 249
rect 1163 215 1263 249
rect 1119 199 1263 215
rect 1032 177 1062 199
rect 1139 177 1169 199
rect 1223 177 1253 199
rect 89 21 119 47
rect 173 21 203 47
rect 381 21 411 47
rect 470 21 500 47
rect 574 21 604 47
rect 678 21 708 47
rect 750 21 780 47
rect 951 21 981 47
rect 1032 21 1062 47
rect 1139 21 1169 47
rect 1223 21 1253 47
<< polycont >>
rect 43 230 77 264
rect 145 230 179 264
rect 303 215 337 249
rect 668 331 702 365
rect 804 323 838 357
rect 557 271 591 305
rect 463 169 497 203
rect 572 163 606 197
rect 842 215 876 249
rect 1033 215 1067 249
rect 1129 215 1163 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 17 477 79 493
rect 17 443 35 477
rect 69 443 79 477
rect 17 409 79 443
rect 113 461 179 527
rect 113 427 129 461
rect 163 427 179 461
rect 213 477 267 493
rect 213 443 223 477
rect 257 443 267 477
rect 17 375 35 409
rect 69 393 79 409
rect 213 409 267 443
rect 69 375 155 393
rect 17 359 155 375
rect 17 264 87 325
rect 17 230 43 264
rect 77 230 87 264
rect 17 197 87 230
rect 121 323 155 359
rect 121 280 155 289
rect 213 357 223 409
rect 257 357 267 409
rect 213 337 267 357
rect 311 483 377 493
rect 311 449 327 483
rect 361 449 377 483
rect 311 415 377 449
rect 311 381 327 415
rect 361 381 377 415
rect 121 264 179 280
rect 121 230 145 264
rect 121 214 179 230
rect 121 161 155 214
rect 45 127 155 161
rect 45 106 79 127
rect 213 106 247 337
rect 311 333 377 381
rect 411 485 465 527
rect 411 451 421 485
rect 455 451 465 485
rect 810 477 927 527
rect 411 417 465 451
rect 604 472 770 477
rect 604 438 620 472
rect 654 438 770 472
rect 604 433 770 438
rect 411 383 421 417
rect 455 383 465 417
rect 411 367 465 383
rect 625 391 702 399
rect 625 357 656 391
rect 690 365 702 391
rect 311 299 423 333
rect 287 249 353 265
rect 287 215 303 249
rect 337 215 353 249
rect 287 191 353 215
rect 389 219 423 299
rect 489 323 591 337
rect 489 289 545 323
rect 579 305 591 323
rect 489 271 557 289
rect 489 253 591 271
rect 625 331 668 357
rect 625 315 702 331
rect 625 219 659 315
rect 736 265 770 433
rect 844 443 892 477
rect 926 443 927 477
rect 810 427 927 443
rect 977 477 1034 493
rect 977 443 991 477
rect 1025 443 1034 477
rect 977 409 1034 443
rect 977 375 991 409
rect 1025 375 1034 409
rect 1069 485 1129 527
rect 1069 451 1085 485
rect 1119 451 1129 485
rect 1163 485 1241 491
rect 1163 451 1179 485
rect 1213 451 1241 485
rect 1069 430 1129 451
rect 1069 411 1135 430
rect 1069 377 1085 411
rect 1119 377 1135 411
rect 1179 417 1241 451
rect 1213 383 1241 417
rect 977 373 1034 375
rect 804 357 1034 373
rect 838 341 1034 357
rect 1179 349 1241 383
rect 838 323 991 341
rect 804 307 991 323
rect 1025 307 1145 341
rect 736 249 876 265
rect 736 233 842 249
rect 389 203 507 219
rect 389 169 463 203
rect 497 169 507 203
rect 389 157 507 169
rect 45 56 79 72
rect 113 59 129 93
rect 163 59 179 93
rect 113 17 179 59
rect 213 56 247 72
rect 332 153 507 157
rect 556 197 659 219
rect 556 163 572 197
rect 606 163 659 197
rect 332 123 423 153
rect 556 147 659 163
rect 698 215 842 233
rect 698 199 876 215
rect 332 119 371 123
rect 332 85 337 119
rect 698 113 732 199
rect 910 165 944 307
rect 1111 265 1145 307
rect 1213 315 1241 349
rect 1179 299 1241 315
rect 1275 485 1316 527
rect 1309 451 1316 485
rect 1275 417 1316 451
rect 1309 383 1316 417
rect 1275 349 1316 383
rect 1309 315 1316 349
rect 1275 299 1316 315
rect 1207 265 1241 299
rect 978 249 1077 265
rect 978 215 1033 249
rect 1067 215 1077 249
rect 978 199 1077 215
rect 1111 249 1173 265
rect 1111 215 1129 249
rect 1163 215 1173 249
rect 1111 199 1173 215
rect 1207 211 1287 265
rect 1207 165 1241 211
rect 891 131 907 165
rect 941 131 957 165
rect 608 106 732 113
rect 332 69 371 85
rect 405 55 421 89
rect 455 55 471 89
rect 608 72 624 106
rect 658 72 732 106
rect 608 56 732 72
rect 774 106 840 122
rect 774 72 790 106
rect 824 72 840 106
rect 405 17 471 55
rect 774 17 840 72
rect 891 93 957 131
rect 891 59 907 93
rect 941 59 957 93
rect 891 51 957 59
rect 1063 131 1079 165
rect 1113 131 1129 165
rect 1063 93 1129 131
rect 1063 59 1079 93
rect 1113 59 1129 93
rect 1063 17 1129 59
rect 1163 161 1241 165
rect 1163 127 1179 161
rect 1213 127 1241 161
rect 1163 93 1241 127
rect 1163 59 1179 93
rect 1213 59 1241 93
rect 1163 51 1241 59
rect 1275 161 1317 177
rect 1309 127 1317 161
rect 1275 93 1317 127
rect 1309 59 1317 93
rect 1275 17 1317 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 121 289 155 323
rect 223 375 257 391
rect 223 357 257 375
rect 656 365 690 391
rect 656 357 668 365
rect 668 357 690 365
rect 545 305 579 323
rect 545 289 557 305
rect 557 289 579 305
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 211 391 269 397
rect 211 357 223 391
rect 257 388 269 391
rect 644 391 702 397
rect 644 388 656 391
rect 257 360 656 388
rect 257 357 269 360
rect 211 351 269 357
rect 644 357 656 360
rect 690 357 702 391
rect 644 351 702 357
rect 109 323 167 329
rect 109 289 121 323
rect 155 320 167 323
rect 533 323 591 329
rect 533 320 545 323
rect 155 292 545 320
rect 155 289 167 292
rect 109 283 167 289
rect 533 289 545 292
rect 579 289 591 323
rect 533 283 591 289
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 1041 221 1075 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 GATE
port 2 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew signal input
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 dlrtp_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 772238
string GDS_START 760736
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string path 0.000 0.000 34.500 0.000 
<< end >>
