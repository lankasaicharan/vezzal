magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 37 49 859 259
rect 0 0 864 49
<< scnmos >>
rect 116 65 146 233
rect 202 65 232 233
rect 288 65 318 233
rect 374 65 404 233
rect 460 65 490 233
rect 546 65 576 233
rect 664 65 694 233
rect 750 65 780 233
<< scpmoshvt >>
rect 116 367 146 619
rect 202 367 232 619
rect 288 367 318 619
rect 374 367 404 619
rect 460 367 490 619
rect 546 367 576 619
rect 664 367 694 619
rect 750 367 780 619
<< ndiff >>
rect 63 221 116 233
rect 63 187 71 221
rect 105 187 116 221
rect 63 111 116 187
rect 63 77 71 111
rect 105 77 116 111
rect 63 65 116 77
rect 146 183 202 233
rect 146 149 157 183
rect 191 149 202 183
rect 146 107 202 149
rect 146 73 157 107
rect 191 73 202 107
rect 146 65 202 73
rect 232 221 288 233
rect 232 187 243 221
rect 277 187 288 221
rect 232 111 288 187
rect 232 77 243 111
rect 277 77 288 111
rect 232 65 288 77
rect 318 183 374 233
rect 318 149 329 183
rect 363 149 374 183
rect 318 111 374 149
rect 318 77 329 111
rect 363 77 374 111
rect 318 65 374 77
rect 404 221 460 233
rect 404 187 415 221
rect 449 187 460 221
rect 404 111 460 187
rect 404 77 415 111
rect 449 77 460 111
rect 404 65 460 77
rect 490 225 546 233
rect 490 191 501 225
rect 535 191 546 225
rect 490 157 546 191
rect 490 123 501 157
rect 535 123 546 157
rect 490 65 546 123
rect 576 181 664 233
rect 576 147 603 181
rect 637 147 664 181
rect 576 107 664 147
rect 576 73 603 107
rect 637 73 664 107
rect 576 65 664 73
rect 694 225 750 233
rect 694 191 705 225
rect 739 191 750 225
rect 694 155 750 191
rect 694 121 705 155
rect 739 121 750 155
rect 694 65 750 121
rect 780 221 833 233
rect 780 187 791 221
rect 825 187 833 221
rect 780 111 833 187
rect 780 77 791 111
rect 825 77 833 111
rect 780 65 833 77
<< pdiff >>
rect 33 607 116 619
rect 33 573 59 607
rect 93 573 116 607
rect 33 515 116 573
rect 33 481 59 515
rect 93 481 116 515
rect 33 411 116 481
rect 33 377 59 411
rect 93 377 116 411
rect 33 367 116 377
rect 146 595 202 619
rect 146 561 157 595
rect 191 561 202 595
rect 146 518 202 561
rect 146 484 157 518
rect 191 484 202 518
rect 146 436 202 484
rect 146 402 157 436
rect 191 402 202 436
rect 146 367 202 402
rect 232 607 288 619
rect 232 573 243 607
rect 277 573 288 607
rect 232 496 288 573
rect 232 462 243 496
rect 277 462 288 496
rect 232 367 288 462
rect 318 595 374 619
rect 318 561 329 595
rect 363 561 374 595
rect 318 518 374 561
rect 318 484 329 518
rect 363 484 374 518
rect 318 436 374 484
rect 318 402 329 436
rect 363 402 374 436
rect 318 367 374 402
rect 404 607 460 619
rect 404 573 415 607
rect 449 573 460 607
rect 404 496 460 573
rect 404 462 415 496
rect 449 462 460 496
rect 404 367 460 462
rect 490 595 546 619
rect 490 561 501 595
rect 535 561 546 595
rect 490 518 546 561
rect 490 484 501 518
rect 535 484 546 518
rect 490 436 546 484
rect 490 402 501 436
rect 535 402 546 436
rect 490 367 546 402
rect 576 607 664 619
rect 576 573 600 607
rect 634 573 664 607
rect 576 496 664 573
rect 576 462 600 496
rect 634 462 664 496
rect 576 367 664 462
rect 694 595 750 619
rect 694 561 705 595
rect 739 561 750 595
rect 694 518 750 561
rect 694 484 705 518
rect 739 484 750 518
rect 694 436 750 484
rect 694 402 705 436
rect 739 402 750 436
rect 694 367 750 402
rect 780 607 833 619
rect 780 573 791 607
rect 825 573 833 607
rect 780 507 833 573
rect 780 473 791 507
rect 825 473 833 507
rect 780 413 833 473
rect 780 379 791 413
rect 825 379 833 413
rect 780 367 833 379
<< ndiffc >>
rect 71 187 105 221
rect 71 77 105 111
rect 157 149 191 183
rect 157 73 191 107
rect 243 187 277 221
rect 243 77 277 111
rect 329 149 363 183
rect 329 77 363 111
rect 415 187 449 221
rect 415 77 449 111
rect 501 191 535 225
rect 501 123 535 157
rect 603 147 637 181
rect 603 73 637 107
rect 705 191 739 225
rect 705 121 739 155
rect 791 187 825 221
rect 791 77 825 111
<< pdiffc >>
rect 59 573 93 607
rect 59 481 93 515
rect 59 377 93 411
rect 157 561 191 595
rect 157 484 191 518
rect 157 402 191 436
rect 243 573 277 607
rect 243 462 277 496
rect 329 561 363 595
rect 329 484 363 518
rect 329 402 363 436
rect 415 573 449 607
rect 415 462 449 496
rect 501 561 535 595
rect 501 484 535 518
rect 501 402 535 436
rect 600 573 634 607
rect 600 462 634 496
rect 705 561 739 595
rect 705 484 739 518
rect 705 402 739 436
rect 791 573 825 607
rect 791 473 825 507
rect 791 379 825 413
<< poly >>
rect 116 619 146 645
rect 202 619 232 645
rect 288 619 318 645
rect 374 619 404 645
rect 460 619 490 645
rect 546 619 576 645
rect 664 619 694 645
rect 750 619 780 645
rect 116 335 146 367
rect 202 335 232 367
rect 288 335 318 367
rect 374 335 404 367
rect 116 319 404 335
rect 116 285 143 319
rect 177 285 211 319
rect 245 285 279 319
rect 313 285 347 319
rect 381 285 404 319
rect 116 269 404 285
rect 116 233 146 269
rect 202 233 232 269
rect 288 233 318 269
rect 374 233 404 269
rect 460 335 490 367
rect 546 335 576 367
rect 664 335 694 367
rect 750 335 780 367
rect 460 319 780 335
rect 460 285 601 319
rect 635 285 669 319
rect 703 285 780 319
rect 460 269 780 285
rect 460 233 490 269
rect 546 233 576 269
rect 664 233 694 269
rect 750 233 780 269
rect 116 39 146 65
rect 202 39 232 65
rect 288 39 318 65
rect 374 39 404 65
rect 460 39 490 65
rect 546 39 576 65
rect 664 39 694 65
rect 750 39 780 65
<< polycont >>
rect 143 285 177 319
rect 211 285 245 319
rect 279 285 313 319
rect 347 285 381 319
rect 601 285 635 319
rect 669 285 703 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 25 607 93 649
rect 25 573 59 607
rect 25 515 93 573
rect 25 481 59 515
rect 25 411 93 481
rect 25 377 59 411
rect 127 595 193 611
rect 127 561 157 595
rect 191 561 193 595
rect 127 518 193 561
rect 127 484 157 518
rect 191 484 193 518
rect 127 436 193 484
rect 227 607 293 649
rect 227 573 243 607
rect 277 573 293 607
rect 227 496 293 573
rect 227 462 243 496
rect 277 462 293 496
rect 327 595 365 611
rect 327 561 329 595
rect 363 561 365 595
rect 327 518 365 561
rect 327 484 329 518
rect 363 484 365 518
rect 127 402 157 436
rect 191 428 193 436
rect 327 436 365 484
rect 399 607 465 649
rect 399 573 415 607
rect 449 573 465 607
rect 399 496 465 573
rect 399 462 415 496
rect 449 462 465 496
rect 499 595 550 611
rect 499 561 501 595
rect 535 561 550 595
rect 499 518 550 561
rect 499 484 501 518
rect 535 484 550 518
rect 327 428 329 436
rect 191 402 329 428
rect 363 428 365 436
rect 499 436 550 484
rect 584 607 650 649
rect 584 573 600 607
rect 634 573 650 607
rect 584 496 650 573
rect 584 462 600 496
rect 634 462 650 496
rect 684 595 754 611
rect 684 561 705 595
rect 739 561 754 595
rect 684 518 754 561
rect 684 484 705 518
rect 739 484 754 518
rect 499 428 501 436
rect 363 402 501 428
rect 535 428 550 436
rect 684 436 754 484
rect 684 428 705 436
rect 535 402 705 428
rect 739 402 754 436
rect 127 386 754 402
rect 788 607 841 649
rect 788 573 791 607
rect 825 573 841 607
rect 788 507 841 573
rect 788 473 791 507
rect 825 473 841 507
rect 788 413 841 473
rect 25 361 93 377
rect 127 319 449 352
rect 127 285 143 319
rect 177 285 211 319
rect 245 285 279 319
rect 313 285 347 319
rect 381 285 449 319
rect 57 221 451 251
rect 57 187 71 221
rect 105 217 243 221
rect 105 187 107 217
rect 57 111 107 187
rect 241 187 243 217
rect 277 217 415 221
rect 277 187 279 217
rect 57 77 71 111
rect 105 77 107 111
rect 57 61 107 77
rect 141 149 157 183
rect 191 149 207 183
rect 141 107 207 149
rect 141 73 157 107
rect 191 73 207 107
rect 141 17 207 73
rect 241 111 279 187
rect 413 187 415 217
rect 449 187 451 221
rect 241 77 243 111
rect 277 77 279 111
rect 241 61 279 77
rect 313 149 329 183
rect 363 149 379 183
rect 313 111 379 149
rect 313 77 329 111
rect 363 77 379 111
rect 313 17 379 77
rect 413 111 451 187
rect 485 249 551 386
rect 788 379 791 413
rect 825 379 841 413
rect 788 363 841 379
rect 585 319 754 352
rect 585 285 601 319
rect 635 285 669 319
rect 703 285 754 319
rect 585 283 754 285
rect 485 225 755 249
rect 485 191 501 225
rect 535 215 705 225
rect 535 191 551 215
rect 485 157 551 191
rect 687 191 705 215
rect 739 191 755 225
rect 485 123 501 157
rect 535 123 551 157
rect 587 147 603 181
rect 637 147 653 181
rect 413 77 415 111
rect 449 87 451 111
rect 587 107 653 147
rect 687 155 755 191
rect 687 121 705 155
rect 739 121 755 155
rect 789 221 841 237
rect 789 187 791 221
rect 825 187 841 221
rect 587 87 603 107
rect 449 77 603 87
rect 413 73 603 77
rect 637 87 653 107
rect 789 111 841 187
rect 789 87 791 111
rect 637 77 791 87
rect 825 77 841 111
rect 637 73 841 77
rect 413 53 841 73
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2_4
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5780140
string GDS_START 5771496
<< end >>
