magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4082 1975
<< nwell >>
rect -38 331 2822 704
rect 2224 291 2441 331
<< pwell >>
rect 1695 229 1809 282
rect 649 222 1809 229
rect 649 191 1941 222
rect 296 185 1941 191
rect 1 178 1941 185
rect 1 157 2289 178
rect 2482 157 2756 269
rect 1 49 2756 157
rect 0 0 2784 49
<< scnmos >>
rect 80 75 110 159
rect 270 75 300 159
rect 372 81 402 165
rect 458 81 488 165
rect 530 81 560 165
rect 630 81 660 165
rect 810 119 840 203
rect 896 119 926 203
rect 1006 119 1036 203
rect 1092 119 1122 203
rect 1314 119 1344 203
rect 1400 119 1430 203
rect 1472 119 1502 203
rect 1544 119 1574 203
rect 1676 68 1706 196
rect 1820 68 1850 196
rect 1930 68 1960 152
rect 2002 68 2032 152
rect 2108 68 2138 152
rect 2180 68 2210 152
rect 2370 47 2400 131
rect 2561 75 2591 243
rect 2647 75 2677 243
<< scpmoshvt >>
rect 179 491 209 619
rect 265 491 295 619
rect 337 491 367 619
rect 423 491 453 619
rect 522 491 552 619
rect 630 491 660 619
rect 908 367 938 619
rect 994 367 1024 619
rect 1216 463 1246 547
rect 1302 463 1332 547
rect 1374 463 1404 547
rect 1506 463 1536 547
rect 1696 379 1726 547
rect 1782 379 1812 547
rect 1923 496 1953 580
rect 2034 496 2064 580
rect 2129 509 2159 593
rect 2215 509 2245 593
rect 2322 327 2352 455
rect 2555 367 2585 619
rect 2641 367 2671 619
<< ndiff >>
rect 675 165 810 203
rect 322 159 372 165
rect 27 147 80 159
rect 27 113 35 147
rect 69 113 80 147
rect 27 75 80 113
rect 110 121 163 159
rect 110 87 121 121
rect 155 87 163 121
rect 110 75 163 87
rect 217 131 270 159
rect 217 97 225 131
rect 259 97 270 131
rect 217 75 270 97
rect 300 81 372 159
rect 402 157 458 165
rect 402 123 413 157
rect 447 123 458 157
rect 402 81 458 123
rect 488 81 530 165
rect 560 125 630 165
rect 560 91 571 125
rect 605 91 630 125
rect 560 81 630 91
rect 660 129 810 165
rect 660 95 671 129
rect 705 119 810 129
rect 840 190 896 203
rect 840 156 851 190
rect 885 156 896 190
rect 840 119 896 156
rect 926 138 1006 203
rect 926 119 949 138
rect 705 95 795 119
rect 660 81 795 95
rect 941 104 949 119
rect 983 119 1006 138
rect 1036 186 1092 203
rect 1036 152 1047 186
rect 1081 152 1092 186
rect 1036 119 1092 152
rect 1122 176 1181 203
rect 1122 142 1133 176
rect 1167 142 1181 176
rect 1122 119 1181 142
rect 1261 190 1314 203
rect 1261 156 1269 190
rect 1303 156 1314 190
rect 1261 119 1314 156
rect 1344 180 1400 203
rect 1344 146 1355 180
rect 1389 146 1400 180
rect 1344 119 1400 146
rect 1430 119 1472 203
rect 1502 119 1544 203
rect 1574 196 1661 203
rect 1721 246 1783 256
rect 1721 212 1733 246
rect 1767 212 1783 246
rect 1721 196 1783 212
rect 1574 119 1676 196
rect 983 104 991 119
rect 941 88 991 104
rect 300 75 350 81
rect 1589 110 1676 119
rect 1589 76 1606 110
rect 1640 76 1676 110
rect 1589 68 1676 76
rect 1706 68 1820 196
rect 1850 152 1915 196
rect 2508 231 2561 243
rect 2508 197 2516 231
rect 2550 197 2561 231
rect 1850 124 1930 152
rect 1850 90 1885 124
rect 1919 90 1930 124
rect 1850 68 1930 90
rect 1960 68 2002 152
rect 2032 118 2108 152
rect 2032 84 2043 118
rect 2077 84 2108 118
rect 2032 68 2108 84
rect 2138 68 2180 152
rect 2210 140 2263 152
rect 2210 106 2221 140
rect 2255 106 2263 140
rect 2210 68 2263 106
rect 2317 105 2370 131
rect 2317 71 2325 105
rect 2359 71 2370 105
rect 2317 47 2370 71
rect 2400 106 2453 131
rect 2400 72 2411 106
rect 2445 72 2453 106
rect 2508 121 2561 197
rect 2508 87 2516 121
rect 2550 87 2561 121
rect 2508 75 2561 87
rect 2591 219 2647 243
rect 2591 185 2602 219
rect 2636 185 2647 219
rect 2591 117 2647 185
rect 2591 83 2602 117
rect 2636 83 2647 117
rect 2591 75 2647 83
rect 2677 219 2730 243
rect 2677 185 2688 219
rect 2722 185 2730 219
rect 2677 121 2730 185
rect 2677 87 2688 121
rect 2722 87 2730 121
rect 2677 75 2730 87
rect 2400 47 2453 72
<< pdiff >>
rect 126 607 179 619
rect 126 573 134 607
rect 168 573 179 607
rect 126 537 179 573
rect 126 503 134 537
rect 168 503 179 537
rect 126 491 179 503
rect 209 611 265 619
rect 209 577 220 611
rect 254 577 265 611
rect 209 537 265 577
rect 209 503 220 537
rect 254 503 265 537
rect 209 491 265 503
rect 295 491 337 619
rect 367 607 423 619
rect 367 573 378 607
rect 412 573 423 607
rect 367 537 423 573
rect 367 503 378 537
rect 412 503 423 537
rect 367 491 423 503
rect 453 491 522 619
rect 552 596 630 619
rect 552 562 571 596
rect 605 562 630 596
rect 552 491 630 562
rect 660 607 713 619
rect 660 573 671 607
rect 705 573 713 607
rect 660 537 713 573
rect 660 503 671 537
rect 705 503 713 537
rect 660 491 713 503
rect 855 433 908 619
rect 855 399 863 433
rect 897 399 908 433
rect 855 367 908 399
rect 938 596 994 619
rect 938 562 949 596
rect 983 562 994 596
rect 938 367 994 562
rect 1024 427 1077 619
rect 1024 393 1035 427
rect 1069 393 1077 427
rect 1024 367 1077 393
rect 1419 575 1477 583
rect 1419 547 1431 575
rect 1147 521 1216 547
rect 1147 487 1171 521
rect 1205 487 1216 521
rect 1147 463 1216 487
rect 1246 536 1302 547
rect 1246 502 1257 536
rect 1291 502 1302 536
rect 1246 463 1302 502
rect 1332 463 1374 547
rect 1404 541 1431 547
rect 1465 547 1477 575
rect 2079 580 2129 593
rect 1832 549 1923 580
rect 1832 547 1854 549
rect 1465 541 1506 547
rect 1404 463 1506 541
rect 1536 521 1589 547
rect 1536 487 1547 521
rect 1581 487 1589 521
rect 1536 463 1589 487
rect 1643 535 1696 547
rect 1643 501 1651 535
rect 1685 501 1696 535
rect 1643 425 1696 501
rect 1643 391 1651 425
rect 1685 391 1696 425
rect 1643 379 1696 391
rect 1726 535 1782 547
rect 1726 501 1737 535
rect 1771 501 1782 535
rect 1726 425 1782 501
rect 1726 391 1737 425
rect 1771 391 1782 425
rect 1726 379 1782 391
rect 1812 515 1854 547
rect 1888 515 1923 549
rect 1812 496 1923 515
rect 1953 496 2034 580
rect 2064 559 2129 580
rect 2064 525 2079 559
rect 2113 525 2129 559
rect 2064 509 2129 525
rect 2159 568 2215 593
rect 2159 534 2170 568
rect 2204 534 2215 568
rect 2159 509 2215 534
rect 2245 577 2305 593
rect 2245 543 2263 577
rect 2297 543 2305 577
rect 2245 509 2305 543
rect 2064 496 2114 509
rect 1812 379 1862 496
rect 2260 443 2322 455
rect 2260 409 2277 443
rect 2311 409 2322 443
rect 2260 327 2322 409
rect 2352 441 2405 455
rect 2352 407 2363 441
rect 2397 407 2405 441
rect 2352 373 2405 407
rect 2352 339 2363 373
rect 2397 339 2405 373
rect 2502 441 2555 619
rect 2502 407 2510 441
rect 2544 407 2555 441
rect 2502 367 2555 407
rect 2585 601 2641 619
rect 2585 567 2596 601
rect 2630 567 2641 601
rect 2585 367 2641 567
rect 2671 599 2724 619
rect 2671 565 2682 599
rect 2716 565 2724 599
rect 2671 510 2724 565
rect 2671 476 2682 510
rect 2716 476 2724 510
rect 2671 421 2724 476
rect 2671 387 2682 421
rect 2716 387 2724 421
rect 2671 367 2724 387
rect 2352 327 2405 339
<< ndiffc >>
rect 35 113 69 147
rect 121 87 155 121
rect 225 97 259 131
rect 413 123 447 157
rect 571 91 605 125
rect 671 95 705 129
rect 851 156 885 190
rect 949 104 983 138
rect 1047 152 1081 186
rect 1133 142 1167 176
rect 1269 156 1303 190
rect 1355 146 1389 180
rect 1733 212 1767 246
rect 1606 76 1640 110
rect 2516 197 2550 231
rect 1885 90 1919 124
rect 2043 84 2077 118
rect 2221 106 2255 140
rect 2325 71 2359 105
rect 2411 72 2445 106
rect 2516 87 2550 121
rect 2602 185 2636 219
rect 2602 83 2636 117
rect 2688 185 2722 219
rect 2688 87 2722 121
<< pdiffc >>
rect 134 573 168 607
rect 134 503 168 537
rect 220 577 254 611
rect 220 503 254 537
rect 378 573 412 607
rect 378 503 412 537
rect 571 562 605 596
rect 671 573 705 607
rect 671 503 705 537
rect 863 399 897 433
rect 949 562 983 596
rect 1035 393 1069 427
rect 1171 487 1205 521
rect 1257 502 1291 536
rect 1431 541 1465 575
rect 1547 487 1581 521
rect 1651 501 1685 535
rect 1651 391 1685 425
rect 1737 501 1771 535
rect 1737 391 1771 425
rect 1854 515 1888 549
rect 2079 525 2113 559
rect 2170 534 2204 568
rect 2263 543 2297 577
rect 2277 409 2311 443
rect 2363 407 2397 441
rect 2363 339 2397 373
rect 2510 407 2544 441
rect 2596 567 2630 601
rect 2682 565 2716 599
rect 2682 476 2716 510
rect 2682 387 2716 421
<< poly >>
rect 179 619 209 645
rect 265 619 295 645
rect 337 619 367 645
rect 423 619 453 645
rect 522 619 552 645
rect 630 619 660 645
rect 908 619 938 645
rect 994 619 1024 645
rect 179 469 209 491
rect 265 469 295 491
rect 179 439 295 469
rect 179 373 209 439
rect 80 357 247 373
rect 80 323 127 357
rect 161 323 197 357
rect 231 323 247 357
rect 80 307 247 323
rect 337 319 367 491
rect 423 459 453 491
rect 409 443 475 459
rect 409 409 425 443
rect 459 409 475 443
rect 409 393 475 409
rect 522 424 552 491
rect 630 456 660 491
rect 630 440 728 456
rect 522 408 588 424
rect 522 374 538 408
rect 572 374 588 408
rect 414 329 480 345
rect 80 159 110 307
rect 295 303 372 319
rect 295 269 311 303
rect 345 269 372 303
rect 414 295 430 329
rect 464 295 480 329
rect 414 279 480 295
rect 522 340 588 374
rect 522 306 538 340
rect 572 306 588 340
rect 522 290 588 306
rect 630 406 678 440
rect 712 406 728 440
rect 630 390 728 406
rect 295 253 372 269
rect 181 231 247 247
rect 181 197 197 231
rect 231 211 247 231
rect 342 231 372 253
rect 450 242 480 279
rect 231 197 300 211
rect 342 201 402 231
rect 450 212 488 242
rect 181 181 300 197
rect 270 159 300 181
rect 372 165 402 201
rect 458 165 488 212
rect 530 165 560 290
rect 630 165 660 390
rect 1092 615 1812 645
rect 908 308 938 367
rect 994 335 1024 367
rect 1092 335 1122 615
rect 1216 547 1246 573
rect 1302 547 1332 615
rect 1374 547 1404 573
rect 1506 547 1536 573
rect 1696 547 1726 573
rect 1782 547 1812 615
rect 1923 580 1953 606
rect 2034 580 2064 606
rect 2129 593 2159 619
rect 2215 615 2460 645
rect 2555 619 2585 645
rect 2641 619 2671 645
rect 2215 593 2245 615
rect 2394 605 2460 615
rect 1216 394 1246 463
rect 1302 437 1332 463
rect 810 292 938 308
rect 810 258 859 292
rect 893 258 938 292
rect 810 242 938 258
rect 980 319 1122 335
rect 980 285 996 319
rect 1030 285 1122 319
rect 1164 378 1246 394
rect 1164 344 1180 378
rect 1214 344 1246 378
rect 1374 431 1404 463
rect 1506 448 1536 463
rect 1374 415 1464 431
rect 1506 429 1611 448
rect 1510 426 1611 429
rect 1515 422 1611 426
rect 1519 418 1611 422
rect 1374 381 1413 415
rect 1447 398 1464 415
rect 1544 415 1611 418
rect 1447 392 1472 398
rect 1447 383 1484 392
rect 1447 381 1495 383
rect 1374 379 1495 381
rect 1544 381 1561 415
rect 1595 381 1611 415
rect 1374 362 1502 379
rect 1446 360 1502 362
rect 1457 353 1502 360
rect 1463 347 1502 353
rect 1164 320 1246 344
rect 1468 339 1502 347
rect 1164 290 1430 320
rect 980 252 1122 285
rect 810 203 840 242
rect 896 203 926 242
rect 1006 203 1036 252
rect 1092 248 1122 252
rect 1092 218 1344 248
rect 1092 203 1122 218
rect 1314 203 1344 218
rect 1400 203 1430 290
rect 1472 203 1502 339
rect 1544 364 1611 381
rect 2394 571 2410 605
rect 2444 571 2460 605
rect 2394 537 2460 571
rect 1923 464 1953 496
rect 1892 448 1960 464
rect 1892 414 1910 448
rect 1944 414 1960 448
rect 1892 398 1960 414
rect 1544 203 1574 364
rect 1696 344 1726 379
rect 1649 328 1726 344
rect 1649 294 1665 328
rect 1699 294 1726 328
rect 1782 356 1812 379
rect 1782 326 1960 356
rect 1649 278 1726 294
rect 810 93 840 119
rect 896 93 926 119
rect 1676 196 1706 278
rect 1820 268 1886 284
rect 1820 234 1836 268
rect 1870 234 1886 268
rect 1820 218 1886 234
rect 1820 196 1850 218
rect 1006 93 1036 119
rect 1092 93 1122 119
rect 1314 93 1344 119
rect 1400 93 1430 119
rect 1472 93 1502 119
rect 80 49 110 75
rect 270 49 300 75
rect 372 55 402 81
rect 458 55 488 81
rect 530 55 560 81
rect 630 51 660 81
rect 1544 51 1574 119
rect 1930 152 1960 326
rect 2034 283 2064 496
rect 2129 440 2159 509
rect 2107 424 2173 440
rect 2107 390 2123 424
rect 2157 390 2173 424
rect 2107 374 2173 390
rect 2108 304 2140 374
rect 2002 267 2068 283
rect 2002 233 2018 267
rect 2052 233 2068 267
rect 2002 217 2068 233
rect 2002 152 2032 217
rect 2110 204 2140 304
rect 2215 295 2245 509
rect 2394 503 2410 537
rect 2444 503 2460 537
rect 2394 487 2460 503
rect 2322 455 2352 481
rect 2108 193 2140 204
rect 2182 279 2252 295
rect 2182 245 2202 279
rect 2236 259 2252 279
rect 2322 259 2352 327
rect 2555 295 2585 367
rect 2641 335 2671 367
rect 2633 319 2699 335
rect 2236 245 2352 259
rect 2182 229 2352 245
rect 2399 279 2591 295
rect 2399 245 2415 279
rect 2449 265 2591 279
rect 2633 285 2649 319
rect 2683 285 2699 319
rect 2633 269 2699 285
rect 2449 245 2465 265
rect 2399 229 2465 245
rect 2561 243 2591 265
rect 2647 243 2677 269
rect 2108 152 2138 193
rect 2182 180 2212 229
rect 2180 167 2212 180
rect 2313 183 2352 229
rect 2180 152 2210 167
rect 2313 153 2400 183
rect 2370 131 2400 153
rect 630 21 1574 51
rect 1676 42 1706 68
rect 1820 42 1850 68
rect 1930 42 1960 68
rect 2002 42 2032 68
rect 2108 42 2138 68
rect 2180 42 2210 68
rect 2561 49 2591 75
rect 2647 49 2677 75
rect 2370 21 2400 47
<< polycont >>
rect 127 323 161 357
rect 197 323 231 357
rect 425 409 459 443
rect 538 374 572 408
rect 311 269 345 303
rect 430 295 464 329
rect 538 306 572 340
rect 678 406 712 440
rect 197 197 231 231
rect 859 258 893 292
rect 996 285 1030 319
rect 1180 344 1214 378
rect 1413 381 1447 415
rect 1561 381 1595 415
rect 2410 571 2444 605
rect 1910 414 1944 448
rect 1665 294 1699 328
rect 1836 234 1870 268
rect 2123 390 2157 424
rect 2018 233 2052 267
rect 2410 503 2444 537
rect 2202 245 2236 279
rect 2415 245 2449 279
rect 2649 285 2683 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 118 607 184 615
rect 118 573 134 607
rect 168 573 184 607
rect 118 537 184 573
rect 118 503 134 537
rect 168 503 184 537
rect 118 443 184 503
rect 218 611 270 649
rect 218 577 220 611
rect 254 577 270 611
rect 218 537 270 577
rect 218 503 220 537
rect 254 503 270 537
rect 218 487 270 503
rect 362 607 428 615
rect 362 573 378 607
rect 412 573 428 607
rect 362 537 428 573
rect 555 596 621 649
rect 555 562 571 596
rect 605 562 621 596
rect 555 558 621 562
rect 655 607 721 615
rect 655 573 671 607
rect 705 573 721 607
rect 362 503 378 537
rect 412 524 428 537
rect 655 537 721 573
rect 933 596 999 649
rect 933 562 949 596
rect 983 562 999 596
rect 933 558 999 562
rect 1415 575 1481 649
rect 655 524 671 537
rect 412 503 671 524
rect 705 524 721 537
rect 1155 524 1207 537
rect 705 521 1207 524
rect 705 503 1171 521
rect 362 490 1171 503
rect 362 483 655 490
rect 1155 487 1171 490
rect 1205 487 1207 521
rect 1241 536 1381 555
rect 1415 541 1431 575
rect 1465 541 1481 575
rect 1415 539 1481 541
rect 1241 502 1257 536
rect 1291 505 1381 536
rect 1517 521 1598 537
rect 1517 505 1547 521
rect 1291 502 1547 505
rect 1241 499 1547 502
rect 362 477 642 483
rect 31 409 425 443
rect 459 409 475 443
rect 31 407 475 409
rect 511 408 572 443
rect 31 247 65 407
rect 511 374 538 408
rect 111 357 477 373
rect 111 323 127 357
rect 161 323 197 357
rect 231 339 477 357
rect 231 323 261 339
rect 111 307 261 323
rect 414 329 477 339
rect 295 303 361 305
rect 295 269 311 303
rect 345 269 361 303
rect 414 295 430 329
rect 464 295 477 329
rect 414 279 477 295
rect 511 340 572 374
rect 511 306 538 340
rect 31 231 247 247
rect 31 197 197 231
rect 231 197 247 231
rect 31 181 247 197
rect 31 147 73 181
rect 295 156 361 269
rect 511 231 572 306
rect 608 197 642 477
rect 1155 465 1207 487
rect 1345 487 1547 499
rect 1581 487 1598 521
rect 1345 467 1598 487
rect 1650 535 1696 649
rect 1650 501 1651 535
rect 1685 501 1696 535
rect 676 440 750 456
rect 676 406 678 440
rect 712 424 750 440
rect 676 390 703 406
rect 737 390 750 424
rect 847 433 999 443
rect 847 399 863 433
rect 897 399 999 433
rect 847 390 999 399
rect 682 292 929 356
rect 682 258 859 292
rect 893 258 929 292
rect 682 240 929 258
rect 965 343 999 390
rect 1033 427 1096 443
rect 1155 431 1303 465
rect 1033 393 1035 427
rect 1069 394 1096 427
rect 1069 393 1235 394
rect 1033 378 1235 393
rect 1033 377 1180 378
rect 1064 348 1180 377
rect 1080 344 1180 348
rect 1214 344 1235 378
rect 965 319 1030 343
rect 965 285 996 319
rect 1030 285 1046 319
rect 965 269 1030 285
rect 965 206 999 269
rect 1080 259 1235 344
rect 1069 247 1235 259
rect 1058 235 1235 247
rect 397 163 642 197
rect 851 190 999 206
rect 397 157 463 163
rect 31 113 35 147
rect 69 113 73 147
rect 31 97 73 113
rect 117 121 159 137
rect 117 87 121 121
rect 155 87 159 121
rect 117 17 159 87
rect 209 131 261 147
rect 209 97 225 131
rect 259 97 261 131
rect 397 123 413 157
rect 447 123 463 157
rect 885 172 999 190
rect 1037 226 1235 235
rect 1037 217 1107 226
rect 1037 186 1097 217
rect 851 134 885 156
rect 1037 152 1047 186
rect 1081 152 1097 186
rect 655 129 721 131
rect 397 119 463 123
rect 555 125 621 129
rect 209 85 261 97
rect 555 91 571 125
rect 605 91 621 125
rect 555 85 621 91
rect 209 51 621 85
rect 655 95 671 129
rect 705 95 721 129
rect 655 17 721 95
rect 933 104 949 138
rect 983 104 999 138
rect 1037 136 1097 152
rect 1131 176 1167 192
rect 1131 142 1133 176
rect 933 17 999 104
rect 1131 17 1167 142
rect 1201 85 1235 226
rect 1269 190 1303 431
rect 1269 140 1303 156
rect 1345 196 1379 467
rect 1413 415 1449 431
rect 1447 381 1449 415
rect 1413 259 1449 381
rect 1485 330 1521 467
rect 1555 424 1616 433
rect 1555 415 1567 424
rect 1555 381 1561 415
rect 1601 390 1616 424
rect 1595 381 1616 390
rect 1555 364 1616 381
rect 1650 425 1696 501
rect 1650 391 1651 425
rect 1685 391 1696 425
rect 1650 375 1696 391
rect 1732 535 1783 584
rect 1732 501 1737 535
rect 1771 501 1783 535
rect 1732 425 1783 501
rect 1838 549 2012 584
rect 1838 515 1854 549
rect 1888 515 2012 549
rect 1838 499 2012 515
rect 2070 559 2122 649
rect 2070 525 2079 559
rect 2113 525 2122 559
rect 2070 509 2122 525
rect 2158 568 2227 584
rect 2158 534 2170 568
rect 2204 534 2227 568
rect 1908 452 1944 464
rect 1732 391 1737 425
rect 1771 391 1783 425
rect 1732 375 1783 391
rect 1485 328 1715 330
rect 1485 294 1665 328
rect 1699 294 1715 328
rect 1485 293 1715 294
rect 1749 259 1783 375
rect 1413 246 1783 259
rect 1413 222 1733 246
rect 1421 212 1733 222
rect 1767 212 1783 246
rect 1817 448 1944 452
rect 1817 414 1910 448
rect 1817 390 1944 414
rect 1817 268 1870 390
rect 1978 345 2012 499
rect 2158 474 2227 534
rect 2046 424 2159 440
rect 2046 390 2047 424
rect 2081 390 2123 424
rect 2157 390 2159 424
rect 2046 374 2159 390
rect 1817 234 1836 268
rect 1817 218 1870 234
rect 1910 337 2012 345
rect 2193 371 2227 474
rect 2261 577 2327 649
rect 2261 543 2263 577
rect 2297 543 2327 577
rect 2261 443 2327 543
rect 2394 605 2460 615
rect 2394 571 2410 605
rect 2444 571 2460 605
rect 2394 537 2460 571
rect 2580 601 2646 649
rect 2580 567 2596 601
rect 2630 567 2646 601
rect 2580 559 2646 567
rect 2680 599 2753 615
rect 2680 565 2682 599
rect 2716 565 2753 599
rect 2394 503 2410 537
rect 2444 525 2460 537
rect 2444 503 2646 525
rect 2394 491 2646 503
rect 2261 409 2277 443
rect 2311 409 2327 443
rect 2261 405 2327 409
rect 2361 441 2461 457
rect 2361 407 2363 441
rect 2397 407 2461 441
rect 2361 373 2461 407
rect 2193 337 2318 371
rect 1910 303 2136 337
rect 1345 180 1389 196
rect 1345 146 1355 180
rect 1817 178 1851 218
rect 1910 187 1966 303
rect 2102 279 2238 303
rect 2102 269 2202 279
rect 2000 267 2068 269
rect 2000 233 2018 267
rect 2052 233 2068 267
rect 2195 245 2202 269
rect 2236 245 2238 279
rect 2000 199 2161 233
rect 2195 229 2238 245
rect 1345 130 1389 146
rect 1522 144 1851 178
rect 1522 85 1556 144
rect 1885 124 1966 187
rect 2127 195 2161 199
rect 2272 195 2318 337
rect 2361 339 2363 373
rect 2397 339 2461 373
rect 2361 323 2461 339
rect 2127 145 2318 195
rect 2409 279 2461 323
rect 2409 245 2415 279
rect 2449 245 2461 279
rect 1201 51 1556 85
rect 1590 76 1606 110
rect 1640 76 1656 110
rect 1590 17 1656 76
rect 1919 90 1966 124
rect 2205 140 2271 145
rect 1885 66 1966 90
rect 2027 118 2093 122
rect 2027 84 2043 118
rect 2077 84 2093 118
rect 2205 106 2221 140
rect 2255 106 2271 140
rect 2205 102 2271 106
rect 2309 105 2375 111
rect 2027 17 2093 84
rect 2309 71 2325 105
rect 2359 71 2375 105
rect 2309 17 2375 71
rect 2409 106 2461 245
rect 2409 72 2411 106
rect 2445 72 2461 106
rect 2409 56 2461 72
rect 2495 441 2564 457
rect 2495 407 2510 441
rect 2544 407 2564 441
rect 2495 231 2564 407
rect 2608 335 2646 491
rect 2680 510 2753 565
rect 2680 476 2682 510
rect 2716 476 2753 510
rect 2680 421 2753 476
rect 2680 387 2682 421
rect 2716 387 2753 421
rect 2680 371 2753 387
rect 2608 319 2683 335
rect 2608 285 2649 319
rect 2608 269 2683 285
rect 2717 235 2753 371
rect 2495 197 2516 231
rect 2550 197 2564 231
rect 2495 121 2564 197
rect 2495 87 2516 121
rect 2550 87 2564 121
rect 2495 71 2564 87
rect 2598 219 2645 235
rect 2598 185 2602 219
rect 2636 185 2645 219
rect 2598 117 2645 185
rect 2598 83 2602 117
rect 2636 83 2645 117
rect 2598 17 2645 83
rect 2679 219 2753 235
rect 2679 185 2688 219
rect 2722 185 2753 219
rect 2679 121 2753 185
rect 2679 87 2688 121
rect 2722 87 2753 121
rect 2679 71 2753 87
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 703 406 712 424
rect 712 406 737 424
rect 703 390 737 406
rect 1567 415 1601 424
rect 1567 390 1595 415
rect 1595 390 1601 415
rect 2047 390 2081 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 691 424 749 430
rect 691 390 703 424
rect 737 421 749 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 737 393 1567 421
rect 737 390 749 393
rect 691 384 749 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2035 424 2093 430
rect 2035 421 2047 424
rect 1601 393 2047 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2035 390 2047 393
rect 2081 390 2093 424
rect 2035 384 2093 390
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfrbp_1
flabel comment s 1477 630 1477 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1106 36 1106 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 2230 418 2230 418 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 2047 390 2081 424 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2527 94 2561 128 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2527 168 2561 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2527 242 2561 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2527 316 2561 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2527 390 2561 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2719 242 2753 276 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2719 316 2753 350 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2719 390 2753 424 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2719 464 2753 498 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2719 538 2753 572 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry R90
string GDS_END 6455802
string GDS_START 6432598
<< end >>
