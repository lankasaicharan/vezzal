magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 860 263 1179 279
rect 328 247 1179 263
rect 1 226 1179 247
rect 1 49 1627 226
rect 0 0 1632 49
<< scnmos >>
rect 83 53 113 221
rect 214 137 244 221
rect 410 109 440 237
rect 510 109 540 237
rect 745 69 775 237
rect 966 125 996 253
rect 1066 125 1096 253
rect 1175 116 1205 200
rect 1293 72 1323 200
rect 1384 72 1414 200
rect 1514 72 1544 200
<< scpmoshvt >>
rect 81 367 111 619
rect 217 367 247 495
rect 410 451 440 619
rect 519 409 549 577
rect 724 367 754 619
rect 951 373 981 541
rect 1060 373 1090 501
rect 1146 373 1176 501
rect 1275 373 1305 541
rect 1407 383 1437 583
rect 1514 383 1544 583
<< ndiff >>
rect 354 225 410 237
rect 27 209 83 221
rect 27 175 38 209
rect 72 175 83 209
rect 27 101 83 175
rect 27 67 38 101
rect 72 67 83 101
rect 27 53 83 67
rect 113 137 214 221
rect 244 209 300 221
rect 244 175 255 209
rect 289 175 300 209
rect 244 137 300 175
rect 354 191 365 225
rect 399 191 410 225
rect 113 73 192 137
rect 354 109 410 191
rect 440 170 510 237
rect 440 136 465 170
rect 499 136 510 170
rect 440 109 510 136
rect 540 170 611 237
rect 540 136 565 170
rect 599 136 611 170
rect 540 109 611 136
rect 665 89 745 237
rect 113 53 146 73
rect 135 39 146 53
rect 180 39 192 73
rect 665 55 677 89
rect 711 69 745 89
rect 775 225 832 237
rect 775 191 786 225
rect 820 191 832 225
rect 775 69 832 191
rect 886 125 966 253
rect 996 225 1066 253
rect 996 191 1007 225
rect 1041 191 1066 225
rect 996 125 1066 191
rect 1096 239 1153 253
rect 1096 205 1107 239
rect 1141 205 1153 239
rect 1096 200 1153 205
rect 1096 125 1175 200
rect 886 89 944 125
rect 711 55 723 69
rect 665 43 723 55
rect 886 55 898 89
rect 932 55 944 89
rect 886 43 944 55
rect 1125 116 1175 125
rect 1205 170 1293 200
rect 1205 136 1239 170
rect 1273 136 1293 170
rect 1205 116 1293 136
rect 1227 72 1293 116
rect 1323 186 1384 200
rect 1323 152 1339 186
rect 1373 152 1384 186
rect 1323 118 1384 152
rect 1323 84 1339 118
rect 1373 84 1384 118
rect 1323 72 1384 84
rect 1414 118 1514 200
rect 1414 84 1439 118
rect 1473 84 1514 118
rect 1414 72 1514 84
rect 1544 188 1601 200
rect 1544 154 1555 188
rect 1589 154 1601 188
rect 1544 118 1601 154
rect 1544 84 1555 118
rect 1589 84 1601 118
rect 1544 72 1601 84
rect 135 27 192 39
<< pdiff >>
rect 27 599 81 619
rect 27 565 36 599
rect 70 565 81 599
rect 27 506 81 565
rect 27 472 36 506
rect 70 472 81 506
rect 27 413 81 472
rect 27 379 36 413
rect 70 379 81 413
rect 27 367 81 379
rect 111 607 168 619
rect 111 573 122 607
rect 156 573 168 607
rect 111 508 168 573
rect 111 474 122 508
rect 156 495 168 508
rect 355 510 410 619
rect 156 474 217 495
rect 111 367 217 474
rect 247 461 301 495
rect 247 427 258 461
rect 292 427 301 461
rect 355 476 365 510
rect 399 476 410 510
rect 355 451 410 476
rect 440 607 497 619
rect 440 573 451 607
rect 485 577 497 607
rect 667 607 724 619
rect 485 573 519 577
rect 440 451 519 573
rect 247 367 301 427
rect 469 409 519 451
rect 549 455 613 577
rect 549 421 567 455
rect 601 421 613 455
rect 549 409 613 421
rect 667 573 679 607
rect 713 573 724 607
rect 667 367 724 573
rect 754 424 811 619
rect 754 390 765 424
rect 799 390 811 424
rect 754 367 811 390
rect 871 576 929 588
rect 871 542 883 576
rect 917 542 929 576
rect 871 541 929 542
rect 871 373 951 541
rect 981 529 1038 541
rect 981 495 992 529
rect 1026 501 1038 529
rect 1327 571 1407 583
rect 1327 541 1339 571
rect 1225 501 1275 541
rect 1026 495 1060 501
rect 981 425 1060 495
rect 981 391 992 425
rect 1026 391 1060 425
rect 981 373 1060 391
rect 1090 489 1146 501
rect 1090 455 1101 489
rect 1135 455 1146 489
rect 1090 419 1146 455
rect 1090 385 1101 419
rect 1135 385 1146 419
rect 1090 373 1146 385
rect 1176 436 1275 501
rect 1176 402 1187 436
rect 1221 402 1275 436
rect 1176 373 1275 402
rect 1305 537 1339 541
rect 1373 537 1407 571
rect 1305 503 1407 537
rect 1305 469 1339 503
rect 1373 469 1407 503
rect 1305 419 1407 469
rect 1305 385 1339 419
rect 1373 385 1407 419
rect 1305 383 1407 385
rect 1437 571 1514 583
rect 1437 537 1448 571
rect 1482 537 1514 571
rect 1437 503 1514 537
rect 1437 469 1448 503
rect 1482 469 1514 503
rect 1437 383 1514 469
rect 1544 571 1601 583
rect 1544 537 1555 571
rect 1589 537 1601 571
rect 1544 500 1601 537
rect 1544 466 1555 500
rect 1589 466 1601 500
rect 1544 429 1601 466
rect 1544 395 1555 429
rect 1589 395 1601 429
rect 1544 383 1601 395
rect 1305 373 1385 383
<< ndiffc >>
rect 38 175 72 209
rect 38 67 72 101
rect 255 175 289 209
rect 365 191 399 225
rect 465 136 499 170
rect 565 136 599 170
rect 146 39 180 73
rect 677 55 711 89
rect 786 191 820 225
rect 1007 191 1041 225
rect 1107 205 1141 239
rect 898 55 932 89
rect 1239 136 1273 170
rect 1339 152 1373 186
rect 1339 84 1373 118
rect 1439 84 1473 118
rect 1555 154 1589 188
rect 1555 84 1589 118
<< pdiffc >>
rect 36 565 70 599
rect 36 472 70 506
rect 36 379 70 413
rect 122 573 156 607
rect 122 474 156 508
rect 258 427 292 461
rect 365 476 399 510
rect 451 573 485 607
rect 567 421 601 455
rect 679 573 713 607
rect 765 390 799 424
rect 883 542 917 576
rect 992 495 1026 529
rect 992 391 1026 425
rect 1101 455 1135 489
rect 1101 385 1135 419
rect 1187 402 1221 436
rect 1339 537 1373 571
rect 1339 469 1373 503
rect 1339 385 1373 419
rect 1448 537 1482 571
rect 1448 469 1482 503
rect 1555 537 1589 571
rect 1555 466 1589 500
rect 1555 395 1589 429
<< poly >>
rect 81 619 111 645
rect 410 619 440 645
rect 724 619 754 645
rect 217 495 247 521
rect 519 577 549 603
rect 81 325 111 367
rect 217 335 247 367
rect 81 309 147 325
rect 81 275 97 309
rect 131 275 147 309
rect 81 259 147 275
rect 205 319 271 335
rect 205 285 221 319
rect 255 299 271 319
rect 410 299 440 451
rect 519 377 549 409
rect 482 361 549 377
rect 826 615 1305 645
rect 482 327 498 361
rect 532 327 549 361
rect 724 335 754 367
rect 826 335 856 615
rect 951 541 981 567
rect 1060 501 1090 615
rect 1275 541 1305 615
rect 1407 583 1437 609
rect 1514 583 1544 609
rect 1146 501 1176 527
rect 951 341 981 373
rect 482 311 549 327
rect 703 319 856 335
rect 255 285 440 299
rect 205 269 440 285
rect 83 221 113 259
rect 214 221 244 269
rect 410 237 440 269
rect 510 237 540 311
rect 703 285 719 319
rect 753 305 856 319
rect 898 325 981 341
rect 753 285 775 305
rect 703 269 775 285
rect 898 291 914 325
rect 948 305 981 325
rect 1060 351 1090 373
rect 1060 321 1096 351
rect 948 291 996 305
rect 898 275 996 291
rect 745 237 775 269
rect 966 253 996 275
rect 1066 253 1096 321
rect 1146 298 1176 373
rect 1275 341 1305 373
rect 1275 311 1323 341
rect 1146 268 1205 298
rect 214 111 244 137
rect 410 83 440 109
rect 510 83 540 109
rect 83 27 113 53
rect 1175 200 1205 268
rect 1293 200 1323 311
rect 1407 302 1437 383
rect 1514 304 1544 383
rect 1371 286 1437 302
rect 1371 252 1387 286
rect 1421 252 1437 286
rect 1371 236 1437 252
rect 1479 288 1551 304
rect 1479 254 1495 288
rect 1529 254 1551 288
rect 1479 238 1551 254
rect 1384 200 1414 236
rect 1514 200 1544 238
rect 745 43 775 69
rect 966 51 996 125
rect 1066 99 1096 125
rect 1175 51 1205 116
rect 966 21 1205 51
rect 1293 46 1323 72
rect 1384 46 1414 72
rect 1514 46 1544 72
<< polycont >>
rect 97 275 131 309
rect 221 285 255 319
rect 498 327 532 361
rect 719 285 753 319
rect 914 291 948 325
rect 1387 252 1421 286
rect 1495 254 1529 288
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 20 599 70 615
rect 20 565 36 599
rect 20 506 70 565
rect 20 472 36 506
rect 20 413 70 472
rect 106 607 156 649
rect 663 607 729 649
rect 106 573 122 607
rect 106 508 156 573
rect 106 474 122 508
rect 106 458 156 474
rect 190 573 451 607
rect 485 573 501 607
rect 663 573 679 607
rect 713 573 729 607
rect 867 579 1389 613
rect 867 576 933 579
rect 190 424 224 573
rect 867 542 883 576
rect 917 542 933 576
rect 1323 571 1389 579
rect 365 510 669 539
rect 20 379 36 413
rect 20 363 70 379
rect 122 390 224 424
rect 258 461 331 499
rect 292 427 331 461
rect 399 508 669 510
rect 976 529 1042 545
rect 1323 537 1339 571
rect 1373 537 1389 571
rect 976 508 992 529
rect 399 505 992 508
rect 399 476 415 505
rect 365 447 415 476
rect 635 495 992 505
rect 1026 495 1042 529
rect 635 474 1042 495
rect 567 455 601 471
rect 258 390 331 427
rect 20 225 54 363
rect 122 325 156 390
rect 297 377 331 390
rect 297 361 533 377
rect 88 309 156 325
rect 88 275 97 309
rect 131 275 156 309
rect 88 259 156 275
rect 205 319 263 356
rect 205 285 221 319
rect 255 285 263 319
rect 205 269 263 285
rect 297 327 498 361
rect 532 327 533 361
rect 297 311 533 327
rect 20 209 88 225
rect 20 175 38 209
rect 72 175 88 209
rect 20 101 88 175
rect 122 141 156 259
rect 297 225 331 311
rect 567 277 601 421
rect 239 209 331 225
rect 239 175 255 209
rect 289 175 331 209
rect 365 276 601 277
rect 365 242 511 276
rect 545 242 601 276
rect 365 236 601 242
rect 365 225 415 236
rect 399 191 415 225
rect 635 202 669 474
rect 749 424 932 440
rect 749 390 765 424
rect 799 406 932 424
rect 799 390 837 406
rect 703 319 769 356
rect 703 285 719 319
rect 753 285 769 319
rect 703 269 769 285
rect 803 225 837 390
rect 898 341 932 406
rect 976 425 1042 474
rect 976 391 992 425
rect 1026 391 1042 425
rect 976 375 1042 391
rect 1085 503 1289 537
rect 1085 498 1151 503
rect 1085 464 1087 498
rect 1121 489 1151 498
rect 1085 455 1101 464
rect 1135 455 1151 489
rect 1085 419 1151 455
rect 1085 385 1101 419
rect 1135 385 1151 419
rect 1085 369 1151 385
rect 1187 436 1221 469
rect 898 325 957 341
rect 1187 325 1221 402
rect 898 291 914 325
rect 948 291 957 325
rect 898 275 957 291
rect 991 291 1221 325
rect 1255 335 1289 503
rect 1323 503 1389 537
rect 1323 469 1339 503
rect 1373 469 1389 503
rect 1432 571 1498 649
rect 1432 537 1448 571
rect 1482 537 1498 571
rect 1432 503 1498 537
rect 1432 469 1448 503
rect 1482 469 1498 503
rect 1539 571 1615 587
rect 1539 537 1555 571
rect 1589 537 1615 571
rect 1539 500 1615 537
rect 1323 435 1389 469
rect 1539 466 1555 500
rect 1589 498 1615 500
rect 1539 464 1567 466
rect 1601 464 1615 498
rect 1323 419 1505 435
rect 1323 385 1339 419
rect 1373 385 1505 419
rect 1323 369 1505 385
rect 1539 429 1615 464
rect 1539 395 1555 429
rect 1589 395 1615 429
rect 1539 379 1615 395
rect 991 276 1057 291
rect 1025 242 1057 276
rect 1255 257 1313 335
rect 1471 304 1505 369
rect 991 241 1057 242
rect 365 175 415 191
rect 449 170 515 202
rect 449 141 465 170
rect 122 136 465 141
rect 499 136 515 170
rect 122 107 515 136
rect 449 105 515 107
rect 549 170 669 202
rect 770 191 786 225
rect 820 191 837 225
rect 985 225 1057 241
rect 985 191 1007 225
rect 1041 191 1057 225
rect 1091 239 1313 257
rect 1091 205 1107 239
rect 1141 223 1313 239
rect 1369 286 1437 302
rect 1369 252 1387 286
rect 1421 252 1437 286
rect 1369 236 1437 252
rect 1471 288 1529 304
rect 1471 254 1495 288
rect 1471 238 1529 254
rect 1141 205 1157 223
rect 1091 187 1157 205
rect 1471 189 1505 238
rect 1567 204 1615 379
rect 549 136 565 170
rect 599 157 669 170
rect 1223 170 1289 188
rect 599 153 1016 157
rect 1223 153 1239 170
rect 599 136 1239 153
rect 1273 136 1289 170
rect 549 123 1289 136
rect 549 105 615 123
rect 982 119 1289 123
rect 1323 186 1505 189
rect 1323 152 1339 186
rect 1373 155 1505 186
rect 1539 188 1615 204
rect 1373 152 1389 155
rect 1323 118 1389 152
rect 1539 154 1555 188
rect 1589 154 1615 188
rect 20 67 38 101
rect 72 67 88 101
rect 20 51 88 67
rect 130 39 146 73
rect 180 39 196 73
rect 130 17 196 39
rect 661 55 677 89
rect 711 55 727 89
rect 661 17 727 55
rect 882 55 898 89
rect 932 85 948 89
rect 1323 85 1339 118
rect 932 84 1339 85
rect 1373 84 1389 118
rect 932 55 1389 84
rect 882 51 1389 55
rect 1423 118 1489 121
rect 1423 84 1439 118
rect 1473 84 1489 118
rect 1423 17 1489 84
rect 1539 118 1615 154
rect 1539 84 1555 118
rect 1589 84 1615 118
rect 1539 68 1615 84
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 511 242 545 276
rect 1087 489 1121 498
rect 1087 464 1101 489
rect 1101 464 1121 489
rect 1567 466 1589 498
rect 1589 466 1601 498
rect 1567 464 1601 466
rect 991 242 1025 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 1075 498 1133 504
rect 1075 464 1087 498
rect 1121 495 1133 498
rect 1555 498 1613 504
rect 1555 495 1567 498
rect 1121 467 1567 495
rect 1121 464 1133 467
rect 1075 458 1133 464
rect 1555 464 1567 467
rect 1601 464 1613 498
rect 1555 458 1613 464
rect 499 276 557 282
rect 499 242 511 276
rect 545 273 557 276
rect 979 276 1037 282
rect 979 273 991 276
rect 545 245 991 273
rect 545 242 557 245
rect 499 236 557 242
rect 979 242 991 245
rect 1025 242 1037 276
rect 979 236 1037 242
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xnor3_1
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 733306
string GDS_START 721414
<< end >>
