magic
tech sky130A
magscale 1 2
timestamp 1627202617
<< checkpaint >>
rect -1298 -1308 2218 1852
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 861 203
rect 30 -17 64 21
<< scnmos >>
rect 80 47 110 177
rect 166 47 196 177
rect 356 47 386 177
rect 428 47 458 177
rect 536 47 566 177
rect 644 47 674 177
rect 752 47 782 177
<< scpmoshvt >>
rect 80 297 110 497
rect 166 297 196 497
rect 342 297 372 497
rect 428 297 458 497
rect 536 297 566 497
rect 644 297 674 497
rect 752 297 782 497
<< ndiff >>
rect 27 161 80 177
rect 27 127 35 161
rect 69 127 80 161
rect 27 93 80 127
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 169 166 177
rect 110 135 121 169
rect 155 135 166 169
rect 110 101 166 135
rect 110 67 121 101
rect 155 67 166 101
rect 110 47 166 67
rect 196 93 249 177
rect 196 59 207 93
rect 241 59 249 93
rect 196 47 249 59
rect 303 165 356 177
rect 303 131 311 165
rect 345 131 356 165
rect 303 97 356 131
rect 303 63 311 97
rect 345 63 356 97
rect 303 47 356 63
rect 386 47 428 177
rect 458 47 536 177
rect 566 165 644 177
rect 566 131 589 165
rect 623 131 644 165
rect 566 97 644 131
rect 566 63 589 97
rect 623 63 644 97
rect 566 47 644 63
rect 674 91 752 177
rect 674 57 693 91
rect 727 57 752 91
rect 674 47 752 57
rect 782 165 835 177
rect 782 131 793 165
rect 827 131 835 165
rect 782 97 835 131
rect 782 63 793 97
rect 827 63 835 97
rect 782 47 835 63
<< pdiff >>
rect 27 485 80 497
rect 27 451 35 485
rect 69 451 80 485
rect 27 417 80 451
rect 27 383 35 417
rect 69 383 80 417
rect 27 349 80 383
rect 27 315 35 349
rect 69 315 80 349
rect 27 297 80 315
rect 110 485 166 497
rect 110 451 121 485
rect 155 451 166 485
rect 110 417 166 451
rect 110 383 121 417
rect 155 383 166 417
rect 110 349 166 383
rect 110 315 121 349
rect 155 315 166 349
rect 110 297 166 315
rect 196 489 342 497
rect 196 455 207 489
rect 241 455 297 489
rect 331 455 342 489
rect 196 297 342 455
rect 372 477 428 497
rect 372 443 383 477
rect 417 443 428 477
rect 372 394 428 443
rect 372 360 383 394
rect 417 360 428 394
rect 372 297 428 360
rect 458 485 536 497
rect 458 451 481 485
rect 515 451 536 485
rect 458 297 536 451
rect 566 485 644 497
rect 566 451 589 485
rect 623 451 644 485
rect 566 394 644 451
rect 566 360 589 394
rect 623 360 644 394
rect 566 297 644 360
rect 674 297 752 497
rect 782 485 835 497
rect 782 451 793 485
rect 827 451 835 485
rect 782 417 835 451
rect 782 383 793 417
rect 827 383 835 417
rect 782 349 835 383
rect 782 315 793 349
rect 827 315 835 349
rect 782 297 835 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 121 135 155 169
rect 121 67 155 101
rect 207 59 241 93
rect 311 131 345 165
rect 311 63 345 97
rect 589 131 623 165
rect 589 63 623 97
rect 693 57 727 91
rect 793 131 827 165
rect 793 63 827 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 121 451 155 485
rect 121 383 155 417
rect 121 315 155 349
rect 207 455 241 489
rect 297 455 331 489
rect 383 443 417 477
rect 383 360 417 394
rect 481 451 515 485
rect 589 451 623 485
rect 589 360 623 394
rect 793 451 827 485
rect 793 383 827 417
rect 793 315 827 349
<< poly >>
rect 80 497 110 523
rect 166 497 196 523
rect 342 497 372 523
rect 428 497 458 523
rect 536 497 566 523
rect 644 497 674 523
rect 752 497 782 523
rect 80 265 110 297
rect 166 265 196 297
rect 342 265 372 297
rect 80 249 250 265
rect 80 215 206 249
rect 240 215 250 249
rect 80 199 250 215
rect 301 249 386 265
rect 301 215 317 249
rect 351 215 386 249
rect 301 199 386 215
rect 80 177 110 199
rect 166 177 196 199
rect 356 177 386 199
rect 428 259 458 297
rect 536 259 566 297
rect 644 259 674 297
rect 752 259 782 297
rect 428 249 494 259
rect 428 215 444 249
rect 478 215 494 249
rect 428 205 494 215
rect 536 249 602 259
rect 536 215 552 249
rect 586 215 602 249
rect 536 205 602 215
rect 644 249 710 259
rect 644 215 660 249
rect 694 215 710 249
rect 644 205 710 215
rect 752 249 843 259
rect 752 215 793 249
rect 827 215 843 249
rect 752 205 843 215
rect 428 177 458 205
rect 536 177 566 205
rect 644 177 674 205
rect 752 177 782 205
rect 80 21 110 47
rect 166 21 196 47
rect 356 21 386 47
rect 428 21 458 47
rect 536 21 566 47
rect 644 21 674 47
rect 752 21 782 47
<< polycont >>
rect 206 215 240 249
rect 317 215 351 249
rect 444 215 478 249
rect 552 215 586 249
rect 660 215 694 249
rect 793 215 827 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 27 485 69 527
rect 27 451 35 485
rect 27 417 69 451
rect 27 383 35 417
rect 27 349 69 383
rect 27 315 35 349
rect 27 299 69 315
rect 103 485 171 493
rect 103 451 121 485
rect 155 451 171 485
rect 103 417 171 451
rect 207 489 331 527
rect 241 455 297 489
rect 207 439 331 455
rect 372 477 428 493
rect 372 443 383 477
rect 417 443 428 477
rect 465 485 531 527
rect 465 451 481 485
rect 515 451 531 485
rect 573 485 639 493
rect 573 451 589 485
rect 623 451 639 485
rect 777 485 828 527
rect 103 383 121 417
rect 155 383 171 417
rect 372 405 428 443
rect 573 405 639 451
rect 103 349 171 383
rect 103 315 121 349
rect 155 315 171 349
rect 27 161 69 177
rect 27 127 35 161
rect 27 93 69 127
rect 27 59 35 93
rect 27 17 69 59
rect 103 169 171 315
rect 103 135 121 169
rect 155 135 171 169
rect 206 394 639 405
rect 206 360 383 394
rect 417 360 589 394
rect 623 360 639 394
rect 206 357 639 360
rect 206 249 261 357
rect 240 215 261 249
rect 301 249 367 323
rect 301 215 317 249
rect 351 215 367 249
rect 401 249 478 323
rect 401 215 444 249
rect 536 249 620 323
rect 674 265 732 474
rect 777 451 793 485
rect 827 451 828 485
rect 777 417 828 451
rect 777 383 793 417
rect 827 383 828 417
rect 777 349 828 383
rect 777 315 793 349
rect 827 315 828 349
rect 777 299 828 315
rect 536 215 552 249
rect 586 215 620 249
rect 660 249 732 265
rect 862 263 903 471
rect 694 215 732 249
rect 206 177 261 215
rect 206 165 361 177
rect 206 143 311 165
rect 103 101 171 135
rect 295 131 311 143
rect 345 131 361 165
rect 103 67 121 101
rect 155 67 171 101
rect 103 51 171 67
rect 207 93 257 109
rect 241 59 257 93
rect 207 17 257 59
rect 295 97 361 131
rect 295 63 311 97
rect 345 63 361 97
rect 295 51 361 63
rect 401 51 478 215
rect 660 199 732 215
rect 766 249 903 263
rect 766 215 793 249
rect 827 215 903 249
rect 766 201 903 215
rect 573 131 589 165
rect 623 131 793 165
rect 827 131 843 165
rect 573 125 843 131
rect 573 97 639 125
rect 573 63 589 97
rect 623 63 639 97
rect 777 97 843 125
rect 573 51 639 63
rect 677 57 693 91
rect 727 57 743 91
rect 677 17 743 57
rect 777 63 793 97
rect 827 63 843 97
rect 777 51 843 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 310 221 344 255 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 402 85 436 119 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 678 425 712 459 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 678 221 712 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 770 221 804 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 586 221 620 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 122 425 156 459 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 122 85 156 119 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 862 221 896 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o2111a_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 2905472
string GDS_START 2897364
string path 0.000 0.000 23.000 0.000 
<< end >>
