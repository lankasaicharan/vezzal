magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3698 1975
<< nwell >>
rect -38 331 2438 704
<< pwell >>
rect 1141 241 1852 243
rect 1141 229 2397 241
rect 422 200 2397 229
rect 1 49 2397 200
rect 0 0 2400 49
<< scnmos >>
rect 80 90 110 174
rect 248 90 278 174
rect 501 119 531 203
rect 573 119 603 203
rect 659 119 689 203
rect 799 119 829 203
rect 875 119 905 203
rect 983 105 1013 189
rect 1115 61 1145 189
rect 1247 61 1277 189
rect 1419 133 1449 217
rect 1527 133 1557 217
rect 1667 133 1697 217
rect 1739 133 1769 217
rect 1944 47 1974 215
rect 2030 47 2060 215
rect 2116 47 2146 215
rect 2202 47 2232 215
rect 2288 47 2318 215
<< scpmoshvt >>
rect 100 462 130 590
rect 186 462 216 590
rect 393 535 423 619
rect 479 535 509 619
rect 565 535 595 619
rect 659 535 689 619
rect 731 535 761 619
rect 832 535 862 619
rect 1139 449 1169 617
rect 1225 449 1255 617
rect 1350 488 1380 572
rect 1475 488 1505 572
rect 1648 488 1678 572
rect 1739 488 1769 572
rect 1944 367 1974 619
rect 2030 367 2060 619
rect 2116 367 2146 619
rect 2202 367 2232 619
rect 2288 367 2318 619
<< ndiff >>
rect 27 149 80 174
rect 27 115 35 149
rect 69 115 80 149
rect 27 90 80 115
rect 110 132 248 174
rect 110 98 123 132
rect 157 98 248 132
rect 110 90 248 98
rect 278 162 335 174
rect 278 128 293 162
rect 327 128 335 162
rect 278 90 335 128
rect 448 167 501 203
rect 448 133 456 167
rect 490 133 501 167
rect 448 119 501 133
rect 531 119 573 203
rect 603 195 659 203
rect 603 161 614 195
rect 648 161 659 195
rect 603 119 659 161
rect 689 193 799 203
rect 689 159 754 193
rect 788 159 799 193
rect 689 119 799 159
rect 829 119 875 203
rect 905 189 955 203
rect 1167 209 1225 217
rect 1167 189 1179 209
rect 905 119 983 189
rect 933 105 983 119
rect 1013 105 1115 189
rect 1035 69 1115 105
rect 1035 35 1047 69
rect 1081 61 1115 69
rect 1145 175 1179 189
rect 1213 189 1225 209
rect 1299 209 1419 217
rect 1299 189 1347 209
rect 1213 175 1247 189
rect 1145 61 1247 175
rect 1277 175 1347 189
rect 1381 175 1419 209
rect 1277 133 1419 175
rect 1449 133 1527 217
rect 1557 180 1667 217
rect 1557 146 1595 180
rect 1629 146 1667 180
rect 1557 133 1667 146
rect 1697 133 1739 217
rect 1769 180 1826 217
rect 1769 146 1784 180
rect 1818 146 1826 180
rect 1769 133 1826 146
rect 1891 203 1944 215
rect 1891 169 1899 203
rect 1933 169 1944 203
rect 1277 61 1397 133
rect 1081 35 1093 61
rect 1891 101 1944 169
rect 1891 67 1899 101
rect 1933 67 1944 101
rect 1891 47 1944 67
rect 1974 203 2030 215
rect 1974 169 1985 203
rect 2019 169 2030 203
rect 1974 89 2030 169
rect 1974 55 1985 89
rect 2019 55 2030 89
rect 1974 47 2030 55
rect 2060 207 2116 215
rect 2060 173 2071 207
rect 2105 173 2116 207
rect 2060 101 2116 173
rect 2060 67 2071 101
rect 2105 67 2116 101
rect 2060 47 2116 67
rect 2146 163 2202 215
rect 2146 129 2157 163
rect 2191 129 2202 163
rect 2146 89 2202 129
rect 2146 55 2157 89
rect 2191 55 2202 89
rect 2146 47 2202 55
rect 2232 207 2288 215
rect 2232 173 2243 207
rect 2277 173 2288 207
rect 2232 101 2288 173
rect 2232 67 2243 101
rect 2277 67 2288 101
rect 2232 47 2288 67
rect 2318 179 2371 215
rect 2318 145 2329 179
rect 2363 145 2371 179
rect 2318 93 2371 145
rect 2318 59 2329 93
rect 2363 59 2371 93
rect 2318 47 2371 59
rect 1035 27 1093 35
<< pdiff >>
rect 1059 631 1117 639
rect 340 594 393 619
rect 47 578 100 590
rect 47 544 55 578
rect 89 544 100 578
rect 47 510 100 544
rect 47 476 55 510
rect 89 476 100 510
rect 47 462 100 476
rect 130 578 186 590
rect 130 544 141 578
rect 175 544 186 578
rect 130 462 186 544
rect 216 576 269 590
rect 216 542 227 576
rect 261 542 269 576
rect 216 508 269 542
rect 340 560 348 594
rect 382 560 393 594
rect 340 535 393 560
rect 423 600 479 619
rect 423 566 434 600
rect 468 566 479 600
rect 423 535 479 566
rect 509 594 565 619
rect 509 560 520 594
rect 554 560 565 594
rect 509 535 565 560
rect 595 599 659 619
rect 595 565 614 599
rect 648 565 659 599
rect 595 535 659 565
rect 689 535 731 619
rect 761 609 832 619
rect 761 575 787 609
rect 821 575 832 609
rect 761 535 832 575
rect 862 594 915 619
rect 862 560 873 594
rect 907 560 915 594
rect 862 535 915 560
rect 1059 597 1071 631
rect 1105 617 1117 631
rect 1105 597 1139 617
rect 216 474 227 508
rect 261 474 269 508
rect 216 462 269 474
rect 1059 449 1139 597
rect 1169 491 1225 617
rect 1169 457 1180 491
rect 1214 457 1225 491
rect 1169 449 1225 457
rect 1255 572 1324 617
rect 1891 599 1944 619
rect 1255 519 1350 572
rect 1255 485 1282 519
rect 1316 488 1350 519
rect 1380 488 1475 572
rect 1505 564 1648 572
rect 1505 530 1559 564
rect 1593 530 1648 564
rect 1505 488 1648 530
rect 1678 547 1739 572
rect 1678 513 1689 547
rect 1723 513 1739 547
rect 1678 488 1739 513
rect 1769 564 1837 572
rect 1769 530 1791 564
rect 1825 530 1837 564
rect 1769 488 1837 530
rect 1891 565 1899 599
rect 1933 565 1944 599
rect 1891 508 1944 565
rect 1316 485 1324 488
rect 1255 471 1324 485
rect 1255 449 1305 471
rect 1891 474 1899 508
rect 1933 474 1944 508
rect 1891 413 1944 474
rect 1891 379 1899 413
rect 1933 379 1944 413
rect 1891 367 1944 379
rect 1974 611 2030 619
rect 1974 577 1985 611
rect 2019 577 2030 611
rect 1974 513 2030 577
rect 1974 479 1985 513
rect 2019 479 2030 513
rect 1974 413 2030 479
rect 1974 379 1985 413
rect 2019 379 2030 413
rect 1974 367 2030 379
rect 2060 599 2116 619
rect 2060 565 2071 599
rect 2105 565 2116 599
rect 2060 508 2116 565
rect 2060 474 2071 508
rect 2105 474 2116 508
rect 2060 409 2116 474
rect 2060 375 2071 409
rect 2105 375 2116 409
rect 2060 367 2116 375
rect 2146 611 2202 619
rect 2146 577 2157 611
rect 2191 577 2202 611
rect 2146 532 2202 577
rect 2146 498 2157 532
rect 2191 498 2202 532
rect 2146 453 2202 498
rect 2146 419 2157 453
rect 2191 419 2202 453
rect 2146 367 2202 419
rect 2232 599 2288 619
rect 2232 565 2243 599
rect 2277 565 2288 599
rect 2232 508 2288 565
rect 2232 474 2243 508
rect 2277 474 2288 508
rect 2232 409 2288 474
rect 2232 375 2243 409
rect 2277 375 2288 409
rect 2232 367 2288 375
rect 2318 607 2371 619
rect 2318 573 2329 607
rect 2363 573 2371 607
rect 2318 532 2371 573
rect 2318 498 2329 532
rect 2363 498 2371 532
rect 2318 453 2371 498
rect 2318 419 2329 453
rect 2363 419 2371 453
rect 2318 367 2371 419
<< ndiffc >>
rect 35 115 69 149
rect 123 98 157 132
rect 293 128 327 162
rect 456 133 490 167
rect 614 161 648 195
rect 754 159 788 193
rect 1047 35 1081 69
rect 1179 175 1213 209
rect 1347 175 1381 209
rect 1595 146 1629 180
rect 1784 146 1818 180
rect 1899 169 1933 203
rect 1899 67 1933 101
rect 1985 169 2019 203
rect 1985 55 2019 89
rect 2071 173 2105 207
rect 2071 67 2105 101
rect 2157 129 2191 163
rect 2157 55 2191 89
rect 2243 173 2277 207
rect 2243 67 2277 101
rect 2329 145 2363 179
rect 2329 59 2363 93
<< pdiffc >>
rect 55 544 89 578
rect 55 476 89 510
rect 141 544 175 578
rect 227 542 261 576
rect 348 560 382 594
rect 434 566 468 600
rect 520 560 554 594
rect 614 565 648 599
rect 787 575 821 609
rect 873 560 907 594
rect 1071 597 1105 631
rect 227 474 261 508
rect 1180 457 1214 491
rect 1282 485 1316 519
rect 1559 530 1593 564
rect 1689 513 1723 547
rect 1791 530 1825 564
rect 1899 565 1933 599
rect 1899 474 1933 508
rect 1899 379 1933 413
rect 1985 577 2019 611
rect 1985 479 2019 513
rect 1985 379 2019 413
rect 2071 565 2105 599
rect 2071 474 2105 508
rect 2071 375 2105 409
rect 2157 577 2191 611
rect 2157 498 2191 532
rect 2157 419 2191 453
rect 2243 565 2277 599
rect 2243 474 2277 508
rect 2243 375 2277 409
rect 2329 573 2363 607
rect 2329 498 2363 532
rect 2329 419 2363 453
<< poly >>
rect 393 619 423 645
rect 479 619 509 645
rect 565 619 595 645
rect 659 619 689 645
rect 731 619 761 645
rect 832 619 862 645
rect 100 590 130 616
rect 186 590 216 616
rect 1139 617 1169 643
rect 1225 617 1255 643
rect 1944 619 1974 645
rect 2030 619 2060 645
rect 2116 619 2146 645
rect 2202 619 2232 645
rect 2288 619 2318 645
rect 100 408 130 462
rect 44 392 130 408
rect 44 358 60 392
rect 94 378 130 392
rect 94 358 110 378
rect 44 324 110 358
rect 186 330 216 462
rect 44 290 60 324
rect 94 290 110 324
rect 44 274 110 290
rect 80 174 110 274
rect 158 314 278 330
rect 158 280 174 314
rect 208 280 278 314
rect 158 246 278 280
rect 158 212 174 246
rect 208 212 278 246
rect 158 196 278 212
rect 248 174 278 196
rect 80 64 110 90
rect 248 64 278 90
rect 393 51 423 535
rect 479 435 509 535
rect 565 471 595 535
rect 473 405 509 435
rect 551 455 617 471
rect 551 421 567 455
rect 601 421 617 455
rect 551 405 617 421
rect 473 357 503 405
rect 473 341 603 357
rect 473 307 489 341
rect 523 307 603 341
rect 473 291 603 307
rect 501 203 531 229
rect 573 203 603 291
rect 659 313 689 535
rect 731 435 761 535
rect 832 507 862 535
rect 832 487 1013 507
rect 832 477 963 487
rect 947 453 963 477
rect 997 453 1013 487
rect 947 437 1013 453
rect 1350 572 1380 598
rect 1475 572 1505 598
rect 1648 572 1678 598
rect 1739 572 1769 598
rect 731 405 905 435
rect 875 363 905 405
rect 767 347 833 363
rect 767 313 783 347
rect 817 313 833 347
rect 659 297 725 313
rect 659 263 675 297
rect 709 263 725 297
rect 659 247 725 263
rect 767 279 833 313
rect 659 203 689 247
rect 767 245 783 279
rect 817 245 833 279
rect 767 229 833 245
rect 875 347 941 363
rect 875 313 891 347
rect 925 313 941 347
rect 875 279 941 313
rect 875 245 891 279
rect 925 245 941 279
rect 875 229 941 245
rect 799 203 829 229
rect 875 203 905 229
rect 983 189 1013 437
rect 1139 417 1169 449
rect 1055 401 1169 417
rect 1055 367 1071 401
rect 1105 387 1169 401
rect 1225 391 1255 449
rect 1350 439 1380 488
rect 1475 456 1505 488
rect 1475 440 1589 456
rect 1341 423 1433 439
rect 1475 426 1539 440
rect 1105 367 1121 387
rect 1055 351 1121 367
rect 1211 375 1277 391
rect 1055 277 1085 351
rect 1211 341 1227 375
rect 1261 341 1277 375
rect 1211 325 1277 341
rect 1341 389 1383 423
rect 1417 389 1433 423
rect 1505 406 1539 426
rect 1573 406 1589 440
rect 1648 424 1678 488
rect 1505 390 1589 406
rect 1631 408 1697 424
rect 1341 373 1433 389
rect 1055 261 1145 277
rect 1341 262 1371 373
rect 1055 227 1071 261
rect 1105 227 1145 261
rect 1055 211 1145 227
rect 1247 232 1371 262
rect 1115 189 1145 211
rect 501 51 531 119
rect 573 93 603 119
rect 659 93 689 119
rect 799 93 829 119
rect 875 93 905 119
rect 983 51 1013 105
rect 393 21 1013 51
rect 1247 189 1277 232
rect 1419 217 1449 243
rect 1527 217 1557 390
rect 1631 374 1647 408
rect 1681 374 1697 408
rect 1631 340 1697 374
rect 1631 306 1647 340
rect 1681 306 1697 340
rect 1631 290 1697 306
rect 1667 217 1697 290
rect 1739 373 1769 488
rect 1739 357 1805 373
rect 1739 323 1755 357
rect 1789 323 1805 357
rect 1739 289 1805 323
rect 1739 255 1755 289
rect 1789 269 1805 289
rect 1944 269 1974 367
rect 1789 255 1974 269
rect 1739 239 1974 255
rect 1739 217 1769 239
rect 1944 215 1974 239
rect 2030 331 2060 367
rect 2116 331 2146 367
rect 2202 331 2232 367
rect 2288 331 2318 367
rect 2030 315 2318 331
rect 2030 281 2046 315
rect 2080 281 2114 315
rect 2148 281 2182 315
rect 2216 281 2250 315
rect 2284 281 2318 315
rect 2030 265 2318 281
rect 2030 215 2060 265
rect 2116 215 2146 265
rect 2202 215 2232 265
rect 2288 215 2318 265
rect 1419 111 1449 133
rect 1419 95 1485 111
rect 1527 107 1557 133
rect 1667 107 1697 133
rect 1739 107 1769 133
rect 1419 61 1435 95
rect 1469 61 1485 95
rect 1115 35 1145 61
rect 1247 35 1277 61
rect 1419 45 1485 61
rect 1944 21 1974 47
rect 2030 21 2060 47
rect 2116 21 2146 47
rect 2202 21 2232 47
rect 2288 21 2318 47
<< polycont >>
rect 60 358 94 392
rect 60 290 94 324
rect 174 280 208 314
rect 174 212 208 246
rect 567 421 601 455
rect 489 307 523 341
rect 963 453 997 487
rect 783 313 817 347
rect 675 263 709 297
rect 783 245 817 279
rect 891 313 925 347
rect 891 245 925 279
rect 1071 367 1105 401
rect 1227 341 1261 375
rect 1383 389 1417 423
rect 1539 406 1573 440
rect 1071 227 1105 261
rect 1647 374 1681 408
rect 1647 306 1681 340
rect 1755 323 1789 357
rect 1755 255 1789 289
rect 2046 281 2080 315
rect 2114 281 2148 315
rect 2182 281 2216 315
rect 2250 281 2284 315
rect 1435 61 1469 95
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 39 578 91 594
rect 39 544 55 578
rect 89 544 91 578
rect 39 510 91 544
rect 125 578 187 649
rect 332 594 384 610
rect 125 544 141 578
rect 175 544 187 578
rect 125 528 187 544
rect 221 576 277 592
rect 221 542 227 576
rect 261 542 277 576
rect 39 476 55 510
rect 89 494 91 510
rect 221 508 277 542
rect 89 476 187 494
rect 39 460 187 476
rect 17 392 94 426
rect 17 358 60 392
rect 17 324 94 358
rect 17 290 60 324
rect 17 240 94 290
rect 153 330 187 460
rect 221 474 227 508
rect 261 474 277 508
rect 332 560 348 594
rect 382 560 384 594
rect 332 525 384 560
rect 418 600 484 649
rect 418 566 434 600
rect 468 566 484 600
rect 418 559 484 566
rect 518 594 564 610
rect 518 560 520 594
rect 554 560 564 594
rect 518 525 564 560
rect 598 599 753 615
rect 598 565 614 599
rect 648 565 753 599
rect 598 559 753 565
rect 787 609 830 649
rect 1055 631 1121 649
rect 821 575 830 609
rect 787 559 830 575
rect 864 594 917 610
rect 1055 597 1071 631
rect 1105 597 1121 631
rect 1055 595 1121 597
rect 864 560 873 594
rect 907 560 917 594
rect 1157 561 1503 591
rect 719 525 753 559
rect 864 525 917 560
rect 979 557 1503 561
rect 979 527 1191 557
rect 332 491 685 525
rect 719 491 909 525
rect 979 504 1013 527
rect 221 457 277 474
rect 221 455 617 457
rect 221 424 567 455
rect 221 390 223 424
rect 257 421 567 424
rect 601 421 617 455
rect 257 417 617 421
rect 257 390 343 417
rect 221 374 343 390
rect 651 383 685 491
rect 153 314 241 330
rect 153 280 174 314
rect 208 280 241 314
rect 153 246 241 280
rect 153 212 174 246
rect 208 212 241 246
rect 153 206 241 212
rect 19 172 241 206
rect 19 149 71 172
rect 19 115 35 149
rect 69 115 71 149
rect 19 99 71 115
rect 105 132 173 138
rect 105 98 123 132
rect 157 98 173 132
rect 105 17 173 98
rect 207 92 241 172
rect 277 162 343 374
rect 395 341 564 370
rect 395 307 489 341
rect 523 307 564 341
rect 395 291 564 307
rect 598 349 685 383
rect 767 424 841 436
rect 767 390 799 424
rect 833 390 841 424
rect 277 128 293 162
rect 327 128 343 162
rect 277 126 343 128
rect 379 217 564 251
rect 379 92 413 217
rect 207 58 413 92
rect 447 167 496 183
rect 447 133 456 167
rect 490 133 496 167
rect 447 17 496 133
rect 530 107 564 217
rect 598 211 639 349
rect 767 347 841 390
rect 875 417 909 491
rect 947 487 1013 504
rect 1266 519 1332 523
rect 947 453 963 487
rect 997 453 1013 487
rect 947 451 1013 453
rect 1157 491 1230 493
rect 1157 457 1180 491
rect 1214 457 1230 491
rect 1266 485 1282 519
rect 1316 485 1332 519
rect 1266 469 1332 485
rect 1157 441 1230 457
rect 875 401 1121 417
rect 875 383 1071 401
rect 1055 367 1071 383
rect 1105 367 1121 401
rect 1055 365 1121 367
rect 767 313 783 347
rect 817 313 841 347
rect 673 297 718 313
rect 673 263 675 297
rect 709 263 718 297
rect 673 247 718 263
rect 598 195 650 211
rect 598 161 614 195
rect 648 161 650 195
rect 598 145 650 161
rect 684 107 718 247
rect 767 279 841 313
rect 767 245 783 279
rect 817 245 841 279
rect 767 243 841 245
rect 875 347 941 349
rect 875 313 891 347
rect 925 331 941 347
rect 1157 331 1191 441
rect 925 313 1191 331
rect 875 297 1191 313
rect 875 279 941 297
rect 875 245 891 279
rect 925 245 941 279
rect 875 243 941 245
rect 1055 261 1121 263
rect 1055 227 1071 261
rect 1105 227 1121 261
rect 1055 209 1121 227
rect 752 193 1121 209
rect 752 159 754 193
rect 788 175 1121 193
rect 1157 213 1191 297
rect 1225 375 1263 391
rect 1225 341 1227 375
rect 1261 341 1263 375
rect 1225 283 1263 341
rect 1297 353 1332 469
rect 1366 424 1433 439
rect 1366 390 1375 424
rect 1409 423 1433 424
rect 1366 389 1383 390
rect 1417 389 1433 423
rect 1366 387 1433 389
rect 1297 319 1369 353
rect 1225 249 1297 283
rect 1157 209 1229 213
rect 1157 175 1179 209
rect 1213 175 1229 209
rect 788 159 792 175
rect 1157 173 1229 175
rect 752 143 792 159
rect 1263 139 1297 249
rect 1331 254 1369 319
rect 1469 324 1503 557
rect 1543 564 1609 649
rect 1543 530 1559 564
rect 1593 530 1609 564
rect 1775 564 1841 649
rect 1543 528 1609 530
rect 1673 547 1739 563
rect 1673 513 1689 547
rect 1723 513 1739 547
rect 1775 530 1791 564
rect 1825 530 1841 564
rect 1775 528 1841 530
rect 1893 599 1942 615
rect 1893 565 1899 599
rect 1933 565 1942 599
rect 1673 494 1739 513
rect 1893 508 1942 565
rect 1537 460 1859 494
rect 1537 440 1589 460
rect 1537 406 1539 440
rect 1573 406 1589 440
rect 1537 390 1589 406
rect 1631 408 1713 424
rect 1631 374 1647 408
rect 1681 374 1713 408
rect 1631 340 1713 374
rect 1631 324 1647 340
rect 1469 306 1647 324
rect 1681 306 1713 340
rect 1469 290 1713 306
rect 1747 357 1791 373
rect 1747 323 1755 357
rect 1789 323 1791 357
rect 1747 289 1791 323
rect 1747 255 1755 289
rect 1789 255 1791 289
rect 1747 254 1791 255
rect 1331 220 1791 254
rect 1331 209 1397 220
rect 1331 175 1347 209
rect 1381 175 1397 209
rect 1825 186 1859 460
rect 1331 173 1397 175
rect 1579 180 1645 186
rect 1579 146 1595 180
rect 1629 146 1645 180
rect 828 107 1485 139
rect 530 105 1485 107
rect 530 73 862 105
rect 1419 95 1485 105
rect 1031 69 1097 71
rect 1031 35 1047 69
rect 1081 35 1097 69
rect 1419 61 1435 95
rect 1469 61 1485 95
rect 1419 51 1485 61
rect 1031 17 1097 35
rect 1579 17 1645 146
rect 1768 180 1859 186
rect 1768 146 1784 180
rect 1818 146 1859 180
rect 1768 130 1859 146
rect 1893 474 1899 508
rect 1933 474 1942 508
rect 1893 413 1942 474
rect 1893 379 1899 413
rect 1933 379 1942 413
rect 1893 317 1942 379
rect 1976 611 2028 649
rect 1976 577 1985 611
rect 2019 577 2028 611
rect 1976 513 2028 577
rect 1976 479 1985 513
rect 2019 479 2028 513
rect 1976 413 2028 479
rect 1976 379 1985 413
rect 2019 379 2028 413
rect 1976 363 2028 379
rect 2062 599 2107 615
rect 2062 565 2071 599
rect 2105 565 2107 599
rect 2062 508 2107 565
rect 2062 474 2071 508
rect 2105 474 2107 508
rect 2062 409 2107 474
rect 2141 611 2207 649
rect 2141 577 2157 611
rect 2191 577 2207 611
rect 2141 532 2207 577
rect 2141 498 2157 532
rect 2191 498 2207 532
rect 2141 453 2207 498
rect 2141 419 2157 453
rect 2191 419 2207 453
rect 2241 599 2279 615
rect 2241 565 2243 599
rect 2277 565 2279 599
rect 2241 508 2279 565
rect 2241 474 2243 508
rect 2277 474 2279 508
rect 2062 375 2071 409
rect 2105 385 2107 409
rect 2241 409 2279 474
rect 2313 607 2379 649
rect 2313 573 2329 607
rect 2363 573 2379 607
rect 2313 532 2379 573
rect 2313 498 2329 532
rect 2363 498 2379 532
rect 2313 453 2379 498
rect 2313 419 2329 453
rect 2363 419 2379 453
rect 2241 385 2243 409
rect 2105 375 2243 385
rect 2277 385 2279 409
rect 2277 375 2370 385
rect 2062 351 2370 375
rect 1893 315 2300 317
rect 1893 281 2046 315
rect 2080 281 2114 315
rect 2148 281 2182 315
rect 2216 281 2250 315
rect 2284 281 2300 315
rect 1893 203 1942 281
rect 2336 247 2370 351
rect 1893 169 1899 203
rect 1933 169 1942 203
rect 1893 101 1942 169
rect 1893 67 1899 101
rect 1933 67 1942 101
rect 1893 51 1942 67
rect 1976 203 2028 219
rect 1976 169 1985 203
rect 2019 169 2028 203
rect 1976 89 2028 169
rect 1976 55 1985 89
rect 2019 55 2028 89
rect 1976 17 2028 55
rect 2062 213 2370 247
rect 2062 207 2107 213
rect 2062 173 2071 207
rect 2105 173 2107 207
rect 2230 207 2279 213
rect 2062 101 2107 173
rect 2062 67 2071 101
rect 2105 67 2107 101
rect 2062 51 2107 67
rect 2141 163 2196 179
rect 2141 129 2157 163
rect 2191 129 2196 163
rect 2141 89 2196 129
rect 2141 55 2157 89
rect 2191 55 2196 89
rect 2141 17 2196 55
rect 2230 173 2243 207
rect 2277 173 2279 207
rect 2230 101 2279 173
rect 2230 67 2243 101
rect 2277 67 2279 101
rect 2230 51 2279 67
rect 2313 145 2329 179
rect 2363 145 2379 179
rect 2313 93 2379 145
rect 2313 59 2329 93
rect 2363 59 2379 93
rect 2313 17 2379 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 223 390 257 424
rect 799 390 833 424
rect 1375 423 1409 424
rect 1375 390 1383 423
rect 1383 390 1409 423
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 787 424 845 430
rect 787 421 799 424
rect 257 393 799 421
rect 257 390 269 393
rect 211 384 269 390
rect 787 390 799 393
rect 833 421 845 424
rect 1363 424 1421 430
rect 1363 421 1375 424
rect 833 393 1375 421
rect 833 390 845 393
rect 787 384 845 390
rect 1363 390 1375 393
rect 1409 390 1421 424
rect 1363 384 1421 390
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< labels >>
flabel pwell s 0 0 2400 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2400 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfrtp_4
flabel comment s 1065 322 1065 322 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 2400 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2400 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1663 390 1697 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2239 168 2273 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2400 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 555228
string GDS_START 537588
<< end >>
