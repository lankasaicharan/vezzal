magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 1 49 1529 247
rect 0 0 1536 49
<< scnmos >>
rect 84 53 114 221
rect 170 53 200 221
rect 256 53 286 221
rect 342 53 372 221
rect 428 53 458 221
rect 514 53 544 221
rect 600 53 630 221
rect 686 53 716 221
rect 772 53 802 221
rect 858 53 888 221
rect 944 53 974 221
rect 1030 53 1060 221
rect 1116 53 1146 221
rect 1216 53 1246 221
rect 1316 53 1346 221
rect 1416 53 1446 221
<< scpmoshvt >>
rect 84 367 114 619
rect 170 367 200 619
rect 256 367 286 619
rect 342 367 372 619
rect 428 367 458 619
rect 514 367 544 619
rect 628 367 658 619
rect 714 367 744 619
rect 800 367 830 619
rect 886 367 916 619
rect 972 367 1002 619
rect 1058 367 1088 619
rect 1144 367 1174 619
rect 1230 367 1260 619
rect 1330 367 1360 619
rect 1416 367 1446 619
<< ndiff >>
rect 27 209 84 221
rect 27 175 39 209
rect 73 175 84 209
rect 27 99 84 175
rect 27 65 39 99
rect 73 65 84 99
rect 27 53 84 65
rect 114 209 170 221
rect 114 175 125 209
rect 159 175 170 209
rect 114 101 170 175
rect 114 67 125 101
rect 159 67 170 101
rect 114 53 170 67
rect 200 99 256 221
rect 200 65 211 99
rect 245 65 256 99
rect 200 53 256 65
rect 286 126 342 221
rect 286 92 297 126
rect 331 92 342 126
rect 286 53 342 92
rect 372 99 428 221
rect 372 65 383 99
rect 417 65 428 99
rect 372 53 428 65
rect 458 126 514 221
rect 458 92 469 126
rect 503 92 514 126
rect 458 53 514 92
rect 544 99 600 221
rect 544 65 555 99
rect 589 65 600 99
rect 544 53 600 65
rect 630 126 686 221
rect 630 92 641 126
rect 675 92 686 126
rect 630 53 686 92
rect 716 189 772 221
rect 716 155 727 189
rect 761 155 772 189
rect 716 53 772 155
rect 802 126 858 221
rect 802 92 813 126
rect 847 92 858 126
rect 802 53 858 92
rect 888 189 944 221
rect 888 155 899 189
rect 933 155 944 189
rect 888 53 944 155
rect 974 126 1030 221
rect 974 92 985 126
rect 1019 92 1030 126
rect 974 53 1030 92
rect 1060 189 1116 221
rect 1060 155 1071 189
rect 1105 155 1116 189
rect 1060 53 1116 155
rect 1146 167 1216 221
rect 1146 133 1171 167
rect 1205 133 1216 167
rect 1146 99 1216 133
rect 1146 65 1171 99
rect 1205 65 1216 99
rect 1146 53 1216 65
rect 1246 181 1316 221
rect 1246 147 1271 181
rect 1305 147 1316 181
rect 1246 53 1316 147
rect 1346 209 1416 221
rect 1346 175 1371 209
rect 1405 175 1416 209
rect 1346 101 1416 175
rect 1346 67 1371 101
rect 1405 67 1416 101
rect 1346 53 1416 67
rect 1446 209 1503 221
rect 1446 175 1457 209
rect 1491 175 1503 209
rect 1446 99 1503 175
rect 1446 65 1457 99
rect 1491 65 1503 99
rect 1446 53 1503 65
<< pdiff >>
rect 27 607 84 619
rect 27 573 39 607
rect 73 573 84 607
rect 27 510 84 573
rect 27 476 39 510
rect 73 476 84 510
rect 27 413 84 476
rect 27 379 39 413
rect 73 379 84 413
rect 27 367 84 379
rect 114 599 170 619
rect 114 565 125 599
rect 159 565 170 599
rect 114 519 170 565
rect 114 485 125 519
rect 159 485 170 519
rect 114 440 170 485
rect 114 406 125 440
rect 159 406 170 440
rect 114 367 170 406
rect 200 591 256 619
rect 200 557 211 591
rect 245 557 256 591
rect 200 367 256 557
rect 286 599 342 619
rect 286 565 297 599
rect 331 565 342 599
rect 286 508 342 565
rect 286 474 297 508
rect 331 474 342 508
rect 286 367 342 474
rect 372 591 428 619
rect 372 557 383 591
rect 417 557 428 591
rect 372 367 428 557
rect 458 599 514 619
rect 458 565 469 599
rect 503 565 514 599
rect 458 508 514 565
rect 458 474 469 508
rect 503 474 514 508
rect 458 367 514 474
rect 544 591 628 619
rect 544 557 569 591
rect 603 557 628 591
rect 544 367 628 557
rect 658 599 714 619
rect 658 565 669 599
rect 703 565 714 599
rect 658 508 714 565
rect 658 474 669 508
rect 703 474 714 508
rect 658 367 714 474
rect 744 531 800 619
rect 744 497 755 531
rect 789 497 800 531
rect 744 419 800 497
rect 744 385 755 419
rect 789 385 800 419
rect 744 367 800 385
rect 830 599 886 619
rect 830 565 841 599
rect 875 565 886 599
rect 830 487 886 565
rect 830 453 841 487
rect 875 453 886 487
rect 830 367 886 453
rect 916 531 972 619
rect 916 497 927 531
rect 961 497 972 531
rect 916 419 972 497
rect 916 385 927 419
rect 961 385 972 419
rect 916 367 972 385
rect 1002 599 1058 619
rect 1002 565 1013 599
rect 1047 565 1058 599
rect 1002 487 1058 565
rect 1002 453 1013 487
rect 1047 453 1058 487
rect 1002 367 1058 453
rect 1088 531 1144 619
rect 1088 497 1099 531
rect 1133 497 1144 531
rect 1088 419 1144 497
rect 1088 385 1099 419
rect 1133 385 1144 419
rect 1088 367 1144 385
rect 1174 599 1230 619
rect 1174 565 1185 599
rect 1219 565 1230 599
rect 1174 471 1230 565
rect 1174 437 1185 471
rect 1219 437 1230 471
rect 1174 367 1230 437
rect 1260 531 1330 619
rect 1260 497 1285 531
rect 1319 497 1330 531
rect 1260 419 1330 497
rect 1260 385 1285 419
rect 1319 385 1330 419
rect 1260 367 1330 385
rect 1360 599 1416 619
rect 1360 565 1371 599
rect 1405 565 1416 599
rect 1360 509 1416 565
rect 1360 475 1371 509
rect 1405 475 1416 509
rect 1360 419 1416 475
rect 1360 385 1371 419
rect 1405 385 1416 419
rect 1360 367 1416 385
rect 1446 607 1503 619
rect 1446 573 1457 607
rect 1491 573 1503 607
rect 1446 513 1503 573
rect 1446 479 1457 513
rect 1491 479 1503 513
rect 1446 419 1503 479
rect 1446 385 1457 419
rect 1491 385 1503 419
rect 1446 367 1503 385
<< ndiffc >>
rect 39 175 73 209
rect 39 65 73 99
rect 125 175 159 209
rect 125 67 159 101
rect 211 65 245 99
rect 297 92 331 126
rect 383 65 417 99
rect 469 92 503 126
rect 555 65 589 99
rect 641 92 675 126
rect 727 155 761 189
rect 813 92 847 126
rect 899 155 933 189
rect 985 92 1019 126
rect 1071 155 1105 189
rect 1171 133 1205 167
rect 1171 65 1205 99
rect 1271 147 1305 181
rect 1371 175 1405 209
rect 1371 67 1405 101
rect 1457 175 1491 209
rect 1457 65 1491 99
<< pdiffc >>
rect 39 573 73 607
rect 39 476 73 510
rect 39 379 73 413
rect 125 565 159 599
rect 125 485 159 519
rect 125 406 159 440
rect 211 557 245 591
rect 297 565 331 599
rect 297 474 331 508
rect 383 557 417 591
rect 469 565 503 599
rect 469 474 503 508
rect 569 557 603 591
rect 669 565 703 599
rect 669 474 703 508
rect 755 497 789 531
rect 755 385 789 419
rect 841 565 875 599
rect 841 453 875 487
rect 927 497 961 531
rect 927 385 961 419
rect 1013 565 1047 599
rect 1013 453 1047 487
rect 1099 497 1133 531
rect 1099 385 1133 419
rect 1185 565 1219 599
rect 1185 437 1219 471
rect 1285 497 1319 531
rect 1285 385 1319 419
rect 1371 565 1405 599
rect 1371 475 1405 509
rect 1371 385 1405 419
rect 1457 573 1491 607
rect 1457 479 1491 513
rect 1457 385 1491 419
<< poly >>
rect 84 619 114 645
rect 170 619 200 645
rect 256 619 286 645
rect 342 619 372 645
rect 428 619 458 645
rect 514 619 544 645
rect 628 619 658 645
rect 714 619 744 645
rect 800 619 830 645
rect 886 619 916 645
rect 972 619 1002 645
rect 1058 619 1088 645
rect 1144 619 1174 645
rect 1230 619 1260 645
rect 1330 619 1360 645
rect 1416 619 1446 645
rect 84 335 114 367
rect 170 335 200 367
rect 256 335 286 367
rect 342 335 372 367
rect 428 335 458 367
rect 514 335 544 367
rect 628 335 658 367
rect 714 335 744 367
rect 800 335 830 367
rect 886 335 916 367
rect 972 335 1002 367
rect 1058 335 1088 367
rect 1144 335 1174 367
rect 1230 335 1260 367
rect 1330 335 1360 367
rect 1416 335 1446 367
rect 84 319 1483 335
rect 84 285 277 319
rect 311 285 345 319
rect 379 285 413 319
rect 447 285 481 319
rect 515 285 549 319
rect 583 285 617 319
rect 651 285 685 319
rect 719 285 753 319
rect 787 285 821 319
rect 855 285 889 319
rect 923 285 957 319
rect 991 285 1025 319
rect 1059 285 1093 319
rect 1127 285 1161 319
rect 1195 285 1229 319
rect 1263 285 1297 319
rect 1331 285 1365 319
rect 1399 285 1433 319
rect 1467 285 1483 319
rect 84 269 1483 285
rect 84 221 114 269
rect 170 221 200 269
rect 256 221 286 269
rect 342 221 372 269
rect 428 221 458 269
rect 514 221 544 269
rect 600 221 630 269
rect 686 221 716 269
rect 772 221 802 269
rect 858 221 888 269
rect 944 221 974 269
rect 1030 221 1060 269
rect 1116 221 1146 269
rect 1216 221 1246 269
rect 1316 221 1346 269
rect 1416 221 1446 269
rect 84 27 114 53
rect 170 27 200 53
rect 256 27 286 53
rect 342 27 372 53
rect 428 27 458 53
rect 514 27 544 53
rect 600 27 630 53
rect 686 27 716 53
rect 772 27 802 53
rect 858 27 888 53
rect 944 27 974 53
rect 1030 27 1060 53
rect 1116 27 1146 53
rect 1216 27 1246 53
rect 1316 27 1346 53
rect 1416 27 1446 53
<< polycont >>
rect 277 285 311 319
rect 345 285 379 319
rect 413 285 447 319
rect 481 285 515 319
rect 549 285 583 319
rect 617 285 651 319
rect 685 285 719 319
rect 753 285 787 319
rect 821 285 855 319
rect 889 285 923 319
rect 957 285 991 319
rect 1025 285 1059 319
rect 1093 285 1127 319
rect 1161 285 1195 319
rect 1229 285 1263 319
rect 1297 285 1331 319
rect 1365 285 1399 319
rect 1433 285 1467 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 23 607 73 649
rect 23 573 39 607
rect 23 510 73 573
rect 23 476 39 510
rect 23 413 73 476
rect 23 379 39 413
rect 109 599 159 615
rect 109 565 125 599
rect 109 519 159 565
rect 195 591 261 649
rect 195 557 211 591
rect 245 557 261 591
rect 195 526 261 557
rect 297 599 331 615
rect 109 485 125 519
rect 297 508 331 565
rect 367 591 417 649
rect 367 557 383 591
rect 367 526 417 557
rect 453 599 519 615
rect 453 565 469 599
rect 503 565 519 599
rect 159 485 297 492
rect 109 474 297 485
rect 453 508 519 565
rect 553 591 619 649
rect 553 557 569 591
rect 603 557 619 591
rect 553 526 619 557
rect 653 599 1405 615
rect 653 565 669 599
rect 703 581 841 599
rect 703 565 719 581
rect 453 492 469 508
rect 331 474 469 492
rect 503 492 519 508
rect 653 508 719 565
rect 825 565 841 581
rect 875 581 1013 599
rect 875 565 891 581
rect 653 492 669 508
rect 503 474 669 492
rect 703 474 719 508
rect 109 458 719 474
rect 755 531 789 547
rect 109 440 159 458
rect 109 406 125 440
rect 755 424 789 497
rect 825 487 891 565
rect 997 565 1013 581
rect 1047 581 1185 599
rect 1047 565 1063 581
rect 825 453 841 487
rect 875 453 891 487
rect 825 437 891 453
rect 927 531 961 547
rect 109 390 159 406
rect 193 419 789 424
rect 193 390 755 419
rect 23 363 73 379
rect 193 356 227 390
rect 927 419 961 497
rect 997 487 1063 565
rect 1169 565 1185 581
rect 1219 581 1371 599
rect 1219 565 1235 581
rect 997 453 1013 487
rect 1047 453 1063 487
rect 997 437 1063 453
rect 1099 531 1133 547
rect 789 385 927 403
rect 1099 419 1133 497
rect 1169 471 1235 565
rect 1169 437 1185 471
rect 1219 437 1235 471
rect 1269 531 1335 547
rect 1269 497 1285 531
rect 1319 497 1335 531
rect 961 385 1099 403
rect 1269 419 1335 497
rect 1269 403 1285 419
rect 1133 385 1285 403
rect 1319 385 1335 419
rect 755 369 1335 385
rect 1371 509 1405 565
rect 1371 419 1405 475
rect 1371 369 1405 385
rect 1441 607 1507 649
rect 1441 573 1457 607
rect 1491 573 1507 607
rect 1441 513 1507 573
rect 1441 479 1457 513
rect 1491 479 1507 513
rect 1441 419 1507 479
rect 1441 385 1457 419
rect 1491 385 1507 419
rect 1441 369 1507 385
rect 121 310 227 356
rect 313 335 647 356
rect 193 235 227 310
rect 261 319 1483 335
rect 261 285 277 319
rect 311 285 345 319
rect 379 285 413 319
rect 447 285 481 319
rect 515 285 549 319
rect 583 285 617 319
rect 651 285 685 319
rect 719 285 753 319
rect 787 285 821 319
rect 855 285 889 319
rect 923 285 957 319
rect 991 285 1025 319
rect 1059 285 1093 319
rect 1127 285 1161 319
rect 1195 285 1229 319
rect 1263 285 1297 319
rect 1331 285 1365 319
rect 1399 285 1433 319
rect 1467 285 1483 319
rect 261 269 1483 285
rect 23 209 73 225
rect 23 175 39 209
rect 23 99 73 175
rect 23 65 39 99
rect 23 17 73 65
rect 109 209 159 225
rect 109 175 125 209
rect 193 201 1321 235
rect 109 167 159 175
rect 711 189 761 201
rect 109 133 675 167
rect 109 101 159 133
rect 109 67 125 101
rect 297 126 331 133
rect 109 51 159 67
rect 195 65 211 99
rect 245 65 261 99
rect 195 17 261 65
rect 469 126 503 133
rect 297 51 331 92
rect 367 65 383 99
rect 417 65 433 99
rect 367 17 433 65
rect 641 126 675 133
rect 469 51 503 92
rect 539 65 555 99
rect 589 65 605 99
rect 539 17 605 65
rect 711 155 727 189
rect 899 189 949 201
rect 711 119 761 155
rect 797 126 863 167
rect 641 85 675 92
rect 797 92 813 126
rect 847 92 863 126
rect 933 155 949 189
rect 1055 189 1121 201
rect 899 119 949 155
rect 985 126 1019 167
rect 797 85 863 92
rect 1055 155 1071 189
rect 1105 155 1121 189
rect 1255 181 1321 201
rect 1055 119 1121 155
rect 1155 133 1171 167
rect 1205 133 1221 167
rect 985 85 1019 92
rect 1155 99 1221 133
rect 1255 147 1271 181
rect 1305 147 1321 181
rect 1255 119 1321 147
rect 1355 209 1421 225
rect 1355 175 1371 209
rect 1405 175 1421 209
rect 1155 85 1171 99
rect 641 65 1171 85
rect 1205 85 1221 99
rect 1355 101 1421 175
rect 1355 85 1371 101
rect 1205 67 1371 85
rect 1405 67 1421 101
rect 1205 65 1421 67
rect 641 51 1421 65
rect 1457 209 1507 225
rect 1491 175 1507 209
rect 1457 99 1507 175
rect 1491 65 1507 99
rect 1457 17 1507 65
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 invlp_8
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6835994
string GDS_START 6824630
<< end >>
