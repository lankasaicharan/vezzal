magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 205 175 855 259
rect 100 49 855 175
rect 0 0 864 49
<< scnmos >>
rect 179 65 209 149
rect 284 65 314 233
rect 370 65 400 233
rect 472 65 502 233
rect 558 65 588 233
rect 660 65 690 233
rect 746 65 776 233
<< scpmoshvt >>
rect 89 500 119 584
rect 284 367 314 619
rect 370 367 400 619
rect 456 367 486 619
rect 574 367 604 619
rect 660 367 690 619
rect 746 367 776 619
<< ndiff >>
rect 231 218 284 233
rect 231 184 239 218
rect 273 184 284 218
rect 231 149 284 184
rect 126 124 179 149
rect 126 90 134 124
rect 168 90 179 124
rect 126 65 179 90
rect 209 111 284 149
rect 209 77 229 111
rect 263 77 284 111
rect 209 65 284 77
rect 314 212 370 233
rect 314 178 325 212
rect 359 178 370 212
rect 314 107 370 178
rect 314 73 325 107
rect 359 73 370 107
rect 314 65 370 73
rect 400 181 472 233
rect 400 147 411 181
rect 445 147 472 181
rect 400 107 472 147
rect 400 73 411 107
rect 445 73 472 107
rect 400 65 472 73
rect 502 181 558 233
rect 502 147 513 181
rect 547 147 558 181
rect 502 107 558 147
rect 502 73 513 107
rect 547 73 558 107
rect 502 65 558 73
rect 588 225 660 233
rect 588 191 615 225
rect 649 191 660 225
rect 588 155 660 191
rect 588 121 615 155
rect 649 121 660 155
rect 588 65 660 121
rect 690 221 746 233
rect 690 187 701 221
rect 735 187 746 221
rect 690 111 746 187
rect 690 77 701 111
rect 735 77 746 111
rect 690 65 746 77
rect 776 221 829 233
rect 776 187 787 221
rect 821 187 829 221
rect 776 111 829 187
rect 776 77 787 111
rect 821 77 829 111
rect 776 65 829 77
<< pdiff >>
rect 231 599 284 619
rect 36 570 89 584
rect 36 536 44 570
rect 78 536 89 570
rect 36 500 89 536
rect 119 559 172 584
rect 119 525 130 559
rect 164 525 172 559
rect 119 500 172 525
rect 231 565 239 599
rect 273 565 284 599
rect 231 507 284 565
rect 231 473 239 507
rect 273 473 284 507
rect 231 416 284 473
rect 231 382 239 416
rect 273 382 284 416
rect 231 367 284 382
rect 314 546 370 619
rect 314 512 325 546
rect 359 512 370 546
rect 314 478 370 512
rect 314 444 325 478
rect 359 444 370 478
rect 314 409 370 444
rect 314 375 325 409
rect 359 375 370 409
rect 314 367 370 375
rect 400 599 456 619
rect 400 565 411 599
rect 445 565 456 599
rect 400 507 456 565
rect 400 473 411 507
rect 445 473 456 507
rect 400 416 456 473
rect 400 382 411 416
rect 445 382 456 416
rect 400 367 456 382
rect 486 573 574 619
rect 486 539 513 573
rect 547 539 574 573
rect 486 367 574 539
rect 604 578 660 619
rect 604 544 615 578
rect 649 544 660 578
rect 604 492 660 544
rect 604 458 615 492
rect 649 458 660 492
rect 604 367 660 458
rect 690 570 746 619
rect 690 536 701 570
rect 735 536 746 570
rect 690 367 746 536
rect 776 599 829 619
rect 776 565 787 599
rect 821 565 829 599
rect 776 507 829 565
rect 776 473 787 507
rect 821 473 829 507
rect 776 413 829 473
rect 776 379 787 413
rect 821 379 829 413
rect 776 367 829 379
<< ndiffc >>
rect 239 184 273 218
rect 134 90 168 124
rect 229 77 263 111
rect 325 178 359 212
rect 325 73 359 107
rect 411 147 445 181
rect 411 73 445 107
rect 513 147 547 181
rect 513 73 547 107
rect 615 191 649 225
rect 615 121 649 155
rect 701 187 735 221
rect 701 77 735 111
rect 787 187 821 221
rect 787 77 821 111
<< pdiffc >>
rect 44 536 78 570
rect 130 525 164 559
rect 239 565 273 599
rect 239 473 273 507
rect 239 382 273 416
rect 325 512 359 546
rect 325 444 359 478
rect 325 375 359 409
rect 411 565 445 599
rect 411 473 445 507
rect 411 382 445 416
rect 513 539 547 573
rect 615 544 649 578
rect 615 458 649 492
rect 701 536 735 570
rect 787 565 821 599
rect 787 473 821 507
rect 787 379 821 413
<< poly >>
rect 284 619 314 645
rect 370 619 400 645
rect 456 619 486 645
rect 574 619 604 645
rect 660 619 690 645
rect 746 619 776 645
rect 89 584 119 610
rect 89 305 119 500
rect 44 289 119 305
rect 44 255 60 289
rect 94 255 119 289
rect 167 305 233 321
rect 167 271 183 305
rect 217 285 233 305
rect 284 285 314 367
rect 370 285 400 367
rect 456 335 486 367
rect 574 335 604 367
rect 660 335 690 367
rect 217 271 400 285
rect 167 255 400 271
rect 450 319 516 335
rect 450 285 466 319
rect 500 285 516 319
rect 450 269 516 285
rect 558 319 690 335
rect 558 285 574 319
rect 608 285 690 319
rect 558 269 690 285
rect 44 221 119 255
rect 284 233 314 255
rect 370 233 400 255
rect 472 233 502 269
rect 558 233 588 269
rect 660 233 690 269
rect 746 335 776 367
rect 746 319 812 335
rect 746 285 762 319
rect 796 285 812 319
rect 746 269 812 285
rect 746 233 776 269
rect 44 187 60 221
rect 94 201 119 221
rect 94 187 209 201
rect 44 171 209 187
rect 179 149 209 171
rect 179 39 209 65
rect 284 39 314 65
rect 370 39 400 65
rect 472 39 502 65
rect 558 39 588 65
rect 660 39 690 65
rect 746 39 776 65
<< polycont >>
rect 60 255 94 289
rect 183 271 217 305
rect 466 285 500 319
rect 574 285 608 319
rect 762 285 796 319
rect 60 187 94 221
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 28 570 94 649
rect 223 599 463 615
rect 28 536 44 570
rect 78 536 94 570
rect 28 532 94 536
rect 128 559 180 575
rect 128 525 130 559
rect 164 525 180 559
rect 17 289 94 498
rect 17 255 60 289
rect 17 221 94 255
rect 17 187 60 221
rect 17 64 94 187
rect 128 321 180 525
rect 223 565 239 599
rect 273 581 411 599
rect 273 565 275 581
rect 223 507 275 565
rect 409 565 411 581
rect 445 565 463 599
rect 223 473 239 507
rect 273 473 275 507
rect 223 416 275 473
rect 223 382 239 416
rect 273 382 275 416
rect 223 366 275 382
rect 309 512 325 546
rect 359 512 375 546
rect 309 478 375 512
rect 309 444 325 478
rect 359 444 375 478
rect 309 409 375 444
rect 309 375 325 409
rect 359 375 375 409
rect 309 364 375 375
rect 409 507 463 565
rect 497 573 563 649
rect 497 539 513 573
rect 547 539 563 573
rect 497 528 563 539
rect 597 578 651 594
rect 597 544 615 578
rect 649 544 651 578
rect 409 473 411 507
rect 445 492 463 507
rect 597 492 651 544
rect 685 570 751 649
rect 685 536 701 570
rect 735 536 751 570
rect 685 526 751 536
rect 785 599 837 615
rect 785 565 787 599
rect 821 565 837 599
rect 785 507 837 565
rect 785 492 787 507
rect 445 473 615 492
rect 409 458 615 473
rect 649 473 787 492
rect 821 473 837 507
rect 649 458 837 473
rect 409 416 449 458
rect 409 382 411 416
rect 445 382 449 416
rect 409 366 449 382
rect 485 385 749 424
rect 128 305 233 321
rect 128 271 183 305
rect 217 271 233 305
rect 128 268 233 271
rect 128 124 184 268
rect 309 249 359 364
rect 485 319 519 385
rect 450 285 466 319
rect 500 285 519 319
rect 558 319 663 350
rect 558 285 574 319
rect 608 285 663 319
rect 703 329 749 385
rect 783 413 837 458
rect 783 379 787 413
rect 821 379 837 413
rect 783 363 837 379
rect 703 319 812 329
rect 703 285 762 319
rect 796 285 812 319
rect 703 271 812 285
rect 128 90 134 124
rect 168 90 184 124
rect 128 74 184 90
rect 223 218 275 234
rect 223 184 239 218
rect 273 184 275 218
rect 223 111 275 184
rect 223 77 229 111
rect 263 77 275 111
rect 223 17 275 77
rect 309 225 665 249
rect 309 215 615 225
rect 309 212 361 215
rect 309 178 325 212
rect 359 178 361 212
rect 599 191 615 215
rect 649 191 665 225
rect 309 107 361 178
rect 309 73 325 107
rect 359 73 361 107
rect 309 57 361 73
rect 395 147 411 181
rect 445 147 461 181
rect 395 107 461 147
rect 395 73 411 107
rect 445 73 461 107
rect 395 17 461 73
rect 497 147 513 181
rect 547 147 563 181
rect 497 107 563 147
rect 599 155 665 191
rect 599 121 615 155
rect 649 121 665 155
rect 699 221 744 237
rect 699 187 701 221
rect 735 187 744 221
rect 497 73 513 107
rect 547 87 563 107
rect 699 111 744 187
rect 699 87 701 111
rect 547 77 701 87
rect 735 77 744 111
rect 547 73 744 77
rect 497 53 744 73
rect 778 221 837 237
rect 778 187 787 221
rect 821 187 837 221
rect 778 111 837 187
rect 778 77 787 111
rect 821 77 837 111
rect 778 17 837 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21boi_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5543476
string GDS_START 5534586
<< end >>
