magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 57 49 669 157
rect 0 0 672 49
<< scnmos >>
rect 140 47 170 131
rect 218 47 248 131
rect 296 47 326 131
rect 398 47 428 131
rect 484 47 514 131
rect 556 47 586 131
<< scpmoshvt >>
rect 84 409 134 609
rect 190 409 240 609
rect 296 409 346 609
rect 406 409 456 609
rect 512 409 562 609
<< ndiff >>
rect 83 101 140 131
rect 83 67 95 101
rect 129 67 140 101
rect 83 47 140 67
rect 170 47 218 131
rect 248 47 296 131
rect 326 47 398 131
rect 428 111 484 131
rect 428 77 439 111
rect 473 77 484 111
rect 428 47 484 77
rect 514 47 556 131
rect 586 97 643 131
rect 586 63 597 97
rect 631 63 643 97
rect 586 47 643 63
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 190 609
rect 134 563 145 597
rect 179 563 190 597
rect 134 514 190 563
rect 134 480 145 514
rect 179 480 190 514
rect 134 409 190 480
rect 240 597 296 609
rect 240 563 251 597
rect 285 563 296 597
rect 240 526 296 563
rect 240 492 251 526
rect 285 492 296 526
rect 240 455 296 492
rect 240 421 251 455
rect 285 421 296 455
rect 240 409 296 421
rect 346 597 406 609
rect 346 563 357 597
rect 391 563 406 597
rect 346 514 406 563
rect 346 480 357 514
rect 391 480 406 514
rect 346 409 406 480
rect 456 597 512 609
rect 456 563 467 597
rect 501 563 512 597
rect 456 526 512 563
rect 456 492 467 526
rect 501 492 512 526
rect 456 455 512 492
rect 456 421 467 455
rect 501 421 512 455
rect 456 409 512 421
rect 562 597 619 609
rect 562 563 573 597
rect 607 563 619 597
rect 562 526 619 563
rect 562 492 573 526
rect 607 492 619 526
rect 562 455 619 492
rect 562 421 573 455
rect 607 421 619 455
rect 562 409 619 421
<< ndiffc >>
rect 95 67 129 101
rect 439 77 473 111
rect 597 63 631 97
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 480 179 514
rect 251 563 285 597
rect 251 492 285 526
rect 251 421 285 455
rect 357 563 391 597
rect 357 480 391 514
rect 467 563 501 597
rect 467 492 501 526
rect 467 421 501 455
rect 573 563 607 597
rect 573 492 607 526
rect 573 421 607 455
<< poly >>
rect 84 609 134 635
rect 190 609 240 635
rect 296 609 346 635
rect 406 609 456 635
rect 512 609 562 635
rect 84 228 134 409
rect 190 356 240 409
rect 296 358 346 409
rect 406 358 456 409
rect 512 358 562 409
rect 182 340 248 356
rect 182 306 198 340
rect 232 306 248 340
rect 182 290 248 306
rect 84 212 170 228
rect 84 178 100 212
rect 134 178 170 212
rect 84 162 170 178
rect 140 131 170 162
rect 218 131 248 290
rect 290 342 356 358
rect 290 308 306 342
rect 340 308 356 342
rect 290 274 356 308
rect 290 240 306 274
rect 340 240 356 274
rect 290 224 356 240
rect 398 342 464 358
rect 398 308 414 342
rect 448 308 464 342
rect 398 274 464 308
rect 398 240 414 274
rect 448 240 464 274
rect 398 224 464 240
rect 512 342 586 358
rect 512 308 528 342
rect 562 308 586 342
rect 512 274 586 308
rect 512 240 528 274
rect 562 240 586 274
rect 512 224 586 240
rect 296 131 326 224
rect 398 131 428 224
rect 556 176 586 224
rect 484 146 586 176
rect 484 131 514 146
rect 556 131 586 146
rect 140 21 170 47
rect 218 21 248 47
rect 296 21 326 47
rect 398 21 428 47
rect 484 21 514 47
rect 556 21 586 47
<< polycont >>
rect 198 306 232 340
rect 100 178 134 212
rect 306 308 340 342
rect 306 240 340 274
rect 414 308 448 342
rect 414 240 448 274
rect 528 308 562 342
rect 528 240 562 274
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 526 89 563
rect 23 492 39 526
rect 73 492 89 526
rect 23 455 89 492
rect 129 597 195 649
rect 129 563 145 597
rect 179 563 195 597
rect 129 514 195 563
rect 129 480 145 514
rect 179 480 195 514
rect 129 464 195 480
rect 235 597 301 613
rect 235 563 251 597
rect 285 563 301 597
rect 235 526 301 563
rect 235 492 251 526
rect 285 492 301 526
rect 23 421 39 455
rect 73 428 89 455
rect 235 455 301 492
rect 341 597 407 649
rect 341 563 357 597
rect 391 563 407 597
rect 341 514 407 563
rect 341 480 357 514
rect 391 480 407 514
rect 341 464 407 480
rect 451 597 517 613
rect 451 563 467 597
rect 501 563 517 597
rect 451 526 517 563
rect 451 492 467 526
rect 501 492 517 526
rect 235 428 251 455
rect 73 421 251 428
rect 285 428 301 455
rect 451 455 517 492
rect 451 428 467 455
rect 285 421 467 428
rect 501 421 517 455
rect 23 394 517 421
rect 557 597 648 613
rect 557 563 573 597
rect 607 563 648 597
rect 557 526 648 563
rect 557 492 573 526
rect 607 492 648 526
rect 557 455 648 492
rect 557 421 573 455
rect 607 421 648 455
rect 557 405 648 421
rect 25 340 248 356
rect 25 306 198 340
rect 232 306 248 340
rect 25 290 248 306
rect 290 342 359 358
rect 290 308 306 342
rect 340 308 359 342
rect 290 274 359 308
rect 290 240 306 274
rect 340 240 359 274
rect 25 212 167 228
rect 25 178 100 212
rect 134 178 167 212
rect 25 162 167 178
rect 79 101 145 126
rect 79 67 95 101
rect 129 67 145 101
rect 290 88 359 240
rect 398 342 464 358
rect 398 308 414 342
rect 448 308 464 342
rect 398 274 464 308
rect 398 240 414 274
rect 448 240 464 274
rect 398 224 464 240
rect 505 342 578 358
rect 505 308 528 342
rect 562 308 578 342
rect 505 274 578 308
rect 505 240 528 274
rect 562 240 578 274
rect 505 224 578 240
rect 614 188 648 405
rect 409 154 648 188
rect 409 111 489 154
rect 79 17 145 67
rect 409 77 439 111
rect 473 77 489 111
rect 409 53 489 77
rect 581 97 647 118
rect 581 63 597 97
rect 631 63 647 97
rect 581 17 647 63
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a41oi_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1346408
string GDS_START 1339252
<< end >>
