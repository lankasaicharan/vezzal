magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 42 49 845 241
rect 0 0 864 49
<< scnmos >>
rect 121 47 151 215
rect 306 47 336 215
rect 448 47 478 215
rect 520 47 550 215
rect 628 47 658 215
rect 736 47 766 215
<< scpmoshvt >>
rect 113 367 143 619
rect 316 367 346 619
rect 402 367 432 619
rect 556 367 586 619
rect 642 367 672 619
rect 736 367 766 619
<< ndiff >>
rect 68 203 121 215
rect 68 169 76 203
rect 110 169 121 203
rect 68 101 121 169
rect 68 67 76 101
rect 110 67 121 101
rect 68 47 121 67
rect 151 132 306 215
rect 151 98 166 132
rect 200 98 261 132
rect 295 98 306 132
rect 151 47 306 98
rect 336 190 448 215
rect 336 156 347 190
rect 381 156 448 190
rect 336 101 448 156
rect 336 67 347 101
rect 381 67 448 101
rect 336 47 448 67
rect 478 47 520 215
rect 550 47 628 215
rect 658 47 736 215
rect 766 187 819 215
rect 766 153 777 187
rect 811 153 819 187
rect 766 93 819 153
rect 766 59 777 93
rect 811 59 819 93
rect 766 47 819 59
<< pdiff >>
rect 60 599 113 619
rect 60 565 68 599
rect 102 565 113 599
rect 60 507 113 565
rect 60 473 68 507
rect 102 473 113 507
rect 60 413 113 473
rect 60 379 68 413
rect 102 379 113 413
rect 60 367 113 379
rect 143 607 196 619
rect 143 573 154 607
rect 188 573 196 607
rect 143 520 196 573
rect 143 486 154 520
rect 188 486 196 520
rect 143 439 196 486
rect 143 405 154 439
rect 188 405 196 439
rect 143 367 196 405
rect 263 599 316 619
rect 263 565 271 599
rect 305 565 316 599
rect 263 510 316 565
rect 263 476 271 510
rect 305 476 316 510
rect 263 413 316 476
rect 263 379 271 413
rect 305 379 316 413
rect 263 367 316 379
rect 346 599 402 619
rect 346 565 357 599
rect 391 565 402 599
rect 346 510 402 565
rect 346 476 357 510
rect 391 476 402 510
rect 346 413 402 476
rect 346 379 357 413
rect 391 379 402 413
rect 346 367 402 379
rect 432 607 556 619
rect 432 573 443 607
rect 477 573 511 607
rect 545 573 556 607
rect 432 524 556 573
rect 432 490 443 524
rect 477 490 511 524
rect 545 490 556 524
rect 432 439 556 490
rect 432 405 443 439
rect 477 405 511 439
rect 545 405 556 439
rect 432 367 556 405
rect 586 599 642 619
rect 586 565 597 599
rect 631 565 642 599
rect 586 510 642 565
rect 586 476 597 510
rect 631 476 642 510
rect 586 413 642 476
rect 586 379 597 413
rect 631 379 642 413
rect 586 367 642 379
rect 672 607 736 619
rect 672 573 687 607
rect 721 573 736 607
rect 672 523 736 573
rect 672 489 687 523
rect 721 489 736 523
rect 672 439 736 489
rect 672 405 687 439
rect 721 405 736 439
rect 672 367 736 405
rect 766 599 819 619
rect 766 565 777 599
rect 811 565 819 599
rect 766 511 819 565
rect 766 477 777 511
rect 811 477 819 511
rect 766 413 819 477
rect 766 379 777 413
rect 811 379 819 413
rect 766 367 819 379
<< ndiffc >>
rect 76 169 110 203
rect 76 67 110 101
rect 166 98 200 132
rect 261 98 295 132
rect 347 156 381 190
rect 347 67 381 101
rect 777 153 811 187
rect 777 59 811 93
<< pdiffc >>
rect 68 565 102 599
rect 68 473 102 507
rect 68 379 102 413
rect 154 573 188 607
rect 154 486 188 520
rect 154 405 188 439
rect 271 565 305 599
rect 271 476 305 510
rect 271 379 305 413
rect 357 565 391 599
rect 357 476 391 510
rect 357 379 391 413
rect 443 573 477 607
rect 511 573 545 607
rect 443 490 477 524
rect 511 490 545 524
rect 443 405 477 439
rect 511 405 545 439
rect 597 565 631 599
rect 597 476 631 510
rect 597 379 631 413
rect 687 573 721 607
rect 687 489 721 523
rect 687 405 721 439
rect 777 565 811 599
rect 777 477 811 511
rect 777 379 811 413
<< poly >>
rect 113 619 143 645
rect 316 619 346 645
rect 402 619 432 645
rect 556 619 586 645
rect 642 619 672 645
rect 736 619 766 645
rect 113 303 143 367
rect 316 303 346 367
rect 402 309 432 367
rect 113 287 200 303
rect 113 253 150 287
rect 184 253 200 287
rect 113 237 200 253
rect 254 287 360 303
rect 254 253 310 287
rect 344 253 360 287
rect 254 237 360 253
rect 402 287 478 309
rect 556 303 586 367
rect 642 303 672 367
rect 736 303 766 367
rect 402 253 428 287
rect 462 253 478 287
rect 402 237 478 253
rect 121 215 151 237
rect 306 215 336 237
rect 448 215 478 237
rect 520 287 586 303
rect 520 253 536 287
rect 570 253 586 287
rect 520 237 586 253
rect 628 287 694 303
rect 628 253 644 287
rect 678 253 694 287
rect 628 237 694 253
rect 736 287 823 303
rect 736 253 773 287
rect 807 253 823 287
rect 736 237 823 253
rect 520 215 550 237
rect 628 215 658 237
rect 736 215 766 237
rect 121 21 151 47
rect 306 21 336 47
rect 448 21 478 47
rect 520 21 550 47
rect 628 21 658 47
rect 736 21 766 47
<< polycont >>
rect 150 253 184 287
rect 310 253 344 287
rect 428 253 462 287
rect 536 253 570 287
rect 644 253 678 287
rect 773 253 807 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 17 599 114 615
rect 17 565 68 599
rect 102 565 114 599
rect 17 507 114 565
rect 17 473 68 507
rect 102 473 114 507
rect 17 413 114 473
rect 17 379 68 413
rect 102 379 114 413
rect 150 607 204 649
rect 150 573 154 607
rect 188 573 204 607
rect 150 520 204 573
rect 150 486 154 520
rect 188 486 204 520
rect 150 439 204 486
rect 150 405 154 439
rect 188 405 204 439
rect 150 389 204 405
rect 255 599 314 615
rect 255 565 271 599
rect 305 565 314 599
rect 255 510 314 565
rect 255 476 271 510
rect 305 476 314 510
rect 255 413 314 476
rect 17 203 114 379
rect 255 379 271 413
rect 305 379 314 413
rect 255 355 314 379
rect 17 169 76 203
rect 110 169 114 203
rect 148 321 314 355
rect 348 599 393 615
rect 348 565 357 599
rect 391 565 393 599
rect 348 510 393 565
rect 348 476 357 510
rect 391 476 393 510
rect 348 413 393 476
rect 348 379 357 413
rect 391 379 393 413
rect 427 607 561 649
rect 427 573 443 607
rect 477 573 511 607
rect 545 573 561 607
rect 427 524 561 573
rect 427 490 443 524
rect 477 490 511 524
rect 545 490 561 524
rect 427 439 561 490
rect 427 405 443 439
rect 477 405 511 439
rect 545 405 561 439
rect 595 599 637 615
rect 595 565 597 599
rect 631 565 637 599
rect 595 510 637 565
rect 595 476 597 510
rect 631 476 637 510
rect 595 413 637 476
rect 348 371 393 379
rect 595 379 597 413
rect 631 379 637 413
rect 671 607 737 649
rect 671 573 687 607
rect 721 573 737 607
rect 671 523 737 573
rect 671 489 687 523
rect 721 489 737 523
rect 671 439 737 489
rect 671 405 687 439
rect 721 405 737 439
rect 771 599 827 615
rect 771 565 777 599
rect 811 565 827 599
rect 771 511 827 565
rect 771 477 777 511
rect 811 477 827 511
rect 771 413 827 477
rect 595 371 637 379
rect 771 379 777 413
rect 811 379 827 413
rect 771 371 827 379
rect 348 337 827 371
rect 148 287 189 321
rect 415 287 469 303
rect 148 253 150 287
rect 184 253 189 287
rect 148 208 189 253
rect 223 253 310 287
rect 344 253 381 287
rect 223 242 381 253
rect 415 253 428 287
rect 462 253 469 287
rect 148 190 381 208
rect 148 174 347 190
rect 17 101 114 169
rect 345 156 347 174
rect 17 67 76 101
rect 110 67 114 101
rect 17 51 114 67
rect 150 132 311 140
rect 150 98 166 132
rect 200 98 261 132
rect 295 98 311 132
rect 150 17 311 98
rect 345 101 381 156
rect 345 67 347 101
rect 415 78 469 253
rect 503 287 570 303
rect 503 253 536 287
rect 503 78 570 253
rect 604 287 737 303
rect 604 253 644 287
rect 678 253 737 287
rect 604 78 737 253
rect 771 287 847 303
rect 771 253 773 287
rect 807 253 847 287
rect 771 237 847 253
rect 771 187 827 203
rect 771 153 777 187
rect 811 153 827 187
rect 771 93 827 153
rect 345 51 381 67
rect 771 59 777 93
rect 811 59 827 93
rect 771 17 827 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a41o_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5528146
string GDS_START 5518658
<< end >>
