magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 1 228 483 248
rect 1 49 856 228
rect 0 0 864 49
<< scnmos >>
rect 84 74 114 222
rect 170 74 200 222
rect 283 74 313 222
rect 370 74 400 222
rect 629 74 659 202
rect 743 74 773 202
<< scpmoshvt >>
rect 92 368 122 592
rect 192 368 222 592
rect 292 368 322 592
rect 416 368 446 592
rect 618 368 648 568
rect 748 368 778 568
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 173 170 222
rect 114 139 125 173
rect 159 139 170 173
rect 114 74 170 139
rect 200 210 283 222
rect 200 176 225 210
rect 259 176 283 210
rect 200 120 283 176
rect 200 86 225 120
rect 259 86 283 120
rect 200 74 283 86
rect 313 142 370 222
rect 313 108 325 142
rect 359 108 370 142
rect 313 74 370 108
rect 400 210 457 222
rect 400 176 411 210
rect 445 176 457 210
rect 400 120 457 176
rect 400 86 411 120
rect 445 86 457 120
rect 400 74 457 86
rect 572 190 629 202
rect 572 156 584 190
rect 618 156 629 190
rect 572 120 629 156
rect 572 86 584 120
rect 618 86 629 120
rect 572 74 629 86
rect 659 190 743 202
rect 659 156 684 190
rect 718 156 743 190
rect 659 120 743 156
rect 659 86 684 120
rect 718 86 743 120
rect 659 74 743 86
rect 773 190 830 202
rect 773 156 784 190
rect 818 156 830 190
rect 773 120 830 156
rect 773 86 784 120
rect 818 86 830 120
rect 773 74 830 86
<< pdiff >>
rect 340 618 398 630
rect 340 592 352 618
rect 33 580 92 592
rect 33 546 45 580
rect 79 546 92 580
rect 33 468 92 546
rect 33 434 45 468
rect 79 434 92 468
rect 33 368 92 434
rect 122 547 192 592
rect 122 513 145 547
rect 179 513 192 547
rect 122 479 192 513
rect 122 445 145 479
rect 179 445 192 479
rect 122 411 192 445
rect 122 377 145 411
rect 179 377 192 411
rect 122 368 192 377
rect 222 584 292 592
rect 222 550 245 584
rect 279 550 292 584
rect 222 505 292 550
rect 222 471 245 505
rect 279 471 292 505
rect 222 368 292 471
rect 322 584 352 592
rect 386 592 398 618
rect 386 584 416 592
rect 322 368 416 584
rect 446 573 505 592
rect 446 539 459 573
rect 493 539 505 573
rect 446 368 505 539
rect 559 414 618 568
rect 559 380 571 414
rect 605 380 618 414
rect 559 368 618 380
rect 648 556 748 568
rect 648 522 676 556
rect 710 522 748 556
rect 648 368 748 522
rect 778 560 837 568
rect 778 526 791 560
rect 825 526 837 560
rect 778 492 837 526
rect 778 458 791 492
rect 825 458 837 492
rect 778 424 837 458
rect 778 390 791 424
rect 825 390 837 424
rect 778 368 837 390
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 139 159 173
rect 225 176 259 210
rect 225 86 259 120
rect 325 108 359 142
rect 411 176 445 210
rect 411 86 445 120
rect 584 156 618 190
rect 584 86 618 120
rect 684 156 718 190
rect 684 86 718 120
rect 784 156 818 190
rect 784 86 818 120
<< pdiffc >>
rect 45 546 79 580
rect 45 434 79 468
rect 145 513 179 547
rect 145 445 179 479
rect 145 377 179 411
rect 245 550 279 584
rect 245 471 279 505
rect 352 584 386 618
rect 459 539 493 573
rect 571 380 605 414
rect 676 522 710 556
rect 791 526 825 560
rect 791 458 825 492
rect 791 390 825 424
<< poly >>
rect 92 592 122 618
rect 192 592 222 618
rect 292 592 322 618
rect 416 592 446 618
rect 618 568 648 594
rect 748 568 778 594
rect 92 353 122 368
rect 192 353 222 368
rect 292 353 322 368
rect 416 353 446 368
rect 618 353 648 368
rect 748 353 778 368
rect 89 326 125 353
rect 189 326 225 353
rect 289 345 325 353
rect 413 345 449 353
rect 615 345 651 353
rect 89 310 241 326
rect 289 315 659 345
rect 745 336 781 353
rect 89 290 191 310
rect 84 276 191 290
rect 225 276 241 310
rect 84 260 241 276
rect 593 314 659 315
rect 593 280 609 314
rect 643 280 659 314
rect 84 222 114 260
rect 170 222 200 260
rect 283 251 545 267
rect 593 264 659 280
rect 707 320 781 336
rect 707 286 723 320
rect 757 286 781 320
rect 707 270 781 286
rect 283 237 495 251
rect 283 222 313 237
rect 370 222 400 237
rect 479 217 495 237
rect 529 217 545 251
rect 479 183 545 217
rect 629 202 659 264
rect 743 202 773 270
rect 479 149 495 183
rect 529 149 545 183
rect 479 115 545 149
rect 479 81 495 115
rect 529 81 545 115
rect 84 48 114 74
rect 170 48 200 74
rect 283 48 313 74
rect 370 48 400 74
rect 479 65 545 81
rect 629 48 659 74
rect 743 48 773 74
<< polycont >>
rect 191 276 225 310
rect 609 280 643 314
rect 723 286 757 320
rect 495 217 529 251
rect 495 149 529 183
rect 495 81 529 115
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 336 618 402 649
rect 29 584 295 615
rect 336 584 352 618
rect 386 584 402 618
rect 29 581 245 584
rect 29 580 95 581
rect 29 546 45 580
rect 79 546 95 580
rect 229 550 245 581
rect 279 550 295 584
rect 443 573 509 596
rect 443 550 459 573
rect 29 468 95 546
rect 29 434 45 468
rect 79 434 95 468
rect 29 428 95 434
rect 129 513 145 547
rect 179 513 195 547
rect 129 479 195 513
rect 129 445 145 479
rect 179 445 195 479
rect 229 539 459 550
rect 493 539 509 573
rect 229 516 509 539
rect 645 556 741 649
rect 645 522 676 556
rect 710 522 741 556
rect 775 560 841 572
rect 775 526 791 560
rect 825 526 841 560
rect 229 505 295 516
rect 229 471 245 505
rect 279 471 295 505
rect 775 492 841 526
rect 775 482 791 492
rect 229 464 295 471
rect 129 430 195 445
rect 393 458 791 482
rect 825 458 841 492
rect 393 448 841 458
rect 129 411 359 430
rect 129 394 145 411
rect 107 377 145 394
rect 179 377 359 411
rect 107 360 359 377
rect 107 226 141 360
rect 393 326 427 448
rect 775 424 841 448
rect 175 310 427 326
rect 175 276 191 310
rect 225 276 427 310
rect 175 260 427 276
rect 479 380 571 414
rect 605 380 621 414
rect 775 390 791 424
rect 825 390 841 424
rect 479 364 621 380
rect 479 251 545 364
rect 23 210 73 226
rect 23 176 39 210
rect 23 120 73 176
rect 107 173 175 226
rect 107 139 125 173
rect 159 139 175 173
rect 107 123 175 139
rect 209 210 445 226
rect 209 176 225 210
rect 259 192 411 210
rect 259 176 275 192
rect 23 86 39 120
rect 23 85 73 86
rect 209 120 275 176
rect 395 176 411 192
rect 209 86 225 120
rect 259 86 275 120
rect 209 85 275 86
rect 23 51 275 85
rect 309 142 359 158
rect 309 108 325 142
rect 309 17 359 108
rect 395 120 445 176
rect 395 86 411 120
rect 395 70 445 86
rect 479 217 495 251
rect 529 217 545 251
rect 593 314 659 330
rect 593 280 609 314
rect 643 280 659 314
rect 593 236 659 280
rect 697 320 773 356
rect 697 286 723 320
rect 757 286 773 320
rect 697 270 773 286
rect 479 202 545 217
rect 807 206 841 390
rect 479 190 634 202
rect 479 183 584 190
rect 479 149 495 183
rect 529 156 584 183
rect 618 156 634 190
rect 529 149 634 156
rect 479 120 634 149
rect 479 115 584 120
rect 479 81 495 115
rect 529 86 584 115
rect 618 86 634 120
rect 529 81 634 86
rect 479 65 634 81
rect 668 190 734 202
rect 668 156 684 190
rect 718 156 734 190
rect 668 120 734 156
rect 668 86 684 120
rect 718 86 734 120
rect 668 17 734 86
rect 768 190 841 206
rect 768 156 784 190
rect 818 156 841 190
rect 768 120 841 156
rect 768 86 784 120
rect 818 86 841 120
rect 768 70 841 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 ebufn_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 1840778
string GDS_START 1833586
<< end >>
