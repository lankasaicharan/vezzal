magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 1140 241 2002 259
rect 4 49 2002 241
rect 0 0 2016 49
<< scnmos >>
rect 83 47 113 215
rect 169 47 199 215
rect 255 47 285 215
rect 341 47 371 215
rect 427 47 457 215
rect 513 47 543 215
rect 599 47 629 215
rect 685 47 715 215
rect 771 47 801 215
rect 857 47 887 215
rect 943 47 973 215
rect 1029 47 1059 215
rect 1223 65 1253 233
rect 1309 65 1339 233
rect 1395 65 1425 233
rect 1493 65 1523 233
rect 1581 65 1611 233
rect 1691 65 1721 233
rect 1781 65 1811 233
rect 1881 65 1911 233
<< scpmoshvt >>
rect 83 367 113 619
rect 169 367 199 619
rect 255 367 285 619
rect 341 367 371 619
rect 427 367 457 619
rect 513 367 543 619
rect 599 367 629 619
rect 685 367 715 619
rect 877 367 907 619
rect 963 367 993 619
rect 1049 367 1079 619
rect 1135 367 1165 619
rect 1221 367 1251 619
rect 1307 367 1337 619
rect 1393 367 1423 619
rect 1479 367 1509 619
rect 1565 367 1595 619
rect 1651 367 1681 619
rect 1737 367 1767 619
rect 1823 367 1853 619
<< ndiff >>
rect 30 193 83 215
rect 30 159 38 193
rect 72 159 83 193
rect 30 93 83 159
rect 30 59 38 93
rect 72 59 83 93
rect 30 47 83 59
rect 113 186 169 215
rect 113 152 124 186
rect 158 152 169 186
rect 113 101 169 152
rect 113 67 124 101
rect 158 67 169 101
rect 113 47 169 67
rect 199 126 255 215
rect 199 92 210 126
rect 244 92 255 126
rect 199 47 255 92
rect 285 202 341 215
rect 285 168 296 202
rect 330 168 341 202
rect 285 101 341 168
rect 285 67 296 101
rect 330 67 341 101
rect 285 47 341 67
rect 371 126 427 215
rect 371 92 382 126
rect 416 92 427 126
rect 371 47 427 92
rect 457 202 513 215
rect 457 168 468 202
rect 502 168 513 202
rect 457 101 513 168
rect 457 67 468 101
rect 502 67 513 101
rect 457 47 513 67
rect 543 126 599 215
rect 543 92 554 126
rect 588 92 599 126
rect 543 47 599 92
rect 629 202 685 215
rect 629 168 640 202
rect 674 168 685 202
rect 629 101 685 168
rect 629 67 640 101
rect 674 67 685 101
rect 629 47 685 67
rect 715 107 771 215
rect 715 73 726 107
rect 760 73 771 107
rect 715 47 771 73
rect 801 183 857 215
rect 801 149 812 183
rect 846 149 857 183
rect 801 101 857 149
rect 801 67 812 101
rect 846 67 857 101
rect 801 47 857 67
rect 887 107 943 215
rect 887 73 898 107
rect 932 73 943 107
rect 887 47 943 73
rect 973 183 1029 215
rect 973 149 984 183
rect 1018 149 1029 183
rect 973 101 1029 149
rect 973 67 984 101
rect 1018 67 1029 101
rect 973 47 1029 67
rect 1059 105 1112 215
rect 1059 71 1070 105
rect 1104 71 1112 105
rect 1059 47 1112 71
rect 1166 107 1223 233
rect 1166 73 1178 107
rect 1212 73 1223 107
rect 1166 65 1223 73
rect 1253 181 1309 233
rect 1253 147 1264 181
rect 1298 147 1309 181
rect 1253 65 1309 147
rect 1339 107 1395 233
rect 1339 73 1350 107
rect 1384 73 1395 107
rect 1339 65 1395 73
rect 1425 181 1493 233
rect 1425 147 1436 181
rect 1470 147 1493 181
rect 1425 65 1493 147
rect 1523 183 1581 233
rect 1523 149 1536 183
rect 1570 149 1581 183
rect 1523 111 1581 149
rect 1523 77 1536 111
rect 1570 77 1581 111
rect 1523 65 1581 77
rect 1611 225 1691 233
rect 1611 191 1636 225
rect 1670 191 1691 225
rect 1611 153 1691 191
rect 1611 119 1636 153
rect 1670 119 1691 153
rect 1611 65 1691 119
rect 1721 183 1781 233
rect 1721 149 1736 183
rect 1770 149 1781 183
rect 1721 110 1781 149
rect 1721 76 1736 110
rect 1770 76 1781 110
rect 1721 65 1781 76
rect 1811 225 1881 233
rect 1811 191 1836 225
rect 1870 191 1881 225
rect 1811 153 1881 191
rect 1811 119 1836 153
rect 1870 119 1881 153
rect 1811 65 1881 119
rect 1911 222 1976 233
rect 1911 188 1922 222
rect 1956 188 1976 222
rect 1911 111 1976 188
rect 1911 77 1922 111
rect 1956 77 1976 111
rect 1911 65 1976 77
<< pdiff >>
rect 30 599 83 619
rect 30 565 38 599
rect 72 565 83 599
rect 30 507 83 565
rect 30 473 38 507
rect 72 473 83 507
rect 30 413 83 473
rect 30 379 38 413
rect 72 379 83 413
rect 30 367 83 379
rect 113 607 169 619
rect 113 573 124 607
rect 158 573 169 607
rect 113 515 169 573
rect 113 481 124 515
rect 158 481 169 515
rect 113 423 169 481
rect 113 389 124 423
rect 158 389 169 423
rect 113 367 169 389
rect 199 599 255 619
rect 199 565 210 599
rect 244 565 255 599
rect 199 507 255 565
rect 199 473 210 507
rect 244 473 255 507
rect 199 413 255 473
rect 199 379 210 413
rect 244 379 255 413
rect 199 367 255 379
rect 285 607 341 619
rect 285 573 296 607
rect 330 573 341 607
rect 285 515 341 573
rect 285 481 296 515
rect 330 481 341 515
rect 285 423 341 481
rect 285 389 296 423
rect 330 389 341 423
rect 285 367 341 389
rect 371 599 427 619
rect 371 565 382 599
rect 416 565 427 599
rect 371 507 427 565
rect 371 473 382 507
rect 416 473 427 507
rect 371 413 427 473
rect 371 379 382 413
rect 416 379 427 413
rect 371 367 427 379
rect 457 607 513 619
rect 457 573 468 607
rect 502 573 513 607
rect 457 515 513 573
rect 457 481 468 515
rect 502 481 513 515
rect 457 423 513 481
rect 457 389 468 423
rect 502 389 513 423
rect 457 367 513 389
rect 543 531 599 619
rect 543 497 554 531
rect 588 497 599 531
rect 543 413 599 497
rect 543 379 554 413
rect 588 379 599 413
rect 543 367 599 379
rect 629 607 685 619
rect 629 573 640 607
rect 674 573 685 607
rect 629 515 685 573
rect 629 481 640 515
rect 674 481 685 515
rect 629 423 685 481
rect 629 389 640 423
rect 674 389 685 423
rect 629 367 685 389
rect 715 531 768 619
rect 715 497 726 531
rect 760 497 768 531
rect 715 413 768 497
rect 715 379 726 413
rect 760 379 768 413
rect 715 367 768 379
rect 824 531 877 619
rect 824 497 832 531
rect 866 497 877 531
rect 824 418 877 497
rect 824 384 832 418
rect 866 384 877 418
rect 824 367 877 384
rect 907 599 963 619
rect 907 565 918 599
rect 952 565 963 599
rect 907 492 963 565
rect 907 458 918 492
rect 952 458 963 492
rect 907 367 963 458
rect 993 531 1049 619
rect 993 497 1004 531
rect 1038 497 1049 531
rect 993 418 1049 497
rect 993 384 1004 418
rect 1038 384 1049 418
rect 993 367 1049 384
rect 1079 599 1135 619
rect 1079 565 1090 599
rect 1124 565 1135 599
rect 1079 492 1135 565
rect 1079 458 1090 492
rect 1124 458 1135 492
rect 1079 367 1135 458
rect 1165 599 1221 619
rect 1165 565 1176 599
rect 1210 565 1221 599
rect 1165 510 1221 565
rect 1165 476 1176 510
rect 1210 476 1221 510
rect 1165 418 1221 476
rect 1165 384 1176 418
rect 1210 384 1221 418
rect 1165 367 1221 384
rect 1251 607 1307 619
rect 1251 573 1262 607
rect 1296 573 1307 607
rect 1251 492 1307 573
rect 1251 458 1262 492
rect 1296 458 1307 492
rect 1251 367 1307 458
rect 1337 599 1393 619
rect 1337 565 1348 599
rect 1382 565 1393 599
rect 1337 510 1393 565
rect 1337 476 1348 510
rect 1382 476 1393 510
rect 1337 418 1393 476
rect 1337 384 1348 418
rect 1382 384 1393 418
rect 1337 367 1393 384
rect 1423 607 1479 619
rect 1423 573 1434 607
rect 1468 573 1479 607
rect 1423 486 1479 573
rect 1423 452 1434 486
rect 1468 452 1479 486
rect 1423 367 1479 452
rect 1509 599 1565 619
rect 1509 565 1520 599
rect 1554 565 1565 599
rect 1509 510 1565 565
rect 1509 476 1520 510
rect 1554 476 1565 510
rect 1509 418 1565 476
rect 1509 384 1520 418
rect 1554 384 1565 418
rect 1509 367 1565 384
rect 1595 607 1651 619
rect 1595 573 1606 607
rect 1640 573 1651 607
rect 1595 486 1651 573
rect 1595 452 1606 486
rect 1640 452 1651 486
rect 1595 367 1651 452
rect 1681 599 1737 619
rect 1681 565 1692 599
rect 1726 565 1737 599
rect 1681 510 1737 565
rect 1681 476 1692 510
rect 1726 476 1737 510
rect 1681 418 1737 476
rect 1681 384 1692 418
rect 1726 384 1737 418
rect 1681 367 1737 384
rect 1767 607 1823 619
rect 1767 573 1778 607
rect 1812 573 1823 607
rect 1767 486 1823 573
rect 1767 452 1778 486
rect 1812 452 1823 486
rect 1767 367 1823 452
rect 1853 599 1906 619
rect 1853 565 1864 599
rect 1898 565 1906 599
rect 1853 510 1906 565
rect 1853 476 1864 510
rect 1898 476 1906 510
rect 1853 418 1906 476
rect 1853 384 1864 418
rect 1898 384 1906 418
rect 1853 367 1906 384
<< ndiffc >>
rect 38 159 72 193
rect 38 59 72 93
rect 124 152 158 186
rect 124 67 158 101
rect 210 92 244 126
rect 296 168 330 202
rect 296 67 330 101
rect 382 92 416 126
rect 468 168 502 202
rect 468 67 502 101
rect 554 92 588 126
rect 640 168 674 202
rect 640 67 674 101
rect 726 73 760 107
rect 812 149 846 183
rect 812 67 846 101
rect 898 73 932 107
rect 984 149 1018 183
rect 984 67 1018 101
rect 1070 71 1104 105
rect 1178 73 1212 107
rect 1264 147 1298 181
rect 1350 73 1384 107
rect 1436 147 1470 181
rect 1536 149 1570 183
rect 1536 77 1570 111
rect 1636 191 1670 225
rect 1636 119 1670 153
rect 1736 149 1770 183
rect 1736 76 1770 110
rect 1836 191 1870 225
rect 1836 119 1870 153
rect 1922 188 1956 222
rect 1922 77 1956 111
<< pdiffc >>
rect 38 565 72 599
rect 38 473 72 507
rect 38 379 72 413
rect 124 573 158 607
rect 124 481 158 515
rect 124 389 158 423
rect 210 565 244 599
rect 210 473 244 507
rect 210 379 244 413
rect 296 573 330 607
rect 296 481 330 515
rect 296 389 330 423
rect 382 565 416 599
rect 382 473 416 507
rect 382 379 416 413
rect 468 573 502 607
rect 468 481 502 515
rect 468 389 502 423
rect 554 497 588 531
rect 554 379 588 413
rect 640 573 674 607
rect 640 481 674 515
rect 640 389 674 423
rect 726 497 760 531
rect 726 379 760 413
rect 832 497 866 531
rect 832 384 866 418
rect 918 565 952 599
rect 918 458 952 492
rect 1004 497 1038 531
rect 1004 384 1038 418
rect 1090 565 1124 599
rect 1090 458 1124 492
rect 1176 565 1210 599
rect 1176 476 1210 510
rect 1176 384 1210 418
rect 1262 573 1296 607
rect 1262 458 1296 492
rect 1348 565 1382 599
rect 1348 476 1382 510
rect 1348 384 1382 418
rect 1434 573 1468 607
rect 1434 452 1468 486
rect 1520 565 1554 599
rect 1520 476 1554 510
rect 1520 384 1554 418
rect 1606 573 1640 607
rect 1606 452 1640 486
rect 1692 565 1726 599
rect 1692 476 1726 510
rect 1692 384 1726 418
rect 1778 573 1812 607
rect 1778 452 1812 486
rect 1864 565 1898 599
rect 1864 476 1898 510
rect 1864 384 1898 418
<< poly >>
rect 83 619 113 645
rect 169 619 199 645
rect 255 619 285 645
rect 341 619 371 645
rect 427 619 457 645
rect 513 619 543 645
rect 599 619 629 645
rect 685 619 715 645
rect 877 619 907 645
rect 963 619 993 645
rect 1049 619 1079 645
rect 1135 619 1165 645
rect 1221 619 1251 645
rect 1307 619 1337 645
rect 1393 619 1423 645
rect 1479 619 1509 645
rect 1565 619 1595 645
rect 1651 619 1681 645
rect 1737 619 1767 645
rect 1823 619 1853 645
rect 83 303 113 367
rect 169 303 199 367
rect 255 303 285 367
rect 341 303 371 367
rect 33 287 371 303
rect 33 253 49 287
rect 83 253 117 287
rect 151 253 185 287
rect 219 253 253 287
rect 287 253 321 287
rect 355 253 371 287
rect 33 237 371 253
rect 83 215 113 237
rect 169 215 199 237
rect 255 215 285 237
rect 341 215 371 237
rect 427 303 457 367
rect 513 303 543 367
rect 599 303 629 367
rect 685 303 715 367
rect 877 335 907 367
rect 963 335 993 367
rect 1049 335 1079 367
rect 1135 335 1165 367
rect 427 287 715 303
rect 857 319 1165 335
rect 857 299 911 319
rect 427 253 443 287
rect 477 253 511 287
rect 545 253 579 287
rect 613 253 647 287
rect 681 253 715 287
rect 427 237 715 253
rect 427 215 457 237
rect 513 215 543 237
rect 599 215 629 237
rect 685 215 715 237
rect 771 285 911 299
rect 945 285 979 319
rect 1013 285 1047 319
rect 1081 285 1115 319
rect 1149 285 1165 319
rect 1221 345 1251 367
rect 1307 345 1337 367
rect 1393 345 1423 367
rect 1479 345 1509 367
rect 1221 335 1509 345
rect 1565 345 1595 367
rect 1651 345 1681 367
rect 1737 345 1767 367
rect 1823 345 1853 367
rect 1565 335 1853 345
rect 1221 319 1523 335
rect 1221 315 1269 319
rect 771 269 1165 285
rect 1223 285 1269 315
rect 1303 285 1337 319
rect 1371 285 1405 319
rect 1439 285 1473 319
rect 1507 285 1523 319
rect 1223 269 1523 285
rect 1565 319 1971 335
rect 1565 285 1581 319
rect 1615 285 1649 319
rect 1683 285 1717 319
rect 1751 285 1785 319
rect 1819 285 1853 319
rect 1887 285 1921 319
rect 1955 285 1971 319
rect 1565 269 1971 285
rect 771 215 801 269
rect 857 215 887 269
rect 943 215 973 269
rect 1029 215 1059 269
rect 1223 233 1253 269
rect 1309 233 1339 269
rect 1395 233 1425 269
rect 1493 233 1523 269
rect 1581 233 1611 269
rect 1691 233 1721 269
rect 1781 233 1811 269
rect 1881 233 1911 269
rect 83 21 113 47
rect 169 21 199 47
rect 255 21 285 47
rect 341 21 371 47
rect 427 21 457 47
rect 513 21 543 47
rect 599 21 629 47
rect 685 21 715 47
rect 771 21 801 47
rect 857 21 887 47
rect 943 21 973 47
rect 1029 21 1059 47
rect 1223 39 1253 65
rect 1309 39 1339 65
rect 1395 39 1425 65
rect 1493 39 1523 65
rect 1581 39 1611 65
rect 1691 39 1721 65
rect 1781 39 1811 65
rect 1881 39 1911 65
<< polycont >>
rect 49 253 83 287
rect 117 253 151 287
rect 185 253 219 287
rect 253 253 287 287
rect 321 253 355 287
rect 443 253 477 287
rect 511 253 545 287
rect 579 253 613 287
rect 647 253 681 287
rect 911 285 945 319
rect 979 285 1013 319
rect 1047 285 1081 319
rect 1115 285 1149 319
rect 1269 285 1303 319
rect 1337 285 1371 319
rect 1405 285 1439 319
rect 1473 285 1507 319
rect 1581 285 1615 319
rect 1649 285 1683 319
rect 1717 285 1751 319
rect 1785 285 1819 319
rect 1853 285 1887 319
rect 1921 285 1955 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 22 599 74 615
rect 22 565 38 599
rect 72 565 74 599
rect 22 507 74 565
rect 22 473 38 507
rect 72 473 74 507
rect 22 413 74 473
rect 22 379 38 413
rect 72 379 74 413
rect 108 607 174 649
rect 108 573 124 607
rect 158 573 174 607
rect 108 515 174 573
rect 108 481 124 515
rect 158 481 174 515
rect 108 423 174 481
rect 108 389 124 423
rect 158 389 174 423
rect 208 599 246 615
rect 208 565 210 599
rect 244 565 246 599
rect 208 507 246 565
rect 208 473 210 507
rect 244 473 246 507
rect 208 413 246 473
rect 22 355 74 379
rect 208 379 210 413
rect 244 379 246 413
rect 280 607 346 649
rect 280 573 296 607
rect 330 573 346 607
rect 280 515 346 573
rect 280 481 296 515
rect 330 481 346 515
rect 280 423 346 481
rect 280 389 296 423
rect 330 389 346 423
rect 380 599 418 615
rect 380 565 382 599
rect 416 565 418 599
rect 380 507 418 565
rect 380 473 382 507
rect 416 473 418 507
rect 380 413 418 473
rect 208 355 246 379
rect 380 379 382 413
rect 416 379 418 413
rect 452 607 1140 615
rect 452 573 468 607
rect 502 581 640 607
rect 502 573 518 581
rect 452 515 518 573
rect 624 573 640 581
rect 674 599 1140 607
rect 674 581 918 599
rect 674 573 690 581
rect 452 481 468 515
rect 502 481 518 515
rect 452 423 518 481
rect 452 389 468 423
rect 502 389 518 423
rect 552 531 590 547
rect 552 497 554 531
rect 588 497 590 531
rect 552 413 590 497
rect 380 355 418 379
rect 552 379 554 413
rect 588 379 590 413
rect 624 515 690 573
rect 902 565 918 581
rect 952 581 1090 599
rect 952 565 968 581
rect 624 481 640 515
rect 674 481 690 515
rect 624 423 690 481
rect 624 389 640 423
rect 674 389 690 423
rect 724 531 776 547
rect 724 497 726 531
rect 760 497 776 531
rect 724 413 776 497
rect 552 355 590 379
rect 724 379 726 413
rect 760 379 776 413
rect 724 355 776 379
rect 22 321 776 355
rect 816 531 868 547
rect 816 497 832 531
rect 866 497 868 531
rect 816 424 868 497
rect 902 492 968 565
rect 1074 565 1090 581
rect 1124 565 1140 599
rect 902 458 918 492
rect 952 458 968 492
rect 1002 531 1040 547
rect 1002 497 1004 531
rect 1038 497 1040 531
rect 1002 424 1040 497
rect 1074 492 1140 565
rect 1074 458 1090 492
rect 1124 458 1140 492
rect 1174 599 1212 615
rect 1174 565 1176 599
rect 1210 565 1212 599
rect 1174 510 1212 565
rect 1174 476 1176 510
rect 1210 476 1212 510
rect 1174 424 1212 476
rect 1246 607 1312 649
rect 1246 573 1262 607
rect 1296 573 1312 607
rect 1246 492 1312 573
rect 1246 458 1262 492
rect 1296 458 1312 492
rect 1346 599 1384 615
rect 1346 565 1348 599
rect 1382 565 1384 599
rect 1346 510 1384 565
rect 1346 476 1348 510
rect 1382 476 1384 510
rect 1346 424 1384 476
rect 1418 607 1484 649
rect 1418 573 1434 607
rect 1468 573 1484 607
rect 1418 486 1484 573
rect 1418 452 1434 486
rect 1468 452 1484 486
rect 1518 599 1556 615
rect 1518 565 1520 599
rect 1554 565 1556 599
rect 1518 510 1556 565
rect 1518 476 1520 510
rect 1554 476 1556 510
rect 816 418 1384 424
rect 1518 418 1556 476
rect 1590 607 1656 649
rect 1590 573 1606 607
rect 1640 573 1656 607
rect 1590 486 1656 573
rect 1590 452 1606 486
rect 1640 452 1656 486
rect 1690 599 1728 615
rect 1690 565 1692 599
rect 1726 565 1728 599
rect 1690 510 1728 565
rect 1690 476 1692 510
rect 1726 476 1728 510
rect 1690 418 1728 476
rect 1762 607 1828 649
rect 1762 573 1778 607
rect 1812 573 1828 607
rect 1762 486 1828 573
rect 1762 452 1778 486
rect 1812 452 1828 486
rect 1862 599 1914 615
rect 1862 565 1864 599
rect 1898 565 1914 599
rect 1862 510 1914 565
rect 1862 476 1864 510
rect 1898 476 1914 510
rect 1862 418 1914 476
rect 816 384 832 418
rect 866 384 1004 418
rect 1038 384 1176 418
rect 1210 384 1348 418
rect 1382 384 1520 418
rect 1554 384 1692 418
rect 1726 384 1864 418
rect 1898 384 1914 418
rect 18 253 49 287
rect 83 253 117 287
rect 151 253 185 287
rect 219 253 253 287
rect 287 253 321 287
rect 355 253 372 287
rect 18 236 372 253
rect 406 253 443 287
rect 477 253 511 287
rect 545 253 579 287
rect 613 253 647 287
rect 681 253 759 287
rect 406 236 759 253
rect 816 251 859 384
rect 893 319 1219 350
rect 893 285 911 319
rect 945 285 979 319
rect 1013 285 1047 319
rect 1081 285 1115 319
rect 1149 285 1219 319
rect 1253 319 1523 350
rect 1253 285 1269 319
rect 1303 285 1337 319
rect 1371 285 1405 319
rect 1439 285 1473 319
rect 1507 285 1523 319
rect 1557 319 1999 350
rect 1557 285 1581 319
rect 1615 285 1649 319
rect 1683 285 1717 319
rect 1751 285 1785 319
rect 1819 285 1853 319
rect 1887 285 1921 319
rect 1955 285 1999 319
rect 816 225 1886 251
rect 816 217 1636 225
rect 22 193 88 202
rect 22 159 38 193
rect 72 159 88 193
rect 22 93 88 159
rect 22 59 38 93
rect 72 59 88 93
rect 22 17 88 59
rect 122 186 296 202
rect 122 152 124 186
rect 158 168 296 186
rect 330 168 468 202
rect 502 168 640 202
rect 674 183 782 202
rect 1620 191 1636 217
rect 1670 217 1836 225
rect 1670 191 1686 217
rect 674 168 812 183
rect 158 152 160 168
rect 122 101 160 152
rect 122 67 124 101
rect 158 67 160 101
rect 122 51 160 67
rect 194 126 260 134
rect 194 92 210 126
rect 244 92 260 126
rect 194 17 260 92
rect 294 101 332 168
rect 294 67 296 101
rect 330 67 332 101
rect 294 51 332 67
rect 366 126 432 134
rect 366 92 382 126
rect 416 92 432 126
rect 366 17 432 92
rect 466 101 504 168
rect 638 149 812 168
rect 846 149 984 183
rect 1018 181 1486 183
rect 1018 149 1264 181
rect 466 67 468 101
rect 502 67 504 101
rect 466 51 504 67
rect 538 126 604 134
rect 538 92 554 126
rect 588 92 604 126
rect 538 17 604 92
rect 638 101 676 149
rect 638 67 640 101
rect 674 67 676 101
rect 638 51 676 67
rect 710 107 776 115
rect 710 73 726 107
rect 760 73 776 107
rect 710 17 776 73
rect 810 101 848 149
rect 982 147 1264 149
rect 1298 147 1436 181
rect 1470 147 1486 181
rect 982 145 1486 147
rect 1520 149 1536 183
rect 1570 149 1586 183
rect 810 67 812 101
rect 846 67 848 101
rect 810 51 848 67
rect 882 107 948 115
rect 882 73 898 107
rect 932 73 948 107
rect 882 17 948 73
rect 982 101 1020 145
rect 1520 111 1586 149
rect 1620 153 1686 191
rect 1820 191 1836 217
rect 1870 191 1886 225
rect 1620 119 1636 153
rect 1670 119 1686 153
rect 1720 149 1736 183
rect 1770 149 1786 183
rect 982 67 984 101
rect 1018 67 1020 101
rect 982 51 1020 67
rect 1054 105 1120 111
rect 1054 71 1070 105
rect 1104 71 1120 105
rect 1054 17 1120 71
rect 1162 107 1536 111
rect 1162 73 1178 107
rect 1212 73 1350 107
rect 1384 77 1536 107
rect 1570 85 1586 111
rect 1720 110 1786 149
rect 1820 153 1886 191
rect 1820 119 1836 153
rect 1870 119 1886 153
rect 1920 222 1972 238
rect 1920 188 1922 222
rect 1956 188 1972 222
rect 1720 85 1736 110
rect 1570 77 1736 85
rect 1384 76 1736 77
rect 1770 85 1786 110
rect 1920 111 1972 188
rect 1920 85 1922 111
rect 1770 77 1922 85
rect 1956 77 1972 111
rect 1770 76 1972 77
rect 1384 73 1972 76
rect 1162 51 1972 73
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o311ai_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1759 316 1793 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1087 390 1121 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1183 390 1217 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1585892
string GDS_START 1568196
<< end >>
