magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 277 241 861 245
rect 1 49 861 241
rect 0 0 864 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 356 51 386 219
rect 428 51 458 219
rect 536 51 566 219
rect 644 51 674 219
rect 752 51 782 219
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 342 367 372 619
rect 428 367 458 619
rect 536 367 566 619
rect 644 367 674 619
rect 752 367 782 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 93 80 169
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 203 166 215
rect 110 169 121 203
rect 155 169 166 203
rect 110 101 166 169
rect 110 67 121 101
rect 155 67 166 101
rect 110 47 166 67
rect 196 161 249 215
rect 196 127 207 161
rect 241 127 249 161
rect 196 93 249 127
rect 196 59 207 93
rect 241 59 249 93
rect 196 47 249 59
rect 303 207 356 219
rect 303 173 311 207
rect 345 173 356 207
rect 303 101 356 173
rect 303 67 311 101
rect 345 67 356 101
rect 303 51 356 67
rect 386 51 428 219
rect 458 51 536 219
rect 566 207 644 219
rect 566 173 589 207
rect 623 173 644 207
rect 566 97 644 173
rect 566 63 589 97
rect 623 63 644 97
rect 566 51 644 63
rect 674 173 752 219
rect 674 139 693 173
rect 727 139 752 173
rect 674 97 752 139
rect 674 63 693 97
rect 727 63 752 97
rect 674 51 752 63
rect 782 207 835 219
rect 782 173 793 207
rect 827 173 835 207
rect 782 97 835 173
rect 782 63 793 97
rect 827 63 835 97
rect 782 51 835 63
<< pdiff >>
rect 27 607 80 619
rect 27 573 35 607
rect 69 573 80 607
rect 27 505 80 573
rect 27 471 35 505
rect 69 471 80 505
rect 27 414 80 471
rect 27 380 35 414
rect 69 380 80 414
rect 27 367 80 380
rect 110 599 166 619
rect 110 565 121 599
rect 155 565 166 599
rect 110 502 166 565
rect 110 468 121 502
rect 155 468 166 502
rect 110 413 166 468
rect 110 379 121 413
rect 155 379 166 413
rect 110 367 166 379
rect 196 607 342 619
rect 196 573 207 607
rect 241 573 297 607
rect 331 573 342 607
rect 196 493 342 573
rect 196 459 211 493
rect 245 459 297 493
rect 331 459 342 493
rect 196 367 342 459
rect 372 599 428 619
rect 372 565 383 599
rect 417 565 428 599
rect 372 510 428 565
rect 372 476 383 510
rect 417 476 428 510
rect 372 425 428 476
rect 372 391 383 425
rect 417 391 428 425
rect 372 367 428 391
rect 458 607 536 619
rect 458 573 481 607
rect 515 573 536 607
rect 458 497 536 573
rect 458 463 481 497
rect 515 463 536 497
rect 458 367 536 463
rect 566 607 644 619
rect 566 573 589 607
rect 623 573 644 607
rect 566 516 644 573
rect 566 482 589 516
rect 623 482 644 516
rect 566 425 644 482
rect 566 391 589 425
rect 623 391 644 425
rect 566 367 644 391
rect 674 367 752 619
rect 782 607 835 619
rect 782 573 793 607
rect 827 573 835 607
rect 782 511 835 573
rect 782 477 793 511
rect 827 477 835 511
rect 782 418 835 477
rect 782 384 793 418
rect 827 384 835 418
rect 782 367 835 384
<< ndiffc >>
rect 35 169 69 203
rect 35 59 69 93
rect 121 169 155 203
rect 121 67 155 101
rect 207 127 241 161
rect 207 59 241 93
rect 311 173 345 207
rect 311 67 345 101
rect 589 173 623 207
rect 589 63 623 97
rect 693 139 727 173
rect 693 63 727 97
rect 793 173 827 207
rect 793 63 827 97
<< pdiffc >>
rect 35 573 69 607
rect 35 471 69 505
rect 35 380 69 414
rect 121 565 155 599
rect 121 468 155 502
rect 121 379 155 413
rect 207 573 241 607
rect 297 573 331 607
rect 211 459 245 493
rect 297 459 331 493
rect 383 565 417 599
rect 383 476 417 510
rect 383 391 417 425
rect 481 573 515 607
rect 481 463 515 497
rect 589 573 623 607
rect 589 482 623 516
rect 589 391 623 425
rect 793 573 827 607
rect 793 477 827 511
rect 793 384 827 418
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 342 619 372 645
rect 428 619 458 645
rect 536 619 566 645
rect 644 619 674 645
rect 752 619 782 645
rect 80 345 110 367
rect 166 345 196 367
rect 80 287 245 345
rect 342 335 372 367
rect 80 253 195 287
rect 229 253 245 287
rect 295 319 386 335
rect 295 285 311 319
rect 345 285 386 319
rect 295 269 386 285
rect 80 237 245 253
rect 80 215 110 237
rect 166 215 196 237
rect 356 219 386 269
rect 428 307 458 367
rect 536 335 566 367
rect 644 335 674 367
rect 536 319 602 335
rect 428 291 494 307
rect 428 257 444 291
rect 478 257 494 291
rect 428 241 494 257
rect 536 285 552 319
rect 586 285 602 319
rect 536 269 602 285
rect 644 319 710 335
rect 644 285 660 319
rect 694 285 710 319
rect 644 269 710 285
rect 752 325 782 367
rect 752 309 843 325
rect 752 275 793 309
rect 827 275 843 309
rect 428 219 458 241
rect 536 219 566 269
rect 644 219 674 269
rect 752 259 843 275
rect 752 219 782 259
rect 80 21 110 47
rect 166 21 196 47
rect 356 25 386 51
rect 428 25 458 51
rect 536 25 566 51
rect 644 25 674 51
rect 752 25 782 51
<< polycont >>
rect 195 253 229 287
rect 311 285 345 319
rect 444 257 478 291
rect 552 285 586 319
rect 660 285 694 319
rect 793 275 827 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 19 607 78 649
rect 19 573 35 607
rect 69 573 78 607
rect 19 505 78 573
rect 19 471 35 505
rect 69 471 78 505
rect 19 414 78 471
rect 19 380 35 414
rect 69 380 78 414
rect 19 364 78 380
rect 112 599 161 615
rect 112 565 121 599
rect 155 565 161 599
rect 112 502 161 565
rect 112 468 121 502
rect 155 468 161 502
rect 112 413 161 468
rect 195 607 347 649
rect 195 573 207 607
rect 241 573 297 607
rect 331 573 347 607
rect 195 493 347 573
rect 195 459 211 493
rect 245 459 297 493
rect 331 459 347 493
rect 381 599 431 615
rect 381 565 383 599
rect 417 565 431 599
rect 381 510 431 565
rect 381 476 383 510
rect 417 476 431 510
rect 381 425 431 476
rect 465 607 531 649
rect 465 573 481 607
rect 515 573 531 607
rect 465 497 531 573
rect 465 463 481 497
rect 515 463 531 497
rect 465 459 531 463
rect 573 607 639 615
rect 573 573 589 607
rect 623 573 639 607
rect 777 607 843 649
rect 573 516 639 573
rect 573 482 589 516
rect 623 482 639 516
rect 573 425 639 482
rect 112 379 121 413
rect 155 379 161 413
rect 19 203 78 219
rect 19 169 35 203
rect 69 169 78 203
rect 19 93 78 169
rect 19 59 35 93
rect 69 59 78 93
rect 19 17 78 59
rect 112 203 161 379
rect 209 391 383 425
rect 417 391 589 425
rect 623 391 639 425
rect 209 303 261 391
rect 195 287 261 303
rect 229 253 261 287
rect 295 319 368 357
rect 295 285 311 319
rect 345 285 368 319
rect 402 307 464 357
rect 511 319 602 357
rect 687 335 743 596
rect 777 573 793 607
rect 827 573 843 607
rect 777 511 843 573
rect 777 477 793 511
rect 827 477 843 511
rect 777 418 843 477
rect 777 384 793 418
rect 827 384 843 418
rect 511 316 552 319
rect 402 291 478 307
rect 195 245 261 253
rect 402 257 444 291
rect 536 285 552 316
rect 586 285 602 319
rect 644 319 743 335
rect 644 285 660 319
rect 694 285 743 319
rect 777 309 847 350
rect 777 275 793 309
rect 827 275 847 309
rect 195 231 315 245
rect 195 211 361 231
rect 286 207 361 211
rect 286 204 311 207
rect 112 169 121 203
rect 155 169 161 203
rect 112 101 161 169
rect 112 67 121 101
rect 155 67 161 101
rect 112 51 161 67
rect 195 161 257 177
rect 195 127 207 161
rect 241 127 257 161
rect 195 93 257 127
rect 195 59 207 93
rect 241 59 257 93
rect 195 17 257 59
rect 291 173 311 204
rect 345 173 361 207
rect 291 101 361 173
rect 291 67 311 101
rect 345 67 361 101
rect 402 72 478 257
rect 573 207 843 241
rect 573 173 589 207
rect 623 173 639 207
rect 777 173 793 207
rect 827 173 843 207
rect 573 97 639 173
rect 291 51 361 67
rect 573 63 589 97
rect 623 63 639 97
rect 573 51 639 63
rect 677 139 693 173
rect 727 139 743 173
rect 677 97 743 139
rect 677 63 693 97
rect 727 63 743 97
rect 677 17 743 63
rect 777 97 843 173
rect 777 63 793 97
rect 827 63 843 97
rect 777 51 843 63
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2111a_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4197216
string GDS_START 4187974
<< end >>
