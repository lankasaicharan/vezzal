magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 19 49 1499 259
rect 0 0 1536 49
<< scnmos >>
rect 100 65 130 233
rect 186 65 216 233
rect 272 65 302 233
rect 358 65 388 233
rect 444 65 474 233
rect 530 65 560 233
rect 616 65 646 233
rect 702 65 732 233
rect 788 65 818 233
rect 874 65 904 233
rect 960 65 990 233
rect 1046 65 1076 233
rect 1132 65 1162 233
rect 1218 65 1248 233
rect 1304 65 1334 233
rect 1390 65 1420 233
<< scpmoshvt >>
rect 100 367 130 619
rect 186 367 216 619
rect 272 367 302 619
rect 358 367 388 619
rect 444 367 474 619
rect 530 367 560 619
rect 616 367 646 619
rect 702 367 732 619
rect 788 367 818 619
rect 874 367 904 619
rect 960 367 990 619
rect 1046 367 1076 619
rect 1132 367 1162 619
rect 1218 367 1248 619
rect 1304 367 1334 619
rect 1390 367 1420 619
<< ndiff >>
rect 45 221 100 233
rect 45 187 53 221
rect 87 187 100 221
rect 45 111 100 187
rect 45 77 53 111
rect 87 77 100 111
rect 45 65 100 77
rect 130 221 186 233
rect 130 187 141 221
rect 175 187 186 221
rect 130 113 186 187
rect 130 79 141 113
rect 175 79 186 113
rect 130 65 186 79
rect 216 181 272 233
rect 216 147 227 181
rect 261 147 272 181
rect 216 107 272 147
rect 216 73 227 107
rect 261 73 272 107
rect 216 65 272 73
rect 302 221 358 233
rect 302 187 313 221
rect 347 187 358 221
rect 302 113 358 187
rect 302 79 313 113
rect 347 79 358 113
rect 302 65 358 79
rect 388 181 444 233
rect 388 147 399 181
rect 433 147 444 181
rect 388 107 444 147
rect 388 73 399 107
rect 433 73 444 107
rect 388 65 444 73
rect 474 221 530 233
rect 474 187 485 221
rect 519 187 530 221
rect 474 111 530 187
rect 474 77 485 111
rect 519 77 530 111
rect 474 65 530 77
rect 560 208 616 233
rect 560 174 571 208
rect 605 174 616 208
rect 560 111 616 174
rect 560 77 571 111
rect 605 77 616 111
rect 560 65 616 77
rect 646 221 702 233
rect 646 187 657 221
rect 691 187 702 221
rect 646 111 702 187
rect 646 77 657 111
rect 691 77 702 111
rect 646 65 702 77
rect 732 208 788 233
rect 732 174 743 208
rect 777 174 788 208
rect 732 111 788 174
rect 732 77 743 111
rect 777 77 788 111
rect 732 65 788 77
rect 818 221 874 233
rect 818 187 829 221
rect 863 187 874 221
rect 818 111 874 187
rect 818 77 829 111
rect 863 77 874 111
rect 818 65 874 77
rect 904 222 960 233
rect 904 188 915 222
rect 949 188 960 222
rect 904 111 960 188
rect 904 77 915 111
rect 949 77 960 111
rect 904 65 960 77
rect 990 221 1046 233
rect 990 187 1001 221
rect 1035 187 1046 221
rect 990 111 1046 187
rect 990 77 1001 111
rect 1035 77 1046 111
rect 990 65 1046 77
rect 1076 183 1132 233
rect 1076 149 1087 183
rect 1121 149 1132 183
rect 1076 111 1132 149
rect 1076 77 1087 111
rect 1121 77 1132 111
rect 1076 65 1132 77
rect 1162 221 1218 233
rect 1162 187 1173 221
rect 1207 187 1218 221
rect 1162 111 1218 187
rect 1162 77 1173 111
rect 1207 77 1218 111
rect 1162 65 1218 77
rect 1248 183 1304 233
rect 1248 149 1259 183
rect 1293 149 1304 183
rect 1248 111 1304 149
rect 1248 77 1259 111
rect 1293 77 1304 111
rect 1248 65 1304 77
rect 1334 221 1390 233
rect 1334 187 1345 221
rect 1379 187 1390 221
rect 1334 111 1390 187
rect 1334 77 1345 111
rect 1379 77 1390 111
rect 1334 65 1390 77
rect 1420 183 1473 233
rect 1420 149 1431 183
rect 1465 149 1473 183
rect 1420 111 1473 149
rect 1420 77 1431 111
rect 1465 77 1473 111
rect 1420 65 1473 77
<< pdiff >>
rect 47 599 100 619
rect 47 565 55 599
rect 89 565 100 599
rect 47 522 100 565
rect 47 488 55 522
rect 89 488 100 522
rect 47 438 100 488
rect 47 404 55 438
rect 89 404 100 438
rect 47 367 100 404
rect 130 607 186 619
rect 130 573 141 607
rect 175 573 186 607
rect 130 490 186 573
rect 130 456 141 490
rect 175 456 186 490
rect 130 367 186 456
rect 216 599 272 619
rect 216 565 227 599
rect 261 565 272 599
rect 216 522 272 565
rect 216 488 227 522
rect 261 488 272 522
rect 216 438 272 488
rect 216 404 227 438
rect 261 404 272 438
rect 216 367 272 404
rect 302 607 358 619
rect 302 573 313 607
rect 347 573 358 607
rect 302 490 358 573
rect 302 456 313 490
rect 347 456 358 490
rect 302 367 358 456
rect 388 599 444 619
rect 388 565 399 599
rect 433 565 444 599
rect 388 522 444 565
rect 388 488 399 522
rect 433 488 444 522
rect 388 438 444 488
rect 388 404 399 438
rect 433 404 444 438
rect 388 367 444 404
rect 474 607 530 619
rect 474 573 485 607
rect 519 573 530 607
rect 474 490 530 573
rect 474 456 485 490
rect 519 456 530 490
rect 474 367 530 456
rect 560 599 616 619
rect 560 565 571 599
rect 605 565 616 599
rect 560 507 616 565
rect 560 473 571 507
rect 605 473 616 507
rect 560 413 616 473
rect 560 379 571 413
rect 605 379 616 413
rect 560 367 616 379
rect 646 607 702 619
rect 646 573 657 607
rect 691 573 702 607
rect 646 529 702 573
rect 646 495 657 529
rect 691 495 702 529
rect 646 453 702 495
rect 646 419 657 453
rect 691 419 702 453
rect 646 367 702 419
rect 732 599 788 619
rect 732 565 743 599
rect 777 565 788 599
rect 732 507 788 565
rect 732 473 743 507
rect 777 473 788 507
rect 732 413 788 473
rect 732 379 743 413
rect 777 379 788 413
rect 732 367 788 379
rect 818 547 874 619
rect 818 513 829 547
rect 863 513 874 547
rect 818 413 874 513
rect 818 379 829 413
rect 863 379 874 413
rect 818 367 874 379
rect 904 597 960 619
rect 904 563 915 597
rect 949 563 960 597
rect 904 502 960 563
rect 904 468 915 502
rect 949 468 960 502
rect 904 367 960 468
rect 990 547 1046 619
rect 990 513 1001 547
rect 1035 513 1046 547
rect 990 413 1046 513
rect 990 379 1001 413
rect 1035 379 1046 413
rect 990 367 1046 379
rect 1076 597 1132 619
rect 1076 563 1087 597
rect 1121 563 1132 597
rect 1076 502 1132 563
rect 1076 468 1087 502
rect 1121 468 1132 502
rect 1076 367 1132 468
rect 1162 545 1218 619
rect 1162 511 1173 545
rect 1207 511 1218 545
rect 1162 425 1218 511
rect 1162 391 1173 425
rect 1207 391 1218 425
rect 1162 367 1218 391
rect 1248 597 1304 619
rect 1248 563 1259 597
rect 1293 563 1304 597
rect 1248 502 1304 563
rect 1248 468 1259 502
rect 1293 468 1304 502
rect 1248 367 1304 468
rect 1334 545 1390 619
rect 1334 511 1345 545
rect 1379 511 1390 545
rect 1334 425 1390 511
rect 1334 391 1345 425
rect 1379 391 1390 425
rect 1334 367 1390 391
rect 1420 599 1473 619
rect 1420 565 1431 599
rect 1465 565 1473 599
rect 1420 502 1473 565
rect 1420 468 1431 502
rect 1465 468 1473 502
rect 1420 367 1473 468
<< ndiffc >>
rect 53 187 87 221
rect 53 77 87 111
rect 141 187 175 221
rect 141 79 175 113
rect 227 147 261 181
rect 227 73 261 107
rect 313 187 347 221
rect 313 79 347 113
rect 399 147 433 181
rect 399 73 433 107
rect 485 187 519 221
rect 485 77 519 111
rect 571 174 605 208
rect 571 77 605 111
rect 657 187 691 221
rect 657 77 691 111
rect 743 174 777 208
rect 743 77 777 111
rect 829 187 863 221
rect 829 77 863 111
rect 915 188 949 222
rect 915 77 949 111
rect 1001 187 1035 221
rect 1001 77 1035 111
rect 1087 149 1121 183
rect 1087 77 1121 111
rect 1173 187 1207 221
rect 1173 77 1207 111
rect 1259 149 1293 183
rect 1259 77 1293 111
rect 1345 187 1379 221
rect 1345 77 1379 111
rect 1431 149 1465 183
rect 1431 77 1465 111
<< pdiffc >>
rect 55 565 89 599
rect 55 488 89 522
rect 55 404 89 438
rect 141 573 175 607
rect 141 456 175 490
rect 227 565 261 599
rect 227 488 261 522
rect 227 404 261 438
rect 313 573 347 607
rect 313 456 347 490
rect 399 565 433 599
rect 399 488 433 522
rect 399 404 433 438
rect 485 573 519 607
rect 485 456 519 490
rect 571 565 605 599
rect 571 473 605 507
rect 571 379 605 413
rect 657 573 691 607
rect 657 495 691 529
rect 657 419 691 453
rect 743 565 777 599
rect 743 473 777 507
rect 743 379 777 413
rect 829 513 863 547
rect 829 379 863 413
rect 915 563 949 597
rect 915 468 949 502
rect 1001 513 1035 547
rect 1001 379 1035 413
rect 1087 563 1121 597
rect 1087 468 1121 502
rect 1173 511 1207 545
rect 1173 391 1207 425
rect 1259 563 1293 597
rect 1259 468 1293 502
rect 1345 511 1379 545
rect 1345 391 1379 425
rect 1431 565 1465 599
rect 1431 468 1465 502
<< poly >>
rect 100 619 130 645
rect 186 619 216 645
rect 272 619 302 645
rect 358 619 388 645
rect 444 619 474 645
rect 530 619 560 645
rect 616 619 646 645
rect 702 619 732 645
rect 788 619 818 645
rect 874 619 904 645
rect 960 619 990 645
rect 1046 619 1076 645
rect 1132 619 1162 645
rect 1218 619 1248 645
rect 1304 619 1334 645
rect 1390 619 1420 645
rect 100 335 130 367
rect 186 335 216 367
rect 272 335 302 367
rect 358 335 388 367
rect 444 335 474 367
rect 530 335 560 367
rect 616 335 646 367
rect 702 335 732 367
rect 100 319 732 335
rect 100 285 116 319
rect 150 285 184 319
rect 218 285 252 319
rect 286 285 320 319
rect 354 285 388 319
rect 422 285 732 319
rect 100 269 732 285
rect 100 233 130 269
rect 186 233 216 269
rect 272 233 302 269
rect 358 233 388 269
rect 444 233 474 269
rect 530 233 560 269
rect 616 233 646 269
rect 702 233 732 269
rect 788 335 818 367
rect 874 335 904 367
rect 960 335 990 367
rect 1046 335 1076 367
rect 1132 335 1162 367
rect 1218 335 1248 367
rect 1304 335 1334 367
rect 1390 335 1420 367
rect 788 319 1420 335
rect 788 285 1112 319
rect 1146 285 1180 319
rect 1214 285 1248 319
rect 1282 285 1316 319
rect 1350 285 1420 319
rect 788 269 1420 285
rect 788 233 818 269
rect 874 233 904 269
rect 960 233 990 269
rect 1046 233 1076 269
rect 1132 233 1162 269
rect 1218 233 1248 269
rect 1304 233 1334 269
rect 1390 233 1420 269
rect 100 39 130 65
rect 186 39 216 65
rect 272 39 302 65
rect 358 39 388 65
rect 444 39 474 65
rect 530 39 560 65
rect 616 39 646 65
rect 702 39 732 65
rect 788 39 818 65
rect 874 39 904 65
rect 960 39 990 65
rect 1046 39 1076 65
rect 1132 39 1162 65
rect 1218 39 1248 65
rect 1304 39 1334 65
rect 1390 39 1420 65
<< polycont >>
rect 116 285 150 319
rect 184 285 218 319
rect 252 285 286 319
rect 320 285 354 319
rect 388 285 422 319
rect 1112 285 1146 319
rect 1180 285 1214 319
rect 1248 285 1282 319
rect 1316 285 1350 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 37 599 91 615
rect 37 565 55 599
rect 89 565 91 599
rect 37 522 91 565
rect 37 488 55 522
rect 89 488 91 522
rect 37 438 91 488
rect 125 607 191 649
rect 125 573 141 607
rect 175 573 191 607
rect 125 490 191 573
rect 125 456 141 490
rect 175 456 191 490
rect 225 599 263 615
rect 225 565 227 599
rect 261 565 263 599
rect 225 522 263 565
rect 225 488 227 522
rect 261 488 263 522
rect 37 404 55 438
rect 89 422 91 438
rect 225 438 263 488
rect 297 607 363 649
rect 297 573 313 607
rect 347 573 363 607
rect 297 490 363 573
rect 297 456 313 490
rect 347 456 363 490
rect 397 599 435 615
rect 397 565 399 599
rect 433 565 435 599
rect 397 522 435 565
rect 397 488 399 522
rect 433 488 435 522
rect 225 422 227 438
rect 89 404 227 422
rect 261 422 263 438
rect 397 438 435 488
rect 469 607 535 649
rect 469 573 485 607
rect 519 573 535 607
rect 469 490 535 573
rect 469 456 485 490
rect 519 456 535 490
rect 569 599 607 615
rect 569 565 571 599
rect 605 565 607 599
rect 569 507 607 565
rect 569 473 571 507
rect 605 473 607 507
rect 397 422 399 438
rect 261 404 399 422
rect 433 422 435 438
rect 569 422 607 473
rect 433 413 607 422
rect 641 607 707 649
rect 641 573 657 607
rect 691 573 707 607
rect 641 529 707 573
rect 641 495 657 529
rect 691 495 707 529
rect 641 453 707 495
rect 641 419 657 453
rect 691 419 707 453
rect 741 599 1481 615
rect 741 565 743 599
rect 777 597 1431 599
rect 777 581 915 597
rect 777 565 779 581
rect 741 507 779 565
rect 913 563 915 581
rect 949 581 1087 597
rect 949 563 951 581
rect 741 473 743 507
rect 777 473 779 507
rect 433 404 571 413
rect 37 388 571 404
rect 566 379 571 388
rect 605 385 607 413
rect 741 413 779 473
rect 741 385 743 413
rect 605 379 743 385
rect 777 379 779 413
rect 100 319 449 354
rect 566 340 779 379
rect 813 513 829 547
rect 863 513 879 547
rect 813 418 879 513
rect 913 502 951 563
rect 1085 563 1087 581
rect 1121 579 1259 597
rect 1121 563 1123 579
rect 913 468 915 502
rect 949 468 951 502
rect 913 452 951 468
rect 985 513 1001 547
rect 1035 513 1051 547
rect 985 418 1051 513
rect 1085 502 1123 563
rect 1257 563 1259 579
rect 1293 579 1431 597
rect 1293 563 1295 579
rect 1085 468 1087 502
rect 1121 468 1123 502
rect 1085 452 1123 468
rect 1157 511 1173 545
rect 1207 511 1223 545
rect 1157 425 1223 511
rect 1257 502 1295 563
rect 1429 565 1431 579
rect 1465 565 1481 599
rect 1257 468 1259 502
rect 1293 468 1295 502
rect 1257 452 1295 468
rect 1329 511 1345 545
rect 1379 511 1395 545
rect 1157 418 1173 425
rect 813 413 1173 418
rect 813 379 829 413
rect 863 379 1001 413
rect 1035 391 1173 413
rect 1207 418 1223 425
rect 1329 425 1395 511
rect 1429 502 1481 565
rect 1429 468 1431 502
rect 1465 468 1481 502
rect 1429 452 1481 468
rect 1329 418 1345 425
rect 1207 391 1345 418
rect 1379 418 1395 425
rect 1379 391 1519 418
rect 1035 384 1519 391
rect 1035 379 1049 384
rect 100 285 116 319
rect 150 285 184 319
rect 218 285 252 319
rect 286 285 320 319
rect 354 285 388 319
rect 422 285 449 319
rect 813 297 1049 379
rect 100 283 449 285
rect 485 272 1049 297
rect 1083 319 1420 350
rect 1083 285 1112 319
rect 1146 285 1180 319
rect 1214 285 1248 319
rect 1282 285 1316 319
rect 1350 285 1420 319
rect 485 249 865 272
rect 136 242 865 249
rect 37 221 102 237
rect 37 187 53 221
rect 87 187 102 221
rect 37 111 102 187
rect 37 77 53 111
rect 87 77 102 111
rect 37 17 102 77
rect 136 221 521 242
rect 136 187 141 221
rect 175 215 313 221
rect 175 187 177 215
rect 136 113 177 187
rect 311 187 313 215
rect 347 215 485 221
rect 347 187 349 215
rect 136 79 141 113
rect 175 79 177 113
rect 136 63 177 79
rect 211 147 227 181
rect 261 147 277 181
rect 211 107 277 147
rect 211 73 227 107
rect 261 73 277 107
rect 211 17 277 73
rect 311 113 349 187
rect 483 187 485 215
rect 519 187 521 221
rect 655 221 693 242
rect 311 79 313 113
rect 347 79 349 113
rect 311 63 349 79
rect 383 147 399 181
rect 433 147 449 181
rect 383 107 449 147
rect 383 73 399 107
rect 433 73 449 107
rect 383 17 449 73
rect 483 111 521 187
rect 483 77 485 111
rect 519 77 521 111
rect 483 61 521 77
rect 555 174 571 208
rect 605 174 621 208
rect 555 111 621 174
rect 555 77 571 111
rect 605 77 621 111
rect 555 17 621 77
rect 655 187 657 221
rect 691 187 693 221
rect 827 221 865 242
rect 999 251 1049 272
rect 1485 251 1519 384
rect 655 111 693 187
rect 655 77 657 111
rect 691 77 693 111
rect 655 61 693 77
rect 727 174 743 208
rect 777 174 793 208
rect 727 111 793 174
rect 727 77 743 111
rect 777 77 793 111
rect 727 17 793 77
rect 827 187 829 221
rect 863 187 865 221
rect 827 111 865 187
rect 827 77 829 111
rect 863 77 865 111
rect 827 61 865 77
rect 899 222 965 238
rect 899 188 915 222
rect 949 188 965 222
rect 899 111 965 188
rect 899 77 915 111
rect 949 77 965 111
rect 899 17 965 77
rect 999 221 1519 251
rect 999 187 1001 221
rect 1035 217 1173 221
rect 1035 187 1037 217
rect 999 111 1037 187
rect 1171 187 1173 217
rect 1207 217 1345 221
rect 1207 187 1209 217
rect 999 77 1001 111
rect 1035 77 1037 111
rect 999 61 1037 77
rect 1071 149 1087 183
rect 1121 149 1137 183
rect 1071 111 1137 149
rect 1071 77 1087 111
rect 1121 77 1137 111
rect 1071 17 1137 77
rect 1171 111 1209 187
rect 1343 187 1345 217
rect 1379 217 1519 221
rect 1379 187 1381 217
rect 1171 77 1173 111
rect 1207 77 1209 111
rect 1171 61 1209 77
rect 1243 149 1259 183
rect 1293 149 1309 183
rect 1243 111 1309 149
rect 1243 77 1259 111
rect 1293 77 1309 111
rect 1243 17 1309 77
rect 1343 111 1381 187
rect 1343 77 1345 111
rect 1379 77 1381 111
rect 1343 61 1381 77
rect 1415 149 1431 183
rect 1465 149 1481 183
rect 1415 111 1481 149
rect 1415 77 1431 111
rect 1465 77 1481 111
rect 1415 17 1481 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor2_8
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5301972
string GDS_START 5289406
<< end >>
