magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 1 193 682 247
rect 1410 235 1602 241
rect 990 193 1602 235
rect 1 49 1602 193
rect 0 0 1632 49
<< scnmos >>
rect 80 53 110 221
rect 237 137 267 221
rect 315 137 345 221
rect 401 137 431 221
rect 487 137 517 221
rect 573 137 603 221
rect 788 83 818 167
rect 875 83 905 167
rect 964 83 994 167
rect 1096 125 1126 209
rect 1182 125 1212 209
rect 1260 125 1290 209
rect 1374 125 1404 209
rect 1489 47 1519 215
<< scpmoshvt >>
rect 82 367 112 619
rect 201 457 231 541
rect 301 457 331 541
rect 387 457 417 541
rect 473 457 503 541
rect 591 457 621 541
rect 824 411 854 495
rect 916 411 946 495
rect 1002 411 1032 495
rect 1088 411 1118 495
rect 1182 411 1212 495
rect 1260 411 1290 495
rect 1374 411 1404 495
rect 1522 367 1552 619
<< ndiff >>
rect 27 209 80 221
rect 27 175 35 209
rect 69 175 80 209
rect 27 101 80 175
rect 27 67 35 101
rect 69 67 80 101
rect 27 53 80 67
rect 110 193 237 221
rect 110 159 121 193
rect 155 159 192 193
rect 226 159 237 193
rect 110 137 237 159
rect 267 137 315 221
rect 345 196 401 221
rect 345 162 356 196
rect 390 162 401 196
rect 345 137 401 162
rect 431 196 487 221
rect 431 162 442 196
rect 476 162 487 196
rect 431 137 487 162
rect 517 196 573 221
rect 517 162 528 196
rect 562 162 573 196
rect 517 137 573 162
rect 603 196 656 221
rect 603 162 614 196
rect 648 162 656 196
rect 603 137 656 162
rect 110 99 163 137
rect 110 65 121 99
rect 155 65 163 99
rect 110 53 163 65
rect 1436 209 1489 215
rect 1016 195 1096 209
rect 1016 167 1049 195
rect 735 143 788 167
rect 735 109 743 143
rect 777 109 788 143
rect 735 83 788 109
rect 818 143 875 167
rect 818 109 829 143
rect 863 109 875 143
rect 818 83 875 109
rect 905 125 964 167
rect 905 91 919 125
rect 953 91 964 125
rect 905 83 964 91
rect 994 161 1049 167
rect 1083 161 1096 195
rect 994 127 1096 161
rect 994 93 1005 127
rect 1039 125 1096 127
rect 1126 183 1182 209
rect 1126 149 1137 183
rect 1171 149 1182 183
rect 1126 125 1182 149
rect 1212 125 1260 209
rect 1290 125 1374 209
rect 1404 127 1489 209
rect 1404 125 1444 127
rect 1039 93 1074 125
rect 994 83 1074 93
rect 1436 93 1444 125
rect 1478 93 1489 127
rect 1436 47 1489 93
rect 1519 188 1576 215
rect 1519 154 1534 188
rect 1568 154 1576 188
rect 1519 101 1576 154
rect 1519 67 1534 101
rect 1568 67 1576 101
rect 1519 47 1576 67
<< pdiff >>
rect 29 599 82 619
rect 29 565 37 599
rect 71 565 82 599
rect 29 503 82 565
rect 29 469 37 503
rect 71 469 82 503
rect 29 413 82 469
rect 29 379 37 413
rect 71 379 82 413
rect 29 367 82 379
rect 112 570 169 619
rect 112 536 127 570
rect 161 541 169 570
rect 518 568 576 576
rect 518 541 530 568
rect 161 536 201 541
rect 112 457 201 536
rect 231 457 301 541
rect 331 515 387 541
rect 331 481 342 515
rect 376 481 387 515
rect 331 457 387 481
rect 417 515 473 541
rect 417 481 428 515
rect 462 481 473 515
rect 417 457 473 481
rect 503 534 530 541
rect 564 541 576 568
rect 564 534 591 541
rect 503 457 591 534
rect 621 516 674 541
rect 621 482 632 516
rect 666 482 674 516
rect 621 457 674 482
rect 112 367 169 457
rect 1465 571 1522 619
rect 1465 537 1473 571
rect 1507 537 1522 571
rect 1465 495 1522 537
rect 771 470 824 495
rect 771 436 779 470
rect 813 436 824 470
rect 771 411 824 436
rect 854 470 916 495
rect 854 436 871 470
rect 905 436 916 470
rect 854 411 916 436
rect 946 478 1002 495
rect 946 444 957 478
rect 991 444 1002 478
rect 946 411 1002 444
rect 1032 470 1088 495
rect 1032 436 1043 470
rect 1077 436 1088 470
rect 1032 411 1088 436
rect 1118 470 1182 495
rect 1118 436 1137 470
rect 1171 436 1182 470
rect 1118 411 1182 436
rect 1212 411 1260 495
rect 1290 411 1374 495
rect 1404 411 1522 495
rect 1465 403 1522 411
rect 1472 367 1522 403
rect 1552 599 1605 619
rect 1552 565 1563 599
rect 1597 565 1605 599
rect 1552 505 1605 565
rect 1552 471 1563 505
rect 1597 471 1605 505
rect 1552 413 1605 471
rect 1552 379 1563 413
rect 1597 379 1605 413
rect 1552 367 1605 379
<< ndiffc >>
rect 35 175 69 209
rect 35 67 69 101
rect 121 159 155 193
rect 192 159 226 193
rect 356 162 390 196
rect 442 162 476 196
rect 528 162 562 196
rect 614 162 648 196
rect 121 65 155 99
rect 743 109 777 143
rect 829 109 863 143
rect 919 91 953 125
rect 1049 161 1083 195
rect 1005 93 1039 127
rect 1137 149 1171 183
rect 1444 93 1478 127
rect 1534 154 1568 188
rect 1534 67 1568 101
<< pdiffc >>
rect 37 565 71 599
rect 37 469 71 503
rect 37 379 71 413
rect 127 536 161 570
rect 342 481 376 515
rect 428 481 462 515
rect 530 534 564 568
rect 632 482 666 516
rect 1473 537 1507 571
rect 779 436 813 470
rect 871 436 905 470
rect 957 444 991 478
rect 1043 436 1077 470
rect 1137 436 1171 470
rect 1563 565 1597 599
rect 1563 471 1597 505
rect 1563 379 1597 413
<< poly >>
rect 82 619 112 645
rect 387 609 739 639
rect 1522 619 1552 645
rect 201 541 231 567
rect 301 541 331 567
rect 387 541 417 609
rect 709 593 739 609
rect 473 541 503 567
rect 591 541 621 567
rect 709 563 1212 593
rect 82 309 112 367
rect 201 325 231 457
rect 301 442 331 457
rect 387 442 417 457
rect 301 412 345 442
rect 387 412 431 442
rect 201 309 267 325
rect 80 293 159 309
rect 80 259 109 293
rect 143 259 159 293
rect 201 275 217 309
rect 251 275 267 309
rect 201 259 267 275
rect 80 243 159 259
rect 80 221 110 243
rect 237 221 267 259
rect 315 221 345 412
rect 401 221 431 412
rect 473 425 503 457
rect 473 409 539 425
rect 473 375 489 409
rect 523 375 539 409
rect 473 359 539 375
rect 487 221 517 359
rect 591 285 621 457
rect 709 425 739 563
rect 824 495 854 521
rect 916 495 946 563
rect 1002 495 1032 521
rect 1088 495 1118 521
rect 1182 495 1212 563
rect 1260 495 1290 521
rect 1374 495 1404 521
rect 673 409 739 425
rect 673 375 689 409
rect 723 375 739 409
rect 824 396 854 411
rect 673 359 739 375
rect 803 366 854 396
rect 803 285 833 366
rect 916 326 946 411
rect 573 269 833 285
rect 573 255 706 269
rect 573 221 603 255
rect 690 235 706 255
rect 740 235 783 269
rect 817 235 833 269
rect 690 219 833 235
rect 875 296 946 326
rect 690 207 818 219
rect 237 111 267 137
rect 315 63 345 137
rect 401 111 431 137
rect 487 111 517 137
rect 573 63 603 137
rect 690 63 720 207
rect 788 167 818 207
rect 875 167 905 296
rect 1002 254 1032 411
rect 1088 355 1118 411
rect 1074 339 1140 355
rect 1074 305 1090 339
rect 1124 305 1140 339
rect 1074 289 1140 305
rect 964 224 1032 254
rect 964 167 994 224
rect 1096 209 1126 289
rect 1182 209 1212 411
rect 1260 365 1290 411
rect 1374 371 1404 411
rect 1260 349 1326 365
rect 1260 315 1276 349
rect 1310 315 1326 349
rect 1260 281 1326 315
rect 1260 247 1276 281
rect 1310 247 1326 281
rect 1260 231 1326 247
rect 1374 355 1440 371
rect 1374 321 1390 355
rect 1424 321 1440 355
rect 1374 287 1440 321
rect 1522 304 1552 367
rect 1374 253 1390 287
rect 1424 253 1440 287
rect 1374 237 1440 253
rect 1482 288 1552 304
rect 1482 254 1498 288
rect 1532 254 1552 288
rect 1482 238 1552 254
rect 1260 209 1290 231
rect 1374 209 1404 237
rect 1489 215 1519 238
rect 1096 99 1126 125
rect 1182 99 1212 125
rect 1260 99 1290 125
rect 80 27 110 53
rect 315 33 720 63
rect 788 57 818 83
rect 875 57 905 83
rect 964 51 994 83
rect 1374 51 1404 125
rect 964 21 1404 51
rect 1489 21 1519 47
<< polycont >>
rect 109 259 143 293
rect 217 275 251 309
rect 489 375 523 409
rect 689 375 723 409
rect 706 235 740 269
rect 783 235 817 269
rect 1090 305 1124 339
rect 1276 315 1310 349
rect 1276 247 1310 281
rect 1390 321 1424 355
rect 1390 253 1424 287
rect 1498 254 1532 288
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 17 599 75 615
rect 17 565 37 599
rect 71 565 75 599
rect 17 503 75 565
rect 111 570 177 649
rect 111 536 127 570
rect 161 536 177 570
rect 111 528 177 536
rect 514 568 580 649
rect 514 534 530 568
rect 564 534 580 568
rect 17 469 37 503
rect 71 469 75 503
rect 326 515 384 531
rect 326 494 342 515
rect 17 413 75 469
rect 17 379 37 413
rect 71 379 75 413
rect 17 363 75 379
rect 111 481 342 494
rect 376 481 384 515
rect 111 460 384 481
rect 418 515 478 532
rect 514 528 580 534
rect 418 481 428 515
rect 462 494 478 515
rect 616 516 667 532
rect 616 494 632 516
rect 462 482 632 494
rect 666 482 667 516
rect 462 481 667 482
rect 418 460 667 481
rect 17 209 73 363
rect 111 309 159 460
rect 107 293 159 309
rect 107 259 109 293
rect 143 259 159 293
rect 201 424 269 426
rect 201 390 223 424
rect 257 390 269 424
rect 201 309 269 390
rect 201 275 217 309
rect 251 275 269 309
rect 201 259 269 275
rect 340 339 384 460
rect 473 424 557 426
rect 701 424 743 588
rect 473 409 511 424
rect 473 375 489 409
rect 545 390 557 424
rect 523 375 557 390
rect 473 373 557 375
rect 673 409 743 424
rect 777 470 824 649
rect 969 494 1007 649
rect 1457 571 1523 649
rect 1457 537 1473 571
rect 1507 537 1523 571
rect 1457 528 1523 537
rect 1559 599 1615 615
rect 1559 565 1563 599
rect 1597 565 1615 599
rect 1559 505 1615 565
rect 777 436 779 470
rect 813 436 824 470
rect 777 420 824 436
rect 858 470 907 486
rect 858 436 871 470
rect 905 436 907 470
rect 941 478 1007 494
rect 941 444 957 478
rect 991 444 1007 478
rect 941 441 1007 444
rect 1041 470 1087 486
rect 673 375 689 409
rect 723 375 743 409
rect 673 373 743 375
rect 858 407 907 436
rect 1041 436 1043 470
rect 1077 436 1087 470
rect 1041 407 1087 436
rect 1121 470 1525 494
rect 1121 436 1137 470
rect 1171 460 1525 470
rect 1171 436 1175 460
rect 1121 420 1175 436
rect 1364 424 1424 426
rect 858 373 1087 407
rect 1364 390 1375 424
rect 1409 390 1424 424
rect 1183 349 1326 365
rect 340 305 1090 339
rect 1124 305 1140 339
rect 1183 315 1276 349
rect 1310 315 1326 349
rect 107 243 159 259
rect 17 175 35 209
rect 69 175 73 209
rect 17 101 73 175
rect 17 67 35 101
rect 69 67 73 101
rect 17 51 73 67
rect 107 193 240 209
rect 107 159 121 193
rect 155 159 192 193
rect 226 159 240 193
rect 107 99 240 159
rect 340 196 397 305
rect 1183 281 1326 315
rect 1183 271 1276 281
rect 340 162 356 196
rect 390 162 397 196
rect 340 146 397 162
rect 431 237 656 271
rect 431 196 478 237
rect 431 162 442 196
rect 476 162 478 196
rect 431 146 478 162
rect 512 196 578 203
rect 512 162 528 196
rect 562 162 578 196
rect 107 65 121 99
rect 155 65 240 99
rect 107 17 240 65
rect 512 17 578 162
rect 612 196 656 237
rect 690 269 1276 271
rect 690 235 706 269
rect 740 235 783 269
rect 817 247 1276 269
rect 1310 247 1326 281
rect 817 237 1326 247
rect 1364 355 1424 390
rect 1364 321 1390 355
rect 1364 287 1424 321
rect 1364 253 1390 287
rect 1364 237 1424 253
rect 1458 304 1525 460
rect 1559 471 1563 505
rect 1597 471 1615 505
rect 1559 413 1615 471
rect 1559 379 1563 413
rect 1597 379 1615 413
rect 1559 363 1615 379
rect 1458 288 1532 304
rect 1458 254 1498 288
rect 1458 238 1532 254
rect 817 235 1099 237
rect 690 233 1099 235
rect 690 219 787 233
rect 1458 203 1494 238
rect 1568 204 1615 363
rect 612 162 614 196
rect 648 162 656 196
rect 612 146 656 162
rect 821 195 1099 199
rect 821 165 1049 195
rect 727 143 787 159
rect 727 109 743 143
rect 777 109 787 143
rect 727 17 787 109
rect 821 143 869 165
rect 821 109 829 143
rect 863 109 869 143
rect 1003 161 1049 165
rect 1083 161 1099 195
rect 821 93 869 109
rect 903 125 969 131
rect 903 91 919 125
rect 953 91 969 125
rect 903 17 969 91
rect 1003 127 1099 161
rect 1133 183 1494 203
rect 1133 149 1137 183
rect 1171 169 1494 183
rect 1528 188 1615 204
rect 1171 149 1394 169
rect 1133 133 1394 149
rect 1528 154 1534 188
rect 1568 154 1615 188
rect 1003 93 1005 127
rect 1039 93 1099 127
rect 1003 77 1099 93
rect 1428 127 1494 135
rect 1428 93 1444 127
rect 1478 93 1494 127
rect 1428 17 1494 93
rect 1528 101 1615 154
rect 1528 67 1534 101
rect 1568 67 1615 101
rect 1528 51 1615 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 223 390 257 424
rect 511 409 545 424
rect 511 390 523 409
rect 523 390 545 409
rect 1375 390 1409 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 499 424 557 430
rect 499 421 511 424
rect 257 393 511 421
rect 257 390 269 393
rect 211 384 269 390
rect 499 390 511 393
rect 545 421 557 424
rect 1363 424 1421 430
rect 1363 421 1375 424
rect 545 393 1375 421
rect 545 390 557 393
rect 499 384 557 390
rect 1363 390 1375 393
rect 1409 390 1421 424
rect 1363 384 1421 390
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fa_1
flabel metal1 s 223 390 257 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1567 94 1601 128 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2457786
string GDS_START 2445194
<< end >>
