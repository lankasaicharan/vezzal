magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1288 -1260 11504 1935
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_0
timestamp 1627201311
transform 1 0 1656 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_1
timestamp 1627201311
transform 1 0 3368 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_2
timestamp 1627201311
transform 1 0 5080 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_3
timestamp 1627201311
transform 1 0 6792 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_4
timestamp 1627201311
transform 1 0 8504 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_0
timestamp 1627201311
transform 1 0 800 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_1
timestamp 1627201311
transform 1 0 2512 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_2
timestamp 1627201311
transform 1 0 4224 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_3
timestamp 1627201311
transform 1 0 5936 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_4
timestamp 1627201311
transform 1 0 7648 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_5
timestamp 1627201311
transform 1 0 9360 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808338  sky130_fd_pr__hvdfl1sd__example_55959141808338_0
timestamp 1627201311
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808338  sky130_fd_pr__hvdfl1sd__example_55959141808338_1
timestamp 1627201311
transform 1 0 10216 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 10244 675 10244 675 0 FreeSans 300 0 0 0 S
flabel comment s 9388 675 9388 675 0 FreeSans 300 0 0 0 D
flabel comment s 8532 675 8532 675 0 FreeSans 300 0 0 0 S
flabel comment s 7676 675 7676 675 0 FreeSans 300 0 0 0 D
flabel comment s 6820 675 6820 675 0 FreeSans 300 0 0 0 S
flabel comment s 5964 675 5964 675 0 FreeSans 300 0 0 0 D
flabel comment s 5108 675 5108 675 0 FreeSans 300 0 0 0 S
flabel comment s 4252 675 4252 675 0 FreeSans 300 0 0 0 D
flabel comment s 3396 675 3396 675 0 FreeSans 300 0 0 0 S
flabel comment s 2540 675 2540 675 0 FreeSans 300 0 0 0 D
flabel comment s 1684 675 1684 675 0 FreeSans 300 0 0 0 S
flabel comment s 828 675 828 675 0 FreeSans 300 0 0 0 D
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 5045048
string GDS_START 5038308
<< end >>
