magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1250 -1208 3090 2438
<< pwell >>
rect 10 100 1768 1172
<< mvnmos >>
rect 89 1062 1689 1146
rect 89 850 1689 934
rect 89 702 1689 786
rect 89 488 1689 572
rect 89 340 1689 424
rect 89 126 1689 210
<< mvndiff >>
rect 36 1134 89 1146
rect 36 1100 44 1134
rect 78 1100 89 1134
rect 36 1062 89 1100
rect 1689 1134 1742 1146
rect 1689 1100 1700 1134
rect 1734 1100 1742 1134
rect 1689 1062 1742 1100
rect 36 896 89 934
rect 36 862 44 896
rect 78 862 89 896
rect 36 850 89 862
rect 1689 896 1742 934
rect 1689 862 1700 896
rect 1734 862 1742 896
rect 1689 850 1742 862
rect 36 774 89 786
rect 36 740 44 774
rect 78 740 89 774
rect 36 702 89 740
rect 1689 774 1742 786
rect 1689 740 1700 774
rect 1734 740 1742 774
rect 1689 702 1742 740
rect 36 534 89 572
rect 36 500 44 534
rect 78 500 89 534
rect 36 488 89 500
rect 1689 534 1742 572
rect 1689 500 1700 534
rect 1734 500 1742 534
rect 1689 488 1742 500
rect 36 412 89 424
rect 36 378 44 412
rect 78 378 89 412
rect 36 340 89 378
rect 1689 412 1742 424
rect 1689 378 1700 412
rect 1734 378 1742 412
rect 1689 340 1742 378
rect 36 172 89 210
rect 36 138 44 172
rect 78 138 89 172
rect 36 126 89 138
rect 1689 172 1742 210
rect 1689 138 1700 172
rect 1734 138 1742 172
rect 1689 126 1742 138
<< mvndiffc >>
rect 44 1100 78 1134
rect 1700 1100 1734 1134
rect 44 862 78 896
rect 1700 862 1734 896
rect 44 740 78 774
rect 1700 740 1734 774
rect 44 500 78 534
rect 1700 500 1734 534
rect 44 378 78 412
rect 1700 378 1734 412
rect 44 138 78 172
rect 1700 138 1734 172
<< poly >>
rect 89 1146 1689 1178
rect 89 1016 1689 1062
rect 89 982 105 1016
rect 139 982 175 1016
rect 209 982 245 1016
rect 279 982 315 1016
rect 349 982 385 1016
rect 419 982 455 1016
rect 489 982 525 1016
rect 559 982 595 1016
rect 629 982 665 1016
rect 699 982 735 1016
rect 769 982 805 1016
rect 839 982 875 1016
rect 909 982 945 1016
rect 979 982 1015 1016
rect 1049 982 1085 1016
rect 1119 982 1155 1016
rect 1189 982 1225 1016
rect 1259 982 1294 1016
rect 1328 982 1363 1016
rect 1397 982 1432 1016
rect 1466 982 1501 1016
rect 1535 982 1570 1016
rect 1604 982 1639 1016
rect 1673 982 1689 1016
rect 89 934 1689 982
rect 89 786 1689 850
rect 89 654 1689 702
rect 89 620 105 654
rect 139 620 175 654
rect 209 620 245 654
rect 279 620 315 654
rect 349 620 385 654
rect 419 620 455 654
rect 489 620 525 654
rect 559 620 595 654
rect 629 620 665 654
rect 699 620 735 654
rect 769 620 805 654
rect 839 620 875 654
rect 909 620 945 654
rect 979 620 1015 654
rect 1049 620 1085 654
rect 1119 620 1155 654
rect 1189 620 1225 654
rect 1259 620 1294 654
rect 1328 620 1363 654
rect 1397 620 1432 654
rect 1466 620 1501 654
rect 1535 620 1570 654
rect 1604 620 1639 654
rect 1673 620 1689 654
rect 89 572 1689 620
rect 89 424 1689 488
rect 89 292 1689 340
rect 89 258 105 292
rect 139 258 174 292
rect 208 258 243 292
rect 277 258 312 292
rect 346 258 380 292
rect 414 258 448 292
rect 482 258 516 292
rect 550 258 584 292
rect 618 258 652 292
rect 686 258 720 292
rect 754 258 788 292
rect 822 258 856 292
rect 890 258 924 292
rect 958 258 992 292
rect 1026 258 1060 292
rect 1094 258 1128 292
rect 1162 258 1196 292
rect 1230 258 1264 292
rect 1298 258 1332 292
rect 1366 258 1400 292
rect 1434 258 1468 292
rect 1502 258 1536 292
rect 1570 258 1604 292
rect 1638 258 1689 292
rect 89 210 1689 258
rect 89 94 1689 126
<< polycont >>
rect 105 982 139 1016
rect 175 982 209 1016
rect 245 982 279 1016
rect 315 982 349 1016
rect 385 982 419 1016
rect 455 982 489 1016
rect 525 982 559 1016
rect 595 982 629 1016
rect 665 982 699 1016
rect 735 982 769 1016
rect 805 982 839 1016
rect 875 982 909 1016
rect 945 982 979 1016
rect 1015 982 1049 1016
rect 1085 982 1119 1016
rect 1155 982 1189 1016
rect 1225 982 1259 1016
rect 1294 982 1328 1016
rect 1363 982 1397 1016
rect 1432 982 1466 1016
rect 1501 982 1535 1016
rect 1570 982 1604 1016
rect 1639 982 1673 1016
rect 105 620 139 654
rect 175 620 209 654
rect 245 620 279 654
rect 315 620 349 654
rect 385 620 419 654
rect 455 620 489 654
rect 525 620 559 654
rect 595 620 629 654
rect 665 620 699 654
rect 735 620 769 654
rect 805 620 839 654
rect 875 620 909 654
rect 945 620 979 654
rect 1015 620 1049 654
rect 1085 620 1119 654
rect 1155 620 1189 654
rect 1225 620 1259 654
rect 1294 620 1328 654
rect 1363 620 1397 654
rect 1432 620 1466 654
rect 1501 620 1535 654
rect 1570 620 1604 654
rect 1639 620 1673 654
rect 105 258 139 292
rect 174 258 208 292
rect 243 258 277 292
rect 312 258 346 292
rect 380 258 414 292
rect 448 258 482 292
rect 516 258 550 292
rect 584 258 618 292
rect 652 258 686 292
rect 720 258 754 292
rect 788 258 822 292
rect 856 258 890 292
rect 924 258 958 292
rect 992 258 1026 292
rect 1060 258 1094 292
rect 1128 258 1162 292
rect 1196 258 1230 292
rect 1264 258 1298 292
rect 1332 258 1366 292
rect 1400 258 1434 292
rect 1468 258 1502 292
rect 1536 258 1570 292
rect 1604 258 1638 292
<< locali >>
rect 78 1116 116 1150
rect 1662 1116 1700 1150
rect 44 1084 78 1100
rect 1700 1084 1734 1100
rect 89 982 105 1016
rect 139 982 175 1016
rect 209 982 245 1016
rect 279 982 315 1016
rect 349 982 385 1016
rect 419 982 455 1016
rect 489 982 525 1016
rect 559 982 595 1016
rect 629 982 665 1016
rect 699 982 735 1016
rect 769 982 805 1016
rect 839 982 875 1016
rect 909 982 945 1016
rect 979 982 1015 1016
rect 1049 982 1085 1016
rect 1119 982 1155 1016
rect 1189 982 1225 1016
rect 1259 982 1294 1016
rect 1328 982 1363 1016
rect 1397 982 1432 1016
rect 1466 982 1501 1016
rect 1535 982 1570 1016
rect 1604 982 1639 1016
rect 1673 982 1689 1016
rect 44 896 78 912
rect 78 846 116 880
rect 78 756 116 790
rect 44 724 78 740
rect 225 654 1558 982
rect 1700 896 1734 912
rect 1662 846 1700 880
rect 1662 756 1700 790
rect 1700 724 1734 740
rect 89 620 105 654
rect 139 620 175 654
rect 209 620 245 654
rect 279 620 315 654
rect 349 620 385 654
rect 419 620 455 654
rect 489 620 525 654
rect 559 620 595 654
rect 629 620 665 654
rect 699 620 735 654
rect 769 620 805 654
rect 839 620 875 654
rect 909 620 945 654
rect 979 620 1015 654
rect 1049 620 1085 654
rect 1119 620 1155 654
rect 1189 620 1225 654
rect 1259 620 1294 654
rect 1328 620 1363 654
rect 1397 620 1432 654
rect 1466 620 1501 654
rect 1535 620 1570 654
rect 1604 620 1639 654
rect 1673 620 1689 654
rect 44 534 78 550
rect 78 484 116 518
rect 78 394 116 428
rect 44 362 78 378
rect 225 292 1558 620
rect 1700 534 1734 550
rect 1662 484 1700 518
rect 1662 394 1700 428
rect 1734 378 1830 426
rect 89 258 105 292
rect 139 258 174 292
rect 208 258 243 292
rect 277 258 312 292
rect 346 258 380 292
rect 414 258 448 292
rect 482 258 516 292
rect 550 258 584 292
rect 618 258 652 292
rect 686 258 720 292
rect 754 258 788 292
rect 822 258 856 292
rect 890 258 924 292
rect 958 258 992 292
rect 1026 258 1060 292
rect 1094 258 1128 292
rect 1162 258 1196 292
rect 1230 258 1264 292
rect 1298 258 1332 292
rect 1366 258 1400 292
rect 1434 258 1468 292
rect 1502 258 1536 292
rect 1570 258 1604 292
rect 1638 258 1654 292
rect 44 172 78 188
rect 1700 172 1830 378
rect 78 122 116 156
rect 1734 138 1830 172
rect 1700 122 1830 138
<< viali >>
rect 44 1134 78 1150
rect 44 1116 78 1134
rect 116 1116 150 1150
rect 1628 1116 1662 1150
rect 1700 1134 1734 1150
rect 1700 1116 1734 1134
rect 44 862 78 880
rect 44 846 78 862
rect 116 846 150 880
rect 44 774 78 790
rect 44 756 78 774
rect 116 756 150 790
rect 1628 846 1662 880
rect 1700 862 1734 880
rect 1700 846 1734 862
rect 1628 756 1662 790
rect 1700 774 1734 790
rect 1700 756 1734 774
rect 44 500 78 518
rect 44 484 78 500
rect 116 484 150 518
rect 44 412 78 428
rect 44 394 78 412
rect 116 394 150 428
rect 1628 484 1662 518
rect 1700 500 1734 518
rect 1700 484 1734 500
rect 1628 394 1662 428
rect 1700 412 1734 428
rect 1700 394 1734 412
rect 44 138 78 156
rect 44 122 78 138
rect 116 122 150 156
<< metal1 >>
rect 38 1156 841 1162
rect 32 1150 841 1156
rect 32 1116 44 1150
rect 78 1116 116 1150
rect 150 1116 841 1150
rect 32 1110 841 1116
rect 38 1104 841 1110
rect 842 1105 843 1161
rect 883 1105 884 1161
rect 885 1156 1740 1162
tri 1740 1156 1746 1162 sw
rect 885 1150 1746 1156
rect 885 1116 1628 1150
rect 1662 1116 1700 1150
rect 1734 1116 1746 1150
rect 885 1110 1746 1116
rect 885 1104 1740 1110
tri 1740 1104 1746 1110 nw
rect 1694 892 1740 1104
rect 38 886 841 892
rect 32 880 841 886
rect 32 846 44 880
rect 78 846 116 880
rect 150 846 841 880
rect 32 840 841 846
rect 38 834 841 840
rect 842 835 843 891
rect 883 835 884 891
rect 885 886 1740 892
tri 1740 886 1746 892 sw
rect 885 880 1746 886
rect 885 846 1628 880
rect 1662 846 1700 880
rect 1734 846 1746 880
rect 885 840 1746 846
rect 885 834 1740 840
tri 1740 834 1746 840 nw
rect 38 802 84 834
rect 38 796 841 802
rect 32 790 841 796
rect 32 756 44 790
rect 78 756 116 790
rect 150 756 841 790
rect 32 750 841 756
rect 38 744 841 750
rect 842 745 843 801
rect 883 745 884 801
rect 885 790 1746 802
rect 885 756 1628 790
rect 1662 756 1700 790
rect 1734 756 1746 790
rect 885 744 1746 756
rect 1694 530 1746 744
rect 32 518 841 530
rect 32 484 44 518
rect 78 484 116 518
rect 150 484 841 518
rect 32 472 841 484
rect 842 473 843 529
rect 883 473 884 529
rect 885 518 1746 530
rect 885 484 1628 518
rect 1662 484 1700 518
rect 1734 484 1746 518
rect 885 472 1746 484
rect 32 440 84 472
rect 32 428 841 440
rect 32 394 44 428
rect 78 394 116 428
rect 150 394 841 428
rect 32 382 841 394
rect 842 383 843 439
rect 883 383 884 439
rect 885 434 1740 440
rect 885 428 1746 434
rect 885 394 1628 428
rect 1662 394 1700 428
rect 1734 394 1746 428
rect 885 388 1746 394
rect 885 382 1740 388
rect 1307 335 1365 382
rect 1308 333 1364 334
rect 1308 292 1364 293
rect 1307 239 1365 291
rect 38 162 221 168
rect 32 156 221 162
rect 32 122 44 156
rect 78 122 116 156
rect 150 122 221 156
rect 32 116 221 122
rect 38 110 221 116
rect 937 110 1694 168
rect 38 52 84 110
<< rmetal1 >>
rect 841 1161 843 1162
rect 841 1105 842 1161
rect 841 1104 843 1105
rect 883 1161 885 1162
rect 884 1105 885 1161
rect 883 1104 885 1105
rect 841 891 843 892
rect 841 835 842 891
rect 841 834 843 835
rect 883 891 885 892
rect 884 835 885 891
rect 883 834 885 835
rect 841 801 843 802
rect 841 745 842 801
rect 841 744 843 745
rect 883 801 885 802
rect 884 745 885 801
rect 883 744 885 745
rect 841 529 843 530
rect 841 473 842 529
rect 841 472 843 473
rect 883 529 885 530
rect 884 473 885 529
rect 883 472 885 473
rect 841 439 843 440
rect 841 383 842 439
rect 841 382 843 383
rect 883 439 885 440
rect 884 383 885 439
rect 883 382 885 383
rect 1307 334 1365 335
rect 1307 333 1308 334
rect 1364 333 1365 334
rect 1307 292 1308 293
rect 1364 292 1365 293
rect 1307 291 1365 292
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1627201311
transform 1 0 1628 0 1 1116
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1627201311
transform 1 0 1628 0 1 846
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1627201311
transform 1 0 44 0 1 1116
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1627201311
transform 1 0 44 0 1 846
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1627201311
transform 1 0 44 0 1 756
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1627201311
transform 1 0 44 0 1 484
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1627201311
transform 1 0 44 0 1 394
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1627201311
transform 1 0 1628 0 1 484
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1627201311
transform 1 0 1628 0 1 394
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1627201311
transform 1 0 1628 0 1 756
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1627201311
transform 1 0 44 0 1 122
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_5595914180895  sky130_fd_pr__nfet_01v8__example_5595914180895_0
timestamp 1627201311
transform 1 0 89 0 -1 424
box -28 0 1628 13
use sky130_fd_pr__nfet_01v8__example_5595914180895  sky130_fd_pr__nfet_01v8__example_5595914180895_1
timestamp 1627201311
transform 1 0 89 0 -1 786
box -28 0 1628 13
use sky130_fd_pr__nfet_01v8__example_5595914180895  sky130_fd_pr__nfet_01v8__example_5595914180895_2
timestamp 1627201311
transform 1 0 89 0 1 488
box -28 0 1628 13
use sky130_fd_pr__nfet_01v8__example_5595914180895  sky130_fd_pr__nfet_01v8__example_5595914180895_3
timestamp 1627201311
transform 1 0 89 0 1 850
box -28 0 1628 13
use sky130_fd_pr__nfet_01v8__example_5595914180895  sky130_fd_pr__nfet_01v8__example_5595914180895_4
timestamp 1627201311
transform 1 0 89 0 -1 1146
box -28 0 1628 13
use sky130_fd_pr__nfet_01v8__example_5595914180892  sky130_fd_pr__nfet_01v8__example_5595914180892_0
timestamp 1627201311
transform 1 0 89 0 1 126
box -28 0 1628 29
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_0
timestamp 1627201311
transform 0 1 1307 1 0 239
box 0 24 148 28
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_1
timestamp 1627201311
transform 1 0 789 0 1 382
box 0 24 148 28
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_2
timestamp 1627201311
transform 1 0 789 0 1 744
box 0 24 148 28
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_3
timestamp 1627201311
transform 1 0 789 0 -1 530
box 0 24 148 28
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_4
timestamp 1627201311
transform 1 0 789 0 1 1104
box 0 24 148 28
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_5
timestamp 1627201311
transform 1 0 789 0 -1 892
box 0 24 148 28
<< labels >>
flabel metal1 s 38 110 221 168 3 FreeSans 520 0 0 0 VGND
port 1 nsew
flabel metal1 s 38 1104 201 1162 3 FreeSans 520 0 0 0 OUT
port 2 nsew
flabel locali s 724 552 891 620 3 FreeSans 520 0 0 0 E_N
port 3 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 40067526
string GDS_START 40058978
<< end >>
