magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4466 1975
<< nwell >>
rect -38 331 3206 704
<< pwell >>
rect 1779 235 2137 279
rect 2612 235 3144 247
rect 37 49 541 229
rect 1489 191 3144 235
rect 1046 167 3144 191
rect 770 49 3144 167
rect 0 0 3168 49
<< scnmos >>
rect 116 119 146 203
rect 188 119 218 203
rect 274 119 304 203
rect 346 119 376 203
rect 432 119 462 203
rect 849 57 879 141
rect 935 57 965 141
rect 1199 81 1229 165
rect 1285 81 1315 165
rect 1357 81 1387 165
rect 1568 125 1598 209
rect 1640 125 1670 209
rect 1858 125 1888 253
rect 1930 125 1960 253
rect 2133 125 2163 209
rect 2218 125 2248 209
rect 2313 125 2343 209
rect 2421 125 2451 209
rect 2691 53 2721 221
rect 2777 53 2807 221
rect 2863 53 2893 221
rect 2949 53 2979 221
rect 3035 53 3065 221
<< scpmoshvt >>
rect 80 479 110 607
rect 166 479 196 607
rect 238 479 268 607
rect 346 479 376 607
rect 634 481 664 609
rect 845 491 875 619
rect 931 491 961 619
rect 1181 463 1211 547
rect 1267 463 1297 547
rect 1339 463 1369 547
rect 1479 463 1509 547
rect 1573 463 1603 547
rect 1721 379 1751 547
rect 1930 463 1960 547
rect 2035 379 2065 547
rect 2231 517 2261 601
rect 2317 517 2347 601
rect 2507 483 2537 567
rect 2697 367 2727 619
rect 2783 367 2813 619
rect 2869 367 2899 619
rect 2955 367 2985 619
rect 3041 367 3071 619
<< ndiff >>
rect 63 178 116 203
rect 63 144 71 178
rect 105 144 116 178
rect 63 119 116 144
rect 146 119 188 203
rect 218 178 274 203
rect 218 144 229 178
rect 263 144 274 178
rect 218 119 274 144
rect 304 119 346 203
rect 376 178 432 203
rect 376 144 387 178
rect 421 144 432 178
rect 376 119 432 144
rect 462 178 515 203
rect 462 144 473 178
rect 507 144 515 178
rect 462 119 515 144
rect 1805 220 1858 253
rect 1805 209 1813 220
rect 1515 197 1568 209
rect 1072 157 1199 165
rect 796 116 849 141
rect 796 82 804 116
rect 838 82 849 116
rect 796 57 849 82
rect 879 116 935 141
rect 879 82 890 116
rect 924 82 935 116
rect 879 57 935 82
rect 965 116 1018 141
rect 965 82 976 116
rect 1010 82 1018 116
rect 965 57 1018 82
rect 1072 123 1086 157
rect 1120 123 1199 157
rect 1072 81 1199 123
rect 1229 157 1285 165
rect 1229 123 1240 157
rect 1274 123 1285 157
rect 1229 81 1285 123
rect 1315 81 1357 165
rect 1387 140 1440 165
rect 1387 106 1398 140
rect 1432 106 1440 140
rect 1515 163 1523 197
rect 1557 163 1568 197
rect 1515 125 1568 163
rect 1598 125 1640 209
rect 1670 201 1813 209
rect 1670 167 1681 201
rect 1715 186 1813 201
rect 1847 186 1858 220
rect 1715 167 1858 186
rect 1670 125 1858 167
rect 1888 125 1930 253
rect 1960 217 2111 253
rect 1960 183 1974 217
rect 2008 183 2069 217
rect 2103 209 2111 217
rect 2638 209 2691 221
rect 2103 183 2133 209
rect 1960 125 2133 183
rect 2163 125 2218 209
rect 2248 125 2313 209
rect 2343 185 2421 209
rect 2343 151 2365 185
rect 2399 151 2421 185
rect 2343 125 2421 151
rect 2451 185 2504 209
rect 2451 151 2462 185
rect 2496 151 2504 185
rect 2451 125 2504 151
rect 2638 175 2646 209
rect 2680 175 2691 209
rect 1387 81 1440 106
rect 2638 101 2691 175
rect 2638 67 2646 101
rect 2680 67 2691 101
rect 2638 53 2691 67
rect 2721 210 2777 221
rect 2721 176 2732 210
rect 2766 176 2777 210
rect 2721 95 2777 176
rect 2721 61 2732 95
rect 2766 61 2777 95
rect 2721 53 2777 61
rect 2807 213 2863 221
rect 2807 179 2818 213
rect 2852 179 2863 213
rect 2807 101 2863 179
rect 2807 67 2818 101
rect 2852 67 2863 101
rect 2807 53 2863 67
rect 2893 181 2949 221
rect 2893 147 2904 181
rect 2938 147 2949 181
rect 2893 95 2949 147
rect 2893 61 2904 95
rect 2938 61 2949 95
rect 2893 53 2949 61
rect 2979 213 3035 221
rect 2979 179 2990 213
rect 3024 179 3035 213
rect 2979 101 3035 179
rect 2979 67 2990 101
rect 3024 67 3035 101
rect 2979 53 3035 67
rect 3065 181 3118 221
rect 3065 147 3076 181
rect 3110 147 3118 181
rect 3065 99 3118 147
rect 3065 65 3076 99
rect 3110 65 3118 99
rect 3065 53 3118 65
<< pdiff >>
rect 27 593 80 607
rect 27 559 35 593
rect 69 559 80 593
rect 27 525 80 559
rect 27 491 35 525
rect 69 491 80 525
rect 27 479 80 491
rect 110 575 166 607
rect 110 541 121 575
rect 155 541 166 575
rect 110 479 166 541
rect 196 479 238 607
rect 268 575 346 607
rect 268 541 290 575
rect 324 541 346 575
rect 268 479 346 541
rect 376 531 429 607
rect 376 497 387 531
rect 421 497 429 531
rect 376 479 429 497
rect 527 595 634 609
rect 527 561 535 595
rect 569 561 634 595
rect 527 481 634 561
rect 664 531 717 609
rect 664 497 675 531
rect 709 497 717 531
rect 664 481 717 497
rect 773 491 845 619
rect 875 609 931 619
rect 875 575 886 609
rect 920 575 931 609
rect 875 491 931 575
rect 961 599 1014 619
rect 961 565 972 599
rect 1006 565 1014 599
rect 961 491 1014 565
rect 773 455 823 491
rect 773 421 781 455
rect 815 421 823 455
rect 773 409 823 421
rect 1858 565 1908 577
rect 1074 509 1181 547
rect 1074 475 1082 509
rect 1116 475 1181 509
rect 1074 463 1181 475
rect 1211 511 1267 547
rect 1211 477 1222 511
rect 1256 477 1267 511
rect 1211 463 1267 477
rect 1297 463 1339 547
rect 1369 537 1479 547
rect 1369 503 1380 537
rect 1414 503 1479 537
rect 1369 463 1479 503
rect 1509 507 1573 547
rect 1509 473 1520 507
rect 1554 473 1573 507
rect 1509 463 1573 473
rect 1603 535 1721 547
rect 1603 501 1676 535
rect 1710 501 1721 535
rect 1603 463 1721 501
rect 1668 461 1721 463
rect 1668 427 1676 461
rect 1710 427 1721 461
rect 1668 379 1721 427
rect 1751 509 1804 547
rect 1751 475 1762 509
rect 1796 475 1804 509
rect 1751 379 1804 475
rect 1858 531 1866 565
rect 1900 547 1908 565
rect 1900 531 1930 547
rect 1858 463 1930 531
rect 1960 463 2035 547
rect 1982 425 2035 463
rect 1982 391 1990 425
rect 2024 391 2035 425
rect 1982 379 2035 391
rect 2065 499 2118 547
rect 2065 465 2076 499
rect 2110 465 2118 499
rect 2065 379 2118 465
rect 2178 589 2231 601
rect 2178 555 2186 589
rect 2220 555 2231 589
rect 2178 517 2231 555
rect 2261 576 2317 601
rect 2261 542 2272 576
rect 2306 542 2317 576
rect 2261 517 2317 542
rect 2347 576 2400 601
rect 2644 599 2697 619
rect 2347 542 2358 576
rect 2392 542 2400 576
rect 2347 517 2400 542
rect 2454 542 2507 567
rect 2454 508 2462 542
rect 2496 508 2507 542
rect 2454 483 2507 508
rect 2537 542 2590 567
rect 2537 508 2548 542
rect 2582 508 2590 542
rect 2537 483 2590 508
rect 2644 565 2652 599
rect 2686 565 2697 599
rect 2644 507 2697 565
rect 2644 473 2652 507
rect 2686 473 2697 507
rect 2644 413 2697 473
rect 2644 379 2652 413
rect 2686 379 2697 413
rect 2644 367 2697 379
rect 2727 611 2783 619
rect 2727 577 2738 611
rect 2772 577 2783 611
rect 2727 510 2783 577
rect 2727 476 2738 510
rect 2772 476 2783 510
rect 2727 413 2783 476
rect 2727 379 2738 413
rect 2772 379 2783 413
rect 2727 367 2783 379
rect 2813 599 2869 619
rect 2813 565 2824 599
rect 2858 565 2869 599
rect 2813 507 2869 565
rect 2813 473 2824 507
rect 2858 473 2869 507
rect 2813 409 2869 473
rect 2813 375 2824 409
rect 2858 375 2869 409
rect 2813 367 2869 375
rect 2899 611 2955 619
rect 2899 577 2910 611
rect 2944 577 2955 611
rect 2899 534 2955 577
rect 2899 500 2910 534
rect 2944 500 2955 534
rect 2899 455 2955 500
rect 2899 421 2910 455
rect 2944 421 2955 455
rect 2899 367 2955 421
rect 2985 599 3041 619
rect 2985 565 2996 599
rect 3030 565 3041 599
rect 2985 507 3041 565
rect 2985 473 2996 507
rect 3030 473 3041 507
rect 2985 409 3041 473
rect 2985 375 2996 409
rect 3030 375 3041 409
rect 2985 367 3041 375
rect 3071 607 3124 619
rect 3071 573 3082 607
rect 3116 573 3124 607
rect 3071 534 3124 573
rect 3071 500 3082 534
rect 3116 500 3124 534
rect 3071 455 3124 500
rect 3071 421 3082 455
rect 3116 421 3124 455
rect 3071 367 3124 421
<< ndiffc >>
rect 71 144 105 178
rect 229 144 263 178
rect 387 144 421 178
rect 473 144 507 178
rect 804 82 838 116
rect 890 82 924 116
rect 976 82 1010 116
rect 1086 123 1120 157
rect 1240 123 1274 157
rect 1398 106 1432 140
rect 1523 163 1557 197
rect 1681 167 1715 201
rect 1813 186 1847 220
rect 1974 183 2008 217
rect 2069 183 2103 217
rect 2365 151 2399 185
rect 2462 151 2496 185
rect 2646 175 2680 209
rect 2646 67 2680 101
rect 2732 176 2766 210
rect 2732 61 2766 95
rect 2818 179 2852 213
rect 2818 67 2852 101
rect 2904 147 2938 181
rect 2904 61 2938 95
rect 2990 179 3024 213
rect 2990 67 3024 101
rect 3076 147 3110 181
rect 3076 65 3110 99
<< pdiffc >>
rect 35 559 69 593
rect 35 491 69 525
rect 121 541 155 575
rect 290 541 324 575
rect 387 497 421 531
rect 535 561 569 595
rect 675 497 709 531
rect 886 575 920 609
rect 972 565 1006 599
rect 781 421 815 455
rect 1082 475 1116 509
rect 1222 477 1256 511
rect 1380 503 1414 537
rect 1520 473 1554 507
rect 1676 501 1710 535
rect 1676 427 1710 461
rect 1762 475 1796 509
rect 1866 531 1900 565
rect 1990 391 2024 425
rect 2076 465 2110 499
rect 2186 555 2220 589
rect 2272 542 2306 576
rect 2358 542 2392 576
rect 2462 508 2496 542
rect 2548 508 2582 542
rect 2652 565 2686 599
rect 2652 473 2686 507
rect 2652 379 2686 413
rect 2738 577 2772 611
rect 2738 476 2772 510
rect 2738 379 2772 413
rect 2824 565 2858 599
rect 2824 473 2858 507
rect 2824 375 2858 409
rect 2910 577 2944 611
rect 2910 500 2944 534
rect 2910 421 2944 455
rect 2996 565 3030 599
rect 2996 473 3030 507
rect 2996 375 3030 409
rect 3082 573 3116 607
rect 3082 500 3116 534
rect 3082 421 3116 455
<< poly >>
rect 80 607 110 633
rect 166 607 196 633
rect 238 607 268 633
rect 346 607 376 633
rect 634 609 664 635
rect 845 619 875 645
rect 931 619 961 645
rect 1029 615 2163 645
rect 80 359 110 479
rect 44 343 110 359
rect 44 309 60 343
rect 94 309 110 343
rect 166 333 196 479
rect 238 447 268 479
rect 238 431 304 447
rect 238 397 254 431
rect 288 397 304 431
rect 238 381 304 397
rect 346 381 376 479
rect 634 459 664 481
rect 634 429 717 459
rect 44 275 110 309
rect 160 303 218 333
rect 44 241 60 275
rect 94 255 110 275
rect 94 241 146 255
rect 44 225 146 241
rect 116 203 146 225
rect 188 203 218 303
rect 268 303 298 381
rect 346 365 605 381
rect 346 351 555 365
rect 268 273 304 303
rect 274 203 304 273
rect 346 203 376 351
rect 539 331 555 351
rect 589 331 605 365
rect 539 297 605 331
rect 539 263 555 297
rect 589 263 605 297
rect 539 247 605 263
rect 432 203 462 229
rect 687 228 717 429
rect 845 302 875 491
rect 931 455 961 491
rect 1029 455 1059 615
rect 1181 547 1211 573
rect 1267 547 1297 615
rect 1339 547 1369 573
rect 1479 547 1509 573
rect 1573 547 1603 573
rect 1721 547 1751 573
rect 931 439 1059 455
rect 931 405 947 439
rect 981 425 1059 439
rect 981 405 997 425
rect 931 389 997 405
rect 1181 393 1211 463
rect 1267 437 1297 463
rect 1339 397 1369 463
rect 827 286 893 302
rect 827 252 843 286
rect 877 252 893 286
rect 687 212 753 228
rect 687 178 703 212
rect 737 178 753 212
rect 687 144 753 178
rect 827 218 893 252
rect 827 184 843 218
rect 877 184 893 218
rect 967 217 997 389
rect 1136 377 1285 393
rect 1136 343 1152 377
rect 1186 343 1285 377
rect 1136 309 1285 343
rect 1339 381 1405 397
rect 1339 347 1355 381
rect 1389 347 1405 381
rect 1339 331 1405 347
rect 1136 275 1152 309
rect 1186 289 1285 309
rect 1186 275 1315 289
rect 1136 259 1315 275
rect 827 168 893 184
rect 935 187 1229 217
rect 116 93 146 119
rect 188 51 218 119
rect 274 93 304 119
rect 346 93 376 119
rect 432 51 462 119
rect 687 110 703 144
rect 737 110 753 144
rect 849 141 879 168
rect 935 141 965 187
rect 1199 165 1229 187
rect 1285 165 1315 259
rect 1375 253 1405 331
rect 1479 323 1509 463
rect 1573 364 1603 463
rect 1930 547 1960 573
rect 2035 547 2065 573
rect 1930 419 1960 463
rect 1872 403 1960 419
rect 1573 334 1670 364
rect 1465 307 1531 323
rect 1465 273 1481 307
rect 1515 286 1531 307
rect 1515 273 1598 286
rect 1465 256 1598 273
rect 1357 237 1423 253
rect 1357 203 1373 237
rect 1407 203 1423 237
rect 1568 209 1598 256
rect 1640 209 1670 334
rect 1721 341 1751 379
rect 1872 369 1888 403
rect 1922 369 1960 403
rect 1872 353 1960 369
rect 1721 325 1787 341
rect 1721 291 1737 325
rect 1771 305 1787 325
rect 1771 291 1888 305
rect 1721 275 1888 291
rect 1858 253 1888 275
rect 1930 253 1960 353
rect 2035 339 2065 379
rect 2133 339 2163 615
rect 2231 601 2261 627
rect 2317 601 2347 627
rect 2697 619 2727 645
rect 2783 619 2813 645
rect 2869 619 2899 645
rect 2955 619 2985 645
rect 3041 619 3071 645
rect 2507 567 2537 593
rect 2035 297 2163 339
rect 2231 297 2261 517
rect 2317 367 2347 517
rect 2507 451 2537 483
rect 2427 435 2537 451
rect 2427 401 2443 435
rect 2477 401 2537 435
rect 2427 367 2537 401
rect 2313 351 2379 367
rect 2313 317 2329 351
rect 2363 317 2379 351
rect 2427 345 2443 367
rect 2313 301 2379 317
rect 2421 333 2443 345
rect 2477 345 2537 367
rect 2697 345 2727 367
rect 2477 333 2727 345
rect 2783 335 2813 367
rect 2869 335 2899 367
rect 2955 335 2985 367
rect 3041 335 3071 367
rect 2421 315 2727 333
rect 2769 319 3071 335
rect 1357 187 1423 203
rect 1357 165 1387 187
rect 687 94 753 110
rect 687 51 717 94
rect 2133 209 2163 297
rect 2205 281 2271 297
rect 2205 247 2221 281
rect 2255 247 2271 281
rect 2205 231 2271 247
rect 2218 209 2248 231
rect 2313 209 2343 301
rect 2421 209 2451 315
rect 2691 221 2721 315
rect 2769 285 2785 319
rect 2819 285 2853 319
rect 2887 285 2921 319
rect 2955 285 3071 319
rect 2769 269 3071 285
rect 2777 221 2807 269
rect 2863 221 2893 269
rect 2949 221 2979 269
rect 3035 221 3065 269
rect 1568 99 1598 125
rect 1640 103 1670 125
rect 1640 87 1729 103
rect 1858 99 1888 125
rect 1930 99 1960 125
rect 2133 99 2163 125
rect 2218 99 2248 125
rect 2313 99 2343 125
rect 2421 99 2451 125
rect 188 21 717 51
rect 849 31 879 57
rect 935 31 965 57
rect 1199 55 1229 81
rect 1285 55 1315 81
rect 1357 55 1387 81
rect 1640 73 1679 87
rect 1663 53 1679 73
rect 1713 53 1729 87
rect 1663 37 1729 53
rect 2691 27 2721 53
rect 2777 27 2807 53
rect 2863 27 2893 53
rect 2949 27 2979 53
rect 3035 27 3065 53
<< polycont >>
rect 60 309 94 343
rect 254 397 288 431
rect 60 241 94 275
rect 555 331 589 365
rect 555 263 589 297
rect 947 405 981 439
rect 843 252 877 286
rect 703 178 737 212
rect 843 184 877 218
rect 1152 343 1186 377
rect 1355 347 1389 381
rect 1152 275 1186 309
rect 703 110 737 144
rect 1481 273 1515 307
rect 1373 203 1407 237
rect 1888 369 1922 403
rect 1737 291 1771 325
rect 2443 401 2477 435
rect 2329 317 2363 351
rect 2443 333 2477 367
rect 2221 247 2255 281
rect 2785 285 2819 319
rect 2853 285 2887 319
rect 2921 285 2955 319
rect 1679 53 1713 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 19 593 71 609
rect 19 559 35 593
rect 69 559 71 593
rect 19 525 71 559
rect 105 575 171 649
rect 105 541 121 575
rect 155 541 171 575
rect 105 533 171 541
rect 274 581 495 615
rect 274 575 340 581
rect 274 541 290 575
rect 324 541 340 575
rect 274 533 340 541
rect 19 491 35 525
rect 69 499 71 525
rect 374 531 427 547
rect 374 499 387 531
rect 69 497 387 499
rect 421 497 427 531
rect 69 491 427 497
rect 19 465 427 491
rect 461 511 495 581
rect 529 595 571 649
rect 529 561 535 595
rect 569 561 571 595
rect 529 545 571 561
rect 605 581 836 615
rect 605 511 639 581
rect 461 477 639 511
rect 673 531 725 547
rect 673 497 675 531
rect 709 497 725 531
rect 17 397 254 431
rect 288 397 451 431
rect 17 387 451 397
rect 144 374 451 387
rect 17 343 110 353
rect 17 309 60 343
rect 94 309 110 343
rect 17 275 110 309
rect 485 308 519 477
rect 673 420 725 497
rect 791 525 836 581
rect 870 609 922 649
rect 870 575 886 609
rect 920 575 922 609
rect 870 559 922 575
rect 956 599 1344 615
rect 956 565 972 599
rect 1006 565 1344 599
rect 956 561 1344 565
rect 956 559 1186 561
rect 791 509 1118 525
rect 791 491 1082 509
rect 1068 475 1082 491
rect 1116 475 1118 509
rect 17 241 60 275
rect 94 241 110 275
rect 17 228 110 241
rect 213 243 519 308
rect 553 386 725 420
rect 765 455 997 457
rect 765 421 781 455
rect 815 439 997 455
rect 815 421 947 439
rect 765 405 947 421
rect 981 405 997 439
rect 773 389 997 405
rect 553 365 605 386
rect 553 331 555 365
rect 589 331 605 365
rect 553 297 605 331
rect 553 263 555 297
rect 589 263 605 297
rect 55 178 121 194
rect 55 144 71 178
rect 105 144 121 178
rect 55 17 121 144
rect 213 178 279 243
rect 553 194 605 263
rect 213 144 229 178
rect 263 144 279 178
rect 213 128 279 144
rect 371 178 437 194
rect 371 144 387 178
rect 421 144 437 178
rect 371 17 437 144
rect 471 178 605 194
rect 471 144 473 178
rect 507 144 605 178
rect 471 128 605 144
rect 687 212 739 352
rect 687 178 703 212
rect 737 178 739 212
rect 687 144 739 178
rect 687 110 703 144
rect 737 110 739 144
rect 687 78 739 110
rect 773 132 807 389
rect 841 286 956 355
rect 841 252 843 286
rect 877 252 956 286
rect 841 218 956 252
rect 841 184 843 218
rect 877 184 956 218
rect 841 166 956 184
rect 1068 161 1118 475
rect 1152 393 1186 559
rect 1220 511 1274 527
rect 1220 477 1222 511
rect 1256 477 1274 511
rect 1220 461 1274 477
rect 1152 377 1204 393
rect 1186 343 1204 377
rect 1152 309 1204 343
rect 1186 275 1204 309
rect 1152 259 1204 275
rect 1068 157 1136 161
rect 773 116 848 132
rect 773 82 804 116
rect 838 82 848 116
rect 773 66 848 82
rect 882 116 932 132
rect 882 82 890 116
rect 924 82 932 116
rect 882 17 932 82
rect 966 116 1014 132
rect 1068 123 1086 157
rect 1120 123 1136 157
rect 1068 119 1136 123
rect 966 82 976 116
rect 1010 85 1014 116
rect 1170 85 1204 259
rect 1238 309 1274 461
rect 1308 453 1344 561
rect 1378 537 1416 649
rect 1378 503 1380 537
rect 1414 503 1416 537
rect 1378 487 1416 503
rect 1450 557 1624 591
rect 1450 453 1484 557
rect 1308 419 1484 453
rect 1518 507 1556 523
rect 1518 473 1520 507
rect 1554 473 1556 507
rect 1518 385 1556 473
rect 1339 381 1556 385
rect 1339 347 1355 381
rect 1389 347 1556 381
rect 1590 393 1624 557
rect 1660 535 1726 649
rect 1660 501 1676 535
rect 1710 501 1726 535
rect 1850 589 2224 605
rect 1850 565 2186 589
rect 1850 531 1866 565
rect 1900 555 2186 565
rect 2220 555 2224 589
rect 1900 539 2224 555
rect 2268 576 2310 649
rect 2268 542 2272 576
rect 2306 542 2310 576
rect 1900 531 1916 539
rect 1850 529 1916 531
rect 1660 461 1726 501
rect 1660 427 1676 461
rect 1710 427 1726 461
rect 1760 509 1800 527
rect 2268 526 2310 542
rect 2354 576 2412 592
rect 2354 542 2358 576
rect 2392 542 2412 576
rect 1760 475 1762 509
rect 1796 495 1800 509
rect 2060 499 2126 505
rect 2060 495 2076 499
rect 1796 475 2076 495
rect 1760 465 2076 475
rect 2110 465 2126 499
rect 1760 459 2126 465
rect 2354 451 2412 542
rect 2446 542 2505 649
rect 2632 599 2696 615
rect 2632 565 2652 599
rect 2686 565 2696 599
rect 2446 508 2462 542
rect 2496 508 2505 542
rect 2446 492 2505 508
rect 2539 542 2598 558
rect 2539 508 2548 542
rect 2582 508 2598 542
rect 2354 435 2493 451
rect 2354 425 2443 435
rect 1872 393 1888 403
rect 1590 369 1888 393
rect 1922 369 1938 403
rect 1590 359 1938 369
rect 1974 391 1990 425
rect 2024 401 2443 425
rect 2477 401 2493 435
rect 2024 391 2493 401
rect 1974 387 2493 391
rect 1339 343 1556 347
rect 1721 309 1737 325
rect 1238 307 1737 309
rect 1238 273 1481 307
rect 1515 291 1737 307
rect 1771 291 1787 325
rect 1515 273 1787 291
rect 1238 271 1787 273
rect 1238 173 1274 271
rect 1357 203 1373 237
rect 1407 203 1557 237
rect 1357 197 1557 203
rect 1357 190 1523 197
rect 1238 157 1290 173
rect 1238 123 1240 157
rect 1274 123 1290 157
rect 1519 163 1523 190
rect 1238 107 1290 123
rect 1382 140 1448 156
rect 1519 147 1557 163
rect 1593 220 1863 237
rect 1593 201 1813 220
rect 1593 167 1681 201
rect 1715 186 1813 201
rect 1847 186 1863 220
rect 1715 167 1863 186
rect 1974 217 2103 387
rect 2422 367 2493 387
rect 2008 183 2069 217
rect 1974 167 2103 183
rect 2137 351 2379 353
rect 2137 317 2329 351
rect 2363 317 2379 351
rect 2422 333 2443 367
rect 2477 333 2493 367
rect 2422 317 2493 333
rect 1010 82 1204 85
rect 966 51 1204 82
rect 1382 106 1398 140
rect 1432 106 1448 140
rect 1382 17 1448 106
rect 1593 17 1627 167
rect 2137 133 2171 317
rect 2539 283 2598 508
rect 2205 281 2598 283
rect 2205 247 2221 281
rect 2255 247 2598 281
rect 2632 507 2696 565
rect 2632 473 2652 507
rect 2686 473 2696 507
rect 2632 413 2696 473
rect 2632 379 2652 413
rect 2686 379 2696 413
rect 2632 319 2696 379
rect 2730 611 2780 649
rect 2730 577 2738 611
rect 2772 577 2780 611
rect 2730 510 2780 577
rect 2730 476 2738 510
rect 2772 476 2780 510
rect 2730 413 2780 476
rect 2730 379 2738 413
rect 2772 379 2780 413
rect 2730 363 2780 379
rect 2814 599 2860 615
rect 2814 565 2824 599
rect 2858 565 2860 599
rect 2814 507 2860 565
rect 2814 473 2824 507
rect 2858 473 2860 507
rect 2814 409 2860 473
rect 2894 611 2960 649
rect 2894 577 2910 611
rect 2944 577 2960 611
rect 2894 534 2960 577
rect 2894 500 2910 534
rect 2944 500 2960 534
rect 2894 455 2960 500
rect 2894 421 2910 455
rect 2944 421 2960 455
rect 2994 599 3032 615
rect 2994 565 2996 599
rect 3030 565 3032 599
rect 2994 507 3032 565
rect 2994 473 2996 507
rect 3030 473 3032 507
rect 2814 375 2824 409
rect 2858 387 2860 409
rect 2994 409 3032 473
rect 3066 607 3132 649
rect 3066 573 3082 607
rect 3116 573 3132 607
rect 3066 534 3132 573
rect 3066 500 3082 534
rect 3116 500 3132 534
rect 3066 455 3132 500
rect 3066 421 3082 455
rect 3116 421 3132 455
rect 2994 387 2996 409
rect 2858 375 2996 387
rect 3030 387 3032 409
rect 3030 375 3137 387
rect 2814 353 3137 375
rect 2632 285 2785 319
rect 2819 285 2853 319
rect 2887 285 2921 319
rect 2955 285 2971 319
rect 2205 235 2512 247
rect 1661 87 2171 133
rect 1661 53 1679 87
rect 1713 53 2171 87
rect 1661 51 2171 53
rect 2349 185 2415 201
rect 2349 151 2365 185
rect 2399 151 2415 185
rect 2349 17 2415 151
rect 2453 185 2512 235
rect 2453 151 2462 185
rect 2496 151 2512 185
rect 2453 135 2512 151
rect 2632 209 2682 285
rect 3007 251 3137 353
rect 2632 175 2646 209
rect 2680 175 2682 209
rect 2632 101 2682 175
rect 2632 67 2646 101
rect 2680 67 2682 101
rect 2632 51 2682 67
rect 2716 210 2782 226
rect 2716 176 2732 210
rect 2766 176 2782 210
rect 2716 95 2782 176
rect 2716 61 2732 95
rect 2766 61 2782 95
rect 2716 17 2782 61
rect 2816 215 3137 251
rect 2816 213 2854 215
rect 2816 179 2818 213
rect 2852 179 2854 213
rect 2988 213 3026 215
rect 2816 101 2854 179
rect 2816 67 2818 101
rect 2852 67 2854 101
rect 2816 51 2854 67
rect 2888 147 2904 181
rect 2938 147 2954 181
rect 2888 95 2954 147
rect 2888 61 2904 95
rect 2938 61 2954 95
rect 2888 17 2954 61
rect 2988 179 2990 213
rect 3024 179 3026 213
rect 2988 101 3026 179
rect 2988 67 2990 101
rect 3024 67 3026 101
rect 2988 51 3026 67
rect 3060 147 3076 181
rect 3110 147 3126 181
rect 3060 99 3126 147
rect 3060 65 3076 99
rect 3110 65 3126 99
rect 3060 17 3126 65
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
<< metal1 >>
rect 0 683 3168 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 0 617 3168 649
rect 0 17 3168 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
rect 0 -49 3168 -17
<< labels >>
flabel pwell s 0 0 3168 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 3168 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfstp_4
flabel comment s 1385 301 1385 301 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 3168 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 3168 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 3007 242 3041 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3103 242 3137 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 1663 94 1697 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 1759 94 1793 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 1855 94 1889 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 1951 94 1985 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 2047 94 2081 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3168 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 132016
string GDS_START 110222
<< end >>
