magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 331 1958 704
<< pwell >>
rect 1 49 1907 157
rect 0 0 1920 49
<< scnmos >>
rect 86 47 116 131
rect 172 47 202 131
rect 258 47 288 131
rect 344 47 374 131
rect 508 47 538 131
rect 594 47 624 131
rect 680 47 710 131
rect 766 47 796 131
rect 852 47 882 131
rect 938 47 968 131
rect 1024 47 1054 131
rect 1110 47 1140 131
rect 1196 47 1226 131
rect 1282 47 1312 131
rect 1368 47 1398 131
rect 1454 47 1484 131
rect 1540 47 1570 131
rect 1626 47 1656 131
rect 1712 47 1742 131
rect 1798 47 1828 131
<< scpmoshvt >>
rect 86 367 116 619
rect 172 367 202 619
rect 258 367 288 619
rect 344 367 374 619
rect 508 367 538 619
rect 594 367 624 619
rect 680 367 710 619
rect 766 367 796 619
rect 852 367 882 619
rect 938 367 968 619
rect 1024 367 1054 619
rect 1110 367 1140 619
rect 1196 367 1226 619
rect 1282 367 1312 619
rect 1368 367 1398 619
rect 1454 367 1484 619
rect 1540 367 1570 619
rect 1626 367 1656 619
rect 1712 367 1742 619
rect 1798 367 1828 619
<< ndiff >>
rect 27 106 86 131
rect 27 72 41 106
rect 75 72 86 106
rect 27 47 86 72
rect 116 106 172 131
rect 116 72 127 106
rect 161 72 172 106
rect 116 47 172 72
rect 202 105 258 131
rect 202 71 213 105
rect 247 71 258 105
rect 202 47 258 71
rect 288 106 344 131
rect 288 72 299 106
rect 333 72 344 106
rect 288 47 344 72
rect 374 105 508 131
rect 374 71 385 105
rect 419 71 463 105
rect 497 71 508 105
rect 374 47 508 71
rect 538 105 594 131
rect 538 71 549 105
rect 583 71 594 105
rect 538 47 594 71
rect 624 105 680 131
rect 624 71 635 105
rect 669 71 680 105
rect 624 47 680 71
rect 710 105 766 131
rect 710 71 721 105
rect 755 71 766 105
rect 710 47 766 71
rect 796 105 852 131
rect 796 71 807 105
rect 841 71 852 105
rect 796 47 852 71
rect 882 105 938 131
rect 882 71 893 105
rect 927 71 938 105
rect 882 47 938 71
rect 968 105 1024 131
rect 968 71 979 105
rect 1013 71 1024 105
rect 968 47 1024 71
rect 1054 105 1110 131
rect 1054 71 1065 105
rect 1099 71 1110 105
rect 1054 47 1110 71
rect 1140 105 1196 131
rect 1140 71 1151 105
rect 1185 71 1196 105
rect 1140 47 1196 71
rect 1226 105 1282 131
rect 1226 71 1237 105
rect 1271 71 1282 105
rect 1226 47 1282 71
rect 1312 105 1368 131
rect 1312 71 1323 105
rect 1357 71 1368 105
rect 1312 47 1368 71
rect 1398 105 1454 131
rect 1398 71 1409 105
rect 1443 71 1454 105
rect 1398 47 1454 71
rect 1484 105 1540 131
rect 1484 71 1495 105
rect 1529 71 1540 105
rect 1484 47 1540 71
rect 1570 105 1626 131
rect 1570 71 1581 105
rect 1615 71 1626 105
rect 1570 47 1626 71
rect 1656 105 1712 131
rect 1656 71 1667 105
rect 1701 71 1712 105
rect 1656 47 1712 71
rect 1742 105 1798 131
rect 1742 71 1753 105
rect 1787 71 1798 105
rect 1742 47 1798 71
rect 1828 105 1881 131
rect 1828 71 1839 105
rect 1873 71 1881 105
rect 1828 47 1881 71
<< pdiff >>
rect 27 595 86 619
rect 27 561 41 595
rect 75 561 86 595
rect 27 509 86 561
rect 27 475 41 509
rect 75 475 86 509
rect 27 425 86 475
rect 27 391 41 425
rect 75 391 86 425
rect 27 367 86 391
rect 116 595 172 619
rect 116 561 127 595
rect 161 561 172 595
rect 116 509 172 561
rect 116 475 127 509
rect 161 475 172 509
rect 116 425 172 475
rect 116 391 127 425
rect 161 391 172 425
rect 116 367 172 391
rect 202 603 258 619
rect 202 569 213 603
rect 247 569 258 603
rect 202 525 258 569
rect 202 491 213 525
rect 247 491 258 525
rect 202 455 258 491
rect 202 421 213 455
rect 247 421 258 455
rect 202 367 258 421
rect 288 595 344 619
rect 288 561 299 595
rect 333 561 344 595
rect 288 509 344 561
rect 288 475 299 509
rect 333 475 344 509
rect 288 425 344 475
rect 288 391 299 425
rect 333 391 344 425
rect 288 367 344 391
rect 374 603 508 619
rect 374 569 385 603
rect 419 569 463 603
rect 497 569 508 603
rect 374 525 508 569
rect 374 491 385 525
rect 419 491 463 525
rect 497 491 508 525
rect 374 455 508 491
rect 374 421 385 455
rect 419 421 463 455
rect 497 421 508 455
rect 374 367 508 421
rect 538 595 594 619
rect 538 561 549 595
rect 583 561 594 595
rect 538 509 594 561
rect 538 475 549 509
rect 583 475 594 509
rect 538 425 594 475
rect 538 391 549 425
rect 583 391 594 425
rect 538 367 594 391
rect 624 595 680 619
rect 624 561 635 595
rect 669 561 680 595
rect 624 509 680 561
rect 624 475 635 509
rect 669 475 680 509
rect 624 425 680 475
rect 624 391 635 425
rect 669 391 680 425
rect 624 367 680 391
rect 710 595 766 619
rect 710 561 721 595
rect 755 561 766 595
rect 710 509 766 561
rect 710 475 721 509
rect 755 475 766 509
rect 710 425 766 475
rect 710 391 721 425
rect 755 391 766 425
rect 710 367 766 391
rect 796 595 852 619
rect 796 561 807 595
rect 841 561 852 595
rect 796 509 852 561
rect 796 475 807 509
rect 841 475 852 509
rect 796 425 852 475
rect 796 391 807 425
rect 841 391 852 425
rect 796 367 852 391
rect 882 595 938 619
rect 882 561 893 595
rect 927 561 938 595
rect 882 509 938 561
rect 882 475 893 509
rect 927 475 938 509
rect 882 425 938 475
rect 882 391 893 425
rect 927 391 938 425
rect 882 367 938 391
rect 968 595 1024 619
rect 968 561 979 595
rect 1013 561 1024 595
rect 968 509 1024 561
rect 968 475 979 509
rect 1013 475 1024 509
rect 968 425 1024 475
rect 968 391 979 425
rect 1013 391 1024 425
rect 968 367 1024 391
rect 1054 595 1110 619
rect 1054 561 1065 595
rect 1099 561 1110 595
rect 1054 509 1110 561
rect 1054 475 1065 509
rect 1099 475 1110 509
rect 1054 425 1110 475
rect 1054 391 1065 425
rect 1099 391 1110 425
rect 1054 367 1110 391
rect 1140 595 1196 619
rect 1140 561 1151 595
rect 1185 561 1196 595
rect 1140 509 1196 561
rect 1140 475 1151 509
rect 1185 475 1196 509
rect 1140 425 1196 475
rect 1140 391 1151 425
rect 1185 391 1196 425
rect 1140 367 1196 391
rect 1226 595 1282 619
rect 1226 561 1237 595
rect 1271 561 1282 595
rect 1226 509 1282 561
rect 1226 475 1237 509
rect 1271 475 1282 509
rect 1226 425 1282 475
rect 1226 391 1237 425
rect 1271 391 1282 425
rect 1226 367 1282 391
rect 1312 595 1368 619
rect 1312 561 1323 595
rect 1357 561 1368 595
rect 1312 509 1368 561
rect 1312 475 1323 509
rect 1357 475 1368 509
rect 1312 425 1368 475
rect 1312 391 1323 425
rect 1357 391 1368 425
rect 1312 367 1368 391
rect 1398 595 1454 619
rect 1398 561 1409 595
rect 1443 561 1454 595
rect 1398 509 1454 561
rect 1398 475 1409 509
rect 1443 475 1454 509
rect 1398 425 1454 475
rect 1398 391 1409 425
rect 1443 391 1454 425
rect 1398 367 1454 391
rect 1484 595 1540 619
rect 1484 561 1495 595
rect 1529 561 1540 595
rect 1484 509 1540 561
rect 1484 475 1495 509
rect 1529 475 1540 509
rect 1484 425 1540 475
rect 1484 391 1495 425
rect 1529 391 1540 425
rect 1484 367 1540 391
rect 1570 595 1626 619
rect 1570 561 1581 595
rect 1615 561 1626 595
rect 1570 509 1626 561
rect 1570 475 1581 509
rect 1615 475 1626 509
rect 1570 425 1626 475
rect 1570 391 1581 425
rect 1615 391 1626 425
rect 1570 367 1626 391
rect 1656 595 1712 619
rect 1656 561 1667 595
rect 1701 561 1712 595
rect 1656 509 1712 561
rect 1656 475 1667 509
rect 1701 475 1712 509
rect 1656 425 1712 475
rect 1656 391 1667 425
rect 1701 391 1712 425
rect 1656 367 1712 391
rect 1742 595 1798 619
rect 1742 561 1753 595
rect 1787 561 1798 595
rect 1742 509 1798 561
rect 1742 475 1753 509
rect 1787 475 1798 509
rect 1742 425 1798 475
rect 1742 391 1753 425
rect 1787 391 1798 425
rect 1742 367 1798 391
rect 1828 595 1881 619
rect 1828 561 1839 595
rect 1873 561 1881 595
rect 1828 509 1881 561
rect 1828 475 1839 509
rect 1873 475 1881 509
rect 1828 425 1881 475
rect 1828 391 1839 425
rect 1873 391 1881 425
rect 1828 367 1881 391
<< ndiffc >>
rect 41 72 75 106
rect 127 72 161 106
rect 213 71 247 105
rect 299 72 333 106
rect 385 71 419 105
rect 463 71 497 105
rect 549 71 583 105
rect 635 71 669 105
rect 721 71 755 105
rect 807 71 841 105
rect 893 71 927 105
rect 979 71 1013 105
rect 1065 71 1099 105
rect 1151 71 1185 105
rect 1237 71 1271 105
rect 1323 71 1357 105
rect 1409 71 1443 105
rect 1495 71 1529 105
rect 1581 71 1615 105
rect 1667 71 1701 105
rect 1753 71 1787 105
rect 1839 71 1873 105
<< pdiffc >>
rect 41 561 75 595
rect 41 475 75 509
rect 41 391 75 425
rect 127 561 161 595
rect 127 475 161 509
rect 127 391 161 425
rect 213 569 247 603
rect 213 491 247 525
rect 213 421 247 455
rect 299 561 333 595
rect 299 475 333 509
rect 299 391 333 425
rect 385 569 419 603
rect 463 569 497 603
rect 385 491 419 525
rect 463 491 497 525
rect 385 421 419 455
rect 463 421 497 455
rect 549 561 583 595
rect 549 475 583 509
rect 549 391 583 425
rect 635 561 669 595
rect 635 475 669 509
rect 635 391 669 425
rect 721 561 755 595
rect 721 475 755 509
rect 721 391 755 425
rect 807 561 841 595
rect 807 475 841 509
rect 807 391 841 425
rect 893 561 927 595
rect 893 475 927 509
rect 893 391 927 425
rect 979 561 1013 595
rect 979 475 1013 509
rect 979 391 1013 425
rect 1065 561 1099 595
rect 1065 475 1099 509
rect 1065 391 1099 425
rect 1151 561 1185 595
rect 1151 475 1185 509
rect 1151 391 1185 425
rect 1237 561 1271 595
rect 1237 475 1271 509
rect 1237 391 1271 425
rect 1323 561 1357 595
rect 1323 475 1357 509
rect 1323 391 1357 425
rect 1409 561 1443 595
rect 1409 475 1443 509
rect 1409 391 1443 425
rect 1495 561 1529 595
rect 1495 475 1529 509
rect 1495 391 1529 425
rect 1581 561 1615 595
rect 1581 475 1615 509
rect 1581 391 1615 425
rect 1667 561 1701 595
rect 1667 475 1701 509
rect 1667 391 1701 425
rect 1753 561 1787 595
rect 1753 475 1787 509
rect 1753 391 1787 425
rect 1839 561 1873 595
rect 1839 475 1873 509
rect 1839 391 1873 425
<< poly >>
rect 86 619 116 645
rect 172 619 202 645
rect 258 619 288 645
rect 344 619 374 645
rect 508 619 538 645
rect 594 619 624 645
rect 680 619 710 645
rect 766 619 796 645
rect 852 619 882 645
rect 938 619 968 645
rect 1024 619 1054 645
rect 1110 619 1140 645
rect 1196 619 1226 645
rect 1282 619 1312 645
rect 1368 619 1398 645
rect 1454 619 1484 645
rect 1540 619 1570 645
rect 1626 619 1656 645
rect 1712 619 1742 645
rect 1798 619 1828 645
rect 86 291 116 367
rect 172 291 202 367
rect 258 291 288 367
rect 344 291 374 367
rect 508 307 538 367
rect 594 307 624 367
rect 680 307 710 367
rect 766 307 796 367
rect 852 307 882 367
rect 938 307 968 367
rect 1024 307 1054 367
rect 1110 307 1140 367
rect 1196 307 1226 367
rect 1282 307 1312 367
rect 1368 307 1398 367
rect 1454 307 1484 367
rect 1540 307 1570 367
rect 1626 307 1656 367
rect 1712 307 1742 367
rect 1798 307 1828 367
rect 86 275 374 291
rect 86 241 118 275
rect 152 241 186 275
rect 220 241 254 275
rect 288 241 322 275
rect 356 241 374 275
rect 86 225 374 241
rect 86 131 116 225
rect 172 131 202 225
rect 258 131 288 225
rect 344 131 374 225
rect 423 291 1828 307
rect 423 257 439 291
rect 473 257 636 291
rect 670 257 808 291
rect 842 257 980 291
rect 1014 257 1152 291
rect 1186 257 1323 291
rect 1357 257 1496 291
rect 1530 257 1668 291
rect 1702 257 1828 291
rect 423 242 1828 257
rect 423 223 538 242
rect 423 189 439 223
rect 473 189 538 223
rect 423 173 538 189
rect 508 131 538 173
rect 594 241 1828 242
rect 594 131 624 241
rect 680 131 710 241
rect 766 131 796 241
rect 852 131 882 241
rect 938 131 968 241
rect 1024 131 1054 241
rect 1110 131 1140 241
rect 1196 131 1226 241
rect 1282 131 1312 241
rect 1368 131 1398 241
rect 1454 131 1484 241
rect 1540 131 1570 241
rect 1626 131 1656 241
rect 1712 131 1742 241
rect 1798 131 1828 241
rect 86 21 116 47
rect 172 21 202 47
rect 258 21 288 47
rect 344 21 374 47
rect 508 21 538 47
rect 594 21 624 47
rect 680 21 710 47
rect 766 21 796 47
rect 852 21 882 47
rect 938 21 968 47
rect 1024 21 1054 47
rect 1110 21 1140 47
rect 1196 21 1226 47
rect 1282 21 1312 47
rect 1368 21 1398 47
rect 1454 21 1484 47
rect 1540 21 1570 47
rect 1626 21 1656 47
rect 1712 21 1742 47
rect 1798 21 1828 47
<< polycont >>
rect 118 241 152 275
rect 186 241 220 275
rect 254 241 288 275
rect 322 241 356 275
rect 439 257 473 291
rect 636 257 670 291
rect 808 257 842 291
rect 980 257 1014 291
rect 1152 257 1186 291
rect 1323 257 1357 291
rect 1496 257 1530 291
rect 1668 257 1702 291
rect 439 189 473 223
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 25 595 84 649
rect 25 561 41 595
rect 75 561 84 595
rect 25 509 84 561
rect 25 475 41 509
rect 75 475 84 509
rect 25 425 84 475
rect 25 391 41 425
rect 75 391 84 425
rect 25 375 84 391
rect 118 595 171 615
rect 118 561 127 595
rect 161 561 171 595
rect 118 509 171 561
rect 118 475 127 509
rect 161 475 171 509
rect 118 425 171 475
rect 118 391 127 425
rect 161 391 171 425
rect 205 603 258 649
rect 205 569 213 603
rect 247 569 258 603
rect 205 525 258 569
rect 205 491 213 525
rect 247 491 258 525
rect 205 455 258 491
rect 205 421 213 455
rect 247 421 258 455
rect 205 405 258 421
rect 292 595 342 615
rect 292 561 299 595
rect 333 561 342 595
rect 292 509 342 561
rect 292 475 299 509
rect 333 475 342 509
rect 292 425 342 475
rect 118 371 171 391
rect 292 391 299 425
rect 333 391 342 425
rect 376 603 510 649
rect 376 569 385 603
rect 419 569 463 603
rect 497 569 510 603
rect 376 525 510 569
rect 376 491 385 525
rect 419 491 463 525
rect 497 491 510 525
rect 376 455 510 491
rect 376 421 385 455
rect 419 421 463 455
rect 497 421 510 455
rect 376 405 510 421
rect 544 595 587 611
rect 544 561 549 595
rect 583 561 587 595
rect 544 509 587 561
rect 544 475 549 509
rect 583 475 587 509
rect 544 425 587 475
rect 292 371 342 391
rect 544 390 549 425
rect 583 390 587 425
rect 118 337 440 371
rect 397 307 440 337
rect 397 291 510 307
rect 86 275 363 291
rect 86 241 118 275
rect 152 241 186 275
rect 220 241 254 275
rect 288 241 322 275
rect 356 241 363 275
rect 86 225 363 241
rect 397 276 439 291
rect 397 242 404 276
rect 438 257 439 276
rect 473 276 510 291
rect 473 257 476 276
rect 438 242 476 257
rect 397 223 510 242
rect 397 189 439 223
rect 473 189 510 223
rect 118 155 510 189
rect 25 106 84 122
rect 25 72 41 106
rect 75 72 84 106
rect 25 17 84 72
rect 118 106 168 155
rect 118 72 127 106
rect 161 72 168 106
rect 118 56 168 72
rect 202 105 258 121
rect 202 71 213 105
rect 247 71 258 105
rect 202 17 258 71
rect 292 106 341 155
rect 292 72 299 106
rect 333 72 341 106
rect 292 56 341 72
rect 375 105 510 121
rect 375 71 385 105
rect 419 71 463 105
rect 497 71 510 105
rect 375 17 510 71
rect 544 105 587 390
rect 621 595 683 649
rect 621 561 635 595
rect 669 561 683 595
rect 621 509 683 561
rect 621 475 635 509
rect 669 475 683 509
rect 621 425 683 475
rect 621 391 635 425
rect 669 391 683 425
rect 621 375 683 391
rect 717 595 759 611
rect 717 561 721 595
rect 755 561 759 595
rect 717 509 759 561
rect 717 475 721 509
rect 755 475 759 509
rect 717 425 759 475
rect 717 390 721 425
rect 755 390 759 425
rect 621 291 683 307
rect 621 242 636 291
rect 670 242 683 291
rect 621 241 683 242
rect 544 71 549 105
rect 583 71 587 105
rect 544 55 587 71
rect 621 105 683 121
rect 621 71 635 105
rect 669 71 683 105
rect 621 17 683 71
rect 717 105 759 390
rect 793 595 855 649
rect 793 561 807 595
rect 841 561 855 595
rect 793 509 855 561
rect 793 475 807 509
rect 841 475 855 509
rect 793 425 855 475
rect 793 391 807 425
rect 841 391 855 425
rect 793 375 855 391
rect 889 595 931 611
rect 889 561 893 595
rect 927 561 931 595
rect 889 509 931 561
rect 889 475 893 509
rect 927 475 931 509
rect 889 425 931 475
rect 889 390 893 425
rect 927 390 931 425
rect 793 291 855 307
rect 793 242 808 291
rect 842 242 855 291
rect 793 241 855 242
rect 717 71 721 105
rect 755 71 759 105
rect 717 55 759 71
rect 793 105 855 121
rect 793 71 807 105
rect 841 71 855 105
rect 793 17 855 71
rect 889 105 931 390
rect 965 595 1027 649
rect 965 561 979 595
rect 1013 561 1027 595
rect 965 509 1027 561
rect 965 475 979 509
rect 1013 475 1027 509
rect 965 425 1027 475
rect 965 391 979 425
rect 1013 391 1027 425
rect 965 375 1027 391
rect 1061 595 1103 611
rect 1061 561 1065 595
rect 1099 561 1103 595
rect 1061 509 1103 561
rect 1061 475 1065 509
rect 1099 475 1103 509
rect 1061 425 1103 475
rect 1061 390 1065 425
rect 1099 390 1103 425
rect 965 291 1027 307
rect 965 242 980 291
rect 1014 242 1027 291
rect 965 241 1027 242
rect 889 71 893 105
rect 927 71 931 105
rect 889 55 931 71
rect 965 105 1027 121
rect 965 71 979 105
rect 1013 71 1027 105
rect 965 17 1027 71
rect 1061 105 1103 390
rect 1137 595 1199 649
rect 1137 561 1151 595
rect 1185 561 1199 595
rect 1137 509 1199 561
rect 1137 475 1151 509
rect 1185 475 1199 509
rect 1137 425 1199 475
rect 1137 391 1151 425
rect 1185 391 1199 425
rect 1137 375 1199 391
rect 1233 595 1275 611
rect 1233 561 1237 595
rect 1271 561 1275 595
rect 1233 509 1275 561
rect 1233 475 1237 509
rect 1271 475 1275 509
rect 1233 425 1275 475
rect 1233 390 1237 425
rect 1271 390 1275 425
rect 1137 291 1199 307
rect 1137 242 1152 291
rect 1186 242 1199 291
rect 1137 241 1199 242
rect 1061 71 1065 105
rect 1099 71 1103 105
rect 1061 55 1103 71
rect 1137 105 1199 121
rect 1137 71 1151 105
rect 1185 71 1199 105
rect 1137 17 1199 71
rect 1233 105 1275 390
rect 1309 595 1370 649
rect 1309 561 1323 595
rect 1357 561 1370 595
rect 1309 509 1370 561
rect 1309 475 1323 509
rect 1357 475 1370 509
rect 1309 425 1370 475
rect 1309 391 1323 425
rect 1357 391 1370 425
rect 1309 375 1370 391
rect 1404 595 1447 611
rect 1404 561 1409 595
rect 1443 561 1447 595
rect 1404 509 1447 561
rect 1404 475 1409 509
rect 1443 475 1447 509
rect 1404 425 1447 475
rect 1404 390 1409 425
rect 1443 390 1447 425
rect 1309 291 1370 307
rect 1309 242 1323 291
rect 1357 242 1370 291
rect 1309 241 1370 242
rect 1233 71 1237 105
rect 1271 71 1275 105
rect 1233 55 1275 71
rect 1309 105 1370 121
rect 1309 71 1323 105
rect 1357 71 1370 105
rect 1309 17 1370 71
rect 1404 105 1447 390
rect 1481 595 1543 649
rect 1481 561 1495 595
rect 1529 561 1543 595
rect 1481 509 1543 561
rect 1481 475 1495 509
rect 1529 475 1543 509
rect 1481 425 1543 475
rect 1481 391 1495 425
rect 1529 391 1543 425
rect 1481 375 1543 391
rect 1577 595 1619 611
rect 1577 561 1581 595
rect 1615 561 1619 595
rect 1577 509 1619 561
rect 1577 475 1581 509
rect 1615 475 1619 509
rect 1577 425 1619 475
rect 1577 390 1581 425
rect 1615 390 1619 425
rect 1481 291 1543 307
rect 1481 242 1496 291
rect 1530 242 1543 291
rect 1481 241 1543 242
rect 1404 71 1409 105
rect 1443 71 1447 105
rect 1404 55 1447 71
rect 1481 105 1543 121
rect 1481 71 1495 105
rect 1529 71 1543 105
rect 1481 17 1543 71
rect 1577 105 1619 390
rect 1653 595 1715 649
rect 1653 561 1667 595
rect 1701 561 1715 595
rect 1653 509 1715 561
rect 1653 475 1667 509
rect 1701 475 1715 509
rect 1653 425 1715 475
rect 1653 391 1667 425
rect 1701 391 1715 425
rect 1653 375 1715 391
rect 1749 595 1791 611
rect 1749 561 1753 595
rect 1787 561 1791 595
rect 1749 509 1791 561
rect 1749 475 1753 509
rect 1787 475 1791 509
rect 1749 425 1791 475
rect 1749 390 1753 425
rect 1787 390 1791 425
rect 1653 291 1715 307
rect 1653 242 1668 291
rect 1702 242 1715 291
rect 1653 241 1715 242
rect 1577 71 1581 105
rect 1615 71 1619 105
rect 1577 55 1619 71
rect 1653 105 1715 121
rect 1653 71 1667 105
rect 1701 71 1715 105
rect 1653 17 1715 71
rect 1749 105 1791 390
rect 1825 595 1889 649
rect 1825 561 1839 595
rect 1873 561 1889 595
rect 1825 509 1889 561
rect 1825 475 1839 509
rect 1873 475 1889 509
rect 1825 425 1889 475
rect 1825 391 1839 425
rect 1873 391 1889 425
rect 1825 375 1889 391
rect 1749 71 1753 105
rect 1787 71 1791 105
rect 1749 55 1791 71
rect 1825 105 1889 121
rect 1825 71 1839 105
rect 1873 71 1889 105
rect 1825 17 1889 71
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 549 391 583 424
rect 549 390 583 391
rect 404 242 438 276
rect 476 242 510 276
rect 721 391 755 424
rect 721 390 755 391
rect 636 257 670 276
rect 636 242 670 257
rect 893 391 927 424
rect 893 390 927 391
rect 808 257 842 276
rect 808 242 842 257
rect 1065 391 1099 424
rect 1065 390 1099 391
rect 980 257 1014 276
rect 980 242 1014 257
rect 1237 391 1271 424
rect 1237 390 1271 391
rect 1152 257 1186 276
rect 1152 242 1186 257
rect 1409 391 1443 424
rect 1409 390 1443 391
rect 1323 257 1357 276
rect 1323 242 1357 257
rect 1581 391 1615 424
rect 1581 390 1615 391
rect 1496 257 1530 276
rect 1496 242 1530 257
rect 1753 391 1787 424
rect 1753 390 1787 391
rect 1668 257 1702 276
rect 1668 242 1702 257
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 537 424 1807 430
rect 537 390 549 424
rect 583 390 721 424
rect 755 390 893 424
rect 927 390 1065 424
rect 1099 390 1237 424
rect 1271 390 1409 424
rect 1443 390 1581 424
rect 1615 390 1753 424
rect 1787 390 1807 424
rect 537 384 1807 390
rect 392 276 1722 282
rect 392 242 404 276
rect 438 242 476 276
rect 510 242 636 276
rect 670 242 808 276
rect 842 242 980 276
rect 1014 242 1152 276
rect 1186 242 1323 276
rect 1357 242 1496 276
rect 1530 242 1668 276
rect 1702 242 1722 276
rect 392 236 1722 242
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel pwell s 1551 24 1551 24 0 FreeSans 200 0 0 0 VNB
port 3 nsew
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkbuf_16
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 537 390 1807 424 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 681728
string GDS_START 666216
<< end >>
