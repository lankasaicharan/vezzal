magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 7 243 507 247
rect 7 49 912 243
rect 0 0 960 49
<< scnmos >>
rect 86 53 116 221
rect 172 53 202 221
rect 326 53 356 221
rect 398 53 428 221
rect 623 49 653 217
rect 709 49 739 217
rect 803 49 833 217
<< scpmoshvt >>
rect 86 367 116 619
rect 172 367 202 619
rect 304 367 334 619
rect 397 367 427 619
rect 623 367 653 619
rect 709 367 739 619
rect 803 367 833 619
<< ndiff >>
rect 33 209 86 221
rect 33 175 41 209
rect 75 175 86 209
rect 33 99 86 175
rect 33 65 41 99
rect 75 65 86 99
rect 33 53 86 65
rect 116 213 172 221
rect 116 179 127 213
rect 161 179 172 213
rect 116 101 172 179
rect 116 67 127 101
rect 161 67 172 101
rect 116 53 172 67
rect 202 163 326 221
rect 202 61 213 163
rect 315 61 326 163
rect 202 53 326 61
rect 356 53 398 221
rect 428 209 481 221
rect 428 175 439 209
rect 473 175 481 209
rect 428 101 481 175
rect 428 67 439 101
rect 473 67 481 101
rect 428 53 481 67
rect 570 181 623 217
rect 570 147 578 181
rect 612 147 623 181
rect 570 95 623 147
rect 570 61 578 95
rect 612 61 623 95
rect 570 49 623 61
rect 653 205 709 217
rect 653 171 664 205
rect 698 171 709 205
rect 653 101 709 171
rect 653 67 664 101
rect 698 67 709 101
rect 653 49 709 67
rect 739 49 803 217
rect 833 205 886 217
rect 833 171 844 205
rect 878 171 886 205
rect 833 95 886 171
rect 833 61 844 95
rect 878 61 886 95
rect 833 49 886 61
<< pdiff >>
rect 33 607 86 619
rect 33 573 41 607
rect 75 573 86 607
rect 33 507 86 573
rect 33 473 41 507
rect 75 473 86 507
rect 33 413 86 473
rect 33 379 41 413
rect 75 379 86 413
rect 33 367 86 379
rect 116 599 172 619
rect 116 565 127 599
rect 161 565 172 599
rect 116 497 172 565
rect 116 463 127 497
rect 161 463 172 497
rect 116 413 172 463
rect 116 379 127 413
rect 161 379 172 413
rect 116 367 172 379
rect 202 607 304 619
rect 202 573 237 607
rect 271 573 304 607
rect 202 512 304 573
rect 202 478 237 512
rect 271 478 304 512
rect 202 418 304 478
rect 202 384 237 418
rect 271 384 304 418
rect 202 367 304 384
rect 334 599 397 619
rect 334 565 345 599
rect 379 565 397 599
rect 334 522 397 565
rect 334 488 345 522
rect 379 488 397 522
rect 334 434 397 488
rect 334 400 345 434
rect 379 400 397 434
rect 334 367 397 400
rect 427 607 480 619
rect 427 573 438 607
rect 472 573 480 607
rect 427 367 480 573
rect 570 436 623 619
rect 570 402 578 436
rect 612 402 623 436
rect 570 367 623 402
rect 653 596 709 619
rect 653 562 664 596
rect 698 562 709 596
rect 653 367 709 562
rect 739 514 803 619
rect 739 480 750 514
rect 784 480 803 514
rect 739 434 803 480
rect 739 400 750 434
rect 784 400 803 434
rect 739 367 803 400
rect 833 599 886 619
rect 833 565 844 599
rect 878 565 886 599
rect 833 516 886 565
rect 833 482 844 516
rect 878 482 886 516
rect 833 434 886 482
rect 833 400 844 434
rect 878 400 886 434
rect 833 367 886 400
<< ndiffc >>
rect 41 175 75 209
rect 41 65 75 99
rect 127 179 161 213
rect 127 67 161 101
rect 213 61 315 163
rect 439 175 473 209
rect 439 67 473 101
rect 578 147 612 181
rect 578 61 612 95
rect 664 171 698 205
rect 664 67 698 101
rect 844 171 878 205
rect 844 61 878 95
<< pdiffc >>
rect 41 573 75 607
rect 41 473 75 507
rect 41 379 75 413
rect 127 565 161 599
rect 127 463 161 497
rect 127 379 161 413
rect 237 573 271 607
rect 237 478 271 512
rect 237 384 271 418
rect 345 565 379 599
rect 345 488 379 522
rect 345 400 379 434
rect 438 573 472 607
rect 578 402 612 436
rect 664 562 698 596
rect 750 480 784 514
rect 750 400 784 434
rect 844 565 878 599
rect 844 482 878 516
rect 844 400 878 434
<< poly >>
rect 86 619 116 645
rect 172 619 202 645
rect 304 619 334 645
rect 397 619 427 645
rect 623 619 653 645
rect 709 619 739 645
rect 803 619 833 645
rect 86 309 116 367
rect 172 309 202 367
rect 304 335 334 367
rect 397 335 427 367
rect 623 335 653 367
rect 709 335 739 367
rect 289 319 355 335
rect 86 293 247 309
rect 86 259 197 293
rect 231 259 247 293
rect 289 285 305 319
rect 339 285 355 319
rect 289 269 355 285
rect 397 319 481 335
rect 397 285 431 319
rect 465 285 481 319
rect 397 269 481 285
rect 587 319 653 335
rect 587 285 603 319
rect 637 285 653 319
rect 587 269 653 285
rect 695 319 761 335
rect 695 285 711 319
rect 745 285 761 319
rect 695 269 761 285
rect 803 305 833 367
rect 803 289 869 305
rect 86 243 247 259
rect 325 258 355 269
rect 325 249 356 258
rect 86 221 116 243
rect 172 221 202 243
rect 326 221 356 249
rect 398 221 428 269
rect 623 217 653 269
rect 709 217 739 269
rect 803 255 819 289
rect 853 255 869 289
rect 803 239 869 255
rect 803 217 833 239
rect 86 27 116 53
rect 172 27 202 53
rect 326 27 356 53
rect 398 27 428 53
rect 623 23 653 49
rect 709 23 739 49
rect 803 23 833 49
<< polycont >>
rect 197 259 231 293
rect 305 285 339 319
rect 431 285 465 319
rect 603 285 637 319
rect 711 285 745 319
rect 819 255 853 289
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 25 607 85 649
rect 25 573 41 607
rect 75 573 85 607
rect 25 507 85 573
rect 25 473 41 507
rect 75 473 85 507
rect 25 413 85 473
rect 25 379 41 413
rect 75 379 85 413
rect 25 363 85 379
rect 119 599 163 615
rect 119 565 127 599
rect 161 565 163 599
rect 119 497 163 565
rect 119 463 127 497
rect 161 463 163 497
rect 119 413 163 463
rect 119 379 127 413
rect 161 379 163 413
rect 221 607 287 649
rect 221 573 237 607
rect 271 573 287 607
rect 221 512 287 573
rect 221 478 237 512
rect 271 478 287 512
rect 221 418 287 478
rect 221 384 237 418
rect 271 384 287 418
rect 329 599 388 615
rect 329 565 345 599
rect 379 565 388 599
rect 422 607 488 649
rect 422 573 438 607
rect 472 573 488 607
rect 422 569 488 573
rect 648 599 894 615
rect 648 596 844 599
rect 329 522 388 565
rect 648 562 664 596
rect 698 565 844 596
rect 878 565 894 599
rect 698 562 894 565
rect 648 554 894 562
rect 329 488 345 522
rect 379 520 388 522
rect 379 514 800 520
rect 379 488 750 514
rect 329 486 750 488
rect 329 434 381 486
rect 734 480 750 486
rect 784 480 800 514
rect 329 400 345 434
rect 379 400 381 434
rect 329 384 381 400
rect 25 209 85 225
rect 25 175 41 209
rect 75 175 85 209
rect 25 99 85 175
rect 25 65 41 99
rect 75 65 85 99
rect 25 17 85 65
rect 119 213 163 379
rect 289 319 367 350
rect 197 293 247 309
rect 231 259 247 293
rect 289 285 305 319
rect 339 285 367 319
rect 415 319 481 452
rect 415 285 431 319
rect 465 285 481 319
rect 517 436 616 452
rect 517 402 578 436
rect 612 402 616 436
rect 517 386 616 402
rect 734 434 800 480
rect 734 400 750 434
rect 784 400 800 434
rect 197 249 247 259
rect 517 251 551 386
rect 734 384 800 400
rect 834 516 894 554
rect 834 482 844 516
rect 878 482 894 516
rect 834 434 894 482
rect 834 400 844 434
rect 878 400 894 434
rect 834 384 894 400
rect 587 319 653 352
rect 587 285 603 319
rect 637 285 653 319
rect 687 319 761 350
rect 687 285 711 319
rect 745 285 761 319
rect 799 289 929 350
rect 799 255 819 289
rect 853 255 929 289
rect 517 249 714 251
rect 197 215 714 249
rect 799 242 929 255
rect 119 179 127 213
rect 161 179 163 213
rect 423 209 489 215
rect 119 101 163 179
rect 119 67 127 101
rect 161 67 163 101
rect 119 51 163 67
rect 197 163 331 181
rect 197 61 213 163
rect 315 61 331 163
rect 197 17 331 61
rect 423 175 439 209
rect 473 175 489 209
rect 662 205 714 215
rect 423 101 489 175
rect 423 67 439 101
rect 473 67 489 101
rect 423 51 489 67
rect 562 147 578 181
rect 612 147 628 181
rect 562 95 628 147
rect 562 61 578 95
rect 612 61 628 95
rect 562 17 628 61
rect 662 171 664 205
rect 698 171 714 205
rect 662 101 714 171
rect 662 67 664 101
rect 698 67 714 101
rect 662 51 714 67
rect 828 205 894 208
rect 828 171 844 205
rect 878 171 894 205
rect 828 95 894 171
rect 828 61 844 95
rect 878 61 894 95
rect 828 17 894 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a221o_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6041596
string GDS_START 6032222
<< end >>
