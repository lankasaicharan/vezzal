magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 1 49 611 157
rect 0 0 672 49
<< scnmos >>
rect 84 47 114 131
rect 156 47 186 131
rect 264 47 294 131
rect 342 47 372 131
rect 420 47 450 131
rect 498 47 528 131
<< scpmoshvt >>
rect 87 409 137 609
rect 200 409 250 609
rect 306 409 356 609
rect 428 409 478 609
rect 534 409 584 609
<< ndiff >>
rect 27 111 84 131
rect 27 77 39 111
rect 73 77 84 111
rect 27 47 84 77
rect 114 47 156 131
rect 186 97 264 131
rect 186 63 197 97
rect 231 63 264 97
rect 186 47 264 63
rect 294 47 342 131
rect 372 47 420 131
rect 450 47 498 131
rect 528 111 585 131
rect 528 77 539 111
rect 573 77 585 111
rect 528 47 585 77
<< pdiff >>
rect 30 597 87 609
rect 30 563 42 597
rect 76 563 87 597
rect 30 526 87 563
rect 30 492 42 526
rect 76 492 87 526
rect 30 455 87 492
rect 30 421 42 455
rect 76 421 87 455
rect 30 409 87 421
rect 137 597 200 609
rect 137 563 148 597
rect 182 563 200 597
rect 137 514 200 563
rect 137 480 148 514
rect 182 480 200 514
rect 137 409 200 480
rect 250 597 306 609
rect 250 563 261 597
rect 295 563 306 597
rect 250 526 306 563
rect 250 492 261 526
rect 295 492 306 526
rect 250 455 306 492
rect 250 421 261 455
rect 295 421 306 455
rect 250 409 306 421
rect 356 597 428 609
rect 356 563 367 597
rect 401 563 428 597
rect 356 514 428 563
rect 356 480 367 514
rect 401 480 428 514
rect 356 409 428 480
rect 478 597 534 609
rect 478 563 489 597
rect 523 563 534 597
rect 478 526 534 563
rect 478 492 489 526
rect 523 492 534 526
rect 478 455 534 492
rect 478 421 489 455
rect 523 421 534 455
rect 478 409 534 421
rect 584 597 641 609
rect 584 563 595 597
rect 629 563 641 597
rect 584 526 641 563
rect 584 492 595 526
rect 629 492 641 526
rect 584 455 641 492
rect 584 421 595 455
rect 629 421 641 455
rect 584 409 641 421
<< ndiffc >>
rect 39 77 73 111
rect 197 63 231 97
rect 539 77 573 111
<< pdiffc >>
rect 42 563 76 597
rect 42 492 76 526
rect 42 421 76 455
rect 148 563 182 597
rect 148 480 182 514
rect 261 563 295 597
rect 261 492 295 526
rect 261 421 295 455
rect 367 563 401 597
rect 367 480 401 514
rect 489 563 523 597
rect 489 492 523 526
rect 489 421 523 455
rect 595 563 629 597
rect 595 492 629 526
rect 595 421 629 455
<< poly >>
rect 87 609 137 635
rect 200 609 250 635
rect 306 609 356 635
rect 428 609 478 635
rect 534 609 584 635
rect 87 322 137 409
rect 200 358 250 409
rect 306 358 356 409
rect 428 358 478 409
rect 534 358 584 409
rect 198 342 264 358
rect 87 306 156 322
rect 87 272 106 306
rect 140 272 156 306
rect 87 238 156 272
rect 87 204 106 238
rect 140 204 156 238
rect 198 308 214 342
rect 248 308 264 342
rect 198 274 264 308
rect 198 240 214 274
rect 248 240 264 274
rect 198 224 264 240
rect 306 342 372 358
rect 306 308 322 342
rect 356 308 372 342
rect 306 274 372 308
rect 306 240 322 274
rect 356 240 372 274
rect 306 224 372 240
rect 87 176 156 204
rect 234 176 264 224
rect 84 146 186 176
rect 234 146 294 176
rect 84 131 114 146
rect 156 131 186 146
rect 264 131 294 146
rect 342 131 372 224
rect 420 342 486 358
rect 420 308 436 342
rect 470 308 486 342
rect 420 274 486 308
rect 420 240 436 274
rect 470 240 486 274
rect 420 224 486 240
rect 534 342 600 358
rect 534 308 550 342
rect 584 308 600 342
rect 534 274 600 308
rect 534 240 550 274
rect 584 240 600 274
rect 534 224 600 240
rect 420 131 450 224
rect 534 176 564 224
rect 498 146 564 176
rect 498 131 528 146
rect 84 21 114 47
rect 156 21 186 47
rect 264 21 294 47
rect 342 21 372 47
rect 420 21 450 47
rect 498 21 528 47
<< polycont >>
rect 106 272 140 306
rect 106 204 140 238
rect 214 308 248 342
rect 214 240 248 274
rect 322 308 356 342
rect 322 240 356 274
rect 436 308 470 342
rect 436 240 470 274
rect 550 308 584 342
rect 550 240 584 274
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 20 597 92 613
rect 20 563 42 597
rect 76 563 92 597
rect 20 526 92 563
rect 20 492 42 526
rect 76 492 92 526
rect 20 455 92 492
rect 132 597 198 649
rect 132 563 148 597
rect 182 563 198 597
rect 132 514 198 563
rect 132 480 148 514
rect 182 480 198 514
rect 132 464 198 480
rect 245 597 311 613
rect 245 563 261 597
rect 295 563 311 597
rect 245 526 311 563
rect 245 492 261 526
rect 295 492 311 526
rect 20 421 42 455
rect 76 421 92 455
rect 245 455 311 492
rect 351 597 417 649
rect 351 563 367 597
rect 401 563 417 597
rect 351 514 417 563
rect 351 480 367 514
rect 401 480 417 514
rect 351 464 417 480
rect 473 597 539 613
rect 473 563 489 597
rect 523 563 539 597
rect 473 526 539 563
rect 473 492 489 526
rect 523 492 539 526
rect 245 428 261 455
rect 20 384 92 421
rect 128 421 261 428
rect 295 428 311 455
rect 473 455 539 492
rect 473 428 489 455
rect 295 421 489 428
rect 523 421 539 455
rect 128 394 539 421
rect 579 597 645 649
rect 579 563 595 597
rect 629 563 645 597
rect 579 526 645 563
rect 579 492 595 526
rect 629 492 645 526
rect 579 455 645 492
rect 579 421 595 455
rect 629 421 645 455
rect 579 405 645 421
rect 20 135 54 384
rect 128 322 162 394
rect 90 306 162 322
rect 90 272 106 306
rect 140 272 162 306
rect 90 238 162 272
rect 90 204 106 238
rect 140 204 162 238
rect 198 342 264 358
rect 198 308 214 342
rect 248 308 264 342
rect 198 274 264 308
rect 198 240 214 274
rect 248 240 264 274
rect 198 224 264 240
rect 306 342 372 358
rect 306 308 322 342
rect 356 308 372 342
rect 306 274 372 308
rect 306 240 322 274
rect 356 240 372 274
rect 306 224 372 240
rect 409 342 486 358
rect 409 308 436 342
rect 470 308 486 342
rect 409 274 486 308
rect 409 240 436 274
rect 470 240 486 274
rect 409 224 486 240
rect 534 342 647 358
rect 534 308 550 342
rect 584 308 647 342
rect 534 274 647 308
rect 534 240 550 274
rect 584 240 647 274
rect 534 224 647 240
rect 90 188 162 204
rect 128 154 589 188
rect 20 111 89 135
rect 20 77 39 111
rect 73 77 89 111
rect 20 53 89 77
rect 181 97 247 118
rect 181 63 197 97
rect 231 63 247 97
rect 181 17 247 63
rect 523 111 589 154
rect 523 77 539 111
rect 573 77 589 111
rect 523 53 589 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4_lp2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6202478
string GDS_START 6195478
<< end >>
