magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 58 242 332 267
rect 58 49 736 242
rect 0 0 768 49
<< scnmos >>
rect 141 73 171 241
rect 219 73 249 241
rect 509 132 539 216
rect 623 132 653 216
<< scpmoshvt >>
rect 135 367 165 619
rect 213 367 243 619
rect 451 426 481 554
rect 623 426 653 554
<< ndiff >>
rect 84 213 141 241
rect 84 179 96 213
rect 130 179 141 213
rect 84 119 141 179
rect 84 85 96 119
rect 130 85 141 119
rect 84 73 141 85
rect 171 73 219 241
rect 249 229 306 241
rect 249 195 260 229
rect 294 195 306 229
rect 249 119 306 195
rect 452 191 509 216
rect 452 157 464 191
rect 498 157 509 191
rect 452 132 509 157
rect 539 191 623 216
rect 539 157 564 191
rect 598 157 623 191
rect 539 132 623 157
rect 653 191 710 216
rect 653 157 664 191
rect 698 157 710 191
rect 653 132 710 157
rect 249 85 260 119
rect 294 85 306 119
rect 249 73 306 85
<< pdiff >>
rect 78 603 135 619
rect 78 569 90 603
rect 124 569 135 603
rect 78 510 135 569
rect 78 476 90 510
rect 124 476 135 510
rect 78 417 135 476
rect 78 383 90 417
rect 124 383 135 417
rect 78 367 135 383
rect 165 367 213 619
rect 243 607 300 619
rect 243 573 254 607
rect 288 573 300 607
rect 243 510 300 573
rect 243 476 254 510
rect 288 476 300 510
rect 243 413 300 476
rect 394 501 451 554
rect 394 467 406 501
rect 440 467 451 501
rect 394 426 451 467
rect 481 541 623 554
rect 481 507 574 541
rect 608 507 623 541
rect 481 426 623 507
rect 653 542 720 554
rect 653 508 674 542
rect 708 508 720 542
rect 653 472 720 508
rect 653 438 674 472
rect 708 438 720 472
rect 653 426 720 438
rect 243 379 254 413
rect 288 379 300 413
rect 243 367 300 379
<< ndiffc >>
rect 96 179 130 213
rect 96 85 130 119
rect 260 195 294 229
rect 464 157 498 191
rect 564 157 598 191
rect 664 157 698 191
rect 260 85 294 119
<< pdiffc >>
rect 90 569 124 603
rect 90 476 124 510
rect 90 383 124 417
rect 254 573 288 607
rect 254 476 288 510
rect 406 467 440 501
rect 574 507 608 541
rect 674 508 708 542
rect 674 438 708 472
rect 254 379 288 413
<< poly >>
rect 135 619 165 645
rect 213 619 243 645
rect 451 554 481 580
rect 623 554 653 580
rect 451 388 481 426
rect 623 388 653 426
rect 451 372 575 388
rect 135 329 165 367
rect 213 341 243 367
rect 451 341 506 372
rect 213 338 506 341
rect 540 338 575 372
rect 105 313 171 329
rect 105 279 121 313
rect 155 279 171 313
rect 213 311 575 338
rect 105 263 171 279
rect 451 304 575 311
rect 451 270 506 304
rect 540 270 575 304
rect 141 241 171 263
rect 219 241 249 267
rect 451 254 575 270
rect 617 372 683 388
rect 617 338 633 372
rect 667 338 683 372
rect 617 304 683 338
rect 617 270 633 304
rect 667 270 683 304
rect 617 254 683 270
rect 509 216 539 254
rect 623 216 653 254
rect 364 101 430 117
rect 509 106 539 132
rect 623 106 653 132
rect 141 47 171 73
rect 219 51 249 73
rect 364 67 380 101
rect 414 67 430 101
rect 364 51 430 67
rect 219 21 430 51
<< polycont >>
rect 506 338 540 372
rect 121 279 155 313
rect 506 270 540 304
rect 633 338 667 372
rect 633 270 667 304
rect 380 67 414 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 25 603 140 615
rect 25 569 90 603
rect 124 569 140 603
rect 25 510 140 569
rect 25 476 90 510
rect 124 476 140 510
rect 25 417 140 476
rect 25 383 90 417
rect 124 383 140 417
rect 25 363 140 383
rect 238 607 304 649
rect 238 573 254 607
rect 288 573 304 607
rect 238 510 304 573
rect 238 476 254 510
rect 288 476 304 510
rect 238 413 304 476
rect 238 379 254 413
rect 288 379 304 413
rect 25 229 71 363
rect 238 359 304 379
rect 338 581 524 615
rect 105 325 171 329
rect 338 325 372 581
rect 105 313 372 325
rect 105 279 121 313
rect 155 291 372 313
rect 406 501 456 547
rect 440 467 456 501
rect 155 279 171 291
rect 105 263 171 279
rect 244 229 310 245
rect 25 213 146 229
rect 25 179 96 213
rect 130 179 146 213
rect 25 119 146 179
rect 25 85 96 119
rect 130 85 146 119
rect 25 69 146 85
rect 244 195 260 229
rect 294 195 310 229
rect 244 119 310 195
rect 244 85 260 119
rect 294 85 310 119
rect 406 220 456 467
rect 490 456 524 581
rect 558 541 624 649
rect 558 507 574 541
rect 608 507 624 541
rect 558 490 624 507
rect 658 542 751 558
rect 658 508 674 542
rect 708 508 751 542
rect 658 472 751 508
rect 658 456 674 472
rect 490 438 674 456
rect 708 438 751 472
rect 490 422 751 438
rect 490 372 556 388
rect 490 338 506 372
rect 540 338 556 372
rect 490 304 556 338
rect 490 270 506 304
rect 540 270 556 304
rect 490 254 556 270
rect 601 372 683 388
rect 601 338 633 372
rect 667 338 683 372
rect 601 304 683 338
rect 601 270 633 304
rect 667 270 683 304
rect 601 254 683 270
rect 717 220 751 422
rect 406 191 514 220
rect 406 157 464 191
rect 498 157 514 191
rect 406 128 514 157
rect 548 191 614 220
rect 548 157 564 191
rect 598 157 614 191
rect 406 117 440 128
rect 244 17 310 85
rect 364 101 440 117
rect 364 67 380 101
rect 414 67 440 101
rect 364 51 440 67
rect 548 17 614 157
rect 648 191 751 220
rect 648 157 664 191
rect 698 186 751 191
rect 698 157 714 186
rect 648 128 714 157
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ebufn_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3338648
string GDS_START 3332026
<< end >>
