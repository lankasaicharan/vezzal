magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 59 49 936 241
rect 0 0 960 49
<< scnmos >>
rect 138 47 168 215
rect 224 47 254 215
rect 402 47 432 215
rect 474 47 504 215
rect 601 47 631 215
rect 709 47 739 215
rect 817 47 847 215
<< scpmoshvt >>
rect 108 367 138 619
rect 194 367 224 619
rect 398 367 428 619
rect 484 367 514 619
rect 626 367 656 619
rect 731 367 761 619
rect 817 367 847 619
<< ndiff >>
rect 85 179 138 215
rect 85 145 93 179
rect 127 145 138 179
rect 85 93 138 145
rect 85 59 93 93
rect 127 59 138 93
rect 85 47 138 59
rect 168 203 224 215
rect 168 169 179 203
rect 213 169 224 203
rect 168 101 224 169
rect 168 67 179 101
rect 213 67 224 101
rect 168 47 224 67
rect 254 167 402 215
rect 254 133 265 167
rect 299 133 357 167
rect 391 133 402 167
rect 254 93 402 133
rect 254 59 265 93
rect 299 59 357 93
rect 391 59 402 93
rect 254 47 402 59
rect 432 47 474 215
rect 504 185 601 215
rect 504 151 530 185
rect 564 151 601 185
rect 504 101 601 151
rect 504 67 530 101
rect 564 67 601 101
rect 504 47 601 67
rect 631 47 709 215
rect 739 47 817 215
rect 847 192 910 215
rect 847 158 868 192
rect 902 158 910 192
rect 847 93 910 158
rect 847 59 868 93
rect 902 59 910 93
rect 847 47 910 59
<< pdiff >>
rect 55 599 108 619
rect 55 565 63 599
rect 97 565 108 599
rect 55 505 108 565
rect 55 471 63 505
rect 97 471 108 505
rect 55 413 108 471
rect 55 379 63 413
rect 97 379 108 413
rect 55 367 108 379
rect 138 611 194 619
rect 138 577 149 611
rect 183 577 194 611
rect 138 534 194 577
rect 138 500 149 534
rect 183 500 194 534
rect 138 457 194 500
rect 138 423 149 457
rect 183 423 194 457
rect 138 367 194 423
rect 224 599 277 619
rect 224 565 235 599
rect 269 565 277 599
rect 224 505 277 565
rect 224 471 235 505
rect 269 471 277 505
rect 224 413 277 471
rect 224 379 235 413
rect 269 379 277 413
rect 224 367 277 379
rect 345 606 398 619
rect 345 572 353 606
rect 387 572 398 606
rect 345 511 398 572
rect 345 477 353 511
rect 387 477 398 511
rect 345 420 398 477
rect 345 386 353 420
rect 387 386 398 420
rect 345 367 398 386
rect 428 531 484 619
rect 428 497 439 531
rect 473 497 484 531
rect 428 413 484 497
rect 428 379 439 413
rect 473 379 484 413
rect 428 367 484 379
rect 514 599 626 619
rect 514 565 525 599
rect 559 565 626 599
rect 514 513 626 565
rect 514 479 581 513
rect 615 479 626 513
rect 514 413 626 479
rect 514 379 581 413
rect 615 379 626 413
rect 514 367 626 379
rect 656 607 731 619
rect 656 573 676 607
rect 710 573 731 607
rect 656 531 731 573
rect 656 497 676 531
rect 710 497 731 531
rect 656 455 731 497
rect 656 421 676 455
rect 710 421 731 455
rect 656 367 731 421
rect 761 599 817 619
rect 761 565 772 599
rect 806 565 817 599
rect 761 506 817 565
rect 761 472 772 506
rect 806 472 817 506
rect 761 413 817 472
rect 761 379 772 413
rect 806 379 817 413
rect 761 367 817 379
rect 847 607 900 619
rect 847 573 858 607
rect 892 573 900 607
rect 847 509 900 573
rect 847 475 858 509
rect 892 475 900 509
rect 847 418 900 475
rect 847 384 858 418
rect 892 384 900 418
rect 847 367 900 384
<< ndiffc >>
rect 93 145 127 179
rect 93 59 127 93
rect 179 169 213 203
rect 179 67 213 101
rect 265 133 299 167
rect 357 133 391 167
rect 265 59 299 93
rect 357 59 391 93
rect 530 151 564 185
rect 530 67 564 101
rect 868 158 902 192
rect 868 59 902 93
<< pdiffc >>
rect 63 565 97 599
rect 63 471 97 505
rect 63 379 97 413
rect 149 577 183 611
rect 149 500 183 534
rect 149 423 183 457
rect 235 565 269 599
rect 235 471 269 505
rect 235 379 269 413
rect 353 572 387 606
rect 353 477 387 511
rect 353 386 387 420
rect 439 497 473 531
rect 439 379 473 413
rect 525 565 559 599
rect 581 479 615 513
rect 581 379 615 413
rect 676 573 710 607
rect 676 497 710 531
rect 676 421 710 455
rect 772 565 806 599
rect 772 472 806 506
rect 772 379 806 413
rect 858 573 892 607
rect 858 475 892 509
rect 858 384 892 418
<< poly >>
rect 108 619 138 645
rect 194 619 224 645
rect 398 619 428 645
rect 484 619 514 645
rect 626 619 656 645
rect 731 619 761 645
rect 817 619 847 645
rect 108 297 138 367
rect 194 333 224 367
rect 398 345 428 367
rect 194 317 283 333
rect 194 297 233 317
rect 108 283 233 297
rect 267 283 283 317
rect 108 267 283 283
rect 331 319 428 345
rect 331 285 347 319
rect 381 299 428 319
rect 484 303 514 367
rect 626 303 656 367
rect 731 303 761 367
rect 817 308 847 367
rect 381 285 432 299
rect 331 269 432 285
rect 138 215 168 267
rect 224 215 254 267
rect 402 215 432 269
rect 484 287 559 303
rect 484 267 509 287
rect 474 253 509 267
rect 543 253 559 287
rect 474 237 559 253
rect 601 287 667 303
rect 601 253 617 287
rect 651 253 667 287
rect 601 237 667 253
rect 709 287 775 303
rect 709 253 725 287
rect 759 253 775 287
rect 709 237 775 253
rect 817 292 919 308
rect 817 258 869 292
rect 903 258 919 292
rect 817 242 919 258
rect 474 215 504 237
rect 601 215 631 237
rect 709 215 739 237
rect 817 215 847 242
rect 138 21 168 47
rect 224 21 254 47
rect 402 21 432 47
rect 474 21 504 47
rect 601 21 631 47
rect 709 21 739 47
rect 817 21 847 47
<< polycont >>
rect 233 283 267 317
rect 347 285 381 319
rect 509 253 543 287
rect 617 253 651 287
rect 725 253 759 287
rect 869 258 903 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 31 599 99 615
rect 31 565 63 599
rect 97 565 99 599
rect 31 505 99 565
rect 31 471 63 505
rect 97 471 99 505
rect 31 413 99 471
rect 133 611 199 649
rect 133 577 149 611
rect 183 577 199 611
rect 133 534 199 577
rect 133 500 149 534
rect 183 500 199 534
rect 133 457 199 500
rect 133 423 149 457
rect 183 423 199 457
rect 233 599 283 615
rect 233 565 235 599
rect 269 565 283 599
rect 233 505 283 565
rect 233 471 235 505
rect 269 471 283 505
rect 31 379 63 413
rect 97 389 99 413
rect 233 413 283 471
rect 233 389 235 413
rect 97 379 235 389
rect 269 379 283 413
rect 337 606 626 615
rect 337 572 353 606
rect 387 599 626 606
rect 387 581 525 599
rect 387 572 403 581
rect 337 511 403 572
rect 513 565 525 581
rect 559 565 626 599
rect 513 549 626 565
rect 337 477 353 511
rect 387 477 403 511
rect 337 420 403 477
rect 337 386 353 420
rect 387 386 403 420
rect 437 531 475 547
rect 437 497 439 531
rect 473 497 475 531
rect 437 413 475 497
rect 31 355 283 379
rect 437 379 439 413
rect 473 379 475 413
rect 31 247 175 355
rect 217 317 283 321
rect 217 283 233 317
rect 267 283 283 317
rect 217 281 283 283
rect 31 213 215 247
rect 177 203 215 213
rect 77 145 93 179
rect 127 145 143 179
rect 77 93 143 145
rect 77 59 93 93
rect 127 59 143 93
rect 77 17 143 59
rect 177 169 179 203
rect 213 169 215 203
rect 249 235 283 281
rect 317 319 403 352
rect 317 285 347 319
rect 381 285 403 319
rect 317 269 403 285
rect 437 235 475 379
rect 509 287 547 515
rect 581 513 626 549
rect 615 479 626 513
rect 581 413 626 479
rect 660 607 726 649
rect 660 573 676 607
rect 710 573 726 607
rect 660 531 726 573
rect 660 497 676 531
rect 710 497 726 531
rect 660 455 726 497
rect 660 421 676 455
rect 710 421 726 455
rect 760 599 808 615
rect 760 565 772 599
rect 806 565 808 599
rect 760 506 808 565
rect 760 472 772 506
rect 806 472 808 506
rect 615 385 626 413
rect 760 413 808 472
rect 760 385 772 413
rect 615 379 772 385
rect 806 379 808 413
rect 842 607 908 649
rect 842 573 858 607
rect 892 573 908 607
rect 842 509 908 573
rect 842 475 858 509
rect 892 475 908 509
rect 842 418 908 475
rect 842 384 858 418
rect 892 384 908 418
rect 581 351 808 379
rect 543 253 547 287
rect 509 237 547 253
rect 607 287 651 303
rect 607 253 617 287
rect 249 201 475 235
rect 177 101 215 169
rect 441 185 573 201
rect 177 67 179 101
rect 213 67 215 101
rect 177 51 215 67
rect 249 133 265 167
rect 299 133 357 167
rect 391 133 407 167
rect 249 93 407 133
rect 249 59 265 93
rect 299 59 357 93
rect 391 59 407 93
rect 249 17 407 59
rect 441 151 530 185
rect 564 151 573 185
rect 441 101 573 151
rect 441 67 530 101
rect 564 67 573 101
rect 607 72 651 253
rect 685 287 833 303
rect 685 253 725 287
rect 759 253 833 287
rect 685 72 833 253
rect 869 292 943 350
rect 903 258 943 292
rect 869 242 943 258
rect 867 192 918 208
rect 867 158 868 192
rect 902 158 918 192
rect 867 93 918 158
rect 441 51 573 67
rect 867 59 868 93
rect 902 59 918 93
rect 867 17 918 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a32o_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2177710
string GDS_START 2168086
<< end >>
