magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 82 49 666 167
rect 0 0 672 49
<< scnmos >>
rect 165 57 195 141
rect 237 57 267 141
rect 323 57 353 141
rect 395 57 425 141
rect 481 57 511 141
rect 553 57 583 141
<< scpmoshvt >>
rect 205 408 255 608
rect 303 408 353 608
rect 533 409 583 609
<< ndiff >>
rect 108 116 165 141
rect 108 82 120 116
rect 154 82 165 116
rect 108 57 165 82
rect 195 57 237 141
rect 267 116 323 141
rect 267 82 278 116
rect 312 82 323 116
rect 267 57 323 82
rect 353 57 395 141
rect 425 108 481 141
rect 425 74 436 108
rect 470 74 481 108
rect 425 57 481 74
rect 511 57 553 141
rect 583 116 640 141
rect 583 82 594 116
rect 628 82 640 116
rect 583 57 640 82
<< pdiff >>
rect 148 596 205 608
rect 148 562 160 596
rect 194 562 205 596
rect 148 525 205 562
rect 148 491 160 525
rect 194 491 205 525
rect 148 454 205 491
rect 148 420 160 454
rect 194 420 205 454
rect 148 408 205 420
rect 255 408 303 608
rect 353 596 410 608
rect 353 562 364 596
rect 398 562 410 596
rect 353 525 410 562
rect 353 491 364 525
rect 398 491 410 525
rect 353 454 410 491
rect 353 420 364 454
rect 398 420 410 454
rect 353 408 410 420
rect 476 597 533 609
rect 476 563 488 597
rect 522 563 533 597
rect 476 526 533 563
rect 476 492 488 526
rect 522 492 533 526
rect 476 455 533 492
rect 476 421 488 455
rect 522 421 533 455
rect 476 409 533 421
rect 583 597 640 609
rect 583 563 594 597
rect 628 563 640 597
rect 583 526 640 563
rect 583 492 594 526
rect 628 492 640 526
rect 583 455 640 492
rect 583 421 594 455
rect 628 421 640 455
rect 583 409 640 421
<< ndiffc >>
rect 120 82 154 116
rect 278 82 312 116
rect 436 74 470 108
rect 594 82 628 116
<< pdiffc >>
rect 160 562 194 596
rect 160 491 194 525
rect 160 420 194 454
rect 364 562 398 596
rect 364 491 398 525
rect 364 420 398 454
rect 488 563 522 597
rect 488 492 522 526
rect 488 421 522 455
rect 594 563 628 597
rect 594 492 628 526
rect 594 421 628 455
<< poly >>
rect 205 608 255 634
rect 303 608 353 634
rect 533 609 583 635
rect 205 356 255 408
rect 165 340 255 356
rect 165 306 181 340
rect 215 306 255 340
rect 165 272 255 306
rect 303 300 353 408
rect 533 369 583 409
rect 165 238 181 272
rect 215 252 255 272
rect 323 264 353 300
rect 395 352 461 368
rect 395 318 411 352
rect 445 318 461 352
rect 395 284 461 318
rect 395 264 411 284
rect 215 238 267 252
rect 165 222 267 238
rect 165 141 195 222
rect 237 141 267 222
rect 323 250 411 264
rect 445 250 461 284
rect 323 234 461 250
rect 509 353 583 369
rect 509 319 525 353
rect 559 319 583 353
rect 509 285 583 319
rect 509 251 525 285
rect 559 251 583 285
rect 509 235 583 251
rect 323 141 353 234
rect 395 141 425 234
rect 553 186 583 235
rect 481 156 583 186
rect 481 141 511 156
rect 553 141 583 156
rect 165 31 195 57
rect 237 31 267 57
rect 323 31 353 57
rect 395 31 425 57
rect 481 31 511 57
rect 553 31 583 57
<< polycont >>
rect 181 306 215 340
rect 181 238 215 272
rect 411 318 445 352
rect 411 250 445 284
rect 525 319 559 353
rect 525 251 559 285
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 144 596 210 649
rect 144 562 160 596
rect 194 562 210 596
rect 144 525 210 562
rect 144 491 160 525
rect 194 491 210 525
rect 144 454 210 491
rect 144 420 160 454
rect 194 420 210 454
rect 144 404 210 420
rect 313 596 414 612
rect 313 562 364 596
rect 398 562 414 596
rect 313 525 414 562
rect 313 491 364 525
rect 398 491 414 525
rect 313 454 414 491
rect 313 420 364 454
rect 398 420 414 454
rect 313 404 414 420
rect 472 597 538 649
rect 472 563 488 597
rect 522 563 538 597
rect 472 526 538 563
rect 472 492 488 526
rect 522 492 538 526
rect 472 455 538 492
rect 472 421 488 455
rect 522 421 538 455
rect 472 405 538 421
rect 578 597 645 613
rect 578 563 594 597
rect 628 563 645 597
rect 578 526 645 563
rect 578 492 594 526
rect 628 492 645 526
rect 578 455 645 492
rect 578 421 594 455
rect 628 421 645 455
rect 578 405 645 421
rect 25 340 263 356
rect 25 306 181 340
rect 215 306 263 340
rect 25 272 263 306
rect 25 238 181 272
rect 215 238 263 272
rect 25 222 263 238
rect 313 145 359 404
rect 395 352 461 368
rect 395 318 411 352
rect 445 318 461 352
rect 395 284 461 318
rect 395 250 411 284
rect 445 250 461 284
rect 395 199 461 250
rect 505 353 575 369
rect 505 319 525 353
rect 559 319 575 353
rect 505 285 575 319
rect 505 251 525 285
rect 559 251 575 285
rect 505 235 575 251
rect 611 199 645 405
rect 395 165 645 199
rect 104 116 170 145
rect 104 82 120 116
rect 154 82 170 116
rect 104 17 170 82
rect 262 116 359 145
rect 262 82 278 116
rect 312 82 359 116
rect 262 53 359 82
rect 420 108 486 129
rect 420 74 436 108
rect 470 74 486 108
rect 420 17 486 74
rect 578 116 645 165
rect 578 82 594 116
rect 628 82 645 116
rect 578 53 645 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor2b_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5271998
string GDS_START 5265098
<< end >>
