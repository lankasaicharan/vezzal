magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 1 190 940 248
rect 1 49 957 190
rect 0 0 960 49
<< scpmos >>
rect 84 368 120 592
rect 182 368 218 592
rect 280 368 316 592
rect 374 368 410 592
rect 536 368 572 592
rect 626 368 662 592
rect 738 368 774 592
rect 828 368 864 592
<< nmoslvt >>
rect 84 74 114 222
rect 188 74 218 222
rect 274 74 304 222
rect 360 74 390 222
rect 572 74 602 222
rect 658 74 688 222
rect 744 74 774 222
rect 834 74 864 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 144 188 222
rect 114 110 139 144
rect 173 110 188 144
rect 114 74 188 110
rect 218 210 274 222
rect 218 176 229 210
rect 263 176 274 210
rect 218 120 274 176
rect 218 86 229 120
rect 263 86 274 120
rect 218 74 274 86
rect 304 189 360 222
rect 304 155 315 189
rect 349 155 360 189
rect 304 74 360 155
rect 390 164 440 222
rect 390 136 461 164
rect 522 150 572 222
rect 390 102 415 136
rect 449 102 461 136
rect 390 74 461 102
rect 515 142 572 150
rect 515 108 527 142
rect 561 108 572 142
rect 515 74 572 108
rect 602 179 658 222
rect 602 145 613 179
rect 647 145 658 179
rect 602 74 658 145
rect 688 210 744 222
rect 688 176 699 210
rect 733 176 744 210
rect 688 120 744 176
rect 688 86 699 120
rect 733 86 744 120
rect 688 74 744 86
rect 774 179 834 222
rect 774 145 785 179
rect 819 145 834 179
rect 774 74 834 145
rect 864 164 914 222
rect 864 136 931 164
rect 864 102 885 136
rect 919 102 931 136
rect 864 74 931 102
<< pdiff >>
rect 27 580 84 592
rect 27 546 39 580
rect 73 546 84 580
rect 27 503 84 546
rect 27 469 39 503
rect 73 469 84 503
rect 27 424 84 469
rect 27 390 39 424
rect 73 390 84 424
rect 27 368 84 390
rect 120 580 182 592
rect 120 546 130 580
rect 164 546 182 580
rect 120 508 182 546
rect 120 474 130 508
rect 164 474 182 508
rect 120 440 182 474
rect 120 406 130 440
rect 164 406 182 440
rect 120 368 182 406
rect 218 580 280 592
rect 218 546 230 580
rect 264 546 280 580
rect 218 499 280 546
rect 218 465 230 499
rect 264 465 280 499
rect 218 368 280 465
rect 316 580 374 592
rect 316 546 330 580
rect 364 546 374 580
rect 316 503 374 546
rect 316 469 330 503
rect 364 469 374 503
rect 316 424 374 469
rect 316 390 330 424
rect 364 390 374 424
rect 316 368 374 390
rect 410 580 536 592
rect 410 546 420 580
rect 454 546 492 580
rect 526 546 536 580
rect 410 508 536 546
rect 410 474 420 508
rect 454 474 492 508
rect 526 474 536 508
rect 410 368 536 474
rect 572 580 626 592
rect 572 546 582 580
rect 616 546 626 580
rect 572 503 626 546
rect 572 469 582 503
rect 616 469 626 503
rect 572 424 626 469
rect 572 390 582 424
rect 616 390 626 424
rect 572 368 626 390
rect 662 580 738 592
rect 662 546 682 580
rect 716 546 738 580
rect 662 499 738 546
rect 662 465 682 499
rect 716 465 738 499
rect 662 368 738 465
rect 774 580 828 592
rect 774 546 784 580
rect 818 546 828 580
rect 774 503 828 546
rect 774 469 784 503
rect 818 469 828 503
rect 774 424 828 469
rect 774 390 784 424
rect 818 390 828 424
rect 774 368 828 390
rect 864 580 924 592
rect 864 546 875 580
rect 909 546 924 580
rect 864 499 924 546
rect 864 465 875 499
rect 909 465 924 499
rect 864 368 924 465
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 110 173 144
rect 229 176 263 210
rect 229 86 263 120
rect 315 155 349 189
rect 415 102 449 136
rect 527 108 561 142
rect 613 145 647 179
rect 699 176 733 210
rect 699 86 733 120
rect 785 145 819 179
rect 885 102 919 136
<< pdiffc >>
rect 39 546 73 580
rect 39 469 73 503
rect 39 390 73 424
rect 130 546 164 580
rect 130 474 164 508
rect 130 406 164 440
rect 230 546 264 580
rect 230 465 264 499
rect 330 546 364 580
rect 330 469 364 503
rect 330 390 364 424
rect 420 546 454 580
rect 492 546 526 580
rect 420 474 454 508
rect 492 474 526 508
rect 582 546 616 580
rect 582 469 616 503
rect 582 390 616 424
rect 682 546 716 580
rect 682 465 716 499
rect 784 546 818 580
rect 784 469 818 503
rect 784 390 818 424
rect 875 546 909 580
rect 875 465 909 499
<< poly >>
rect 84 592 120 618
rect 182 592 218 618
rect 280 592 316 618
rect 374 592 410 618
rect 536 592 572 618
rect 626 592 662 618
rect 738 592 774 618
rect 828 592 864 618
rect 84 336 120 368
rect 182 336 218 368
rect 84 320 218 336
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 218 320
rect 280 336 316 368
rect 374 336 410 368
rect 536 336 572 368
rect 626 336 662 368
rect 738 336 774 368
rect 828 336 864 368
rect 280 320 488 336
rect 280 300 302 320
rect 84 270 218 286
rect 84 222 114 270
rect 188 222 218 270
rect 274 286 302 300
rect 336 286 370 320
rect 404 286 438 320
rect 472 286 488 320
rect 274 270 488 286
rect 536 320 688 336
rect 536 286 552 320
rect 586 286 638 320
rect 672 286 688 320
rect 536 270 688 286
rect 274 222 304 270
rect 360 222 390 270
rect 572 222 602 270
rect 658 222 688 270
rect 744 320 864 336
rect 744 286 793 320
rect 827 286 864 320
rect 744 270 864 286
rect 744 222 774 270
rect 834 222 864 270
rect 84 48 114 74
rect 188 48 218 74
rect 274 48 304 74
rect 360 48 390 74
rect 572 48 602 74
rect 658 48 688 74
rect 744 48 774 74
rect 834 48 864 74
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 302 286 336 320
rect 370 286 404 320
rect 438 286 472 320
rect 552 286 586 320
rect 638 286 672 320
rect 793 286 827 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 580 90 649
rect 23 546 39 580
rect 73 546 90 580
rect 23 503 90 546
rect 23 469 39 503
rect 73 469 90 503
rect 23 424 90 469
rect 23 390 39 424
rect 73 390 90 424
rect 127 580 180 596
rect 127 546 130 580
rect 164 546 180 580
rect 127 508 180 546
rect 127 474 130 508
rect 164 474 180 508
rect 127 440 180 474
rect 214 580 280 649
rect 214 546 230 580
rect 264 546 280 580
rect 214 499 280 546
rect 214 465 230 499
rect 264 465 280 499
rect 214 458 280 465
rect 314 580 380 596
rect 314 546 330 580
rect 364 546 380 580
rect 314 503 380 546
rect 314 469 330 503
rect 364 469 380 503
rect 127 406 130 440
rect 164 424 180 440
rect 314 424 380 469
rect 416 580 530 649
rect 416 546 420 580
rect 454 546 492 580
rect 526 546 530 580
rect 416 508 530 546
rect 416 474 420 508
rect 454 474 492 508
rect 526 474 530 508
rect 416 458 530 474
rect 566 580 632 596
rect 566 546 582 580
rect 616 546 632 580
rect 566 503 632 546
rect 566 469 582 503
rect 616 469 632 503
rect 566 424 632 469
rect 666 580 732 649
rect 666 546 682 580
rect 716 546 732 580
rect 666 499 732 546
rect 666 465 682 499
rect 716 465 732 499
rect 666 458 732 465
rect 768 580 825 596
rect 768 546 784 580
rect 818 546 825 580
rect 768 503 825 546
rect 768 469 784 503
rect 818 469 825 503
rect 768 430 825 469
rect 859 580 925 649
rect 859 546 875 580
rect 909 546 925 580
rect 859 499 925 546
rect 859 465 875 499
rect 909 465 925 499
rect 859 464 925 465
rect 768 424 935 430
rect 164 406 330 424
rect 127 390 330 406
rect 364 390 582 424
rect 616 390 784 424
rect 818 390 935 424
rect 25 320 218 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 218 320
rect 25 270 218 286
rect 286 320 488 356
rect 286 286 302 320
rect 336 286 370 320
rect 404 286 438 320
rect 472 286 488 320
rect 286 270 488 286
rect 536 320 743 356
rect 536 286 552 320
rect 586 286 638 320
rect 672 286 743 320
rect 536 270 743 286
rect 777 320 843 356
rect 777 286 793 320
rect 827 286 843 320
rect 777 270 843 286
rect 889 236 935 390
rect 23 210 263 236
rect 23 176 39 210
rect 73 202 229 210
rect 73 176 89 202
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 144 189 168
rect 123 110 139 144
rect 173 110 189 144
rect 123 17 189 110
rect 229 120 263 176
rect 299 202 663 236
rect 299 189 365 202
rect 299 155 315 189
rect 349 155 365 189
rect 597 179 663 202
rect 299 119 365 155
rect 399 136 465 168
rect 229 85 263 86
rect 399 102 415 136
rect 449 102 465 136
rect 399 85 465 102
rect 229 51 465 85
rect 511 142 563 168
rect 511 108 527 142
rect 561 108 563 142
rect 597 145 613 179
rect 647 145 663 179
rect 597 129 663 145
rect 697 210 735 226
rect 697 176 699 210
rect 733 176 735 210
rect 511 85 563 108
rect 697 120 735 176
rect 769 202 935 236
rect 769 179 835 202
rect 769 145 785 179
rect 819 145 835 179
rect 769 129 835 145
rect 869 136 935 168
rect 697 86 699 120
rect 733 86 735 120
rect 697 85 735 86
rect 869 102 885 136
rect 919 102 935 136
rect 869 85 935 102
rect 511 51 935 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 2625174
string GDS_START 2616492
<< end >>
