magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 214 165 762 183
rect 1 49 762 165
rect 0 0 768 49
<< scnmos >>
rect 80 55 110 139
rect 293 73 323 157
rect 365 73 395 157
rect 437 73 467 157
rect 545 73 575 157
rect 653 73 683 157
<< scpmoshvt >>
rect 185 397 215 481
rect 277 397 307 481
rect 365 397 395 481
rect 454 397 484 481
rect 545 397 575 481
rect 653 397 683 481
<< ndiff >>
rect 27 127 80 139
rect 27 93 35 127
rect 69 93 80 127
rect 27 55 80 93
rect 110 101 163 139
rect 110 67 121 101
rect 155 67 163 101
rect 110 55 163 67
rect 240 145 293 157
rect 240 111 248 145
rect 282 111 293 145
rect 240 73 293 111
rect 323 73 365 157
rect 395 73 437 157
rect 467 73 545 157
rect 575 119 653 157
rect 575 85 586 119
rect 620 85 653 119
rect 575 73 653 85
rect 683 144 736 157
rect 683 110 694 144
rect 728 110 736 144
rect 683 73 736 110
<< pdiff >>
rect 132 443 185 481
rect 132 409 140 443
rect 174 409 185 443
rect 132 397 185 409
rect 215 469 277 481
rect 215 435 226 469
rect 260 435 277 469
rect 215 397 277 435
rect 307 443 365 481
rect 307 409 318 443
rect 352 409 365 443
rect 307 397 365 409
rect 395 469 454 481
rect 395 435 408 469
rect 442 435 454 469
rect 395 397 454 435
rect 484 443 545 481
rect 484 409 500 443
rect 534 409 545 443
rect 484 397 545 409
rect 575 469 653 481
rect 575 435 602 469
rect 636 435 653 469
rect 575 397 653 435
rect 683 443 736 481
rect 683 409 694 443
rect 728 409 736 443
rect 683 397 736 409
<< ndiffc >>
rect 35 93 69 127
rect 121 67 155 101
rect 248 111 282 145
rect 586 85 620 119
rect 694 110 728 144
<< pdiffc >>
rect 140 409 174 443
rect 226 435 260 469
rect 318 409 352 443
rect 408 435 442 469
rect 500 409 534 443
rect 602 435 636 469
rect 694 409 728 443
<< poly >>
rect 496 605 562 621
rect 496 571 512 605
rect 546 585 562 605
rect 546 571 683 585
rect 496 555 683 571
rect 185 481 215 507
rect 277 481 307 507
rect 365 481 395 507
rect 454 481 484 507
rect 545 481 575 507
rect 653 481 683 555
rect 185 373 215 397
rect 277 375 307 397
rect 44 343 215 373
rect 257 345 307 375
rect 44 313 110 343
rect 44 279 60 313
rect 94 279 110 313
rect 257 295 287 345
rect 365 297 395 397
rect 454 313 484 397
rect 545 313 575 397
rect 44 245 110 279
rect 44 211 60 245
rect 94 211 110 245
rect 44 195 110 211
rect 80 139 110 195
rect 152 279 287 295
rect 152 245 168 279
rect 202 265 287 279
rect 329 281 395 297
rect 202 245 218 265
rect 152 211 218 245
rect 329 247 345 281
rect 379 247 395 281
rect 329 231 395 247
rect 152 177 168 211
rect 202 177 218 211
rect 152 161 218 177
rect 80 29 110 55
rect 188 51 218 161
rect 293 157 323 183
rect 365 157 395 231
rect 437 297 503 313
rect 437 263 453 297
rect 487 263 503 297
rect 437 229 503 263
rect 437 195 453 229
rect 487 195 503 229
rect 437 179 503 195
rect 545 297 611 313
rect 545 263 561 297
rect 595 263 611 297
rect 545 229 611 263
rect 545 195 561 229
rect 595 195 611 229
rect 545 179 611 195
rect 437 157 467 179
rect 545 157 575 179
rect 653 157 683 397
rect 293 51 323 73
rect 188 21 323 51
rect 365 47 395 73
rect 437 47 467 73
rect 545 47 575 73
rect 653 47 683 73
<< polycont >>
rect 512 571 546 605
rect 60 279 94 313
rect 60 211 94 245
rect 168 245 202 279
rect 345 247 379 281
rect 168 177 202 211
rect 453 263 487 297
rect 453 195 487 229
rect 561 263 595 297
rect 561 195 595 229
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 222 469 264 649
rect 136 443 178 459
rect 136 409 140 443
rect 174 409 178 443
rect 222 435 226 469
rect 260 435 264 469
rect 392 469 458 649
rect 222 419 264 435
rect 314 443 356 459
rect 136 383 178 409
rect 314 409 318 443
rect 352 409 356 443
rect 392 435 408 469
rect 442 435 458 469
rect 392 431 458 435
rect 496 571 512 605
rect 546 571 562 605
rect 496 443 538 571
rect 314 383 356 409
rect 496 409 500 443
rect 534 409 538 443
rect 598 469 640 649
rect 598 435 602 469
rect 636 435 640 469
rect 598 419 640 435
rect 690 443 737 572
rect 496 383 538 409
rect 136 349 202 383
rect 31 279 60 313
rect 94 279 110 313
rect 31 245 110 279
rect 31 211 60 245
rect 94 211 110 245
rect 168 279 202 349
rect 168 211 202 245
rect 168 175 202 177
rect 31 141 202 175
rect 244 349 538 383
rect 690 409 694 443
rect 728 409 737 443
rect 244 145 282 349
rect 415 297 487 313
rect 31 127 69 141
rect 31 93 35 127
rect 244 111 248 145
rect 31 77 69 93
rect 105 101 171 105
rect 105 67 121 101
rect 155 67 171 101
rect 244 95 282 111
rect 319 281 379 297
rect 319 247 345 281
rect 319 94 379 247
rect 415 263 453 297
rect 415 229 487 263
rect 415 195 453 229
rect 415 94 487 195
rect 561 297 641 313
rect 595 263 641 297
rect 561 229 641 263
rect 595 195 641 229
rect 561 168 641 195
rect 690 144 737 409
rect 570 119 636 123
rect 105 17 171 67
rect 570 85 586 119
rect 620 85 636 119
rect 690 110 694 144
rect 728 110 737 144
rect 690 94 737 110
rect 570 17 636 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4b_m
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5329506
string GDS_START 5321906
<< end >>
