magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 37 49 854 241
rect 0 0 864 49
<< scnmos >>
rect 116 131 146 215
rect 188 131 218 215
rect 274 131 304 215
rect 446 131 476 215
rect 532 131 562 215
rect 637 47 667 215
rect 723 47 753 215
<< scpmoshvt >>
rect 80 481 110 609
rect 174 481 204 609
rect 260 481 290 609
rect 450 367 480 495
rect 522 367 552 495
rect 637 367 667 619
rect 723 367 753 619
<< ndiff >>
rect 63 190 116 215
rect 63 156 71 190
rect 105 156 116 190
rect 63 131 116 156
rect 146 131 188 215
rect 218 187 274 215
rect 218 153 229 187
rect 263 153 274 187
rect 218 131 274 153
rect 304 136 446 215
rect 304 131 338 136
rect 326 102 338 131
rect 372 131 446 136
rect 476 190 532 215
rect 476 156 487 190
rect 521 156 532 190
rect 476 131 532 156
rect 562 161 637 215
rect 562 131 592 161
rect 372 102 384 131
rect 584 127 592 131
rect 626 127 637 161
rect 326 94 384 102
rect 584 93 637 127
rect 584 59 592 93
rect 626 59 637 93
rect 584 47 637 59
rect 667 203 723 215
rect 667 169 678 203
rect 712 169 723 203
rect 667 101 723 169
rect 667 67 678 101
rect 712 67 723 101
rect 667 47 723 67
rect 753 203 828 215
rect 753 169 782 203
rect 816 169 828 203
rect 753 93 828 169
rect 753 59 782 93
rect 816 59 828 93
rect 753 47 828 59
<< pdiff >>
rect 27 597 80 609
rect 27 563 35 597
rect 69 563 80 597
rect 27 527 80 563
rect 27 493 35 527
rect 69 493 80 527
rect 27 481 80 493
rect 110 587 174 609
rect 110 553 125 587
rect 159 553 174 587
rect 110 481 174 553
rect 204 597 260 609
rect 204 563 215 597
rect 249 563 260 597
rect 204 529 260 563
rect 204 495 215 529
rect 249 495 260 529
rect 204 481 260 495
rect 290 595 343 609
rect 290 561 301 595
rect 335 561 343 595
rect 290 527 343 561
rect 290 493 301 527
rect 335 493 343 527
rect 584 573 637 619
rect 584 539 592 573
rect 626 539 637 573
rect 584 495 637 539
rect 290 481 343 493
rect 397 418 450 495
rect 397 384 405 418
rect 439 384 450 418
rect 397 367 450 384
rect 480 367 522 495
rect 552 367 637 495
rect 667 599 723 619
rect 667 565 678 599
rect 712 565 723 599
rect 667 512 723 565
rect 667 478 678 512
rect 712 478 723 512
rect 667 420 723 478
rect 667 386 678 420
rect 712 386 723 420
rect 667 367 723 386
rect 753 607 828 619
rect 753 573 782 607
rect 816 573 828 607
rect 753 506 828 573
rect 753 472 782 506
rect 816 472 828 506
rect 753 413 828 472
rect 753 379 782 413
rect 816 379 828 413
rect 753 367 828 379
<< ndiffc >>
rect 71 156 105 190
rect 229 153 263 187
rect 338 102 372 136
rect 487 156 521 190
rect 592 127 626 161
rect 592 59 626 93
rect 678 169 712 203
rect 678 67 712 101
rect 782 169 816 203
rect 782 59 816 93
<< pdiffc >>
rect 35 563 69 597
rect 35 493 69 527
rect 125 553 159 587
rect 215 563 249 597
rect 215 495 249 529
rect 301 561 335 595
rect 301 493 335 527
rect 592 539 626 573
rect 405 384 439 418
rect 678 565 712 599
rect 678 478 712 512
rect 678 386 712 420
rect 782 573 816 607
rect 782 472 816 506
rect 782 379 816 413
<< poly >>
rect 80 609 110 635
rect 174 609 204 635
rect 260 609 290 635
rect 637 619 667 645
rect 723 619 753 645
rect 450 495 480 521
rect 522 495 552 521
rect 80 303 110 481
rect 174 443 204 481
rect 152 427 218 443
rect 152 393 168 427
rect 202 393 218 427
rect 152 359 218 393
rect 152 325 168 359
rect 202 325 218 359
rect 260 371 290 481
rect 260 355 358 371
rect 260 341 308 355
rect 152 309 218 325
rect 21 287 110 303
rect 21 253 37 287
rect 71 267 110 287
rect 71 253 146 267
rect 21 237 146 253
rect 116 215 146 237
rect 188 215 218 309
rect 274 321 308 341
rect 342 321 358 355
rect 274 287 358 321
rect 450 303 480 367
rect 274 253 308 287
rect 342 253 358 287
rect 274 237 358 253
rect 409 287 480 303
rect 409 253 425 287
rect 459 273 480 287
rect 522 308 552 367
rect 637 334 667 367
rect 723 334 753 367
rect 630 318 753 334
rect 522 292 588 308
rect 459 253 476 273
rect 409 237 476 253
rect 522 258 538 292
rect 572 258 588 292
rect 630 284 646 318
rect 680 284 753 318
rect 630 268 753 284
rect 522 242 588 258
rect 274 215 304 237
rect 446 215 476 237
rect 532 215 562 242
rect 637 215 667 268
rect 723 215 753 268
rect 116 105 146 131
rect 188 105 218 131
rect 274 105 304 131
rect 446 105 476 131
rect 532 105 562 131
rect 637 21 667 47
rect 723 21 753 47
<< polycont >>
rect 168 393 202 427
rect 168 325 202 359
rect 37 253 71 287
rect 308 321 342 355
rect 308 253 342 287
rect 425 253 459 287
rect 538 258 572 292
rect 646 284 680 318
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 19 597 73 615
rect 19 563 35 597
rect 69 563 73 597
rect 19 527 73 563
rect 109 587 175 649
rect 109 553 125 587
rect 159 553 175 587
rect 109 545 175 553
rect 211 597 258 613
rect 211 563 215 597
rect 249 563 258 597
rect 19 493 35 527
rect 69 511 73 527
rect 211 529 258 563
rect 211 511 215 529
rect 69 495 215 511
rect 249 495 258 529
rect 69 493 258 495
rect 19 477 258 493
rect 292 595 351 611
rect 292 561 301 595
rect 335 561 351 595
rect 292 527 351 561
rect 576 573 642 649
rect 576 539 592 573
rect 626 539 642 573
rect 576 528 642 539
rect 676 599 748 615
rect 676 565 678 599
rect 712 565 748 599
rect 292 493 301 527
rect 335 494 351 527
rect 676 512 748 565
rect 335 493 642 494
rect 292 460 642 493
rect 292 443 339 460
rect 17 287 79 443
rect 17 253 37 287
rect 71 253 79 287
rect 17 237 79 253
rect 113 427 204 443
rect 113 393 168 427
rect 202 393 204 427
rect 113 359 204 393
rect 113 325 168 359
rect 202 325 204 359
rect 113 237 204 325
rect 238 409 339 443
rect 389 418 455 426
rect 238 203 272 409
rect 389 384 405 418
rect 439 384 455 418
rect 389 371 455 384
rect 55 190 121 203
rect 55 156 71 190
rect 105 156 121 190
rect 55 17 121 156
rect 213 187 272 203
rect 213 153 229 187
rect 263 153 272 187
rect 306 355 455 371
rect 306 321 308 355
rect 342 337 455 355
rect 342 321 358 337
rect 306 287 358 321
rect 509 292 574 426
rect 306 253 308 287
rect 342 253 358 287
rect 306 206 358 253
rect 392 253 425 287
rect 459 253 475 287
rect 392 242 475 253
rect 509 258 538 292
rect 572 258 574 292
rect 608 334 642 460
rect 676 478 678 512
rect 712 478 748 512
rect 676 420 748 478
rect 676 386 678 420
rect 712 386 748 420
rect 676 370 748 386
rect 608 318 680 334
rect 608 284 646 318
rect 608 268 680 284
rect 509 242 574 258
rect 714 219 748 370
rect 782 607 824 649
rect 816 573 824 607
rect 782 506 824 573
rect 816 472 824 506
rect 782 413 824 472
rect 816 379 824 413
rect 782 363 824 379
rect 306 190 525 206
rect 306 172 487 190
rect 213 137 272 153
rect 483 156 487 172
rect 521 156 525 190
rect 674 203 748 219
rect 483 140 525 156
rect 588 161 626 177
rect 322 102 338 136
rect 372 102 388 136
rect 322 17 388 102
rect 588 127 592 161
rect 588 93 626 127
rect 588 59 592 93
rect 588 17 626 59
rect 674 169 678 203
rect 712 169 748 203
rect 674 101 748 169
rect 674 67 678 101
rect 712 67 748 101
rect 674 51 748 67
rect 782 203 824 219
rect 816 169 824 203
rect 782 93 824 169
rect 816 59 824 93
rect 782 17 824 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2bb2o_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5911858
string GDS_START 5903446
<< end >>
