magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 41 49 764 263
rect 0 0 768 49
<< scnmos >>
rect 124 69 154 237
rect 220 69 250 237
rect 306 69 336 237
rect 460 69 490 237
rect 546 69 576 237
rect 646 69 676 237
<< scpmoshvt >>
rect 123 367 153 619
rect 234 367 264 619
rect 328 367 358 619
rect 420 367 450 619
rect 574 367 604 619
rect 646 367 676 619
<< ndiff >>
rect 67 219 124 237
rect 67 185 79 219
rect 113 185 124 219
rect 67 115 124 185
rect 67 81 79 115
rect 113 81 124 115
rect 67 69 124 81
rect 154 192 220 237
rect 154 158 170 192
rect 204 158 220 192
rect 154 111 220 158
rect 154 77 170 111
rect 204 77 220 111
rect 154 69 220 77
rect 250 192 306 237
rect 250 158 261 192
rect 295 158 306 192
rect 250 111 306 158
rect 250 77 261 111
rect 295 77 306 111
rect 250 69 306 77
rect 336 133 460 237
rect 336 99 347 133
rect 381 99 415 133
rect 449 99 460 133
rect 336 69 460 99
rect 490 192 546 237
rect 490 158 501 192
rect 535 158 546 192
rect 490 111 546 158
rect 490 77 501 111
rect 535 77 546 111
rect 490 69 546 77
rect 576 229 646 237
rect 576 195 596 229
rect 630 195 646 229
rect 576 161 646 195
rect 576 127 596 161
rect 630 127 646 161
rect 576 69 646 127
rect 676 192 738 237
rect 676 158 692 192
rect 726 158 738 192
rect 676 111 738 158
rect 676 77 692 111
rect 726 77 738 111
rect 676 69 738 77
<< pdiff >>
rect 66 599 123 619
rect 66 565 74 599
rect 108 565 123 599
rect 66 510 123 565
rect 66 476 74 510
rect 108 476 123 510
rect 66 413 123 476
rect 66 379 74 413
rect 108 379 123 413
rect 66 367 123 379
rect 153 607 234 619
rect 153 573 176 607
rect 210 573 234 607
rect 153 496 234 573
rect 153 462 176 496
rect 210 462 234 496
rect 153 367 234 462
rect 264 367 328 619
rect 358 367 420 619
rect 450 607 574 619
rect 450 573 461 607
rect 495 573 529 607
rect 563 573 574 607
rect 450 513 574 573
rect 450 479 461 513
rect 495 479 529 513
rect 563 479 574 513
rect 450 420 574 479
rect 450 386 461 420
rect 495 386 529 420
rect 563 386 574 420
rect 450 367 574 386
rect 604 367 646 619
rect 676 607 729 619
rect 676 573 687 607
rect 721 573 729 607
rect 676 497 729 573
rect 676 463 687 497
rect 721 463 729 497
rect 676 367 729 463
<< ndiffc >>
rect 79 185 113 219
rect 79 81 113 115
rect 170 158 204 192
rect 170 77 204 111
rect 261 158 295 192
rect 261 77 295 111
rect 347 99 381 133
rect 415 99 449 133
rect 501 158 535 192
rect 501 77 535 111
rect 596 195 630 229
rect 596 127 630 161
rect 692 158 726 192
rect 692 77 726 111
<< pdiffc >>
rect 74 565 108 599
rect 74 476 108 510
rect 74 379 108 413
rect 176 573 210 607
rect 176 462 210 496
rect 461 573 495 607
rect 529 573 563 607
rect 461 479 495 513
rect 529 479 563 513
rect 461 386 495 420
rect 529 386 563 420
rect 687 573 721 607
rect 687 463 721 497
<< poly >>
rect 123 619 153 645
rect 234 619 264 645
rect 328 619 358 645
rect 420 619 450 645
rect 574 619 604 645
rect 646 619 676 645
rect 123 335 153 367
rect 88 319 154 335
rect 234 325 264 367
rect 328 325 358 367
rect 420 325 450 367
rect 574 335 604 367
rect 88 285 104 319
rect 138 285 154 319
rect 88 269 154 285
rect 124 237 154 269
rect 196 309 264 325
rect 196 275 214 309
rect 248 275 264 309
rect 196 259 264 275
rect 306 309 378 325
rect 306 275 328 309
rect 362 275 378 309
rect 306 259 378 275
rect 420 309 490 325
rect 420 275 440 309
rect 474 275 490 309
rect 420 259 490 275
rect 532 319 604 335
rect 532 285 548 319
rect 582 285 604 319
rect 532 269 604 285
rect 646 325 676 367
rect 646 309 738 325
rect 646 275 688 309
rect 722 275 738 309
rect 220 237 250 259
rect 306 237 336 259
rect 460 237 490 259
rect 546 237 576 269
rect 646 259 738 275
rect 646 237 676 259
rect 124 43 154 69
rect 220 43 250 69
rect 306 43 336 69
rect 460 43 490 69
rect 546 43 576 69
rect 646 43 676 69
<< polycont >>
rect 104 285 138 319
rect 214 275 248 309
rect 328 275 362 309
rect 440 275 474 309
rect 548 285 582 319
rect 688 275 722 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 599 112 615
rect 17 565 74 599
rect 108 565 112 599
rect 17 510 112 565
rect 17 476 74 510
rect 108 476 112 510
rect 17 413 112 476
rect 160 607 226 649
rect 160 573 176 607
rect 210 573 226 607
rect 160 496 226 573
rect 160 462 176 496
rect 210 462 226 496
rect 160 454 226 462
rect 443 607 582 615
rect 443 573 461 607
rect 495 573 529 607
rect 563 573 582 607
rect 443 513 582 573
rect 443 479 461 513
rect 495 479 529 513
rect 563 479 582 513
rect 443 420 582 479
rect 671 607 737 649
rect 671 573 687 607
rect 721 573 737 607
rect 671 497 737 573
rect 671 463 687 497
rect 721 463 737 497
rect 671 458 737 463
rect 17 379 74 413
rect 108 379 112 413
rect 17 363 112 379
rect 146 386 461 420
rect 495 386 529 420
rect 563 386 652 420
rect 17 235 53 363
rect 146 329 180 386
rect 88 319 180 329
rect 88 285 104 319
rect 138 285 180 319
rect 88 269 180 285
rect 214 309 271 351
rect 248 275 271 309
rect 214 242 271 275
rect 305 309 369 352
rect 305 275 328 309
rect 362 275 369 309
rect 305 242 369 275
rect 403 309 474 352
rect 403 275 440 309
rect 403 242 474 275
rect 508 319 584 352
rect 508 285 548 319
rect 582 285 584 319
rect 508 269 584 285
rect 618 235 652 386
rect 688 309 751 424
rect 722 275 751 309
rect 688 242 751 275
rect 17 219 120 235
rect 17 185 79 219
rect 113 185 120 219
rect 580 229 652 235
rect 17 115 120 185
rect 17 81 79 115
rect 113 81 120 115
rect 17 65 120 81
rect 154 192 220 208
rect 154 158 170 192
rect 204 158 220 192
rect 154 111 220 158
rect 154 77 170 111
rect 204 77 220 111
rect 154 17 220 77
rect 254 192 546 208
rect 254 158 261 192
rect 295 174 501 192
rect 295 158 297 174
rect 254 111 297 158
rect 499 158 501 174
rect 535 158 546 192
rect 254 77 261 111
rect 295 77 297 111
rect 254 61 297 77
rect 331 133 465 140
rect 331 99 347 133
rect 381 99 415 133
rect 449 99 465 133
rect 331 17 465 99
rect 499 111 546 158
rect 580 195 596 229
rect 630 195 652 229
rect 580 161 652 195
rect 580 127 596 161
rect 630 127 652 161
rect 580 119 652 127
rect 686 192 742 208
rect 686 158 692 192
rect 726 158 742 192
rect 499 77 501 111
rect 535 85 546 111
rect 686 111 742 158
rect 686 85 692 111
rect 535 77 692 85
rect 726 77 742 111
rect 499 51 742 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o32a_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1773022
string GDS_START 1765370
<< end >>
