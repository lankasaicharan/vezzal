magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 6 241 660 259
rect 6 49 1512 241
rect 0 0 1536 49
<< scnmos >>
rect 87 65 117 233
rect 173 65 203 233
rect 259 65 289 233
rect 359 65 389 233
rect 445 65 475 233
rect 531 65 561 233
rect 789 47 819 215
rect 875 47 905 215
rect 961 47 991 215
rect 1047 47 1077 215
rect 1141 47 1171 215
rect 1227 47 1257 215
rect 1313 47 1343 215
rect 1399 47 1429 215
<< scpmoshvt >>
rect 85 367 115 619
rect 171 367 201 619
rect 257 367 287 619
rect 359 367 389 619
rect 445 367 475 619
rect 531 367 561 619
rect 711 367 741 619
rect 797 367 827 619
rect 883 367 913 619
rect 969 367 999 619
rect 1164 367 1194 619
rect 1250 367 1280 619
rect 1336 367 1366 619
rect 1422 367 1452 619
<< ndiff >>
rect 32 192 87 233
rect 32 158 42 192
rect 76 158 87 192
rect 32 111 87 158
rect 32 77 42 111
rect 76 77 87 111
rect 32 65 87 77
rect 117 225 173 233
rect 117 191 128 225
rect 162 191 173 225
rect 117 153 173 191
rect 117 119 128 153
rect 162 119 173 153
rect 117 65 173 119
rect 203 225 259 233
rect 203 191 214 225
rect 248 191 259 225
rect 203 111 259 191
rect 203 77 214 111
rect 248 77 259 111
rect 203 65 259 77
rect 289 175 359 233
rect 289 141 300 175
rect 334 141 359 175
rect 289 107 359 141
rect 289 73 300 107
rect 334 73 359 107
rect 289 65 359 73
rect 389 107 445 233
rect 389 73 400 107
rect 434 73 445 107
rect 389 65 445 73
rect 475 179 531 233
rect 475 145 486 179
rect 520 145 531 179
rect 475 65 531 145
rect 561 225 634 233
rect 561 191 586 225
rect 620 191 634 225
rect 561 157 634 191
rect 561 123 586 157
rect 620 123 634 157
rect 561 65 634 123
rect 736 93 789 215
rect 736 59 744 93
rect 778 59 789 93
rect 736 47 789 59
rect 819 181 875 215
rect 819 147 830 181
rect 864 147 875 181
rect 819 101 875 147
rect 819 67 830 101
rect 864 67 875 101
rect 819 47 875 67
rect 905 106 961 215
rect 905 72 916 106
rect 950 72 961 106
rect 905 47 961 72
rect 991 181 1047 215
rect 991 147 1002 181
rect 1036 147 1047 181
rect 991 101 1047 147
rect 991 67 1002 101
rect 1036 67 1047 101
rect 991 47 1047 67
rect 1077 170 1141 215
rect 1077 136 1092 170
rect 1126 136 1141 170
rect 1077 93 1141 136
rect 1077 59 1092 93
rect 1126 59 1141 93
rect 1077 47 1141 59
rect 1171 203 1227 215
rect 1171 169 1182 203
rect 1216 169 1227 203
rect 1171 101 1227 169
rect 1171 67 1182 101
rect 1216 67 1227 101
rect 1171 47 1227 67
rect 1257 175 1313 215
rect 1257 141 1268 175
rect 1302 141 1313 175
rect 1257 89 1313 141
rect 1257 55 1268 89
rect 1302 55 1313 89
rect 1257 47 1313 55
rect 1343 203 1399 215
rect 1343 169 1354 203
rect 1388 169 1399 203
rect 1343 101 1399 169
rect 1343 67 1354 101
rect 1388 67 1399 101
rect 1343 47 1399 67
rect 1429 175 1486 215
rect 1429 141 1440 175
rect 1474 141 1486 175
rect 1429 89 1486 141
rect 1429 55 1440 89
rect 1474 55 1486 89
rect 1429 47 1486 55
<< pdiff >>
rect 32 599 85 619
rect 32 565 40 599
rect 74 565 85 599
rect 32 510 85 565
rect 32 476 40 510
rect 74 476 85 510
rect 32 413 85 476
rect 32 379 40 413
rect 74 379 85 413
rect 32 367 85 379
rect 115 607 171 619
rect 115 573 126 607
rect 160 573 171 607
rect 115 534 171 573
rect 115 500 126 534
rect 160 500 171 534
rect 115 465 171 500
rect 115 431 126 465
rect 160 431 171 465
rect 115 367 171 431
rect 201 599 257 619
rect 201 565 212 599
rect 246 565 257 599
rect 201 510 257 565
rect 201 476 212 510
rect 246 476 257 510
rect 201 413 257 476
rect 201 379 212 413
rect 246 379 257 413
rect 201 367 257 379
rect 287 566 359 619
rect 287 532 305 566
rect 339 532 359 566
rect 287 367 359 532
rect 389 599 445 619
rect 389 565 400 599
rect 434 565 445 599
rect 389 492 445 565
rect 389 458 400 492
rect 434 458 445 492
rect 389 367 445 458
rect 475 572 531 619
rect 475 538 486 572
rect 520 538 531 572
rect 475 367 531 538
rect 561 599 711 619
rect 561 565 572 599
rect 606 565 666 599
rect 700 565 711 599
rect 561 516 711 565
rect 561 482 572 516
rect 606 512 711 516
rect 606 482 666 512
rect 561 478 666 482
rect 700 478 711 512
rect 561 436 711 478
rect 561 402 581 436
rect 615 420 711 436
rect 615 402 666 420
rect 561 386 666 402
rect 700 386 711 420
rect 561 367 711 386
rect 741 599 797 619
rect 741 565 752 599
rect 786 565 797 599
rect 741 506 797 565
rect 741 472 752 506
rect 786 472 797 506
rect 741 367 797 472
rect 827 566 883 619
rect 827 532 838 566
rect 872 532 883 566
rect 827 367 883 532
rect 913 599 969 619
rect 913 565 924 599
rect 958 565 969 599
rect 913 506 969 565
rect 913 472 924 506
rect 958 472 969 506
rect 913 367 969 472
rect 999 599 1052 619
rect 999 565 1010 599
rect 1044 565 1052 599
rect 999 508 1052 565
rect 999 474 1010 508
rect 1044 474 1052 508
rect 999 413 1052 474
rect 999 379 1010 413
rect 1044 379 1052 413
rect 999 367 1052 379
rect 1111 607 1164 619
rect 1111 573 1119 607
rect 1153 573 1164 607
rect 1111 534 1164 573
rect 1111 500 1119 534
rect 1153 500 1164 534
rect 1111 455 1164 500
rect 1111 421 1119 455
rect 1153 421 1164 455
rect 1111 367 1164 421
rect 1194 599 1250 619
rect 1194 565 1205 599
rect 1239 565 1250 599
rect 1194 508 1250 565
rect 1194 474 1205 508
rect 1239 474 1250 508
rect 1194 413 1250 474
rect 1194 379 1205 413
rect 1239 379 1250 413
rect 1194 367 1250 379
rect 1280 607 1336 619
rect 1280 573 1291 607
rect 1325 573 1336 607
rect 1280 532 1336 573
rect 1280 498 1291 532
rect 1325 498 1336 532
rect 1280 453 1336 498
rect 1280 419 1291 453
rect 1325 419 1336 453
rect 1280 367 1336 419
rect 1366 599 1422 619
rect 1366 565 1377 599
rect 1411 565 1422 599
rect 1366 508 1422 565
rect 1366 474 1377 508
rect 1411 474 1422 508
rect 1366 413 1422 474
rect 1366 379 1377 413
rect 1411 379 1422 413
rect 1366 367 1422 379
rect 1452 607 1505 619
rect 1452 573 1463 607
rect 1497 573 1505 607
rect 1452 532 1505 573
rect 1452 498 1463 532
rect 1497 498 1505 532
rect 1452 453 1505 498
rect 1452 419 1463 453
rect 1497 419 1505 453
rect 1452 367 1505 419
<< ndiffc >>
rect 42 158 76 192
rect 42 77 76 111
rect 128 191 162 225
rect 128 119 162 153
rect 214 191 248 225
rect 214 77 248 111
rect 300 141 334 175
rect 300 73 334 107
rect 400 73 434 107
rect 486 145 520 179
rect 586 191 620 225
rect 586 123 620 157
rect 744 59 778 93
rect 830 147 864 181
rect 830 67 864 101
rect 916 72 950 106
rect 1002 147 1036 181
rect 1002 67 1036 101
rect 1092 136 1126 170
rect 1092 59 1126 93
rect 1182 169 1216 203
rect 1182 67 1216 101
rect 1268 141 1302 175
rect 1268 55 1302 89
rect 1354 169 1388 203
rect 1354 67 1388 101
rect 1440 141 1474 175
rect 1440 55 1474 89
<< pdiffc >>
rect 40 565 74 599
rect 40 476 74 510
rect 40 379 74 413
rect 126 573 160 607
rect 126 500 160 534
rect 126 431 160 465
rect 212 565 246 599
rect 212 476 246 510
rect 212 379 246 413
rect 305 532 339 566
rect 400 565 434 599
rect 400 458 434 492
rect 486 538 520 572
rect 572 565 606 599
rect 666 565 700 599
rect 572 482 606 516
rect 666 478 700 512
rect 581 402 615 436
rect 666 386 700 420
rect 752 565 786 599
rect 752 472 786 506
rect 838 532 872 566
rect 924 565 958 599
rect 924 472 958 506
rect 1010 565 1044 599
rect 1010 474 1044 508
rect 1010 379 1044 413
rect 1119 573 1153 607
rect 1119 500 1153 534
rect 1119 421 1153 455
rect 1205 565 1239 599
rect 1205 474 1239 508
rect 1205 379 1239 413
rect 1291 573 1325 607
rect 1291 498 1325 532
rect 1291 419 1325 453
rect 1377 565 1411 599
rect 1377 474 1411 508
rect 1377 379 1411 413
rect 1463 573 1497 607
rect 1463 498 1497 532
rect 1463 419 1497 453
<< poly >>
rect 85 619 115 645
rect 171 619 201 645
rect 257 619 287 645
rect 359 619 389 645
rect 445 619 475 645
rect 531 619 561 645
rect 711 619 741 645
rect 797 619 827 645
rect 883 619 913 645
rect 969 619 999 645
rect 1164 619 1194 645
rect 1250 619 1280 645
rect 1336 619 1366 645
rect 1422 619 1452 645
rect 85 321 115 367
rect 171 321 201 367
rect 257 335 287 367
rect 359 335 389 367
rect 445 335 475 367
rect 24 305 201 321
rect 24 271 40 305
rect 74 271 201 305
rect 24 269 201 271
rect 245 319 311 335
rect 245 285 261 319
rect 295 285 311 319
rect 245 269 311 285
rect 359 319 475 335
rect 359 285 399 319
rect 433 285 475 319
rect 359 269 475 285
rect 24 255 203 269
rect 87 233 117 255
rect 173 233 203 255
rect 259 233 289 269
rect 359 233 389 269
rect 445 233 475 269
rect 531 335 561 367
rect 531 319 616 335
rect 531 285 547 319
rect 581 285 616 319
rect 711 303 741 367
rect 797 345 827 367
rect 883 345 913 367
rect 969 345 999 367
rect 797 319 927 345
rect 797 315 877 319
rect 531 269 616 285
rect 689 287 755 303
rect 531 233 561 269
rect 689 253 705 287
rect 739 267 755 287
rect 861 285 877 315
rect 911 285 927 319
rect 969 315 1099 345
rect 1164 331 1194 367
rect 1250 331 1280 367
rect 1336 331 1366 367
rect 1422 331 1452 367
rect 861 267 927 285
rect 1033 281 1049 315
rect 1083 281 1099 315
rect 739 253 819 267
rect 689 237 819 253
rect 861 237 991 267
rect 1033 265 1099 281
rect 1141 315 1452 331
rect 1141 281 1157 315
rect 1191 281 1225 315
rect 1259 281 1293 315
rect 1327 281 1361 315
rect 1395 281 1452 315
rect 1141 265 1452 281
rect 789 215 819 237
rect 875 215 905 237
rect 961 215 991 237
rect 1047 215 1077 265
rect 1141 215 1171 265
rect 1227 215 1257 265
rect 1313 215 1343 265
rect 1399 215 1429 265
rect 87 39 117 65
rect 173 39 203 65
rect 259 39 289 65
rect 359 39 389 65
rect 445 39 475 65
rect 531 39 561 65
rect 789 21 819 47
rect 875 21 905 47
rect 961 21 991 47
rect 1047 21 1077 47
rect 1141 21 1171 47
rect 1227 21 1257 47
rect 1313 21 1343 47
rect 1399 21 1429 47
<< polycont >>
rect 40 271 74 305
rect 261 285 295 319
rect 399 285 433 319
rect 547 285 581 319
rect 705 253 739 287
rect 877 285 911 319
rect 1049 281 1083 315
rect 1157 281 1191 315
rect 1225 281 1259 315
rect 1293 281 1327 315
rect 1361 281 1395 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 24 599 76 615
rect 24 565 40 599
rect 74 565 76 599
rect 24 510 76 565
rect 24 476 40 510
rect 74 476 76 510
rect 24 413 76 476
rect 110 607 176 649
rect 110 573 126 607
rect 160 573 176 607
rect 110 534 176 573
rect 110 500 126 534
rect 160 500 176 534
rect 110 465 176 500
rect 110 431 126 465
rect 160 431 176 465
rect 210 599 255 615
rect 210 565 212 599
rect 246 565 255 599
rect 210 510 255 565
rect 289 566 355 649
rect 289 532 305 566
rect 339 532 355 566
rect 289 526 355 532
rect 389 599 436 615
rect 389 565 400 599
rect 434 565 436 599
rect 210 476 212 510
rect 246 492 255 510
rect 389 494 436 565
rect 470 572 536 649
rect 470 538 486 572
rect 520 538 536 572
rect 470 528 536 538
rect 570 599 709 615
rect 570 565 572 599
rect 606 565 666 599
rect 700 565 709 599
rect 570 516 709 565
rect 570 494 572 516
rect 389 492 572 494
rect 246 476 400 492
rect 210 458 400 476
rect 434 482 572 492
rect 606 512 709 516
rect 606 482 666 512
rect 434 478 666 482
rect 700 478 709 512
rect 434 458 709 478
rect 24 379 40 413
rect 74 397 76 413
rect 210 413 250 458
rect 581 436 709 458
rect 743 599 788 615
rect 743 565 752 599
rect 786 565 788 599
rect 743 506 788 565
rect 822 566 888 649
rect 822 532 838 566
rect 872 532 888 566
rect 822 524 888 532
rect 922 599 968 615
rect 922 565 924 599
rect 958 565 968 599
rect 743 472 752 506
rect 786 490 788 506
rect 922 506 968 565
rect 922 490 924 506
rect 786 472 924 490
rect 958 472 968 506
rect 743 456 968 472
rect 1002 599 1060 615
rect 1002 565 1010 599
rect 1044 565 1060 599
rect 1002 508 1060 565
rect 1002 474 1010 508
rect 1044 474 1060 508
rect 210 397 212 413
rect 74 379 212 397
rect 246 379 250 413
rect 24 363 250 379
rect 286 390 547 424
rect 17 305 78 321
rect 17 271 40 305
rect 74 271 78 305
rect 17 242 78 271
rect 112 225 178 363
rect 286 329 320 390
rect 245 319 320 329
rect 245 285 261 319
rect 295 285 320 319
rect 354 319 475 356
rect 354 285 399 319
rect 433 285 475 319
rect 511 285 547 390
rect 615 420 709 436
rect 1002 420 1060 474
rect 1103 607 1169 649
rect 1103 573 1119 607
rect 1153 573 1169 607
rect 1103 534 1169 573
rect 1103 500 1119 534
rect 1153 500 1169 534
rect 1103 455 1169 500
rect 1103 421 1119 455
rect 1153 421 1169 455
rect 1203 599 1241 615
rect 1203 565 1205 599
rect 1239 565 1241 599
rect 1203 508 1241 565
rect 1203 474 1205 508
rect 1239 474 1241 508
rect 615 402 666 420
rect 581 386 666 402
rect 700 413 1060 420
rect 700 386 1010 413
rect 994 379 1010 386
rect 1044 385 1060 413
rect 1203 413 1241 474
rect 1275 607 1341 649
rect 1275 573 1291 607
rect 1325 573 1341 607
rect 1275 532 1341 573
rect 1275 498 1291 532
rect 1325 498 1341 532
rect 1275 453 1341 498
rect 1275 419 1291 453
rect 1325 419 1341 453
rect 1375 599 1413 615
rect 1375 565 1377 599
rect 1411 565 1413 599
rect 1375 508 1413 565
rect 1375 474 1377 508
rect 1411 474 1413 508
rect 1044 379 1169 385
rect 581 285 597 319
rect 674 287 755 350
rect 674 253 705 287
rect 739 253 755 287
rect 789 319 956 352
rect 994 351 1169 379
rect 1203 379 1205 413
rect 1239 385 1241 413
rect 1375 413 1413 474
rect 1447 607 1513 649
rect 1447 573 1463 607
rect 1497 573 1513 607
rect 1447 532 1513 573
rect 1447 498 1463 532
rect 1497 498 1513 532
rect 1447 453 1513 498
rect 1447 419 1463 453
rect 1497 419 1513 453
rect 1375 385 1377 413
rect 1239 379 1377 385
rect 1411 385 1413 413
rect 1411 379 1519 385
rect 1203 351 1519 379
rect 789 285 877 319
rect 911 285 956 319
rect 1135 317 1169 351
rect 789 283 956 285
rect 1033 315 1099 317
rect 26 192 78 208
rect 26 158 42 192
rect 76 158 78 192
rect 26 111 78 158
rect 112 191 128 225
rect 162 191 178 225
rect 112 153 178 191
rect 112 119 128 153
rect 162 119 178 153
rect 212 225 636 251
rect 212 191 214 225
rect 248 217 586 225
rect 248 191 250 217
rect 26 77 42 111
rect 76 85 78 111
rect 212 111 250 191
rect 570 191 586 217
rect 620 191 636 225
rect 674 249 755 253
rect 1033 281 1049 315
rect 1083 281 1099 315
rect 1135 315 1411 317
rect 1135 281 1157 315
rect 1191 281 1225 315
rect 1259 281 1293 315
rect 1327 281 1361 315
rect 1395 281 1411 315
rect 1033 265 1099 281
rect 1033 249 1067 265
rect 674 215 1067 249
rect 1447 247 1519 351
rect 212 85 214 111
rect 76 77 214 85
rect 248 77 250 111
rect 26 51 250 77
rect 284 179 536 183
rect 284 175 486 179
rect 284 141 300 175
rect 334 145 486 175
rect 520 145 536 179
rect 334 141 350 145
rect 284 107 350 141
rect 475 136 536 145
rect 570 157 636 191
rect 1173 213 1519 247
rect 1173 203 1218 213
rect 570 123 586 157
rect 620 123 636 157
rect 570 119 636 123
rect 670 147 830 181
rect 864 147 1002 181
rect 1036 147 1052 181
rect 670 145 866 147
rect 284 73 300 107
rect 334 73 350 107
rect 284 57 350 73
rect 384 107 450 111
rect 384 73 400 107
rect 434 85 450 107
rect 670 85 704 145
rect 434 73 704 85
rect 384 51 704 73
rect 738 93 787 109
rect 738 59 744 93
rect 778 59 787 93
rect 738 17 787 59
rect 821 101 866 145
rect 821 67 830 101
rect 864 67 866 101
rect 821 51 866 67
rect 900 106 966 113
rect 900 72 916 106
rect 950 72 966 106
rect 900 17 966 72
rect 1000 101 1052 147
rect 1000 67 1002 101
rect 1036 67 1052 101
rect 1000 51 1052 67
rect 1086 170 1139 186
rect 1086 136 1092 170
rect 1126 136 1139 170
rect 1086 93 1139 136
rect 1086 59 1092 93
rect 1126 59 1139 93
rect 1086 17 1139 59
rect 1173 169 1182 203
rect 1216 169 1218 203
rect 1352 203 1390 213
rect 1173 101 1218 169
rect 1173 67 1182 101
rect 1216 67 1218 101
rect 1173 51 1218 67
rect 1252 175 1318 179
rect 1252 141 1268 175
rect 1302 141 1318 175
rect 1252 89 1318 141
rect 1252 55 1268 89
rect 1302 55 1318 89
rect 1252 17 1318 55
rect 1352 169 1354 203
rect 1388 169 1390 203
rect 1352 101 1390 169
rect 1352 67 1354 101
rect 1388 67 1390 101
rect 1352 51 1390 67
rect 1424 175 1490 179
rect 1424 141 1440 175
rect 1474 141 1490 175
rect 1424 89 1490 141
rect 1424 55 1440 89
rect 1474 55 1490 89
rect 1424 17 1490 55
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2111a_4
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4152892
string GDS_START 4139776
<< end >>
