magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
rect 427 299 1530 331
<< pwell >>
rect 1 159 427 222
rect 1588 159 2014 184
rect 1 49 2014 159
rect 0 0 2016 49
<< scnmos >>
rect 84 112 114 196
rect 156 112 186 196
rect 242 112 272 196
rect 314 112 344 196
rect 512 49 542 133
rect 584 49 614 133
rect 670 49 700 133
rect 748 49 778 133
rect 914 49 944 133
rect 1028 49 1058 133
rect 1243 49 1273 133
rect 1315 49 1345 133
rect 1401 49 1431 133
rect 1473 49 1503 133
rect 1671 74 1701 158
rect 1743 74 1773 158
rect 1829 74 1859 158
rect 1901 74 1931 158
<< scpmoshvt >>
rect 116 419 166 619
rect 222 419 272 619
rect 520 335 570 535
rect 642 367 692 567
rect 740 367 790 567
rect 905 367 955 567
rect 1028 367 1078 567
rect 1142 367 1192 567
rect 1280 347 1330 547
rect 1387 347 1437 547
rect 1723 374 1773 574
rect 1829 374 1879 574
<< ndiff >>
rect 27 171 84 196
rect 27 137 39 171
rect 73 137 84 171
rect 27 112 84 137
rect 114 112 156 196
rect 186 171 242 196
rect 186 137 197 171
rect 231 137 242 171
rect 186 112 242 137
rect 272 112 314 196
rect 344 171 401 196
rect 344 137 355 171
rect 389 137 401 171
rect 344 112 401 137
rect 1614 133 1671 158
rect 455 112 512 133
rect 455 78 467 112
rect 501 78 512 112
rect 455 49 512 78
rect 542 49 584 133
rect 614 100 670 133
rect 614 66 625 100
rect 659 66 670 100
rect 614 49 670 66
rect 700 49 748 133
rect 778 112 914 133
rect 778 78 860 112
rect 894 78 914 112
rect 778 49 914 78
rect 944 49 1028 133
rect 1058 108 1132 133
rect 1058 74 1086 108
rect 1120 74 1132 108
rect 1058 49 1132 74
rect 1186 108 1243 133
rect 1186 74 1198 108
rect 1232 74 1243 108
rect 1186 49 1243 74
rect 1273 49 1315 133
rect 1345 108 1401 133
rect 1345 74 1356 108
rect 1390 74 1401 108
rect 1345 49 1401 74
rect 1431 49 1473 133
rect 1503 112 1560 133
rect 1503 78 1514 112
rect 1548 78 1560 112
rect 1503 49 1560 78
rect 1614 99 1626 133
rect 1660 99 1671 133
rect 1614 74 1671 99
rect 1701 74 1743 158
rect 1773 133 1829 158
rect 1773 99 1784 133
rect 1818 99 1829 133
rect 1773 74 1829 99
rect 1859 74 1901 158
rect 1931 133 1988 158
rect 1931 99 1942 133
rect 1976 99 1988 133
rect 1931 74 1988 99
<< pdiff >>
rect 59 597 116 619
rect 59 563 71 597
rect 105 563 116 597
rect 59 465 116 563
rect 59 431 71 465
rect 105 431 116 465
rect 59 419 116 431
rect 166 607 222 619
rect 166 573 177 607
rect 211 573 222 607
rect 166 419 222 573
rect 272 466 329 619
rect 585 554 642 567
rect 585 535 597 554
rect 272 432 283 466
rect 317 432 329 466
rect 272 419 329 432
rect 463 381 520 535
rect 463 347 475 381
rect 509 347 520 381
rect 463 335 520 347
rect 570 520 597 535
rect 631 520 642 554
rect 570 367 642 520
rect 692 367 740 567
rect 790 527 905 567
rect 790 493 852 527
rect 886 493 905 527
rect 790 413 905 493
rect 790 379 852 413
rect 886 379 905 413
rect 790 367 905 379
rect 955 367 1028 567
rect 1078 555 1142 567
rect 1078 521 1089 555
rect 1123 521 1142 555
rect 1078 463 1142 521
rect 1078 429 1089 463
rect 1123 429 1142 463
rect 1078 367 1142 429
rect 1192 555 1265 567
rect 1192 521 1219 555
rect 1253 547 1265 555
rect 1253 521 1280 547
rect 1192 474 1280 521
rect 1192 440 1219 474
rect 1253 440 1280 474
rect 1192 393 1280 440
rect 1192 367 1219 393
rect 570 335 620 367
rect 1207 359 1219 367
rect 1253 359 1280 393
rect 1207 347 1280 359
rect 1330 535 1387 547
rect 1330 501 1341 535
rect 1375 501 1387 535
rect 1330 464 1387 501
rect 1330 430 1341 464
rect 1375 430 1387 464
rect 1330 393 1387 430
rect 1330 359 1341 393
rect 1375 359 1387 393
rect 1330 347 1387 359
rect 1437 535 1494 547
rect 1437 501 1448 535
rect 1482 501 1494 535
rect 1437 464 1494 501
rect 1437 430 1448 464
rect 1482 430 1494 464
rect 1666 562 1723 574
rect 1666 528 1678 562
rect 1712 528 1723 562
rect 1666 491 1723 528
rect 1666 457 1678 491
rect 1712 457 1723 491
rect 1437 393 1494 430
rect 1437 359 1448 393
rect 1482 359 1494 393
rect 1666 420 1723 457
rect 1666 386 1678 420
rect 1712 386 1723 420
rect 1666 374 1723 386
rect 1773 562 1829 574
rect 1773 528 1784 562
rect 1818 528 1829 562
rect 1773 491 1829 528
rect 1773 457 1784 491
rect 1818 457 1829 491
rect 1773 420 1829 457
rect 1773 386 1784 420
rect 1818 386 1829 420
rect 1773 374 1829 386
rect 1879 562 1936 574
rect 1879 528 1890 562
rect 1924 528 1936 562
rect 1879 491 1936 528
rect 1879 457 1890 491
rect 1924 457 1936 491
rect 1879 420 1936 457
rect 1879 386 1890 420
rect 1924 386 1936 420
rect 1879 374 1936 386
rect 1437 347 1494 359
<< ndiffc >>
rect 39 137 73 171
rect 197 137 231 171
rect 355 137 389 171
rect 467 78 501 112
rect 625 66 659 100
rect 860 78 894 112
rect 1086 74 1120 108
rect 1198 74 1232 108
rect 1356 74 1390 108
rect 1514 78 1548 112
rect 1626 99 1660 133
rect 1784 99 1818 133
rect 1942 99 1976 133
<< pdiffc >>
rect 71 563 105 597
rect 71 431 105 465
rect 177 573 211 607
rect 283 432 317 466
rect 475 347 509 381
rect 597 520 631 554
rect 852 493 886 527
rect 852 379 886 413
rect 1089 521 1123 555
rect 1089 429 1123 463
rect 1219 521 1253 555
rect 1219 440 1253 474
rect 1219 359 1253 393
rect 1341 501 1375 535
rect 1341 430 1375 464
rect 1341 359 1375 393
rect 1448 501 1482 535
rect 1448 430 1482 464
rect 1678 528 1712 562
rect 1678 457 1712 491
rect 1448 359 1482 393
rect 1678 386 1712 420
rect 1784 528 1818 562
rect 1784 457 1818 491
rect 1784 386 1818 420
rect 1890 528 1924 562
rect 1890 457 1924 491
rect 1890 386 1924 420
<< poly >>
rect 116 619 166 645
rect 222 619 272 645
rect 365 609 692 639
rect 365 597 431 609
rect 365 563 381 597
rect 415 563 431 597
rect 642 567 692 609
rect 1280 615 1589 645
rect 740 567 790 593
rect 905 567 955 593
rect 1028 567 1078 593
rect 1142 567 1192 593
rect 365 547 431 563
rect 520 535 570 561
rect 116 370 166 419
rect 84 354 166 370
rect 84 320 116 354
rect 150 320 166 354
rect 222 370 272 419
rect 222 354 344 370
rect 222 340 285 354
rect 84 286 166 320
rect 84 252 116 286
rect 150 266 166 286
rect 242 320 285 340
rect 319 320 344 354
rect 1280 547 1330 615
rect 1559 578 1589 615
rect 1387 547 1437 573
rect 1559 562 1625 578
rect 1723 574 1773 600
rect 1829 574 1879 600
rect 642 341 692 367
rect 242 286 344 320
rect 520 293 570 335
rect 150 252 186 266
rect 84 236 186 252
rect 84 196 114 236
rect 156 196 186 236
rect 242 252 285 286
rect 319 252 344 286
rect 242 236 344 252
rect 242 196 272 236
rect 314 196 344 236
rect 512 277 614 293
rect 512 243 545 277
rect 579 243 614 277
rect 512 227 614 243
rect 512 133 542 227
rect 584 133 614 227
rect 662 221 692 341
rect 740 335 790 367
rect 734 319 800 335
rect 734 285 750 319
rect 784 285 800 319
rect 905 317 955 367
rect 734 269 800 285
rect 842 287 955 317
rect 1028 335 1078 367
rect 1028 319 1094 335
rect 842 221 872 287
rect 1028 285 1044 319
rect 1078 285 1094 319
rect 1028 269 1094 285
rect 1142 307 1192 367
rect 1559 528 1575 562
rect 1609 528 1625 562
rect 1559 494 1625 528
rect 1559 460 1575 494
rect 1609 460 1625 494
rect 1559 444 1625 460
rect 1142 291 1208 307
rect 662 191 700 221
rect 670 133 700 191
rect 742 205 872 221
rect 742 171 758 205
rect 792 191 872 205
rect 914 223 980 239
rect 792 171 808 191
rect 742 155 808 171
rect 914 189 930 223
rect 964 189 980 223
rect 914 173 980 189
rect 748 133 778 155
rect 914 133 944 173
rect 1028 133 1058 269
rect 1142 257 1158 291
rect 1192 257 1208 291
rect 1280 305 1330 347
rect 1387 307 1437 347
rect 1280 275 1345 305
rect 1142 223 1208 257
rect 1142 189 1158 223
rect 1192 203 1208 223
rect 1192 189 1273 203
rect 1142 173 1273 189
rect 1243 133 1273 173
rect 1315 133 1345 275
rect 1387 291 1453 307
rect 1387 257 1403 291
rect 1437 257 1453 291
rect 1387 223 1453 257
rect 1387 189 1403 223
rect 1437 203 1453 223
rect 1723 203 1773 374
rect 1437 189 1773 203
rect 1387 173 1773 189
rect 1401 133 1431 173
rect 1473 133 1503 173
rect 1671 158 1701 173
rect 1743 158 1773 173
rect 1829 332 1879 374
rect 1829 316 1895 332
rect 1829 282 1845 316
rect 1879 282 1895 316
rect 1829 248 1895 282
rect 1829 214 1845 248
rect 1879 228 1895 248
rect 1879 214 1931 228
rect 1829 198 1931 214
rect 1829 158 1859 198
rect 1901 158 1931 198
rect 84 86 114 112
rect 156 86 186 112
rect 242 86 272 112
rect 314 86 344 112
rect 512 23 542 49
rect 584 23 614 49
rect 670 23 700 49
rect 748 23 778 49
rect 914 23 944 49
rect 1028 23 1058 49
rect 1243 23 1273 49
rect 1315 23 1345 49
rect 1401 23 1431 49
rect 1473 23 1503 49
rect 1671 48 1701 74
rect 1743 48 1773 74
rect 1829 48 1859 74
rect 1901 48 1931 74
<< polycont >>
rect 381 563 415 597
rect 116 320 150 354
rect 116 252 150 286
rect 285 320 319 354
rect 285 252 319 286
rect 545 243 579 277
rect 750 285 784 319
rect 1044 285 1078 319
rect 1575 528 1609 562
rect 1575 460 1609 494
rect 758 171 792 205
rect 930 189 964 223
rect 1158 257 1192 291
rect 1158 189 1192 223
rect 1403 257 1437 291
rect 1403 189 1437 223
rect 1845 282 1879 316
rect 1845 214 1879 248
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 597 121 613
rect 23 563 71 597
rect 105 563 121 597
rect 161 607 227 649
rect 161 573 177 607
rect 211 573 227 607
rect 365 597 431 613
rect 23 537 121 563
rect 365 563 381 597
rect 415 563 431 597
rect 365 537 431 563
rect 23 503 431 537
rect 581 554 647 649
rect 581 520 597 554
rect 631 520 647 554
rect 581 503 647 520
rect 734 579 980 613
rect 23 465 121 503
rect 23 431 71 465
rect 105 431 121 465
rect 23 415 121 431
rect 267 466 595 467
rect 267 432 283 466
rect 317 433 595 466
rect 317 432 333 433
rect 267 415 333 432
rect 23 200 57 415
rect 100 354 167 370
rect 100 320 116 354
rect 150 320 167 354
rect 100 286 167 320
rect 100 252 116 286
rect 150 252 167 286
rect 100 236 167 252
rect 217 354 335 370
rect 217 320 285 354
rect 319 320 335 354
rect 217 286 335 320
rect 217 252 285 286
rect 319 252 335 286
rect 217 236 335 252
rect 371 200 405 433
rect 23 171 89 200
rect 23 137 39 171
rect 73 137 89 171
rect 23 108 89 137
rect 181 171 247 200
rect 181 137 197 171
rect 231 137 247 171
rect 181 17 247 137
rect 339 171 405 200
rect 339 137 355 171
rect 389 137 405 171
rect 339 108 405 137
rect 451 381 525 397
rect 451 347 475 381
rect 509 347 525 381
rect 451 331 525 347
rect 561 335 595 433
rect 734 335 800 579
rect 836 527 902 543
rect 836 493 852 527
rect 886 493 902 527
rect 836 413 902 493
rect 836 379 852 413
rect 886 379 902 413
rect 836 363 902 379
rect 451 191 485 331
rect 561 319 800 335
rect 561 293 750 319
rect 529 285 750 293
rect 784 285 800 319
rect 529 277 800 285
rect 529 243 545 277
rect 579 269 800 277
rect 579 243 595 269
rect 529 227 595 243
rect 742 205 808 221
rect 742 191 758 205
rect 451 171 758 191
rect 792 171 808 205
rect 451 157 808 171
rect 451 112 517 157
rect 742 155 808 157
rect 844 137 878 363
rect 946 239 980 579
rect 1073 555 1139 649
rect 1073 521 1089 555
rect 1123 521 1139 555
rect 1073 463 1139 521
rect 1073 429 1089 463
rect 1123 429 1139 463
rect 1073 413 1139 429
rect 1203 555 1278 571
rect 1203 521 1219 555
rect 1253 521 1278 555
rect 1203 474 1278 521
rect 1203 440 1219 474
rect 1253 440 1278 474
rect 1203 393 1278 440
rect 1203 377 1219 393
rect 1028 359 1219 377
rect 1253 359 1278 393
rect 1028 343 1278 359
rect 1325 535 1391 649
rect 1325 501 1341 535
rect 1375 501 1391 535
rect 1325 464 1391 501
rect 1325 430 1341 464
rect 1375 430 1391 464
rect 1325 393 1391 430
rect 1325 359 1341 393
rect 1375 359 1391 393
rect 1325 343 1391 359
rect 1432 535 1523 578
rect 1432 501 1448 535
rect 1482 501 1523 535
rect 1432 464 1523 501
rect 1432 430 1448 464
rect 1482 430 1523 464
rect 1432 393 1523 430
rect 1432 359 1448 393
rect 1482 359 1523 393
rect 1559 562 1625 578
rect 1559 528 1575 562
rect 1609 528 1625 562
rect 1559 494 1625 528
rect 1559 460 1575 494
rect 1609 460 1625 494
rect 1559 384 1625 460
rect 1662 562 1728 578
rect 1662 528 1678 562
rect 1712 528 1728 562
rect 1662 491 1728 528
rect 1662 457 1678 491
rect 1712 457 1728 491
rect 1662 420 1728 457
rect 1662 386 1678 420
rect 1712 386 1728 420
rect 1432 343 1523 359
rect 1028 319 1094 343
rect 1028 285 1044 319
rect 1078 285 1094 319
rect 1244 307 1278 343
rect 1028 269 1094 285
rect 1142 291 1208 307
rect 914 223 980 239
rect 914 189 930 223
rect 964 189 980 223
rect 1142 257 1158 291
rect 1192 257 1208 291
rect 1142 223 1208 257
rect 1142 207 1158 223
rect 914 173 980 189
rect 1016 189 1158 207
rect 1192 189 1208 223
rect 1016 173 1208 189
rect 1244 291 1453 307
rect 1244 273 1403 291
rect 1016 137 1050 173
rect 1244 137 1278 273
rect 1387 257 1403 273
rect 1437 257 1453 291
rect 1387 223 1453 257
rect 1387 189 1403 223
rect 1437 189 1453 223
rect 1387 173 1453 189
rect 1489 137 1523 343
rect 1662 232 1728 386
rect 1768 562 1834 649
rect 1768 528 1784 562
rect 1818 528 1834 562
rect 1768 491 1834 528
rect 1768 457 1784 491
rect 1818 457 1834 491
rect 1768 420 1834 457
rect 1768 386 1784 420
rect 1818 386 1834 420
rect 1768 370 1834 386
rect 1874 562 1992 578
rect 1874 528 1890 562
rect 1924 528 1992 562
rect 1874 491 1992 528
rect 1874 457 1890 491
rect 1924 457 1992 491
rect 1874 420 1992 457
rect 1874 386 1890 420
rect 1924 386 1992 420
rect 1874 370 1992 386
rect 1829 316 1895 332
rect 1829 282 1845 316
rect 1879 282 1895 316
rect 1829 248 1895 282
rect 1829 232 1845 248
rect 1610 214 1845 232
rect 1879 214 1895 248
rect 1610 198 1895 214
rect 451 78 467 112
rect 501 78 517 112
rect 451 53 517 78
rect 609 100 675 121
rect 609 66 625 100
rect 659 66 675 100
rect 609 17 675 66
rect 844 112 1050 137
rect 844 78 860 112
rect 894 103 1050 112
rect 1086 108 1136 137
rect 894 78 910 103
rect 844 53 910 78
rect 1120 74 1136 108
rect 1086 17 1136 74
rect 1182 108 1278 137
rect 1182 74 1198 108
rect 1232 74 1278 108
rect 1182 61 1278 74
rect 1340 108 1406 137
rect 1340 74 1356 108
rect 1390 74 1406 108
rect 1340 17 1406 74
rect 1489 112 1564 137
rect 1489 78 1514 112
rect 1548 78 1564 112
rect 1489 53 1564 78
rect 1610 133 1676 198
rect 1945 162 1992 370
rect 1610 99 1626 133
rect 1660 99 1676 133
rect 1610 70 1676 99
rect 1768 133 1834 162
rect 1768 99 1784 133
rect 1818 99 1834 133
rect 1768 17 1834 99
rect 1926 133 1992 162
rect 1926 99 1942 133
rect 1976 99 1992 133
rect 1926 70 1992 99
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrbp_lp
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1471 390 1505 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 464 1505 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 538 1505 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1951 94 1985 128 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1951 168 1985 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1951 390 1985 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1951 464 1985 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1951 538 1985 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4320518
string GDS_START 4305862
<< end >>
