magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
rect 277 329 790 331
<< pwell >>
rect 129 49 1140 241
rect 0 0 1248 49
<< scnmos >>
rect 208 47 238 215
rect 294 47 324 215
rect 380 47 410 215
rect 499 47 529 215
rect 585 47 615 215
rect 683 47 713 215
rect 769 47 799 215
rect 855 47 885 215
rect 941 47 971 215
rect 1027 47 1057 215
<< scpmoshvt >>
rect 90 367 120 619
rect 176 367 206 619
rect 366 365 396 617
rect 452 365 482 617
rect 585 365 615 617
rect 671 365 701 617
rect 861 367 891 619
rect 947 367 977 619
rect 1033 367 1063 619
rect 1119 367 1149 619
<< ndiff >>
rect 155 169 208 215
rect 155 135 163 169
rect 197 135 208 169
rect 155 95 208 135
rect 155 61 163 95
rect 197 61 208 95
rect 155 47 208 61
rect 238 169 294 215
rect 238 135 249 169
rect 283 135 294 169
rect 238 47 294 135
rect 324 203 380 215
rect 324 169 335 203
rect 369 169 380 203
rect 324 101 380 169
rect 324 67 335 101
rect 369 67 380 101
rect 324 47 380 67
rect 410 165 499 215
rect 410 131 436 165
rect 470 131 499 165
rect 410 89 499 131
rect 410 55 436 89
rect 470 55 499 89
rect 410 47 499 55
rect 529 203 585 215
rect 529 169 540 203
rect 574 169 585 203
rect 529 101 585 169
rect 529 67 540 101
rect 574 67 585 101
rect 529 47 585 67
rect 615 165 683 215
rect 615 131 630 165
rect 664 131 683 165
rect 615 89 683 131
rect 615 55 630 89
rect 664 55 683 89
rect 615 47 683 55
rect 713 203 769 215
rect 713 169 724 203
rect 758 169 769 203
rect 713 101 769 169
rect 713 67 724 101
rect 758 67 769 101
rect 713 47 769 67
rect 799 165 855 215
rect 799 131 810 165
rect 844 131 855 165
rect 799 89 855 131
rect 799 55 810 89
rect 844 55 855 89
rect 799 47 855 55
rect 885 203 941 215
rect 885 169 896 203
rect 930 169 941 203
rect 885 101 941 169
rect 885 67 896 101
rect 930 67 941 101
rect 885 47 941 67
rect 971 165 1027 215
rect 971 131 982 165
rect 1016 131 1027 165
rect 971 89 1027 131
rect 971 55 982 89
rect 1016 55 1027 89
rect 971 47 1027 55
rect 1057 203 1114 215
rect 1057 169 1072 203
rect 1106 169 1114 203
rect 1057 101 1114 169
rect 1057 67 1072 101
rect 1106 67 1114 101
rect 1057 47 1114 67
<< pdiff >>
rect 37 607 90 619
rect 37 573 45 607
rect 79 573 90 607
rect 37 505 90 573
rect 37 471 45 505
rect 79 471 90 505
rect 37 413 90 471
rect 37 379 45 413
rect 79 379 90 413
rect 37 367 90 379
rect 120 599 176 619
rect 120 565 131 599
rect 165 565 176 599
rect 120 505 176 565
rect 120 471 131 505
rect 165 471 176 505
rect 120 413 176 471
rect 120 379 131 413
rect 165 379 176 413
rect 120 367 176 379
rect 206 607 259 619
rect 206 573 217 607
rect 251 573 259 607
rect 206 523 259 573
rect 206 489 217 523
rect 251 489 259 523
rect 206 443 259 489
rect 206 409 217 443
rect 251 409 259 443
rect 206 367 259 409
rect 313 599 366 617
rect 313 565 321 599
rect 355 565 366 599
rect 313 529 366 565
rect 313 495 321 529
rect 355 495 366 529
rect 313 459 366 495
rect 313 425 321 459
rect 355 425 366 459
rect 313 365 366 425
rect 396 543 452 617
rect 396 509 407 543
rect 441 509 452 543
rect 396 475 452 509
rect 396 441 407 475
rect 441 441 452 475
rect 396 407 452 441
rect 396 373 407 407
rect 441 373 452 407
rect 396 365 452 373
rect 482 607 585 617
rect 482 573 518 607
rect 552 573 585 607
rect 482 509 585 573
rect 482 475 518 509
rect 552 475 585 509
rect 482 418 585 475
rect 482 384 518 418
rect 552 384 585 418
rect 482 365 585 384
rect 615 597 671 617
rect 615 563 626 597
rect 660 563 671 597
rect 615 490 671 563
rect 615 456 626 490
rect 660 456 671 490
rect 615 365 671 456
rect 701 531 754 617
rect 701 497 712 531
rect 746 497 754 531
rect 701 418 754 497
rect 701 384 712 418
rect 746 384 754 418
rect 701 365 754 384
rect 808 531 861 619
rect 808 497 816 531
rect 850 497 861 531
rect 808 418 861 497
rect 808 384 816 418
rect 850 384 861 418
rect 808 367 861 384
rect 891 597 947 619
rect 891 563 902 597
rect 936 563 947 597
rect 891 490 947 563
rect 891 456 902 490
rect 936 456 947 490
rect 891 367 947 456
rect 977 599 1033 619
rect 977 565 988 599
rect 1022 565 1033 599
rect 977 504 1033 565
rect 977 470 988 504
rect 1022 470 1033 504
rect 977 418 1033 470
rect 977 384 988 418
rect 1022 384 1033 418
rect 977 367 1033 384
rect 1063 607 1119 619
rect 1063 573 1074 607
rect 1108 573 1119 607
rect 1063 490 1119 573
rect 1063 456 1074 490
rect 1108 456 1119 490
rect 1063 367 1119 456
rect 1149 599 1202 619
rect 1149 565 1160 599
rect 1194 565 1202 599
rect 1149 504 1202 565
rect 1149 470 1160 504
rect 1194 470 1202 504
rect 1149 418 1202 470
rect 1149 384 1160 418
rect 1194 384 1202 418
rect 1149 367 1202 384
<< ndiffc >>
rect 163 135 197 169
rect 163 61 197 95
rect 249 135 283 169
rect 335 169 369 203
rect 335 67 369 101
rect 436 131 470 165
rect 436 55 470 89
rect 540 169 574 203
rect 540 67 574 101
rect 630 131 664 165
rect 630 55 664 89
rect 724 169 758 203
rect 724 67 758 101
rect 810 131 844 165
rect 810 55 844 89
rect 896 169 930 203
rect 896 67 930 101
rect 982 131 1016 165
rect 982 55 1016 89
rect 1072 169 1106 203
rect 1072 67 1106 101
<< pdiffc >>
rect 45 573 79 607
rect 45 471 79 505
rect 45 379 79 413
rect 131 565 165 599
rect 131 471 165 505
rect 131 379 165 413
rect 217 573 251 607
rect 217 489 251 523
rect 217 409 251 443
rect 321 565 355 599
rect 321 495 355 529
rect 321 425 355 459
rect 407 509 441 543
rect 407 441 441 475
rect 407 373 441 407
rect 518 573 552 607
rect 518 475 552 509
rect 518 384 552 418
rect 626 563 660 597
rect 626 456 660 490
rect 712 497 746 531
rect 712 384 746 418
rect 816 497 850 531
rect 816 384 850 418
rect 902 563 936 597
rect 902 456 936 490
rect 988 565 1022 599
rect 988 470 1022 504
rect 988 384 1022 418
rect 1074 573 1108 607
rect 1074 456 1108 490
rect 1160 565 1194 599
rect 1160 470 1194 504
rect 1160 384 1194 418
<< poly >>
rect 90 619 120 645
rect 176 619 206 645
rect 366 617 396 643
rect 452 617 482 643
rect 585 617 615 643
rect 671 617 701 643
rect 861 619 891 645
rect 947 619 977 645
rect 1033 619 1063 645
rect 1119 619 1149 645
rect 90 321 120 367
rect 176 321 206 367
rect 366 333 396 365
rect 452 333 482 365
rect 67 305 324 321
rect 67 271 83 305
rect 117 271 163 305
rect 197 271 324 305
rect 67 237 324 271
rect 366 317 543 333
rect 366 283 493 317
rect 527 283 543 317
rect 366 267 543 283
rect 585 331 615 365
rect 671 333 701 365
rect 861 345 891 367
rect 947 345 977 367
rect 661 331 727 333
rect 585 317 727 331
rect 585 283 677 317
rect 711 283 727 317
rect 585 267 727 283
rect 769 319 977 345
rect 769 285 811 319
rect 845 315 977 319
rect 1033 317 1063 367
rect 1119 317 1149 367
rect 845 285 885 315
rect 769 269 885 285
rect 67 203 83 237
rect 117 203 133 237
rect 208 215 238 237
rect 294 215 324 237
rect 380 215 410 267
rect 499 215 529 267
rect 585 215 615 267
rect 683 215 713 267
rect 769 215 799 269
rect 855 215 885 269
rect 1033 301 1223 317
rect 1033 267 1080 301
rect 1114 267 1173 301
rect 1207 267 1223 301
rect 941 237 1223 267
rect 941 215 971 237
rect 1027 215 1057 237
rect 67 187 133 203
rect 208 21 238 47
rect 294 21 324 47
rect 380 21 410 47
rect 499 21 529 47
rect 585 21 615 47
rect 683 21 713 47
rect 769 21 799 47
rect 855 21 885 47
rect 941 21 971 47
rect 1027 21 1057 47
<< polycont >>
rect 83 271 117 305
rect 163 271 197 305
rect 493 283 527 317
rect 677 283 711 317
rect 811 285 845 319
rect 83 203 117 237
rect 1080 267 1114 301
rect 1173 267 1207 301
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 29 607 89 649
rect 29 573 45 607
rect 79 573 89 607
rect 29 505 89 573
rect 29 471 45 505
rect 79 471 89 505
rect 29 413 89 471
rect 29 379 45 413
rect 79 379 89 413
rect 29 363 89 379
rect 123 599 167 615
rect 123 565 131 599
rect 165 565 167 599
rect 123 505 167 565
rect 123 471 131 505
rect 165 471 167 505
rect 123 413 167 471
rect 123 379 131 413
rect 165 379 167 413
rect 201 607 267 649
rect 201 573 217 607
rect 251 573 267 607
rect 201 523 267 573
rect 201 489 217 523
rect 251 489 267 523
rect 201 443 267 489
rect 201 409 217 443
rect 251 409 267 443
rect 305 607 568 615
rect 305 599 518 607
rect 305 565 321 599
rect 355 579 518 599
rect 355 565 357 579
rect 305 529 357 565
rect 502 573 518 579
rect 552 573 568 607
rect 305 495 321 529
rect 355 495 357 529
rect 305 459 357 495
rect 305 425 321 459
rect 355 425 357 459
rect 305 409 357 425
rect 391 509 407 543
rect 441 509 457 543
rect 391 475 457 509
rect 391 441 407 475
rect 441 441 457 475
rect 123 375 167 379
rect 391 407 457 441
rect 391 375 407 407
rect 123 373 407 375
rect 441 373 457 407
rect 502 509 568 573
rect 502 475 518 509
rect 552 475 568 509
rect 502 418 568 475
rect 610 597 952 615
rect 610 563 626 597
rect 660 581 902 597
rect 660 563 676 581
rect 610 490 676 563
rect 886 563 902 581
rect 936 563 952 597
rect 610 456 626 490
rect 660 456 676 490
rect 610 452 676 456
rect 710 531 762 547
rect 710 497 712 531
rect 746 497 762 531
rect 710 418 762 497
rect 502 384 518 418
rect 552 384 712 418
rect 746 384 762 418
rect 800 531 852 547
rect 800 497 816 531
rect 850 497 852 531
rect 800 418 852 497
rect 886 490 952 563
rect 886 456 902 490
rect 936 456 952 490
rect 886 452 952 456
rect 986 599 1024 615
rect 986 565 988 599
rect 1022 565 1024 599
rect 986 504 1024 565
rect 986 470 988 504
rect 1022 470 1024 504
rect 986 418 1024 470
rect 1058 607 1124 649
rect 1058 573 1074 607
rect 1108 573 1124 607
rect 1058 490 1124 573
rect 1058 456 1074 490
rect 1108 456 1124 490
rect 1058 452 1124 456
rect 1158 599 1210 615
rect 1158 565 1160 599
rect 1194 565 1210 599
rect 1158 504 1210 565
rect 1158 470 1160 504
rect 1194 470 1210 504
rect 1158 418 1210 470
rect 800 384 816 418
rect 850 384 988 418
rect 1022 384 1160 418
rect 1194 384 1210 418
rect 123 341 457 373
rect 31 271 83 305
rect 117 271 163 305
rect 197 271 213 305
rect 31 237 213 271
rect 31 203 83 237
rect 117 203 213 237
rect 247 267 457 341
rect 491 317 643 350
rect 491 283 493 317
rect 527 283 643 317
rect 491 267 643 283
rect 677 317 752 350
rect 711 283 752 317
rect 677 267 752 283
rect 786 319 1030 350
rect 786 285 811 319
rect 845 285 1030 319
rect 786 267 1030 285
rect 1064 301 1223 350
rect 1064 267 1080 301
rect 1114 267 1173 301
rect 1207 267 1223 301
rect 247 169 297 267
rect 147 135 163 169
rect 197 135 213 169
rect 147 95 213 135
rect 247 135 249 169
rect 283 135 297 169
rect 247 119 297 135
rect 331 203 1122 233
rect 331 169 335 203
rect 369 199 540 203
rect 369 169 385 199
rect 147 61 163 95
rect 197 85 213 95
rect 331 101 385 169
rect 524 169 540 199
rect 574 199 724 203
rect 574 169 580 199
rect 331 85 335 101
rect 197 67 335 85
rect 369 67 385 101
rect 197 61 385 67
rect 147 51 385 61
rect 420 131 436 165
rect 470 131 486 165
rect 420 89 486 131
rect 420 55 436 89
rect 470 55 486 89
rect 420 17 486 55
rect 524 101 580 169
rect 714 169 724 199
rect 758 199 896 203
rect 758 169 760 199
rect 524 67 540 101
rect 574 67 580 101
rect 524 51 580 67
rect 614 131 630 165
rect 664 131 680 165
rect 614 89 680 131
rect 614 55 630 89
rect 664 55 680 89
rect 614 17 680 55
rect 714 101 760 169
rect 894 169 896 199
rect 930 199 1072 203
rect 930 169 932 199
rect 714 67 724 101
rect 758 67 760 101
rect 714 51 760 67
rect 794 131 810 165
rect 844 131 860 165
rect 794 89 860 131
rect 794 55 810 89
rect 844 55 860 89
rect 794 17 860 55
rect 894 101 932 169
rect 1068 169 1072 199
rect 1106 169 1122 203
rect 894 67 896 101
rect 930 67 932 101
rect 894 51 932 67
rect 966 131 982 165
rect 1016 131 1032 165
rect 966 89 1032 131
rect 966 55 982 89
rect 1016 55 1032 89
rect 966 17 1032 55
rect 1068 101 1122 169
rect 1068 67 1072 101
rect 1106 67 1122 101
rect 1068 51 1122 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o41ai_2
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6594652
string GDS_START 6583510
<< end >>
