magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 122 210 666 248
rect 1 49 666 210
rect 0 0 672 49
<< scnmos >>
rect 84 74 114 184
rect 198 74 228 222
rect 284 74 314 222
rect 475 74 505 222
rect 553 74 583 222
<< scpmoshvt >>
rect 86 368 116 536
rect 210 368 240 592
rect 300 368 330 592
rect 466 378 496 578
rect 556 378 586 578
<< ndiff >>
rect 148 184 198 222
rect 27 146 84 184
rect 27 112 39 146
rect 73 112 84 146
rect 27 74 84 112
rect 114 144 198 184
rect 114 110 139 144
rect 173 110 198 144
rect 114 74 198 110
rect 228 210 284 222
rect 228 176 239 210
rect 273 176 284 210
rect 228 120 284 176
rect 228 86 239 120
rect 273 86 284 120
rect 228 74 284 86
rect 314 120 475 222
rect 314 86 339 120
rect 373 86 430 120
rect 464 86 475 120
rect 314 74 475 86
rect 505 74 553 222
rect 583 210 640 222
rect 583 176 594 210
rect 628 176 640 210
rect 583 120 640 176
rect 583 86 594 120
rect 628 86 640 120
rect 583 74 640 86
<< pdiff >>
rect 134 592 192 594
rect 134 582 210 592
rect 134 548 146 582
rect 180 548 210 582
rect 134 536 210 548
rect 27 524 86 536
rect 27 490 39 524
rect 73 490 86 524
rect 27 440 86 490
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 368 210 536
rect 240 414 300 592
rect 240 380 253 414
rect 287 380 300 414
rect 240 368 300 380
rect 330 578 448 592
rect 330 566 466 578
rect 330 532 372 566
rect 406 532 466 566
rect 330 378 466 532
rect 496 427 556 578
rect 496 393 509 427
rect 543 393 556 427
rect 496 378 556 393
rect 586 566 645 578
rect 586 532 599 566
rect 633 532 645 566
rect 586 378 645 532
rect 330 368 383 378
<< ndiffc >>
rect 39 112 73 146
rect 139 110 173 144
rect 239 176 273 210
rect 239 86 273 120
rect 339 86 373 120
rect 430 86 464 120
rect 594 176 628 210
rect 594 86 628 120
<< pdiffc >>
rect 146 548 180 582
rect 39 490 73 524
rect 39 406 73 440
rect 253 380 287 414
rect 372 532 406 566
rect 509 393 543 427
rect 599 532 633 566
<< poly >>
rect 210 592 240 618
rect 300 592 330 618
rect 86 536 116 562
rect 466 578 496 604
rect 556 578 586 604
rect 86 353 116 368
rect 210 353 240 368
rect 300 353 330 368
rect 466 363 496 378
rect 556 363 586 378
rect 83 336 119 353
rect 44 320 119 336
rect 44 286 60 320
rect 94 286 119 320
rect 207 326 243 353
rect 297 326 333 353
rect 207 310 357 326
rect 463 310 499 363
rect 553 326 589 363
rect 553 310 619 326
rect 207 290 307 310
rect 44 270 119 286
rect 198 276 307 290
rect 341 276 357 310
rect 84 184 114 270
rect 198 260 357 276
rect 439 294 505 310
rect 439 260 455 294
rect 489 260 505 294
rect 198 222 228 260
rect 284 222 314 260
rect 439 244 505 260
rect 475 222 505 244
rect 553 276 569 310
rect 603 276 619 310
rect 553 260 619 276
rect 553 222 583 260
rect 84 48 114 74
rect 198 48 228 74
rect 284 48 314 74
rect 475 48 505 74
rect 553 48 583 74
<< polycont >>
rect 60 286 94 320
rect 307 276 341 310
rect 455 260 489 294
rect 569 276 603 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 130 582 196 649
rect 130 548 146 582
rect 180 548 196 582
rect 23 524 89 540
rect 130 532 196 548
rect 327 566 452 649
rect 327 532 372 566
rect 406 532 452 566
rect 583 566 649 649
rect 583 532 599 566
rect 633 532 649 566
rect 23 490 39 524
rect 73 498 89 524
rect 73 490 627 498
rect 23 464 627 490
rect 23 440 178 464
rect 23 406 39 440
rect 73 406 178 440
rect 23 390 178 406
rect 25 320 110 356
rect 25 286 60 320
rect 94 286 110 320
rect 25 270 110 286
rect 144 236 178 390
rect 217 414 303 430
rect 217 380 253 414
rect 287 380 303 414
rect 217 364 303 380
rect 337 427 559 430
rect 337 393 509 427
rect 543 393 559 427
rect 337 374 559 393
rect 23 202 178 236
rect 223 226 257 364
rect 337 326 371 374
rect 593 326 627 464
rect 291 310 371 326
rect 553 310 627 326
rect 291 276 307 310
rect 341 276 371 310
rect 291 260 371 276
rect 223 210 289 226
rect 23 146 89 202
rect 223 176 239 210
rect 273 176 289 210
rect 23 112 39 146
rect 73 112 89 146
rect 23 70 89 112
rect 123 144 189 168
rect 123 110 139 144
rect 173 110 189 144
rect 123 17 189 110
rect 223 120 289 176
rect 337 202 371 260
rect 409 294 505 310
rect 409 260 455 294
rect 489 260 505 294
rect 553 276 569 310
rect 603 276 627 310
rect 553 260 627 276
rect 409 236 505 260
rect 578 210 644 226
rect 578 202 594 210
rect 337 176 594 202
rect 628 176 644 210
rect 337 168 644 176
rect 578 120 644 168
rect 223 86 239 120
rect 273 86 289 120
rect 223 70 289 86
rect 323 86 339 120
rect 373 86 430 120
rect 464 86 480 120
rect 323 17 480 86
rect 578 86 594 120
rect 628 86 644 120
rect 578 70 644 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and2b_2
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 3077010
string GDS_START 3071560
<< end >>
