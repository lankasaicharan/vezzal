magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 40 49 596 192
rect 0 0 672 49
<< scnmos >>
rect 135 82 165 166
rect 221 82 251 166
rect 307 82 337 166
rect 401 82 431 166
rect 487 82 517 166
<< scpmoshvt >>
rect 149 535 179 619
rect 221 535 251 619
rect 307 535 337 619
rect 401 535 431 619
rect 473 535 503 619
<< ndiff >>
rect 66 128 135 166
rect 66 94 74 128
rect 108 94 135 128
rect 66 82 135 94
rect 165 158 221 166
rect 165 124 176 158
rect 210 124 221 158
rect 165 82 221 124
rect 251 128 307 166
rect 251 94 262 128
rect 296 94 307 128
rect 251 82 307 94
rect 337 128 401 166
rect 337 94 352 128
rect 386 94 401 128
rect 337 82 401 94
rect 431 154 487 166
rect 431 120 442 154
rect 476 120 487 154
rect 431 82 487 120
rect 517 128 570 166
rect 517 94 528 128
rect 562 94 570 128
rect 517 82 570 94
<< pdiff >>
rect 49 607 149 619
rect 49 573 57 607
rect 91 573 149 607
rect 49 535 149 573
rect 179 535 221 619
rect 251 584 307 619
rect 251 550 262 584
rect 296 550 307 584
rect 251 535 307 550
rect 337 535 401 619
rect 431 535 473 619
rect 503 607 623 619
rect 503 573 581 607
rect 615 573 623 607
rect 503 535 623 573
<< ndiffc >>
rect 74 94 108 128
rect 176 124 210 158
rect 262 94 296 128
rect 352 94 386 128
rect 442 120 476 154
rect 528 94 562 128
<< pdiffc >>
rect 57 573 91 607
rect 262 550 296 584
rect 581 573 615 607
<< poly >>
rect 149 619 179 645
rect 221 619 251 645
rect 307 619 337 645
rect 401 619 431 645
rect 473 619 503 645
rect 149 478 179 535
rect 57 448 179 478
rect 57 322 87 448
rect 221 400 251 535
rect 21 306 87 322
rect 21 272 37 306
rect 71 272 87 306
rect 21 238 87 272
rect 185 384 251 400
rect 185 350 201 384
rect 235 350 251 384
rect 307 376 337 535
rect 401 400 431 535
rect 473 478 503 535
rect 473 448 592 478
rect 401 384 467 400
rect 185 316 251 350
rect 185 282 201 316
rect 235 282 251 316
rect 185 266 251 282
rect 21 204 37 238
rect 71 218 87 238
rect 71 204 165 218
rect 21 188 165 204
rect 135 166 165 188
rect 221 166 251 266
rect 293 360 359 376
rect 293 326 309 360
rect 343 326 359 360
rect 293 292 359 326
rect 293 258 309 292
rect 343 258 359 292
rect 293 242 359 258
rect 401 350 417 384
rect 451 350 467 384
rect 401 316 467 350
rect 401 282 417 316
rect 451 282 467 316
rect 401 266 467 282
rect 562 322 592 448
rect 562 306 628 322
rect 562 272 578 306
rect 612 272 628 306
rect 307 166 337 242
rect 401 166 431 266
rect 562 238 628 272
rect 562 218 578 238
rect 487 204 578 218
rect 612 204 628 238
rect 487 188 628 204
rect 487 166 517 188
rect 135 56 165 82
rect 221 56 251 82
rect 307 56 337 82
rect 401 56 431 82
rect 487 56 517 82
<< polycont >>
rect 37 272 71 306
rect 201 350 235 384
rect 201 282 235 316
rect 37 204 71 238
rect 309 326 343 360
rect 309 258 343 292
rect 417 350 451 384
rect 417 282 451 316
rect 578 272 612 306
rect 578 204 612 238
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 53 607 91 649
rect 53 573 57 607
rect 581 607 619 649
rect 53 557 91 573
rect 127 584 545 600
rect 127 550 262 584
rect 296 550 545 584
rect 615 573 619 607
rect 581 557 619 573
rect 127 534 545 550
rect 31 306 71 498
rect 31 272 37 306
rect 31 238 71 272
rect 31 204 37 238
rect 31 168 71 204
rect 131 202 165 534
rect 201 384 257 498
rect 235 350 257 384
rect 201 316 257 350
rect 235 282 257 316
rect 201 242 257 282
rect 309 360 353 498
rect 343 326 353 360
rect 309 292 353 326
rect 343 258 353 292
rect 309 242 353 258
rect 415 384 451 498
rect 415 350 417 384
rect 415 316 451 350
rect 415 282 417 316
rect 415 242 451 282
rect 578 306 641 498
rect 612 272 641 306
rect 578 238 641 272
rect 612 204 641 238
rect 131 168 226 202
rect 160 158 226 168
rect 58 128 124 132
rect 58 94 74 128
rect 108 94 124 128
rect 160 124 176 158
rect 210 124 226 158
rect 262 164 476 198
rect 578 168 641 204
rect 262 128 300 164
rect 438 154 476 164
rect 58 88 124 94
rect 296 94 300 128
rect 262 88 300 94
rect 58 54 300 88
rect 336 94 352 128
rect 386 94 402 128
rect 438 120 442 154
rect 438 104 476 120
rect 512 128 578 132
rect 336 17 402 94
rect 512 94 528 128
rect 562 94 578 128
rect 512 17 578 94
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o32ai_m
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2020070
string GDS_START 2011630
<< end >>
