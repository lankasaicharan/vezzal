magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 1 248 211 258
rect 1 49 1151 248
rect 0 0 1152 49
<< scpmos >>
rect 86 368 116 592
rect 186 368 216 592
rect 286 368 316 592
rect 434 368 464 592
rect 524 368 554 592
rect 634 368 664 592
rect 724 368 754 592
rect 834 368 864 592
rect 941 368 971 592
rect 1031 368 1061 592
<< nmoslvt >>
rect 98 84 128 232
rect 296 74 326 222
rect 382 74 412 222
rect 482 74 512 222
rect 568 74 598 222
rect 766 74 796 222
rect 852 74 882 222
rect 938 74 968 222
rect 1034 74 1064 222
<< ndiff >>
rect 27 220 98 232
rect 27 186 39 220
rect 73 186 98 220
rect 27 130 98 186
rect 27 96 39 130
rect 73 96 98 130
rect 27 84 98 96
rect 128 220 185 232
rect 128 186 139 220
rect 173 186 185 220
rect 128 130 185 186
rect 128 96 139 130
rect 173 96 185 130
rect 128 84 185 96
rect 239 152 296 222
rect 239 118 251 152
rect 285 118 296 152
rect 239 74 296 118
rect 326 169 382 222
rect 326 135 337 169
rect 371 135 382 169
rect 326 74 382 135
rect 412 184 482 222
rect 412 150 437 184
rect 471 150 482 184
rect 412 116 482 150
rect 412 82 437 116
rect 471 82 482 116
rect 412 74 482 82
rect 512 116 568 222
rect 512 82 523 116
rect 557 82 568 116
rect 512 74 568 82
rect 598 200 655 222
rect 598 166 609 200
rect 643 166 655 200
rect 598 74 655 166
rect 709 207 766 222
rect 709 173 721 207
rect 755 173 766 207
rect 709 74 766 173
rect 796 120 852 222
rect 796 86 807 120
rect 841 86 852 120
rect 796 74 852 86
rect 882 210 938 222
rect 882 176 893 210
rect 927 176 938 210
rect 882 120 938 176
rect 882 86 893 120
rect 927 86 938 120
rect 882 74 938 86
rect 968 152 1034 222
rect 968 118 979 152
rect 1013 118 1034 152
rect 968 74 1034 118
rect 1064 210 1125 222
rect 1064 176 1079 210
rect 1113 176 1125 210
rect 1064 120 1125 176
rect 1064 86 1079 120
rect 1113 86 1125 120
rect 1064 74 1125 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 504 86 546
rect 27 470 39 504
rect 73 470 86 504
rect 27 425 86 470
rect 27 391 39 425
rect 73 391 86 425
rect 27 368 86 391
rect 116 539 186 592
rect 116 505 139 539
rect 173 505 186 539
rect 116 440 186 505
rect 116 406 139 440
rect 173 406 186 440
rect 116 368 186 406
rect 216 580 286 592
rect 216 546 239 580
rect 273 546 286 580
rect 216 499 286 546
rect 216 465 239 499
rect 273 465 286 499
rect 216 368 286 465
rect 316 573 434 592
rect 316 539 358 573
rect 392 539 434 573
rect 316 368 434 539
rect 464 580 524 592
rect 464 546 477 580
rect 511 546 524 580
rect 464 497 524 546
rect 464 463 477 497
rect 511 463 524 497
rect 464 414 524 463
rect 464 380 477 414
rect 511 380 524 414
rect 464 368 524 380
rect 554 580 634 592
rect 554 546 577 580
rect 611 546 634 580
rect 554 499 634 546
rect 554 465 577 499
rect 611 465 634 499
rect 554 368 634 465
rect 664 580 724 592
rect 664 546 677 580
rect 711 546 724 580
rect 664 510 724 546
rect 664 476 677 510
rect 711 476 724 510
rect 664 440 724 476
rect 664 406 677 440
rect 711 406 724 440
rect 664 368 724 406
rect 754 580 834 592
rect 754 546 777 580
rect 811 546 834 580
rect 754 499 834 546
rect 754 465 777 499
rect 811 465 834 499
rect 754 368 834 465
rect 864 584 941 592
rect 864 550 880 584
rect 914 550 941 584
rect 864 505 941 550
rect 864 471 880 505
rect 914 471 941 505
rect 864 424 941 471
rect 864 390 880 424
rect 914 390 941 424
rect 864 368 941 390
rect 971 584 1031 592
rect 971 550 984 584
rect 1018 550 1031 584
rect 971 499 1031 550
rect 971 465 984 499
rect 1018 465 1031 499
rect 971 368 1031 465
rect 1061 584 1125 592
rect 1061 550 1076 584
rect 1110 550 1125 584
rect 1061 505 1125 550
rect 1061 471 1076 505
rect 1110 471 1125 505
rect 1061 424 1125 471
rect 1061 390 1076 424
rect 1110 390 1125 424
rect 1061 368 1125 390
<< ndiffc >>
rect 39 186 73 220
rect 39 96 73 130
rect 139 186 173 220
rect 139 96 173 130
rect 251 118 285 152
rect 337 135 371 169
rect 437 150 471 184
rect 437 82 471 116
rect 523 82 557 116
rect 609 166 643 200
rect 721 173 755 207
rect 807 86 841 120
rect 893 176 927 210
rect 893 86 927 120
rect 979 118 1013 152
rect 1079 176 1113 210
rect 1079 86 1113 120
<< pdiffc >>
rect 39 546 73 580
rect 39 470 73 504
rect 39 391 73 425
rect 139 505 173 539
rect 139 406 173 440
rect 239 546 273 580
rect 239 465 273 499
rect 358 539 392 573
rect 477 546 511 580
rect 477 463 511 497
rect 477 380 511 414
rect 577 546 611 580
rect 577 465 611 499
rect 677 546 711 580
rect 677 476 711 510
rect 677 406 711 440
rect 777 546 811 580
rect 777 465 811 499
rect 880 550 914 584
rect 880 471 914 505
rect 880 390 914 424
rect 984 550 1018 584
rect 984 465 1018 499
rect 1076 550 1110 584
rect 1076 471 1110 505
rect 1076 390 1110 424
<< poly >>
rect 86 592 116 618
rect 186 592 216 618
rect 286 592 316 618
rect 434 592 464 618
rect 524 592 554 618
rect 634 592 664 618
rect 724 592 754 618
rect 834 592 864 618
rect 941 592 971 618
rect 1031 592 1061 618
rect 86 353 116 368
rect 186 353 216 368
rect 286 353 316 368
rect 434 353 464 368
rect 524 353 554 368
rect 634 353 664 368
rect 724 353 754 368
rect 834 353 864 368
rect 941 353 971 368
rect 1031 353 1061 368
rect 83 336 119 353
rect 183 336 219 353
rect 83 320 219 336
rect 83 286 99 320
rect 133 286 167 320
rect 201 286 219 320
rect 83 270 219 286
rect 283 345 319 353
rect 431 345 467 353
rect 283 320 467 345
rect 283 286 299 320
rect 333 315 467 320
rect 521 326 557 353
rect 631 326 667 353
rect 333 286 412 315
rect 283 270 412 286
rect 98 232 128 270
rect 296 222 326 270
rect 382 222 412 270
rect 521 310 667 326
rect 521 276 549 310
rect 583 276 617 310
rect 651 276 667 310
rect 521 267 667 276
rect 721 300 757 353
rect 831 336 867 353
rect 938 336 974 353
rect 1028 336 1064 353
rect 816 320 882 336
rect 816 300 832 320
rect 721 286 832 300
rect 866 286 882 320
rect 721 270 882 286
rect 482 237 667 267
rect 482 222 512 237
rect 568 222 598 237
rect 766 222 796 270
rect 852 222 882 270
rect 938 320 1064 336
rect 938 286 1001 320
rect 1035 286 1064 320
rect 938 270 1064 286
rect 938 222 968 270
rect 1034 222 1064 270
rect 98 58 128 84
rect 296 48 326 74
rect 382 48 412 74
rect 482 48 512 74
rect 568 48 598 74
rect 766 48 796 74
rect 852 48 882 74
rect 938 48 968 74
rect 1034 48 1064 74
<< polycont >>
rect 99 286 133 320
rect 167 286 201 320
rect 299 286 333 320
rect 549 276 583 310
rect 617 276 651 310
rect 832 286 866 320
rect 1001 286 1035 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 581 289 615
rect 23 580 89 581
rect 23 546 39 580
rect 73 546 89 580
rect 223 580 289 581
rect 23 504 89 546
rect 23 470 39 504
rect 73 470 89 504
rect 23 425 89 470
rect 23 391 39 425
rect 73 391 89 425
rect 23 390 89 391
rect 123 539 189 547
rect 123 505 139 539
rect 173 505 189 539
rect 123 440 189 505
rect 223 546 239 580
rect 273 546 289 580
rect 223 499 289 546
rect 323 573 427 649
rect 323 539 358 573
rect 392 539 427 573
rect 323 530 427 539
rect 461 580 527 596
rect 461 546 477 580
rect 511 546 527 580
rect 223 465 239 499
rect 273 492 289 499
rect 461 497 527 546
rect 461 492 477 497
rect 273 465 477 492
rect 223 463 477 465
rect 511 463 527 497
rect 223 458 527 463
rect 561 580 627 649
rect 561 546 577 580
rect 611 546 627 580
rect 561 499 627 546
rect 561 465 577 499
rect 611 465 627 499
rect 561 458 627 465
rect 661 580 727 596
rect 661 546 677 580
rect 711 546 727 580
rect 661 510 727 546
rect 661 476 677 510
rect 711 476 727 510
rect 123 406 139 440
rect 173 424 189 440
rect 461 424 527 458
rect 661 440 727 476
rect 761 580 827 649
rect 761 546 777 580
rect 811 546 827 580
rect 761 499 827 546
rect 761 465 777 499
rect 811 465 827 499
rect 761 458 827 465
rect 861 584 934 600
rect 861 550 880 584
rect 914 550 934 584
rect 861 505 934 550
rect 861 471 880 505
rect 914 471 934 505
rect 661 424 677 440
rect 173 406 427 424
rect 123 390 427 406
rect 25 320 217 356
rect 25 286 99 320
rect 133 286 167 320
rect 201 286 217 320
rect 283 320 359 356
rect 283 286 299 320
rect 333 286 359 320
rect 393 330 427 390
rect 461 414 677 424
rect 461 380 477 414
rect 511 406 677 414
rect 711 424 727 440
rect 861 424 934 471
rect 968 584 1034 649
rect 968 550 984 584
rect 1018 550 1034 584
rect 968 499 1034 550
rect 968 465 984 499
rect 1018 465 1034 499
rect 968 458 1034 465
rect 1068 584 1129 600
rect 1068 550 1076 584
rect 1110 550 1129 584
rect 1068 505 1129 550
rect 1068 471 1076 505
rect 1110 471 1129 505
rect 1068 424 1129 471
rect 711 406 880 424
rect 511 390 880 406
rect 914 390 1076 424
rect 1110 390 1129 424
rect 511 380 527 390
rect 461 364 527 380
rect 25 270 217 286
rect 393 252 455 330
rect 601 326 743 356
rect 533 310 743 326
rect 533 276 549 310
rect 583 276 617 310
rect 651 276 743 310
rect 533 260 743 276
rect 793 320 935 356
rect 793 286 832 320
rect 866 286 935 320
rect 793 270 935 286
rect 985 320 1127 356
rect 985 286 1001 320
rect 1035 286 1127 320
rect 985 270 1127 286
rect 337 236 455 252
rect 23 220 89 236
rect 23 186 39 220
rect 73 186 89 220
rect 23 130 89 186
rect 23 96 39 130
rect 73 96 89 130
rect 23 17 89 96
rect 123 220 455 236
rect 893 226 1129 236
rect 123 186 139 220
rect 173 218 455 220
rect 173 202 387 218
rect 173 186 189 202
rect 123 130 189 186
rect 337 169 387 202
rect 593 200 659 216
rect 593 184 609 200
rect 123 96 139 130
rect 173 96 189 130
rect 123 80 189 96
rect 235 152 301 168
rect 235 118 251 152
rect 285 118 301 152
rect 371 135 387 169
rect 337 119 387 135
rect 421 150 437 184
rect 471 166 609 184
rect 643 166 659 200
rect 705 210 1129 226
rect 705 207 893 210
rect 705 173 721 207
rect 755 176 893 207
rect 927 202 1079 210
rect 755 173 927 176
rect 705 170 927 173
rect 471 150 659 166
rect 235 85 301 118
rect 421 116 471 150
rect 791 120 857 136
rect 791 116 807 120
rect 421 85 437 116
rect 235 82 437 85
rect 235 51 471 82
rect 507 82 523 116
rect 557 86 807 116
rect 841 86 857 120
rect 557 82 857 86
rect 507 66 857 82
rect 893 120 927 170
rect 1063 176 1079 202
rect 1113 176 1129 210
rect 893 70 927 86
rect 963 152 1029 168
rect 963 118 979 152
rect 1013 118 1029 152
rect 963 17 1029 118
rect 1063 120 1129 176
rect 1063 86 1079 120
rect 1113 86 1129 120
rect 1063 70 1129 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a41oi_2
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 582174
string GDS_START 572020
<< end >>
