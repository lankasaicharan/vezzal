magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3890 1975
<< nwell >>
rect -38 331 2630 704
<< pwell >>
rect 1 235 208 289
rect 887 269 1252 279
rect 887 235 1566 269
rect 2316 241 2590 273
rect 1 201 1566 235
rect 1830 201 2590 241
rect 1 49 2590 201
rect 0 0 2592 49
<< scnmos >>
rect 99 179 129 263
rect 305 125 335 209
rect 477 125 507 209
rect 563 125 593 209
rect 649 125 679 209
rect 721 125 751 209
rect 966 169 996 253
rect 1038 169 1068 253
rect 1143 125 1173 253
rect 1333 159 1363 243
rect 1438 115 1468 243
rect 1647 91 1677 175
rect 1719 91 1749 175
rect 1909 131 1939 215
rect 2014 47 2044 215
rect 2100 47 2130 215
rect 2205 131 2235 215
rect 2395 79 2425 247
rect 2481 79 2511 247
<< scpmoshvt >>
rect 99 395 129 523
rect 357 465 387 593
rect 491 535 521 619
rect 577 535 607 619
rect 671 535 701 619
rect 743 535 773 619
rect 930 535 960 619
rect 1153 535 1183 619
rect 1258 451 1288 619
rect 1330 451 1360 619
rect 1438 451 1468 535
rect 1533 451 1563 535
rect 1619 451 1649 535
rect 1901 367 1931 451
rect 2006 367 2036 619
rect 2092 367 2122 619
rect 2197 367 2227 495
rect 2395 367 2425 619
rect 2481 367 2511 619
<< ndiff >>
rect 27 238 99 263
rect 27 204 53 238
rect 87 204 99 238
rect 27 179 99 204
rect 129 245 182 263
rect 129 211 140 245
rect 174 211 182 245
rect 129 179 182 211
rect 913 228 966 253
rect 248 167 305 209
rect 248 133 260 167
rect 294 133 305 167
rect 248 125 305 133
rect 335 167 477 209
rect 335 133 362 167
rect 396 133 477 167
rect 335 125 477 133
rect 507 184 563 209
rect 507 150 518 184
rect 552 150 563 184
rect 507 125 563 150
rect 593 184 649 209
rect 593 150 604 184
rect 638 150 649 184
rect 593 125 649 150
rect 679 125 721 209
rect 751 175 823 209
rect 751 141 763 175
rect 797 141 823 175
rect 913 194 921 228
rect 955 194 966 228
rect 913 169 966 194
rect 996 169 1038 253
rect 1068 191 1143 253
rect 1068 169 1098 191
rect 1090 157 1098 169
rect 1132 157 1143 191
rect 751 125 823 141
rect 1090 125 1143 157
rect 1173 183 1226 253
rect 1173 149 1184 183
rect 1218 149 1226 183
rect 1280 218 1333 243
rect 1280 184 1288 218
rect 1322 184 1333 218
rect 1280 159 1333 184
rect 1363 231 1438 243
rect 1363 197 1383 231
rect 1417 197 1438 231
rect 1363 159 1438 197
rect 1173 125 1226 149
rect 1385 115 1438 159
rect 1468 115 1540 243
rect 2342 219 2395 247
rect 1856 190 1909 215
rect 1490 91 1540 115
rect 1594 150 1647 175
rect 1594 116 1602 150
rect 1636 116 1647 150
rect 1594 91 1647 116
rect 1677 91 1719 175
rect 1749 150 1802 175
rect 1749 116 1760 150
rect 1794 116 1802 150
rect 1856 156 1864 190
rect 1898 156 1909 190
rect 1856 131 1909 156
rect 1939 163 2014 215
rect 1939 131 1969 163
rect 1749 91 1802 116
rect 1961 129 1969 131
rect 2003 129 2014 163
rect 1961 93 2014 129
rect 1490 57 1498 91
rect 1532 57 1540 91
rect 1490 45 1540 57
rect 1961 59 1969 93
rect 2003 59 2014 93
rect 1961 47 2014 59
rect 2044 207 2100 215
rect 2044 173 2055 207
rect 2089 173 2100 207
rect 2044 101 2100 173
rect 2044 67 2055 101
rect 2089 67 2100 101
rect 2044 47 2100 67
rect 2130 203 2205 215
rect 2130 169 2160 203
rect 2194 169 2205 203
rect 2130 131 2205 169
rect 2235 190 2288 215
rect 2235 156 2246 190
rect 2280 156 2288 190
rect 2235 131 2288 156
rect 2342 185 2350 219
rect 2384 185 2395 219
rect 2130 93 2183 131
rect 2342 125 2395 185
rect 2130 59 2141 93
rect 2175 59 2183 93
rect 2342 91 2350 125
rect 2384 91 2395 125
rect 2342 79 2395 91
rect 2425 235 2481 247
rect 2425 201 2436 235
rect 2470 201 2481 235
rect 2425 125 2481 201
rect 2425 91 2436 125
rect 2470 91 2481 125
rect 2425 79 2481 91
rect 2511 235 2564 247
rect 2511 201 2522 235
rect 2556 201 2564 235
rect 2511 125 2564 201
rect 2511 91 2522 125
rect 2556 91 2564 125
rect 2511 79 2564 91
rect 2130 47 2183 59
<< pdiff >>
rect 437 593 491 619
rect 304 579 357 593
rect 304 545 312 579
rect 346 545 357 579
rect 46 499 99 523
rect 46 465 54 499
rect 88 465 99 499
rect 46 395 99 465
rect 129 508 182 523
rect 129 474 140 508
rect 174 474 182 508
rect 129 395 182 474
rect 304 511 357 545
rect 304 477 312 511
rect 346 477 357 511
rect 304 465 357 477
rect 387 581 491 593
rect 387 547 422 581
rect 456 547 491 581
rect 387 535 491 547
rect 521 589 577 619
rect 521 555 532 589
rect 566 555 577 589
rect 521 535 577 555
rect 607 593 671 619
rect 607 559 625 593
rect 659 559 671 593
rect 607 535 671 559
rect 701 535 743 619
rect 773 606 930 619
rect 773 572 784 606
rect 818 572 885 606
rect 919 572 930 606
rect 773 535 930 572
rect 960 594 1153 619
rect 960 560 971 594
rect 1005 560 1108 594
rect 1142 560 1153 594
rect 960 535 1153 560
rect 1183 582 1258 619
rect 1183 548 1213 582
rect 1247 548 1258 582
rect 1183 535 1258 548
rect 387 465 437 535
rect 1205 451 1258 535
rect 1288 451 1330 619
rect 1360 535 1415 619
rect 1953 607 2006 619
rect 1953 573 1961 607
rect 1995 573 2006 607
rect 1953 536 2006 573
rect 1360 531 1438 535
rect 1360 497 1373 531
rect 1407 497 1438 531
rect 1360 451 1438 497
rect 1468 451 1533 535
rect 1563 505 1619 535
rect 1563 471 1574 505
rect 1608 471 1619 505
rect 1563 451 1619 471
rect 1649 505 1702 535
rect 1649 471 1660 505
rect 1694 471 1702 505
rect 1953 502 1961 536
rect 1995 502 2006 536
rect 1649 451 1702 471
rect 1953 465 2006 502
rect 1953 451 1961 465
rect 1848 426 1901 451
rect 1848 392 1856 426
rect 1890 392 1901 426
rect 1848 367 1901 392
rect 1931 431 1961 451
rect 1995 431 2006 465
rect 1931 367 2006 431
rect 2036 599 2092 619
rect 2036 565 2047 599
rect 2081 565 2092 599
rect 2036 501 2092 565
rect 2036 467 2047 501
rect 2081 467 2092 501
rect 2036 420 2092 467
rect 2036 386 2047 420
rect 2081 386 2092 420
rect 2036 367 2092 386
rect 2122 607 2175 619
rect 2122 573 2133 607
rect 2167 573 2175 607
rect 2122 509 2175 573
rect 2342 607 2395 619
rect 2342 573 2350 607
rect 2384 573 2395 607
rect 2122 475 2133 509
rect 2167 495 2175 509
rect 2342 512 2395 573
rect 2167 475 2197 495
rect 2122 413 2197 475
rect 2122 379 2152 413
rect 2186 379 2197 413
rect 2122 367 2197 379
rect 2227 481 2280 495
rect 2227 447 2238 481
rect 2272 447 2280 481
rect 2227 413 2280 447
rect 2227 379 2238 413
rect 2272 379 2280 413
rect 2227 367 2280 379
rect 2342 478 2350 512
rect 2384 478 2395 512
rect 2342 419 2395 478
rect 2342 385 2350 419
rect 2384 385 2395 419
rect 2342 367 2395 385
rect 2425 599 2481 619
rect 2425 565 2436 599
rect 2470 565 2481 599
rect 2425 502 2481 565
rect 2425 468 2436 502
rect 2470 468 2481 502
rect 2425 409 2481 468
rect 2425 375 2436 409
rect 2470 375 2481 409
rect 2425 367 2481 375
rect 2511 607 2564 619
rect 2511 573 2522 607
rect 2556 573 2564 607
rect 2511 509 2564 573
rect 2511 475 2522 509
rect 2556 475 2564 509
rect 2511 413 2564 475
rect 2511 379 2522 413
rect 2556 379 2564 413
rect 2511 367 2564 379
<< ndiffc >>
rect 53 204 87 238
rect 140 211 174 245
rect 260 133 294 167
rect 362 133 396 167
rect 518 150 552 184
rect 604 150 638 184
rect 763 141 797 175
rect 921 194 955 228
rect 1098 157 1132 191
rect 1184 149 1218 183
rect 1288 184 1322 218
rect 1383 197 1417 231
rect 1602 116 1636 150
rect 1760 116 1794 150
rect 1864 156 1898 190
rect 1969 129 2003 163
rect 1498 57 1532 91
rect 1969 59 2003 93
rect 2055 173 2089 207
rect 2055 67 2089 101
rect 2160 169 2194 203
rect 2246 156 2280 190
rect 2350 185 2384 219
rect 2141 59 2175 93
rect 2350 91 2384 125
rect 2436 201 2470 235
rect 2436 91 2470 125
rect 2522 201 2556 235
rect 2522 91 2556 125
<< pdiffc >>
rect 312 545 346 579
rect 54 465 88 499
rect 140 474 174 508
rect 312 477 346 511
rect 422 547 456 581
rect 532 555 566 589
rect 625 559 659 593
rect 784 572 818 606
rect 885 572 919 606
rect 971 560 1005 594
rect 1108 560 1142 594
rect 1213 548 1247 582
rect 1961 573 1995 607
rect 1373 497 1407 531
rect 1574 471 1608 505
rect 1660 471 1694 505
rect 1961 502 1995 536
rect 1856 392 1890 426
rect 1961 431 1995 465
rect 2047 565 2081 599
rect 2047 467 2081 501
rect 2047 386 2081 420
rect 2133 573 2167 607
rect 2350 573 2384 607
rect 2133 475 2167 509
rect 2152 379 2186 413
rect 2238 447 2272 481
rect 2238 379 2272 413
rect 2350 478 2384 512
rect 2350 385 2384 419
rect 2436 565 2470 599
rect 2436 468 2470 502
rect 2436 375 2470 409
rect 2522 573 2556 607
rect 2522 475 2556 509
rect 2522 379 2556 413
<< poly >>
rect 177 615 387 645
rect 491 619 521 645
rect 577 619 607 645
rect 671 619 701 645
rect 743 619 773 645
rect 930 619 960 645
rect 1153 619 1183 645
rect 1258 619 1288 645
rect 1330 619 1360 645
rect 2006 619 2036 645
rect 2092 619 2122 645
rect 2395 619 2425 645
rect 2481 619 2511 645
rect 177 605 243 615
rect 177 571 193 605
rect 227 571 243 605
rect 357 593 387 615
rect 177 555 243 571
rect 99 523 129 549
rect 491 503 521 535
rect 469 487 535 503
rect 357 439 387 465
rect 469 453 485 487
rect 519 453 535 487
rect 469 437 535 453
rect 243 395 309 411
rect 577 395 607 535
rect 99 363 129 395
rect 243 375 259 395
rect 58 347 129 363
rect 58 313 74 347
rect 108 313 129 347
rect 58 297 129 313
rect 99 263 129 297
rect 197 361 259 375
rect 293 365 607 395
rect 671 437 701 535
rect 743 509 773 535
rect 743 487 885 509
rect 743 479 835 487
rect 819 453 835 479
rect 869 453 885 487
rect 819 437 885 453
rect 930 483 960 535
rect 1153 485 1183 535
rect 930 465 996 483
rect 671 421 745 437
rect 671 387 695 421
rect 729 387 745 421
rect 293 361 309 365
rect 197 345 309 361
rect 671 353 745 387
rect 99 153 129 179
rect 197 103 227 345
rect 671 333 695 353
rect 383 307 449 323
rect 649 319 695 333
rect 729 319 745 353
rect 819 343 849 437
rect 930 431 946 465
rect 980 431 996 465
rect 1139 455 1183 485
rect 1139 435 1169 455
rect 1438 535 1468 561
rect 1533 535 1563 561
rect 1619 535 1649 561
rect 1901 451 1931 477
rect 930 397 996 431
rect 930 363 946 397
rect 980 363 996 397
rect 649 313 745 319
rect 269 281 335 297
rect 269 247 285 281
rect 319 247 335 281
rect 383 273 399 307
rect 433 287 449 307
rect 563 303 745 313
rect 793 327 859 343
rect 433 273 507 287
rect 383 257 507 273
rect 269 231 335 247
rect 305 209 335 231
rect 477 209 507 257
rect 563 283 679 303
rect 793 293 809 327
rect 843 293 859 327
rect 930 321 996 363
rect 563 209 593 283
rect 793 261 859 293
rect 649 209 679 235
rect 721 231 859 261
rect 966 253 996 321
rect 1038 419 1169 435
rect 1038 385 1065 419
rect 1099 385 1169 419
rect 1258 407 1288 451
rect 1038 369 1169 385
rect 1216 391 1288 407
rect 1038 253 1068 369
rect 1216 357 1232 391
rect 1266 357 1288 391
rect 1216 341 1288 357
rect 1330 405 1360 451
rect 1330 389 1396 405
rect 1330 355 1346 389
rect 1380 355 1396 389
rect 1216 305 1246 341
rect 1143 275 1246 305
rect 1330 321 1396 355
rect 1330 287 1346 321
rect 1380 287 1396 321
rect 1143 253 1173 275
rect 1330 271 1396 287
rect 721 209 751 231
rect 966 143 996 169
rect 1038 143 1068 169
rect 1333 243 1363 271
rect 1438 243 1468 451
rect 1533 288 1563 451
rect 1619 419 1649 451
rect 1619 403 1685 419
rect 1619 369 1635 403
rect 1669 383 1685 403
rect 1669 369 1749 383
rect 1619 353 1749 369
rect 2197 495 2227 521
rect 1533 258 1677 288
rect 1605 247 1677 258
rect 1333 133 1363 159
rect 191 87 257 103
rect 305 99 335 125
rect 477 99 507 125
rect 563 99 593 125
rect 191 53 207 87
rect 241 53 257 87
rect 191 51 257 53
rect 649 51 679 125
rect 721 99 751 125
rect 1143 99 1173 125
rect 1605 213 1621 247
rect 1655 213 1677 247
rect 1605 197 1677 213
rect 1647 175 1677 197
rect 1719 175 1749 353
rect 1901 333 1931 367
rect 1865 317 1931 333
rect 1865 283 1881 317
rect 1915 297 1931 317
rect 2006 297 2036 367
rect 2092 297 2122 367
rect 2197 297 2227 367
rect 2395 335 2425 367
rect 2345 319 2425 335
rect 1915 283 2235 297
rect 1865 267 2235 283
rect 2345 285 2361 319
rect 2395 299 2425 319
rect 2481 299 2511 367
rect 2395 285 2511 299
rect 2345 269 2511 285
rect 1909 215 1939 267
rect 2014 215 2044 267
rect 2100 215 2130 267
rect 2205 215 2235 267
rect 2395 247 2425 269
rect 2481 247 2511 269
rect 1438 51 1468 115
rect 191 21 1468 51
rect 1909 105 1939 131
rect 1647 65 1677 91
rect 1719 65 1749 91
rect 2205 105 2235 131
rect 2395 53 2425 79
rect 2481 53 2511 79
rect 2014 21 2044 47
rect 2100 21 2130 47
<< polycont >>
rect 193 571 227 605
rect 485 453 519 487
rect 74 313 108 347
rect 259 361 293 395
rect 835 453 869 487
rect 695 387 729 421
rect 695 319 729 353
rect 946 431 980 465
rect 946 363 980 397
rect 285 247 319 281
rect 399 273 433 307
rect 809 293 843 327
rect 1065 385 1099 419
rect 1232 357 1266 391
rect 1346 355 1380 389
rect 1346 287 1380 321
rect 1635 369 1669 403
rect 207 53 241 87
rect 1621 213 1655 247
rect 1881 283 1915 317
rect 2361 285 2395 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 38 499 104 649
rect 144 605 243 615
rect 144 571 193 605
rect 227 571 243 605
rect 144 555 243 571
rect 296 579 349 595
rect 144 526 190 555
rect 38 465 54 499
rect 88 465 104 499
rect 38 458 104 465
rect 138 508 190 526
rect 138 474 140 508
rect 174 474 190 508
rect 296 545 312 579
rect 346 545 349 579
rect 296 511 349 545
rect 406 581 472 649
rect 406 547 422 581
rect 456 547 472 581
rect 406 537 472 547
rect 528 589 589 605
rect 528 555 532 589
rect 566 555 589 589
rect 528 539 589 555
rect 296 495 312 511
rect 138 458 190 474
rect 17 347 108 424
rect 17 313 74 347
rect 17 297 108 313
rect 144 297 190 458
rect 243 477 312 495
rect 346 477 349 511
rect 243 461 349 477
rect 383 487 519 503
rect 243 395 309 461
rect 243 361 259 395
rect 293 361 309 395
rect 383 453 485 487
rect 383 321 519 453
rect 383 307 449 321
rect 144 281 335 297
rect 144 261 285 281
rect 37 238 90 254
rect 37 204 53 238
rect 87 204 90 238
rect 37 17 90 204
rect 124 247 285 261
rect 319 247 335 281
rect 383 273 399 307
rect 433 273 449 307
rect 553 287 589 539
rect 124 245 335 247
rect 124 211 140 245
rect 174 239 335 245
rect 516 253 589 287
rect 623 593 675 609
rect 623 559 625 593
rect 659 559 675 593
rect 768 606 935 649
rect 768 572 784 606
rect 818 572 885 606
rect 919 572 935 606
rect 768 567 935 572
rect 969 594 1146 615
rect 623 507 675 559
rect 969 560 971 594
rect 1005 560 1108 594
rect 1142 560 1146 594
rect 969 544 1146 560
rect 1197 582 1253 649
rect 1197 548 1213 582
rect 1247 548 1253 582
rect 969 533 1029 544
rect 623 473 799 507
rect 174 211 482 239
rect 124 203 482 211
rect 191 167 310 169
rect 191 133 260 167
rect 294 133 310 167
rect 191 87 310 133
rect 191 53 207 87
rect 241 53 310 87
rect 191 51 310 53
rect 346 167 412 169
rect 346 133 362 167
rect 396 133 412 167
rect 346 17 412 133
rect 448 85 482 203
rect 516 184 563 253
rect 623 200 659 473
rect 516 150 518 184
rect 552 150 563 184
rect 516 134 563 150
rect 597 184 659 200
rect 597 150 604 184
rect 638 150 659 184
rect 597 134 659 150
rect 693 421 731 437
rect 693 387 695 421
rect 729 387 731 421
rect 693 353 731 387
rect 765 397 799 473
rect 835 499 1029 533
rect 1197 532 1253 548
rect 1287 581 1524 615
rect 835 487 869 499
rect 1287 498 1321 581
rect 835 437 869 453
rect 930 431 946 465
rect 980 431 1029 465
rect 930 397 1029 431
rect 765 363 946 397
rect 980 363 1029 397
rect 1063 441 1321 498
rect 1357 531 1450 547
rect 1357 497 1373 531
rect 1407 497 1450 531
rect 1357 481 1450 497
rect 1063 419 1101 441
rect 1063 385 1065 419
rect 1099 385 1101 419
rect 1063 369 1101 385
rect 1135 391 1282 407
rect 693 319 695 353
rect 729 319 731 353
rect 995 335 1029 363
rect 1135 357 1232 391
rect 1266 357 1282 391
rect 1135 341 1282 357
rect 1330 389 1382 405
rect 1330 355 1346 389
rect 1380 355 1382 389
rect 1135 335 1169 341
rect 693 259 731 319
rect 793 327 959 329
rect 793 293 809 327
rect 843 293 959 327
rect 995 301 1169 335
rect 1330 321 1382 355
rect 1330 305 1346 321
rect 693 225 885 259
rect 693 85 729 225
rect 448 51 729 85
rect 763 175 815 191
rect 797 141 815 175
rect 763 17 815 141
rect 851 144 885 225
rect 919 228 959 293
rect 1205 287 1346 305
rect 1380 287 1382 321
rect 1205 271 1382 287
rect 1416 317 1450 481
rect 1486 419 1524 581
rect 1558 505 1617 649
rect 1945 607 2011 649
rect 1945 573 1961 607
rect 1995 573 2011 607
rect 1945 536 2011 573
rect 1558 471 1574 505
rect 1608 471 1617 505
rect 1558 455 1617 471
rect 1651 505 1739 521
rect 1651 471 1660 505
rect 1694 471 1739 505
rect 1651 455 1739 471
rect 1486 403 1669 419
rect 1486 369 1635 403
rect 1486 353 1669 369
rect 1705 329 1739 455
rect 1945 502 1961 536
rect 1995 502 2011 536
rect 1945 465 2011 502
rect 1840 426 1906 442
rect 1945 431 1961 465
rect 1995 431 2011 465
rect 2045 599 2093 615
rect 2045 565 2047 599
rect 2081 565 2093 599
rect 2045 501 2093 565
rect 2045 467 2047 501
rect 2081 467 2093 501
rect 1840 392 1856 426
rect 1890 397 1906 426
rect 2045 420 2093 467
rect 1890 392 2001 397
rect 1840 363 2001 392
rect 1705 317 1931 329
rect 1416 283 1881 317
rect 1915 283 1931 317
rect 1416 281 1931 283
rect 1205 267 1239 271
rect 919 194 921 228
rect 955 194 959 228
rect 919 178 959 194
rect 995 233 1239 267
rect 1416 235 1450 281
rect 1967 247 2001 363
rect 995 144 1029 233
rect 1273 218 1333 234
rect 851 103 1029 144
rect 1082 191 1148 199
rect 1082 157 1098 191
rect 1132 157 1148 191
rect 1082 17 1148 157
rect 1182 183 1234 199
rect 1182 149 1184 183
rect 1218 149 1234 183
rect 1182 93 1234 149
rect 1273 184 1288 218
rect 1322 184 1333 218
rect 1367 231 1450 235
rect 1367 197 1383 231
rect 1417 197 1450 231
rect 1605 213 1621 247
rect 1655 213 2001 247
rect 2045 386 2047 420
rect 2081 386 2093 420
rect 1605 197 1914 213
rect 1367 195 1450 197
rect 1273 161 1333 184
rect 1848 190 1914 197
rect 1273 150 1652 161
rect 1273 127 1602 150
rect 1586 116 1602 127
rect 1636 116 1652 150
rect 1586 100 1652 116
rect 1744 150 1810 163
rect 1744 116 1760 150
rect 1794 116 1810 150
rect 1848 156 1864 190
rect 1898 156 1914 190
rect 2045 207 2093 386
rect 2129 607 2196 649
rect 2129 573 2133 607
rect 2167 573 2196 607
rect 2129 509 2196 573
rect 2129 475 2133 509
rect 2167 475 2196 509
rect 2334 607 2395 649
rect 2334 573 2350 607
rect 2384 573 2395 607
rect 2334 512 2395 573
rect 2129 413 2196 475
rect 2129 379 2152 413
rect 2186 379 2196 413
rect 2129 363 2196 379
rect 2230 481 2293 497
rect 2230 447 2238 481
rect 2272 447 2293 481
rect 2230 413 2293 447
rect 2230 379 2238 413
rect 2272 379 2293 413
rect 2230 335 2293 379
rect 2334 478 2350 512
rect 2384 478 2395 512
rect 2334 419 2395 478
rect 2334 385 2350 419
rect 2384 385 2395 419
rect 2334 369 2395 385
rect 2429 599 2478 615
rect 2429 565 2436 599
rect 2470 565 2478 599
rect 2429 502 2478 565
rect 2429 468 2436 502
rect 2470 468 2478 502
rect 2429 409 2478 468
rect 2429 375 2436 409
rect 2470 375 2478 409
rect 2230 319 2395 335
rect 2230 285 2361 319
rect 2230 269 2395 285
rect 1848 140 1914 156
rect 1953 163 2011 179
rect 1182 91 1548 93
rect 1182 57 1498 91
rect 1532 57 1548 91
rect 1182 53 1548 57
rect 1744 17 1810 116
rect 1953 129 1969 163
rect 2003 129 2011 163
rect 1953 93 2011 129
rect 1953 59 1969 93
rect 2003 59 2011 93
rect 1953 17 2011 59
rect 2045 173 2055 207
rect 2089 173 2093 207
rect 2045 101 2093 173
rect 2045 67 2055 101
rect 2089 67 2093 101
rect 2045 51 2093 67
rect 2127 203 2196 219
rect 2127 169 2160 203
rect 2194 169 2196 203
rect 2127 93 2196 169
rect 2230 190 2296 269
rect 2429 235 2478 375
rect 2512 607 2572 649
rect 2512 573 2522 607
rect 2556 573 2572 607
rect 2512 509 2572 573
rect 2512 475 2522 509
rect 2556 475 2572 509
rect 2512 413 2572 475
rect 2512 379 2522 413
rect 2556 379 2572 413
rect 2512 363 2572 379
rect 2230 156 2246 190
rect 2280 156 2296 190
rect 2230 140 2296 156
rect 2334 219 2395 235
rect 2334 185 2350 219
rect 2384 185 2395 219
rect 2127 59 2141 93
rect 2175 59 2196 93
rect 2127 17 2196 59
rect 2334 125 2395 185
rect 2334 91 2350 125
rect 2384 91 2395 125
rect 2334 17 2395 91
rect 2429 201 2436 235
rect 2470 201 2478 235
rect 2429 125 2478 201
rect 2429 91 2436 125
rect 2470 91 2478 125
rect 2429 75 2478 91
rect 2512 235 2572 251
rect 2512 201 2522 235
rect 2556 201 2572 235
rect 2512 125 2572 201
rect 2512 91 2522 125
rect 2556 91 2572 125
rect 2512 17 2572 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
flabel pwell s 0 0 2592 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2592 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfsbp_2
flabel comment s 210 224 210 224 0 FreeSans 200 90 0 0 no_jumper_check
flabel comment s 830 368 830 368 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 2592 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2592 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 2431 242 2465 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1087 464 1121 498 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2047 94 2081 128 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2047 168 2081 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2047 464 2081 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2047 538 2081 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2592 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2363656
string GDS_START 2344784
<< end >>
