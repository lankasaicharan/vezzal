magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 332 1382 704
<< pwell >>
rect 213 248 681 252
rect 213 228 1343 248
rect 1 49 1343 228
rect 0 0 1344 49
<< scpmos >>
rect 158 368 188 568
rect 268 368 298 568
rect 358 368 388 568
rect 468 368 498 568
rect 558 368 588 568
rect 680 368 710 568
rect 770 368 800 568
rect 887 368 917 592
rect 977 368 1007 592
rect 1087 368 1117 592
rect 1177 368 1207 592
<< nmoslvt >>
rect 84 74 114 202
rect 296 98 326 226
rect 382 98 412 226
rect 468 98 498 226
rect 568 98 598 226
rect 766 94 796 222
rect 852 94 882 222
rect 954 74 984 222
rect 1054 74 1084 222
rect 1144 74 1174 222
rect 1230 74 1260 222
<< ndiff >>
rect 239 214 296 226
rect 27 194 84 202
rect 27 160 39 194
rect 73 160 84 194
rect 27 116 84 160
rect 27 82 39 116
rect 73 82 84 116
rect 27 74 84 82
rect 114 186 173 202
rect 114 152 125 186
rect 159 152 173 186
rect 114 116 173 152
rect 114 82 125 116
rect 159 82 173 116
rect 239 180 251 214
rect 285 180 296 214
rect 239 144 296 180
rect 239 110 251 144
rect 285 110 296 144
rect 239 98 296 110
rect 326 191 382 226
rect 326 157 337 191
rect 371 157 382 191
rect 326 98 382 157
rect 412 214 468 226
rect 412 180 423 214
rect 457 180 468 214
rect 412 144 468 180
rect 412 110 423 144
rect 457 110 468 144
rect 412 98 468 110
rect 498 213 568 226
rect 498 179 523 213
rect 557 179 568 213
rect 498 98 568 179
rect 598 144 655 226
rect 598 110 609 144
rect 643 110 655 144
rect 598 98 655 110
rect 709 152 766 222
rect 709 118 721 152
rect 755 118 766 152
rect 114 74 173 82
rect 709 94 766 118
rect 796 210 852 222
rect 796 176 807 210
rect 841 176 852 210
rect 796 140 852 176
rect 796 106 807 140
rect 841 106 852 140
rect 796 94 852 106
rect 882 210 954 222
rect 882 176 909 210
rect 943 176 954 210
rect 882 120 954 176
rect 882 94 909 120
rect 897 86 909 94
rect 943 86 954 120
rect 897 74 954 86
rect 984 210 1054 222
rect 984 176 1009 210
rect 1043 176 1054 210
rect 984 120 1054 176
rect 984 86 1009 120
rect 1043 86 1054 120
rect 984 74 1054 86
rect 1084 142 1144 222
rect 1084 108 1095 142
rect 1129 108 1144 142
rect 1084 74 1144 108
rect 1174 210 1230 222
rect 1174 176 1185 210
rect 1219 176 1230 210
rect 1174 120 1230 176
rect 1174 86 1185 120
rect 1219 86 1230 120
rect 1174 74 1230 86
rect 1260 210 1317 222
rect 1260 176 1271 210
rect 1305 176 1317 210
rect 1260 120 1317 176
rect 1260 86 1271 120
rect 1305 86 1317 120
rect 1260 74 1317 86
<< pdiff >>
rect 818 580 887 592
rect 818 568 830 580
rect 99 556 158 568
rect 99 522 111 556
rect 145 522 158 556
rect 99 485 158 522
rect 99 451 111 485
rect 145 451 158 485
rect 99 414 158 451
rect 99 380 111 414
rect 145 380 158 414
rect 99 368 158 380
rect 188 556 268 568
rect 188 522 211 556
rect 245 522 268 556
rect 188 447 268 522
rect 188 413 211 447
rect 245 413 268 447
rect 188 368 268 413
rect 298 556 358 568
rect 298 522 311 556
rect 345 522 358 556
rect 298 485 358 522
rect 298 451 311 485
rect 345 451 358 485
rect 298 414 358 451
rect 298 380 311 414
rect 345 380 358 414
rect 298 368 358 380
rect 388 560 468 568
rect 388 526 411 560
rect 445 526 468 560
rect 388 492 468 526
rect 388 458 411 492
rect 445 458 468 492
rect 388 368 468 458
rect 498 560 558 568
rect 498 526 511 560
rect 545 526 558 560
rect 498 492 558 526
rect 498 458 511 492
rect 545 458 558 492
rect 498 424 558 458
rect 498 390 511 424
rect 545 390 558 424
rect 498 368 558 390
rect 588 560 680 568
rect 588 526 611 560
rect 645 526 680 560
rect 588 492 680 526
rect 588 458 611 492
rect 645 458 680 492
rect 588 368 680 458
rect 710 560 770 568
rect 710 526 723 560
rect 757 526 770 560
rect 710 492 770 526
rect 710 458 723 492
rect 757 458 770 492
rect 710 424 770 458
rect 710 390 723 424
rect 757 390 770 424
rect 710 368 770 390
rect 800 546 830 568
rect 864 546 887 580
rect 800 497 887 546
rect 800 463 830 497
rect 864 463 887 497
rect 800 414 887 463
rect 800 380 830 414
rect 864 380 887 414
rect 800 368 887 380
rect 917 580 977 592
rect 917 546 930 580
rect 964 546 977 580
rect 917 497 977 546
rect 917 463 930 497
rect 964 463 977 497
rect 917 414 977 463
rect 917 380 930 414
rect 964 380 977 414
rect 917 368 977 380
rect 1007 580 1087 592
rect 1007 546 1030 580
rect 1064 546 1087 580
rect 1007 467 1087 546
rect 1007 433 1030 467
rect 1064 433 1087 467
rect 1007 368 1087 433
rect 1117 580 1177 592
rect 1117 546 1130 580
rect 1164 546 1177 580
rect 1117 497 1177 546
rect 1117 463 1130 497
rect 1164 463 1177 497
rect 1117 414 1177 463
rect 1117 380 1130 414
rect 1164 380 1177 414
rect 1117 368 1177 380
rect 1207 580 1276 592
rect 1207 546 1230 580
rect 1264 546 1276 580
rect 1207 467 1276 546
rect 1207 433 1230 467
rect 1264 433 1276 467
rect 1207 368 1276 433
<< ndiffc >>
rect 39 160 73 194
rect 39 82 73 116
rect 125 152 159 186
rect 125 82 159 116
rect 251 180 285 214
rect 251 110 285 144
rect 337 157 371 191
rect 423 180 457 214
rect 423 110 457 144
rect 523 179 557 213
rect 609 110 643 144
rect 721 118 755 152
rect 807 176 841 210
rect 807 106 841 140
rect 909 176 943 210
rect 909 86 943 120
rect 1009 176 1043 210
rect 1009 86 1043 120
rect 1095 108 1129 142
rect 1185 176 1219 210
rect 1185 86 1219 120
rect 1271 176 1305 210
rect 1271 86 1305 120
<< pdiffc >>
rect 111 522 145 556
rect 111 451 145 485
rect 111 380 145 414
rect 211 522 245 556
rect 211 413 245 447
rect 311 522 345 556
rect 311 451 345 485
rect 311 380 345 414
rect 411 526 445 560
rect 411 458 445 492
rect 511 526 545 560
rect 511 458 545 492
rect 511 390 545 424
rect 611 526 645 560
rect 611 458 645 492
rect 723 526 757 560
rect 723 458 757 492
rect 723 390 757 424
rect 830 546 864 580
rect 830 463 864 497
rect 830 380 864 414
rect 930 546 964 580
rect 930 463 964 497
rect 930 380 964 414
rect 1030 546 1064 580
rect 1030 433 1064 467
rect 1130 546 1164 580
rect 1130 463 1164 497
rect 1130 380 1164 414
rect 1230 546 1264 580
rect 1230 433 1264 467
<< poly >>
rect 158 568 188 594
rect 268 568 298 594
rect 358 568 388 594
rect 468 568 498 594
rect 558 568 588 594
rect 680 568 710 594
rect 770 568 800 594
rect 887 592 917 618
rect 977 592 1007 618
rect 1087 592 1117 618
rect 1177 592 1207 618
rect 158 353 188 368
rect 268 353 298 368
rect 358 353 388 368
rect 468 353 498 368
rect 558 353 588 368
rect 680 353 710 368
rect 770 353 800 368
rect 887 353 917 368
rect 977 353 1007 368
rect 1087 353 1117 368
rect 1177 353 1207 368
rect 155 302 191 353
rect 265 330 301 353
rect 355 330 391 353
rect 239 314 391 330
rect 84 286 185 302
rect 84 252 117 286
rect 151 252 185 286
rect 239 280 255 314
rect 289 294 391 314
rect 465 336 501 353
rect 555 336 591 353
rect 677 336 713 353
rect 767 336 803 353
rect 465 320 591 336
rect 289 280 412 294
rect 239 264 412 280
rect 465 286 481 320
rect 515 300 591 320
rect 646 320 803 336
rect 515 286 598 300
rect 465 270 598 286
rect 84 236 185 252
rect 84 202 114 236
rect 296 226 326 264
rect 382 226 412 264
rect 468 226 498 270
rect 568 226 598 270
rect 646 286 662 320
rect 696 286 803 320
rect 884 349 920 353
rect 974 349 1010 353
rect 1084 349 1120 353
rect 1174 349 1210 353
rect 884 319 1210 349
rect 646 271 803 286
rect 951 310 1210 319
rect 951 276 967 310
rect 1001 276 1035 310
rect 1069 276 1103 310
rect 1137 290 1210 310
rect 1137 276 1260 290
rect 646 241 882 271
rect 951 260 1260 276
rect 766 222 796 241
rect 852 222 882 241
rect 954 222 984 260
rect 1054 222 1084 260
rect 1144 222 1174 260
rect 1230 222 1260 260
rect 84 48 114 74
rect 296 72 326 98
rect 382 72 412 98
rect 468 72 498 98
rect 568 72 598 98
rect 766 68 796 94
rect 852 68 882 94
rect 954 48 984 74
rect 1054 48 1084 74
rect 1144 48 1174 74
rect 1230 48 1260 74
<< polycont >>
rect 117 252 151 286
rect 255 280 289 314
rect 481 286 515 320
rect 662 286 696 320
rect 967 276 1001 310
rect 1035 276 1069 310
rect 1103 276 1137 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 95 556 161 572
rect 95 522 111 556
rect 145 522 161 556
rect 95 485 161 522
rect 95 451 111 485
rect 145 451 161 485
rect 95 414 161 451
rect 95 380 111 414
rect 145 380 161 414
rect 195 556 261 649
rect 195 522 211 556
rect 245 522 261 556
rect 195 447 261 522
rect 195 413 211 447
rect 245 413 261 447
rect 195 404 261 413
rect 295 556 361 572
rect 295 522 311 556
rect 345 522 361 556
rect 295 485 361 522
rect 295 451 311 485
rect 345 451 361 485
rect 395 560 461 649
rect 395 526 411 560
rect 445 526 461 560
rect 395 492 461 526
rect 395 458 411 492
rect 445 458 461 492
rect 495 560 561 572
rect 495 526 511 560
rect 545 526 561 560
rect 495 492 561 526
rect 495 458 511 492
rect 545 458 561 492
rect 595 560 661 649
rect 814 580 880 649
rect 595 526 611 560
rect 645 526 661 560
rect 595 492 661 526
rect 595 458 611 492
rect 645 458 661 492
rect 707 560 780 572
rect 707 526 723 560
rect 757 526 780 560
rect 707 492 780 526
rect 707 458 723 492
rect 757 458 780 492
rect 295 424 361 451
rect 495 424 561 458
rect 707 424 780 458
rect 295 414 511 424
rect 95 370 161 380
rect 295 380 311 414
rect 345 390 511 414
rect 545 390 723 424
rect 757 390 780 424
rect 345 380 373 390
rect 23 336 261 370
rect 295 364 373 380
rect 23 202 57 336
rect 227 330 261 336
rect 227 314 305 330
rect 101 286 167 302
rect 101 252 117 286
rect 151 252 167 286
rect 227 280 255 314
rect 289 280 305 314
rect 227 264 305 280
rect 101 236 167 252
rect 339 230 373 364
rect 409 320 551 356
rect 409 286 481 320
rect 515 286 551 320
rect 409 270 551 286
rect 601 320 712 356
rect 601 286 662 320
rect 696 286 712 320
rect 746 326 780 390
rect 814 546 830 580
rect 864 546 880 580
rect 814 497 880 546
rect 814 463 830 497
rect 864 463 880 497
rect 814 414 880 463
rect 814 380 830 414
rect 864 380 880 414
rect 814 364 880 380
rect 914 580 980 596
rect 914 546 930 580
rect 964 546 980 580
rect 914 497 980 546
rect 914 463 930 497
rect 964 463 980 497
rect 914 414 980 463
rect 1014 580 1080 649
rect 1014 546 1030 580
rect 1064 546 1080 580
rect 1014 467 1080 546
rect 1014 433 1030 467
rect 1064 433 1080 467
rect 1014 428 1080 433
rect 1114 580 1180 596
rect 1114 546 1130 580
rect 1164 546 1180 580
rect 1114 497 1180 546
rect 1114 463 1130 497
rect 1164 463 1180 497
rect 914 380 930 414
rect 964 394 980 414
rect 1114 414 1180 463
rect 1214 580 1280 649
rect 1214 546 1230 580
rect 1264 546 1280 580
rect 1214 467 1280 546
rect 1214 433 1230 467
rect 1264 433 1280 467
rect 1214 428 1280 433
rect 1114 394 1130 414
rect 964 380 1130 394
rect 1164 394 1180 414
rect 1164 380 1319 394
rect 914 360 1319 380
rect 746 310 1153 326
rect 746 292 967 310
rect 601 270 712 286
rect 951 276 967 292
rect 1001 276 1035 310
rect 1069 276 1103 310
rect 1137 276 1153 310
rect 951 260 1153 276
rect 235 214 301 230
rect 23 194 89 202
rect 23 160 39 194
rect 73 160 89 194
rect 23 116 89 160
rect 23 82 39 116
rect 73 82 89 116
rect 23 70 89 82
rect 123 186 175 202
rect 123 152 125 186
rect 159 152 175 186
rect 123 116 175 152
rect 123 82 125 116
rect 159 82 175 116
rect 123 17 175 82
rect 235 180 251 214
rect 285 180 301 214
rect 235 144 301 180
rect 235 110 251 144
rect 285 110 301 144
rect 337 191 373 230
rect 371 157 373 191
rect 337 119 373 157
rect 407 214 473 230
rect 407 180 423 214
rect 457 180 473 214
rect 407 144 473 180
rect 507 213 857 236
rect 1187 226 1221 360
rect 1273 310 1319 360
rect 507 179 523 213
rect 557 210 857 213
rect 557 202 807 210
rect 557 179 573 202
rect 507 178 573 179
rect 841 176 857 210
rect 705 152 771 168
rect 235 85 301 110
rect 407 110 423 144
rect 457 110 609 144
rect 643 110 659 144
rect 407 94 659 110
rect 705 118 721 152
rect 755 118 771 152
rect 407 85 473 94
rect 235 51 473 85
rect 705 17 771 118
rect 807 140 857 176
rect 841 106 857 140
rect 807 90 857 106
rect 893 210 959 226
rect 893 176 909 210
rect 943 176 959 210
rect 893 120 959 176
rect 893 86 909 120
rect 943 86 959 120
rect 893 17 959 86
rect 993 210 1221 226
rect 993 176 1009 210
rect 1043 192 1185 210
rect 993 120 1043 176
rect 1219 176 1221 210
rect 993 86 1009 120
rect 993 70 1043 86
rect 1079 142 1145 158
rect 1079 108 1095 142
rect 1129 108 1145 142
rect 1079 17 1145 108
rect 1185 120 1221 176
rect 1219 86 1221 120
rect 1185 70 1221 86
rect 1255 210 1321 226
rect 1255 176 1271 210
rect 1305 176 1321 210
rect 1255 120 1321 176
rect 1255 86 1271 120
rect 1305 86 1321 120
rect 1255 17 1321 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and3b_4
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 3533766
string GDS_START 3523040
<< end >>
