magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 157 394 241
rect 1 49 757 157
rect 0 0 768 49
<< scnmos >>
rect 80 47 110 215
rect 207 131 237 215
rect 285 131 315 215
rect 476 47 506 131
rect 562 47 592 131
rect 648 47 678 131
<< scpmoshvt >>
rect 80 367 110 619
rect 256 492 286 576
rect 342 492 372 576
rect 476 492 506 576
rect 562 492 592 576
rect 640 492 670 576
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 101 80 169
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 131 207 215
rect 237 131 285 215
rect 315 190 368 215
rect 315 156 326 190
rect 360 156 368 190
rect 315 131 368 156
rect 110 129 163 131
rect 110 95 121 129
rect 155 95 163 129
rect 423 106 476 131
rect 110 47 163 95
rect 423 72 431 106
rect 465 72 476 106
rect 423 47 476 72
rect 506 106 562 131
rect 506 72 517 106
rect 551 72 562 106
rect 506 47 562 72
rect 592 106 648 131
rect 592 72 603 106
rect 637 72 648 106
rect 592 47 648 72
rect 678 106 731 131
rect 678 72 689 106
rect 723 72 731 106
rect 678 47 731 72
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 504 80 565
rect 27 470 35 504
rect 69 470 80 504
rect 27 413 80 470
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 607 163 619
rect 110 573 121 607
rect 155 576 163 607
rect 155 573 256 576
rect 110 551 256 573
rect 110 517 209 551
rect 243 517 256 551
rect 110 504 256 517
rect 110 470 121 504
rect 155 492 256 504
rect 286 551 342 576
rect 286 517 297 551
rect 331 517 342 551
rect 286 492 342 517
rect 372 568 476 576
rect 372 534 410 568
rect 444 534 476 568
rect 372 492 476 534
rect 506 568 562 576
rect 506 534 517 568
rect 551 534 562 568
rect 506 492 562 534
rect 592 492 640 576
rect 670 552 723 576
rect 670 518 681 552
rect 715 518 723 552
rect 670 492 723 518
rect 155 470 163 492
rect 110 413 163 470
rect 110 379 121 413
rect 155 379 163 413
rect 110 367 163 379
<< ndiffc >>
rect 35 169 69 203
rect 35 67 69 101
rect 326 156 360 190
rect 121 95 155 129
rect 431 72 465 106
rect 517 72 551 106
rect 603 72 637 106
rect 689 72 723 106
<< pdiffc >>
rect 35 565 69 599
rect 35 470 69 504
rect 35 379 69 413
rect 121 573 155 607
rect 209 517 243 551
rect 121 470 155 504
rect 297 517 331 551
rect 410 534 444 568
rect 517 534 551 568
rect 681 518 715 552
rect 121 379 155 413
<< poly >>
rect 80 619 110 645
rect 256 576 286 602
rect 342 576 372 602
rect 476 576 506 602
rect 562 576 592 602
rect 640 576 670 602
rect 256 449 286 492
rect 207 433 286 449
rect 342 440 372 492
rect 207 399 223 433
rect 257 399 286 433
rect 80 303 110 367
rect 207 365 286 399
rect 207 331 223 365
rect 257 331 286 365
rect 207 315 286 331
rect 334 424 400 440
rect 334 390 350 424
rect 384 390 400 424
rect 476 415 506 492
rect 334 374 400 390
rect 448 399 514 415
rect 80 287 159 303
rect 80 253 109 287
rect 143 253 159 287
rect 80 237 159 253
rect 80 215 110 237
rect 207 215 237 315
rect 334 267 364 374
rect 448 365 464 399
rect 498 365 514 399
rect 448 331 514 365
rect 448 297 464 331
rect 498 297 514 331
rect 448 281 514 297
rect 562 326 592 492
rect 640 440 670 492
rect 640 424 732 440
rect 640 390 656 424
rect 690 390 732 424
rect 640 374 732 390
rect 562 310 654 326
rect 285 237 364 267
rect 285 215 315 237
rect 476 131 506 281
rect 562 276 604 310
rect 638 276 654 310
rect 562 260 654 276
rect 562 131 592 260
rect 702 212 732 374
rect 648 182 732 212
rect 648 131 678 182
rect 207 105 237 131
rect 285 105 315 131
rect 80 21 110 47
rect 476 21 506 47
rect 562 21 592 47
rect 648 21 678 47
<< polycont >>
rect 223 399 257 433
rect 223 331 257 365
rect 350 390 384 424
rect 109 253 143 287
rect 464 365 498 399
rect 464 297 498 331
rect 656 390 690 424
rect 604 276 638 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 19 599 71 615
rect 19 565 35 599
rect 69 565 71 599
rect 19 504 71 565
rect 19 470 35 504
rect 69 470 71 504
rect 19 413 71 470
rect 19 379 35 413
rect 69 379 71 413
rect 19 203 71 379
rect 105 607 253 649
rect 105 573 121 607
rect 155 573 253 607
rect 105 551 253 573
rect 394 568 460 649
rect 105 517 209 551
rect 243 517 253 551
rect 105 504 253 517
rect 105 470 121 504
rect 155 501 253 504
rect 287 551 335 567
rect 287 517 297 551
rect 331 517 335 551
rect 394 534 410 568
rect 444 534 460 568
rect 394 530 460 534
rect 501 568 568 584
rect 501 534 517 568
rect 551 534 568 568
rect 501 530 568 534
rect 155 470 171 501
rect 287 496 335 517
rect 287 470 500 496
rect 105 413 171 470
rect 297 462 500 470
rect 105 379 121 413
rect 155 379 171 413
rect 105 363 171 379
rect 207 399 223 433
rect 257 399 276 433
rect 207 365 276 399
rect 207 331 223 365
rect 257 331 276 365
rect 310 424 400 428
rect 310 390 350 424
rect 384 390 400 424
rect 310 351 400 390
rect 448 399 500 462
rect 448 365 464 399
rect 498 365 500 399
rect 19 169 35 203
rect 69 169 71 203
rect 105 287 173 303
rect 105 253 109 287
rect 143 253 173 287
rect 105 206 173 253
rect 207 242 276 331
rect 448 331 500 365
rect 448 315 464 331
rect 310 297 464 315
rect 498 297 500 331
rect 310 281 500 297
rect 105 172 264 206
rect 19 101 71 169
rect 19 67 35 101
rect 69 67 71 101
rect 19 51 71 67
rect 105 129 175 138
rect 105 95 121 129
rect 155 95 175 129
rect 105 17 175 95
rect 209 106 264 172
rect 310 190 376 281
rect 534 245 568 530
rect 665 552 731 649
rect 665 518 681 552
rect 715 518 731 552
rect 665 502 731 518
rect 607 424 737 442
rect 607 390 656 424
rect 690 390 737 424
rect 607 384 737 390
rect 310 156 326 190
rect 360 156 376 190
rect 310 140 376 156
rect 435 211 568 245
rect 602 310 751 350
rect 602 276 604 310
rect 638 276 751 310
rect 602 222 751 276
rect 435 124 474 211
rect 415 106 474 124
rect 209 72 431 106
rect 465 72 474 106
rect 209 56 474 72
rect 508 143 739 177
rect 508 106 553 143
rect 508 72 517 106
rect 551 72 553 106
rect 508 56 553 72
rect 587 106 653 109
rect 587 72 603 106
rect 637 72 653 106
rect 587 17 653 72
rect 687 106 739 143
rect 687 72 689 106
rect 723 72 739 106
rect 687 56 739 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2bb2a_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3625414
string GDS_START 3617138
<< end >>
