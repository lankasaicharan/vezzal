magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 4370 1975
<< nwell >>
rect -38 343 3110 704
rect -38 332 1411 343
rect 1680 332 3110 343
rect 283 326 1411 332
<< pwell >>
rect 618 268 897 284
rect 1453 279 1638 301
rect 285 248 897 268
rect 1272 275 1638 279
rect 1272 274 1881 275
rect 1272 256 3071 274
rect 1157 248 3071 256
rect 285 228 3071 248
rect 1 49 3071 228
rect 0 0 3072 49
<< scnmos >>
rect 84 74 114 202
rect 170 74 200 202
rect 411 94 441 242
rect 506 114 536 242
rect 592 114 622 242
rect 694 130 724 258
rect 788 130 818 258
rect 990 74 1020 222
rect 1248 102 1278 230
rect 1348 125 1378 253
rect 1434 125 1464 253
rect 1532 147 1562 275
rect 1870 120 1900 248
rect 2070 100 2100 248
rect 2156 100 2186 248
rect 2266 100 2296 248
rect 2352 100 2382 248
rect 2566 120 2596 248
rect 2686 100 2716 248
rect 2772 100 2802 248
rect 2858 100 2888 248
rect 2944 100 2974 248
<< scpmoshvt >>
rect 86 392 116 592
rect 176 392 206 592
rect 397 362 427 586
rect 498 362 528 530
rect 589 362 619 530
rect 713 362 743 530
rect 803 362 833 530
rect 1128 368 1158 592
rect 1235 379 1265 547
rect 1354 379 1384 547
rect 1482 423 1512 591
rect 1672 423 1702 591
rect 1779 368 1809 568
rect 1951 368 1981 592
rect 2041 368 2071 592
rect 2165 368 2195 592
rect 2255 368 2285 592
rect 2540 368 2570 568
rect 2657 368 2687 592
rect 2747 368 2777 592
rect 2855 368 2885 592
rect 2947 368 2977 592
<< ndiff >>
rect 644 242 694 258
rect 27 190 84 202
rect 27 156 39 190
rect 73 156 84 190
rect 27 120 84 156
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 184 170 202
rect 114 150 125 184
rect 159 150 170 184
rect 114 116 170 150
rect 114 82 125 116
rect 159 82 170 116
rect 114 74 170 82
rect 200 188 257 202
rect 200 154 211 188
rect 245 154 257 188
rect 200 120 257 154
rect 200 86 211 120
rect 245 86 257 120
rect 200 74 257 86
rect 311 108 411 242
rect 311 74 324 108
rect 358 94 411 108
rect 441 196 506 242
rect 441 162 461 196
rect 495 162 506 196
rect 441 114 506 162
rect 536 234 592 242
rect 536 200 547 234
rect 581 200 592 234
rect 536 166 592 200
rect 536 132 547 166
rect 581 132 592 166
rect 536 114 592 132
rect 622 184 694 242
rect 622 150 633 184
rect 667 150 694 184
rect 622 130 694 150
rect 724 246 788 258
rect 724 212 743 246
rect 777 212 788 246
rect 724 176 788 212
rect 724 142 743 176
rect 777 142 788 176
rect 724 130 788 142
rect 818 244 871 258
rect 818 210 829 244
rect 863 210 871 244
rect 1479 253 1532 275
rect 1298 230 1348 253
rect 818 130 871 210
rect 622 114 679 130
rect 441 94 491 114
rect 358 74 371 94
rect 311 62 371 74
rect 925 91 990 222
rect 925 57 933 91
rect 967 74 990 91
rect 1020 184 1073 222
rect 1183 221 1248 230
rect 1020 150 1031 184
rect 1065 150 1073 184
rect 1020 148 1073 150
rect 1183 187 1195 221
rect 1229 187 1248 221
rect 1183 153 1248 187
rect 1020 116 1077 148
rect 1020 82 1031 116
rect 1065 82 1077 116
rect 1183 119 1191 153
rect 1225 119 1248 153
rect 1183 102 1248 119
rect 1278 153 1348 230
rect 1278 119 1291 153
rect 1325 125 1348 153
rect 1378 239 1434 253
rect 1378 205 1389 239
rect 1423 205 1434 239
rect 1378 125 1434 205
rect 1464 239 1532 253
rect 1464 205 1487 239
rect 1521 205 1532 239
rect 1464 147 1532 205
rect 1562 228 1612 275
rect 1797 248 1855 249
rect 1797 237 1870 248
rect 1562 147 1635 228
rect 1464 125 1514 147
rect 1325 119 1333 125
rect 1278 102 1333 119
rect 1020 74 1077 82
rect 967 57 975 74
rect 925 45 975 57
rect 1582 93 1635 147
rect 1797 203 1809 237
rect 1843 203 1870 237
rect 1797 120 1870 203
rect 1900 120 2070 248
rect 2001 100 2070 120
rect 2100 236 2156 248
rect 2100 202 2111 236
rect 2145 202 2156 236
rect 2100 100 2156 202
rect 2186 100 2266 248
rect 2296 236 2352 248
rect 2296 202 2307 236
rect 2341 202 2352 236
rect 2296 100 2352 202
rect 2382 100 2455 248
rect 2509 236 2566 248
rect 2509 202 2521 236
rect 2555 202 2566 236
rect 2509 120 2566 202
rect 2596 120 2686 248
rect 1577 85 1635 93
rect 1577 51 1589 85
rect 1623 51 1635 85
rect 1577 39 1635 51
rect 2001 84 2055 100
rect 2001 50 2013 84
rect 2047 50 2055 84
rect 2201 84 2251 100
rect 2001 38 2055 50
rect 2201 50 2209 84
rect 2243 50 2251 84
rect 2397 84 2455 100
rect 2611 100 2686 120
rect 2716 220 2772 248
rect 2716 186 2727 220
rect 2761 186 2772 220
rect 2716 146 2772 186
rect 2716 112 2727 146
rect 2761 112 2772 146
rect 2716 100 2772 112
rect 2802 157 2858 248
rect 2802 123 2813 157
rect 2847 123 2858 157
rect 2802 100 2858 123
rect 2888 236 2944 248
rect 2888 202 2899 236
rect 2933 202 2944 236
rect 2888 146 2944 202
rect 2888 112 2899 146
rect 2933 112 2944 146
rect 2888 100 2944 112
rect 2974 236 3045 248
rect 2974 202 2999 236
rect 3033 202 3045 236
rect 2974 146 3045 202
rect 2974 112 2999 146
rect 3033 112 3045 146
rect 2974 100 3045 112
rect 2201 38 2251 50
rect 2397 50 2409 84
rect 2443 50 2455 84
rect 2397 38 2455 50
rect 2611 84 2671 100
rect 2611 50 2624 84
rect 2658 50 2671 84
rect 2611 38 2671 50
<< pdiff >>
rect 319 628 379 639
rect 319 594 332 628
rect 366 594 379 628
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 512 86 546
rect 27 478 39 512
rect 73 478 86 512
rect 27 444 86 478
rect 27 410 39 444
rect 73 410 86 444
rect 27 392 86 410
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 512 176 546
rect 116 478 129 512
rect 163 478 176 512
rect 116 444 176 478
rect 116 410 129 444
rect 163 410 176 444
rect 116 392 176 410
rect 206 580 265 592
rect 206 546 219 580
rect 253 546 265 580
rect 206 512 265 546
rect 206 478 219 512
rect 253 478 265 512
rect 206 444 265 478
rect 206 410 219 444
rect 253 410 265 444
rect 206 392 265 410
rect 319 586 379 594
rect 319 362 397 586
rect 427 530 480 586
rect 637 576 695 588
rect 637 542 649 576
rect 683 542 695 576
rect 1827 624 1933 636
rect 637 530 695 542
rect 427 488 498 530
rect 427 454 451 488
rect 485 454 498 488
rect 427 408 498 454
rect 427 374 451 408
rect 485 374 498 408
rect 427 362 498 374
rect 528 408 589 530
rect 528 374 541 408
rect 575 374 589 408
rect 528 362 589 374
rect 619 362 713 530
rect 743 422 803 530
rect 743 388 756 422
rect 790 388 803 422
rect 743 362 803 388
rect 833 518 892 530
rect 833 484 846 518
rect 880 484 892 518
rect 833 437 892 484
rect 833 403 846 437
rect 880 403 892 437
rect 833 362 892 403
rect 1069 580 1128 592
rect 1069 546 1081 580
rect 1115 546 1128 580
rect 1069 494 1128 546
rect 1069 460 1081 494
rect 1115 460 1128 494
rect 1069 368 1128 460
rect 1158 580 1217 592
rect 1158 546 1171 580
rect 1205 547 1217 580
rect 1402 579 1482 591
rect 1402 547 1424 579
rect 1205 546 1235 547
rect 1158 512 1235 546
rect 1158 478 1171 512
rect 1205 478 1235 512
rect 1158 440 1235 478
rect 1158 406 1171 440
rect 1205 406 1235 440
rect 1158 379 1235 406
rect 1265 522 1354 547
rect 1265 488 1307 522
rect 1341 488 1354 522
rect 1265 379 1354 488
rect 1384 545 1424 547
rect 1458 545 1482 579
rect 1384 423 1482 545
rect 1512 547 1672 591
rect 1512 513 1625 547
rect 1659 513 1672 547
rect 1512 469 1672 513
rect 1512 435 1625 469
rect 1659 435 1672 469
rect 1512 423 1672 435
rect 1702 568 1755 591
rect 1827 590 1863 624
rect 1897 592 1933 624
rect 2089 625 2147 639
rect 2089 592 2101 625
rect 1897 590 1951 592
rect 1827 568 1951 590
rect 1702 423 1779 568
rect 1384 379 1437 423
rect 1720 417 1779 423
rect 1158 368 1211 379
rect 1720 383 1732 417
rect 1766 383 1779 417
rect 1720 368 1779 383
rect 1809 368 1951 568
rect 1981 420 2041 592
rect 1981 386 1994 420
rect 2028 386 2041 420
rect 1981 368 2041 386
rect 2071 591 2101 592
rect 2135 592 2147 625
rect 2303 624 2421 636
rect 2303 592 2345 624
rect 2135 591 2165 592
rect 2071 368 2165 591
rect 2195 420 2255 592
rect 2195 386 2208 420
rect 2242 386 2255 420
rect 2195 368 2255 386
rect 2285 590 2345 592
rect 2379 590 2421 624
rect 2285 368 2421 590
rect 2588 580 2657 592
rect 2588 568 2600 580
rect 2481 560 2540 568
rect 2481 526 2493 560
rect 2527 526 2540 560
rect 2481 492 2540 526
rect 2481 458 2493 492
rect 2527 458 2540 492
rect 2481 424 2540 458
rect 2481 390 2493 424
rect 2527 390 2540 424
rect 2481 368 2540 390
rect 2570 546 2600 568
rect 2634 546 2657 580
rect 2570 503 2657 546
rect 2570 469 2600 503
rect 2634 469 2657 503
rect 2570 424 2657 469
rect 2570 390 2600 424
rect 2634 390 2657 424
rect 2570 368 2657 390
rect 2687 580 2747 592
rect 2687 546 2700 580
rect 2734 546 2747 580
rect 2687 500 2747 546
rect 2687 466 2700 500
rect 2734 466 2747 500
rect 2687 420 2747 466
rect 2687 386 2700 420
rect 2734 386 2747 420
rect 2687 368 2747 386
rect 2777 580 2855 592
rect 2777 546 2800 580
rect 2834 546 2855 580
rect 2777 488 2855 546
rect 2777 454 2800 488
rect 2834 454 2855 488
rect 2777 368 2855 454
rect 2885 580 2947 592
rect 2885 546 2900 580
rect 2934 546 2947 580
rect 2885 500 2947 546
rect 2885 466 2900 500
rect 2934 466 2947 500
rect 2885 420 2947 466
rect 2885 386 2900 420
rect 2934 386 2947 420
rect 2885 368 2947 386
rect 2977 580 3036 592
rect 2977 546 2990 580
rect 3024 546 3036 580
rect 2977 497 3036 546
rect 2977 463 2990 497
rect 3024 463 3036 497
rect 2977 414 3036 463
rect 2977 380 2990 414
rect 3024 380 3036 414
rect 2977 368 3036 380
<< ndiffc >>
rect 39 156 73 190
rect 39 86 73 120
rect 125 150 159 184
rect 125 82 159 116
rect 211 154 245 188
rect 211 86 245 120
rect 324 74 358 108
rect 461 162 495 196
rect 547 200 581 234
rect 547 132 581 166
rect 633 150 667 184
rect 743 212 777 246
rect 743 142 777 176
rect 829 210 863 244
rect 933 57 967 91
rect 1031 150 1065 184
rect 1195 187 1229 221
rect 1031 82 1065 116
rect 1191 119 1225 153
rect 1291 119 1325 153
rect 1389 205 1423 239
rect 1487 205 1521 239
rect 1809 203 1843 237
rect 2111 202 2145 236
rect 2307 202 2341 236
rect 2521 202 2555 236
rect 1589 51 1623 85
rect 2013 50 2047 84
rect 2209 50 2243 84
rect 2727 186 2761 220
rect 2727 112 2761 146
rect 2813 123 2847 157
rect 2899 202 2933 236
rect 2899 112 2933 146
rect 2999 202 3033 236
rect 2999 112 3033 146
rect 2409 50 2443 84
rect 2624 50 2658 84
<< pdiffc >>
rect 332 594 366 628
rect 39 546 73 580
rect 39 478 73 512
rect 39 410 73 444
rect 129 546 163 580
rect 129 478 163 512
rect 129 410 163 444
rect 219 546 253 580
rect 219 478 253 512
rect 219 410 253 444
rect 649 542 683 576
rect 451 454 485 488
rect 451 374 485 408
rect 541 374 575 408
rect 756 388 790 422
rect 846 484 880 518
rect 846 403 880 437
rect 1081 546 1115 580
rect 1081 460 1115 494
rect 1171 546 1205 580
rect 1171 478 1205 512
rect 1171 406 1205 440
rect 1307 488 1341 522
rect 1424 545 1458 579
rect 1625 513 1659 547
rect 1625 435 1659 469
rect 1863 590 1897 624
rect 1732 383 1766 417
rect 1994 386 2028 420
rect 2101 591 2135 625
rect 2208 386 2242 420
rect 2345 590 2379 624
rect 2493 526 2527 560
rect 2493 458 2527 492
rect 2493 390 2527 424
rect 2600 546 2634 580
rect 2600 469 2634 503
rect 2600 390 2634 424
rect 2700 546 2734 580
rect 2700 466 2734 500
rect 2700 386 2734 420
rect 2800 546 2834 580
rect 2800 454 2834 488
rect 2900 546 2934 580
rect 2900 466 2934 500
rect 2900 386 2934 420
rect 2990 546 3024 580
rect 2990 463 3024 497
rect 2990 380 3024 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 397 586 427 612
rect 495 604 957 634
rect 86 377 116 392
rect 176 377 206 392
rect 83 360 119 377
rect 173 360 209 377
rect 495 545 531 604
rect 498 530 528 545
rect 589 530 619 556
rect 710 545 746 604
rect 927 582 957 604
rect 1128 592 1158 618
rect 1232 615 1515 645
rect 927 566 1020 582
rect 713 530 743 545
rect 803 530 833 556
rect 927 532 943 566
rect 977 532 1020 566
rect 927 498 1020 532
rect 927 464 943 498
rect 977 464 1020 498
rect 927 430 1020 464
rect 927 396 943 430
rect 977 396 1020 430
rect 927 362 1020 396
rect 1232 562 1268 615
rect 1479 606 1515 615
rect 1482 591 1512 606
rect 1672 591 1702 617
rect 1235 547 1265 562
rect 1354 547 1384 573
rect 1779 568 1809 594
rect 1951 592 1981 618
rect 2041 592 2071 618
rect 1482 408 1512 423
rect 1672 408 1702 423
rect 1479 398 1515 408
rect 83 344 219 360
rect 397 347 427 362
rect 498 347 528 362
rect 589 347 619 362
rect 713 347 743 362
rect 803 347 833 362
rect 83 324 101 344
rect 84 310 101 324
rect 135 310 169 344
rect 203 310 219 344
rect 84 294 219 310
rect 267 314 333 330
rect 84 202 114 294
rect 170 202 200 294
rect 267 280 283 314
rect 317 294 333 314
rect 394 294 430 347
rect 495 320 531 347
rect 317 280 441 294
rect 495 290 536 320
rect 267 264 441 280
rect 411 242 441 264
rect 506 242 536 290
rect 586 257 622 347
rect 694 317 746 347
rect 694 258 724 317
rect 800 303 836 347
rect 788 273 836 303
rect 927 328 943 362
rect 977 353 1020 362
rect 1128 353 1158 368
rect 1235 364 1265 379
rect 1354 364 1384 379
rect 1452 368 1515 398
rect 1563 378 1705 408
rect 1452 364 1482 368
rect 977 328 1161 353
rect 927 323 1161 328
rect 927 294 1020 323
rect 788 258 818 273
rect 927 260 943 294
rect 977 260 1020 294
rect 1232 275 1268 364
rect 1351 347 1387 364
rect 1326 331 1392 347
rect 1326 297 1342 331
rect 1376 297 1392 331
rect 1326 281 1392 297
rect 1434 334 1482 364
rect 592 242 622 257
rect 927 244 1020 260
rect 990 222 1020 244
rect 1095 259 1278 275
rect 1095 225 1111 259
rect 1145 245 1278 259
rect 1348 253 1378 281
rect 1434 253 1464 334
rect 1563 320 1593 378
rect 2165 592 2195 618
rect 2255 592 2285 618
rect 2540 568 2570 594
rect 2657 592 2687 618
rect 2747 592 2777 618
rect 2855 592 2885 618
rect 2947 592 2977 618
rect 1779 353 1809 368
rect 1951 353 1981 368
rect 2041 353 2071 368
rect 2165 353 2195 368
rect 2255 353 2285 368
rect 2540 353 2570 368
rect 2657 353 2687 368
rect 2747 353 2777 368
rect 2855 353 2885 368
rect 2947 353 2977 368
rect 1776 330 1812 353
rect 1532 290 1593 320
rect 1641 314 1812 330
rect 1532 275 1562 290
rect 1641 280 1657 314
rect 1691 280 1725 314
rect 1759 294 1812 314
rect 1948 336 1984 353
rect 2038 336 2074 353
rect 2162 336 2198 353
rect 2252 337 2288 353
rect 2252 336 2382 337
rect 2537 336 2573 353
rect 2654 336 2690 353
rect 2744 336 2780 353
rect 2852 336 2888 353
rect 2944 336 2980 353
rect 1948 320 2382 336
rect 1759 280 1900 294
rect 1145 225 1161 245
rect 1248 230 1278 245
rect 84 48 114 74
rect 170 48 200 74
rect 411 68 441 94
rect 506 88 536 114
rect 592 56 622 114
rect 694 104 724 130
rect 788 108 818 130
rect 788 92 877 108
rect 788 58 827 92
rect 861 58 877 92
rect 788 56 877 58
rect 592 26 877 56
rect 1095 209 1161 225
rect 1641 264 1900 280
rect 1948 286 1964 320
rect 1998 286 2032 320
rect 2066 286 2100 320
rect 2134 286 2382 320
rect 1948 270 2382 286
rect 2530 320 2596 336
rect 2530 286 2546 320
rect 2580 286 2596 320
rect 2530 270 2596 286
rect 2654 320 2980 336
rect 2654 286 2679 320
rect 2713 286 2747 320
rect 2781 286 2815 320
rect 2849 286 2980 320
rect 2654 274 2980 286
rect 2654 270 2974 274
rect 1870 248 1900 264
rect 2070 248 2100 270
rect 2156 248 2186 270
rect 2266 248 2296 270
rect 2352 248 2382 270
rect 2566 248 2596 270
rect 2686 248 2716 270
rect 2772 248 2802 270
rect 2858 248 2888 270
rect 2944 248 2974 270
rect 1248 76 1278 102
rect 990 48 1020 74
rect 1348 51 1378 125
rect 1434 99 1464 125
rect 1532 51 1562 147
rect 1870 94 1900 120
rect 1348 21 1562 51
rect 2070 74 2100 100
rect 2156 74 2186 100
rect 2266 74 2296 100
rect 2352 74 2382 100
rect 2566 94 2596 120
rect 2686 74 2716 100
rect 2772 74 2802 100
rect 2858 74 2888 100
rect 2944 74 2974 100
<< polycont >>
rect 943 532 977 566
rect 943 464 977 498
rect 943 396 977 430
rect 101 310 135 344
rect 169 310 203 344
rect 283 280 317 314
rect 943 328 977 362
rect 943 260 977 294
rect 1342 297 1376 331
rect 1111 225 1145 259
rect 1657 280 1691 314
rect 1725 280 1759 314
rect 827 58 861 92
rect 1964 286 1998 320
rect 2032 286 2066 320
rect 2100 286 2134 320
rect 2546 286 2580 320
rect 2679 286 2713 320
rect 2747 286 2781 320
rect 2815 286 2849 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 17 580 73 596
rect 17 546 39 580
rect 17 512 73 546
rect 17 478 39 512
rect 17 444 73 478
rect 17 410 39 444
rect 17 394 73 410
rect 113 580 163 649
rect 315 628 383 649
rect 113 546 129 580
rect 113 512 163 546
rect 113 478 129 512
rect 113 444 163 478
rect 113 410 129 444
rect 113 394 163 410
rect 203 580 269 596
rect 315 594 332 628
rect 366 594 383 628
rect 203 546 219 580
rect 253 560 269 580
rect 633 576 699 592
rect 633 560 649 576
rect 253 546 649 560
rect 203 542 649 546
rect 683 542 699 576
rect 203 526 699 542
rect 935 566 1031 582
rect 203 512 269 526
rect 203 478 219 512
rect 253 478 269 512
rect 203 444 269 478
rect 203 410 219 444
rect 253 410 269 444
rect 203 394 269 410
rect 17 268 51 394
rect 85 344 219 360
rect 85 310 101 344
rect 135 310 169 344
rect 203 310 219 344
rect 85 302 219 310
rect 267 314 333 330
rect 267 280 283 314
rect 317 280 333 314
rect 267 268 333 280
rect 17 234 333 268
rect 17 190 73 234
rect 367 200 401 526
rect 846 518 901 534
rect 435 488 846 492
rect 435 454 451 488
rect 485 484 846 488
rect 880 484 901 518
rect 485 458 901 484
rect 485 454 501 458
rect 435 408 501 454
rect 846 437 901 458
rect 435 374 451 408
rect 485 374 501 408
rect 435 358 501 374
rect 541 408 592 424
rect 575 374 592 408
rect 17 156 39 190
rect 17 120 73 156
rect 17 86 39 120
rect 17 70 73 86
rect 109 184 159 200
rect 109 150 125 184
rect 109 116 159 150
rect 109 82 125 116
rect 109 17 159 82
rect 195 192 401 200
rect 461 196 495 358
rect 541 356 592 374
rect 675 390 703 424
rect 737 422 806 424
rect 737 390 756 422
rect 675 388 756 390
rect 790 388 806 422
rect 675 387 806 388
rect 880 403 901 437
rect 846 387 901 403
rect 541 350 641 356
rect 541 316 607 350
rect 541 310 641 316
rect 675 276 709 387
rect 195 188 427 192
rect 195 154 211 188
rect 245 158 427 188
rect 245 154 261 158
rect 195 120 261 154
rect 195 86 211 120
rect 245 86 261 120
rect 195 70 261 86
rect 307 108 359 124
rect 307 74 324 108
rect 358 74 359 108
rect 307 17 359 74
rect 393 85 427 158
rect 461 125 495 162
rect 531 242 709 276
rect 743 350 833 353
rect 743 316 799 350
rect 743 310 833 316
rect 743 246 777 310
rect 867 262 901 387
rect 531 234 597 242
rect 531 200 547 234
rect 581 200 597 234
rect 531 166 597 200
rect 531 132 547 166
rect 581 132 597 166
rect 531 125 597 132
rect 631 184 683 208
rect 631 150 633 184
rect 667 150 683 184
rect 631 85 683 150
rect 743 176 777 212
rect 813 244 901 262
rect 935 532 943 566
rect 977 532 1031 566
rect 935 498 1031 532
rect 935 464 943 498
rect 977 464 1031 498
rect 935 458 1031 464
rect 1065 580 1131 649
rect 1823 624 1937 649
rect 1065 546 1081 580
rect 1115 546 1131 580
rect 1065 494 1131 546
rect 1065 460 1081 494
rect 1115 460 1131 494
rect 1065 458 1131 460
rect 1171 580 1205 596
rect 1171 512 1205 546
rect 935 430 985 458
rect 935 396 943 430
rect 977 396 985 430
rect 1171 440 1205 478
rect 935 362 985 396
rect 935 328 943 362
rect 977 328 985 362
rect 935 294 985 328
rect 935 260 943 294
rect 977 260 985 294
rect 935 244 985 260
rect 1019 406 1171 424
rect 1019 390 1205 406
rect 1239 581 1743 615
rect 1823 590 1863 624
rect 1897 590 1937 624
rect 2085 625 2151 649
rect 2085 591 2101 625
rect 2135 591 2151 625
rect 2085 590 2151 591
rect 2299 624 2425 649
rect 2299 590 2345 624
rect 2379 590 2425 624
rect 1239 430 1273 581
rect 1398 579 1575 581
rect 1307 522 1357 547
rect 1398 545 1424 579
rect 1458 545 1575 579
rect 1709 556 1743 581
rect 2584 580 2650 649
rect 2459 560 2543 572
rect 2459 556 2493 560
rect 1341 498 1357 522
rect 1341 488 1507 498
rect 1307 464 1507 488
rect 1239 396 1297 430
rect 813 210 829 244
rect 863 210 901 244
rect 813 209 901 210
rect 1019 184 1053 390
rect 1087 350 1127 356
rect 1121 316 1127 350
rect 1087 275 1127 316
rect 1177 350 1229 356
rect 1177 316 1183 350
rect 1217 316 1229 350
rect 1177 310 1229 316
rect 1087 259 1161 275
rect 1087 225 1111 259
rect 1145 225 1161 259
rect 1087 218 1161 225
rect 1195 221 1229 310
rect 1263 243 1297 396
rect 1331 424 1415 430
rect 1331 390 1375 424
rect 1409 390 1415 424
rect 1331 331 1415 390
rect 1331 297 1342 331
rect 1376 297 1415 331
rect 1331 281 1415 297
rect 1473 257 1507 464
rect 1541 330 1575 545
rect 1609 513 1625 547
rect 1659 513 1675 547
rect 1709 526 2493 556
rect 2527 526 2543 560
rect 1709 522 2543 526
rect 1609 488 1675 513
rect 2459 492 2543 522
rect 1609 469 2425 488
rect 1609 435 1625 469
rect 1659 454 2425 469
rect 1659 435 1675 454
rect 1609 419 1675 435
rect 1716 417 1843 420
rect 1716 383 1732 417
rect 1766 383 1843 417
rect 1716 380 1843 383
rect 1809 355 1843 380
rect 1978 386 1994 420
rect 2028 386 2208 420
rect 2242 386 2279 420
rect 1978 370 2279 386
rect 1809 350 1895 355
rect 1541 314 1775 330
rect 1541 296 1657 314
rect 1641 280 1657 296
rect 1691 280 1725 314
rect 1759 280 1775 314
rect 1641 264 1775 280
rect 1809 316 1855 350
rect 1889 316 1895 350
rect 1809 310 1895 316
rect 1956 320 2142 336
rect 1263 239 1439 243
rect 1263 209 1389 239
rect 1373 205 1389 209
rect 1423 205 1439 239
rect 1373 203 1439 205
rect 1473 239 1537 257
rect 1473 205 1487 239
rect 1521 221 1537 239
rect 1809 237 1843 310
rect 1521 205 1775 221
rect 1473 187 1775 205
rect 1956 286 1964 320
rect 1998 286 2032 320
rect 2066 286 2100 320
rect 2134 286 2142 320
rect 1956 270 2142 286
rect 1956 236 1990 270
rect 2192 252 2279 370
rect 2192 236 2357 252
rect 1809 187 1843 203
rect 1877 202 1990 236
rect 2095 202 2111 236
rect 2145 202 2307 236
rect 2341 202 2357 236
rect 1019 175 1031 184
rect 743 126 777 142
rect 811 150 1031 175
rect 1065 150 1081 184
rect 1195 175 1229 187
rect 811 141 1081 150
rect 393 51 683 85
rect 811 92 877 141
rect 1019 116 1081 141
rect 1175 153 1241 175
rect 1175 119 1191 153
rect 1225 119 1241 153
rect 1275 153 1341 169
rect 1741 153 1775 187
rect 1877 153 1911 202
rect 2391 168 2425 454
rect 2459 458 2493 492
rect 2527 458 2543 492
rect 2459 424 2543 458
rect 2459 236 2493 424
rect 2527 390 2543 424
rect 2584 546 2600 580
rect 2634 546 2650 580
rect 2584 503 2650 546
rect 2584 469 2600 503
rect 2634 469 2650 503
rect 2584 424 2650 469
rect 2584 390 2600 424
rect 2634 390 2650 424
rect 2684 580 2750 596
rect 2684 546 2700 580
rect 2734 546 2750 580
rect 2684 500 2750 546
rect 2684 466 2700 500
rect 2734 466 2750 500
rect 2684 420 2750 466
rect 2784 580 2850 649
rect 2784 546 2800 580
rect 2834 546 2850 580
rect 2784 488 2850 546
rect 2784 454 2800 488
rect 2834 454 2850 488
rect 2784 438 2850 454
rect 2884 580 2951 596
rect 2884 546 2900 580
rect 2934 546 2951 580
rect 2884 500 2951 546
rect 2884 466 2900 500
rect 2934 466 2951 500
rect 2684 386 2700 420
rect 2734 404 2750 420
rect 2884 420 2951 466
rect 2884 404 2900 420
rect 2734 386 2900 404
rect 2934 386 2951 420
rect 2684 370 2951 386
rect 2990 580 3040 649
rect 3024 546 3040 580
rect 2990 497 3040 546
rect 3024 463 3040 497
rect 2990 414 3040 463
rect 3024 380 3040 414
rect 2527 320 2596 356
rect 2527 286 2546 320
rect 2580 286 2596 320
rect 2527 270 2596 286
rect 2643 320 2865 336
rect 2643 286 2679 320
rect 2713 286 2747 320
rect 2781 286 2815 320
rect 2849 286 2865 320
rect 2643 270 2865 286
rect 2459 202 2521 236
rect 2555 202 2571 236
rect 2643 168 2677 270
rect 2899 236 2949 370
rect 2990 364 3040 380
rect 1275 119 1291 153
rect 1325 119 1707 153
rect 1741 119 1911 153
rect 1945 134 2677 168
rect 2711 220 2899 236
rect 2711 186 2727 220
rect 2761 202 2899 220
rect 2933 202 2949 236
rect 2711 146 2761 186
rect 811 58 827 92
rect 861 58 877 92
rect 811 51 877 58
rect 917 91 983 107
rect 917 57 933 91
rect 967 57 983 91
rect 917 17 983 57
rect 1019 82 1031 116
rect 1065 85 1081 116
rect 1673 85 1707 119
rect 1945 85 1979 134
rect 2711 112 2727 146
rect 1065 82 1589 85
rect 1019 51 1589 82
rect 1623 51 1639 85
rect 1673 51 1979 85
rect 2013 84 2063 100
rect 2047 50 2063 84
rect 2013 17 2063 50
rect 2193 84 2259 100
rect 2193 50 2209 84
rect 2243 50 2259 84
rect 2193 17 2259 50
rect 2393 84 2459 100
rect 2393 50 2409 84
rect 2443 50 2459 84
rect 2393 17 2459 50
rect 2607 84 2675 100
rect 2711 96 2761 112
rect 2797 157 2863 168
rect 2797 123 2813 157
rect 2847 123 2863 157
rect 2607 50 2624 84
rect 2658 50 2675 84
rect 2607 17 2675 50
rect 2797 17 2863 123
rect 2899 146 2949 202
rect 2933 112 2949 146
rect 2899 96 2949 112
rect 2983 236 3049 252
rect 2983 202 2999 236
rect 3033 202 3049 236
rect 2983 146 3049 202
rect 2983 112 2999 146
rect 3033 112 3049 146
rect 2983 17 3049 112
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 703 390 737 424
rect 607 316 641 350
rect 799 316 833 350
rect 1087 316 1121 350
rect 1183 316 1217 350
rect 1375 390 1409 424
rect 1855 316 1889 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 683 3072 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 0 617 3072 649
rect 691 424 749 430
rect 691 390 703 424
rect 737 421 749 424
rect 1363 424 1421 430
rect 1363 421 1375 424
rect 737 393 1375 421
rect 737 390 749 393
rect 691 384 749 390
rect 1363 390 1375 393
rect 1409 390 1421 424
rect 1363 384 1421 390
rect 595 350 653 356
rect 595 316 607 350
rect 641 347 653 350
rect 787 350 845 356
rect 787 347 799 350
rect 641 319 799 347
rect 641 316 653 319
rect 595 310 653 316
rect 787 316 799 319
rect 833 347 845 350
rect 1075 350 1133 356
rect 1075 347 1087 350
rect 833 319 1087 347
rect 833 316 845 319
rect 787 310 845 316
rect 1075 316 1087 319
rect 1121 316 1133 350
rect 1075 310 1133 316
rect 1171 350 1229 356
rect 1171 316 1183 350
rect 1217 347 1229 350
rect 1843 350 1901 356
rect 1843 347 1855 350
rect 1217 319 1855 347
rect 1217 316 1229 319
rect 1171 310 1229 316
rect 1843 316 1855 319
rect 1889 316 1901 350
rect 1843 310 1901 316
rect 0 17 3072 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
rect 0 -49 3072 -17
<< labels >>
rlabel comment s 0 0 0 0 4 fah_4
flabel pwell s 0 0 3072 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 3072 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 0 617 3072 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 0 0 3072 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel locali s 2911 390 2945 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2911 464 2945 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2911 538 2945 572 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2239 316 2273 350 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 991 464 1025 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 991 538 1025 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 2527 316 2561 350 0 FreeSans 340 0 0 0 CI
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3072 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 3403038
string GDS_START 3380906
<< end >>
