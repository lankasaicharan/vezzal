magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4178 1975
<< nwell >>
rect -38 331 2918 704
<< pwell >>
rect 15 157 527 238
rect 1741 235 2047 279
rect 2572 235 2862 263
rect 952 167 1082 191
rect 1393 167 2862 235
rect 952 157 2862 167
rect 15 49 2862 157
rect 0 0 2880 49
<< scnmos >>
rect 94 128 124 212
rect 166 128 196 212
rect 252 128 282 212
rect 324 128 354 212
rect 418 128 448 212
rect 755 47 785 131
rect 841 47 871 131
rect 1105 57 1135 141
rect 1191 57 1221 141
rect 1263 57 1293 141
rect 1472 125 1502 209
rect 1574 125 1604 209
rect 1817 125 1847 253
rect 1889 125 1919 253
rect 2086 125 2116 209
rect 2194 125 2224 209
rect 2266 125 2296 209
rect 2374 125 2404 209
rect 2651 153 2681 237
rect 2753 69 2783 237
<< scpmoshvt >>
rect 80 408 110 536
rect 166 408 196 536
rect 238 408 268 536
rect 346 408 376 536
rect 606 481 636 609
rect 823 483 853 611
rect 909 483 939 611
rect 1105 463 1135 547
rect 1191 463 1221 547
rect 1263 463 1293 547
rect 1415 463 1445 547
rect 1504 463 1534 547
rect 1673 379 1703 547
rect 1882 463 1912 547
rect 1991 379 2021 547
rect 2187 483 2217 567
rect 2273 483 2303 567
rect 2463 483 2493 567
rect 2653 367 2683 495
rect 2770 367 2800 619
<< ndiff >>
rect 41 187 94 212
rect 41 153 49 187
rect 83 153 94 187
rect 41 128 94 153
rect 124 128 166 212
rect 196 187 252 212
rect 196 153 207 187
rect 241 153 252 187
rect 196 128 252 153
rect 282 128 324 212
rect 354 187 418 212
rect 354 153 365 187
rect 399 153 418 187
rect 354 128 418 153
rect 448 198 501 212
rect 448 164 459 198
rect 493 164 501 198
rect 448 128 501 164
rect 978 157 1056 165
rect 702 106 755 131
rect 702 72 710 106
rect 744 72 755 106
rect 702 47 755 72
rect 785 106 841 131
rect 785 72 796 106
rect 830 72 841 106
rect 785 47 841 72
rect 871 106 924 131
rect 871 72 882 106
rect 916 72 924 106
rect 871 47 924 72
rect 978 123 990 157
rect 1024 141 1056 157
rect 1767 209 1817 253
rect 1419 182 1472 209
rect 1419 148 1427 182
rect 1461 148 1472 182
rect 1024 123 1105 141
rect 978 57 1105 123
rect 1135 115 1191 141
rect 1135 81 1146 115
rect 1180 81 1191 115
rect 1135 57 1191 81
rect 1221 57 1263 141
rect 1293 117 1346 141
rect 1419 125 1472 148
rect 1502 125 1574 209
rect 1604 198 1817 209
rect 1604 164 1721 198
rect 1755 164 1817 198
rect 1604 125 1817 164
rect 1847 125 1889 253
rect 1919 245 2021 253
rect 1919 211 1930 245
rect 1964 211 2021 245
rect 1919 209 2021 211
rect 2598 212 2651 237
rect 1919 201 2086 209
rect 1919 167 2006 201
rect 2040 167 2086 201
rect 1919 125 2086 167
rect 2116 125 2194 209
rect 2224 125 2266 209
rect 2296 183 2374 209
rect 2296 149 2315 183
rect 2349 149 2374 183
rect 2296 125 2374 149
rect 2404 183 2457 209
rect 2404 149 2415 183
rect 2449 149 2457 183
rect 2598 178 2606 212
rect 2640 178 2651 212
rect 2598 153 2651 178
rect 2681 225 2753 237
rect 2681 191 2696 225
rect 2730 191 2753 225
rect 2681 153 2753 191
rect 2404 125 2457 149
rect 1293 83 1304 117
rect 1338 83 1346 117
rect 1293 57 1346 83
rect 2700 115 2753 153
rect 2700 81 2708 115
rect 2742 81 2753 115
rect 2700 69 2753 81
rect 2783 209 2836 237
rect 2783 175 2794 209
rect 2828 175 2836 209
rect 2783 115 2836 175
rect 2783 81 2794 115
rect 2828 81 2836 115
rect 2783 69 2836 81
<< pdiff >>
rect 483 609 557 610
rect 483 598 606 609
rect 483 564 491 598
rect 525 564 606 598
rect 27 524 80 536
rect 27 490 35 524
rect 69 490 80 524
rect 27 454 80 490
rect 27 420 35 454
rect 69 420 80 454
rect 27 408 80 420
rect 110 520 166 536
rect 110 486 121 520
rect 155 486 166 520
rect 110 408 166 486
rect 196 408 238 536
rect 268 511 346 536
rect 268 477 290 511
rect 324 477 346 511
rect 268 408 346 477
rect 376 456 429 536
rect 483 481 606 564
rect 636 529 689 609
rect 636 495 647 529
rect 681 495 689 529
rect 636 481 689 495
rect 743 483 823 611
rect 853 603 909 611
rect 853 569 864 603
rect 898 569 909 603
rect 853 483 909 569
rect 939 589 992 611
rect 939 555 950 589
rect 984 555 992 589
rect 939 483 992 555
rect 376 422 387 456
rect 421 422 429 456
rect 376 408 429 422
rect 743 463 801 483
rect 743 429 755 463
rect 789 429 801 463
rect 743 421 801 429
rect 1810 559 1860 573
rect 1052 522 1105 547
rect 1052 488 1060 522
rect 1094 488 1105 522
rect 1052 463 1105 488
rect 1135 522 1191 547
rect 1135 488 1146 522
rect 1180 488 1191 522
rect 1135 463 1191 488
rect 1221 463 1263 547
rect 1293 524 1415 547
rect 1293 490 1304 524
rect 1338 490 1415 524
rect 1293 463 1415 490
rect 1445 518 1504 547
rect 1445 484 1456 518
rect 1490 484 1504 518
rect 1445 463 1504 484
rect 1534 535 1673 547
rect 1534 501 1599 535
rect 1633 501 1673 535
rect 1534 467 1673 501
rect 1534 463 1612 467
rect 1604 433 1612 463
rect 1646 433 1673 467
rect 1604 379 1673 433
rect 1703 535 1756 547
rect 1703 501 1714 535
rect 1748 501 1756 535
rect 1703 467 1756 501
rect 1703 433 1714 467
rect 1748 433 1756 467
rect 1810 525 1818 559
rect 1852 547 1860 559
rect 1852 525 1882 547
rect 1810 463 1882 525
rect 1912 463 1991 547
rect 1703 379 1756 433
rect 1934 421 1991 463
rect 1934 387 1946 421
rect 1980 387 1991 421
rect 1934 379 1991 387
rect 2021 503 2074 547
rect 2021 469 2032 503
rect 2066 469 2074 503
rect 2021 390 2074 469
rect 2021 379 2071 390
rect 2717 607 2770 619
rect 2717 573 2725 607
rect 2759 573 2770 607
rect 2134 543 2187 567
rect 2134 509 2142 543
rect 2176 509 2187 543
rect 2134 483 2187 509
rect 2217 543 2273 567
rect 2217 509 2228 543
rect 2262 509 2273 543
rect 2217 483 2273 509
rect 2303 543 2356 567
rect 2303 509 2314 543
rect 2348 509 2356 543
rect 2303 483 2356 509
rect 2410 543 2463 567
rect 2410 509 2418 543
rect 2452 509 2463 543
rect 2410 483 2463 509
rect 2493 543 2546 567
rect 2493 509 2504 543
rect 2538 509 2546 543
rect 2493 483 2546 509
rect 2717 507 2770 573
rect 2717 495 2725 507
rect 2600 483 2653 495
rect 2600 449 2608 483
rect 2642 449 2653 483
rect 2600 413 2653 449
rect 2600 379 2608 413
rect 2642 379 2653 413
rect 2600 367 2653 379
rect 2683 473 2725 495
rect 2759 473 2770 507
rect 2683 413 2770 473
rect 2683 379 2694 413
rect 2728 379 2770 413
rect 2683 367 2770 379
rect 2800 599 2853 619
rect 2800 565 2811 599
rect 2845 565 2853 599
rect 2800 505 2853 565
rect 2800 471 2811 505
rect 2845 471 2853 505
rect 2800 420 2853 471
rect 2800 386 2811 420
rect 2845 386 2853 420
rect 2800 367 2853 386
<< ndiffc >>
rect 49 153 83 187
rect 207 153 241 187
rect 365 153 399 187
rect 459 164 493 198
rect 710 72 744 106
rect 796 72 830 106
rect 882 72 916 106
rect 990 123 1024 157
rect 1427 148 1461 182
rect 1146 81 1180 115
rect 1721 164 1755 198
rect 1930 211 1964 245
rect 2006 167 2040 201
rect 2315 149 2349 183
rect 2415 149 2449 183
rect 2606 178 2640 212
rect 2696 191 2730 225
rect 1304 83 1338 117
rect 2708 81 2742 115
rect 2794 175 2828 209
rect 2794 81 2828 115
<< pdiffc >>
rect 491 564 525 598
rect 35 490 69 524
rect 35 420 69 454
rect 121 486 155 520
rect 290 477 324 511
rect 647 495 681 529
rect 864 569 898 603
rect 950 555 984 589
rect 387 422 421 456
rect 755 429 789 463
rect 1060 488 1094 522
rect 1146 488 1180 522
rect 1304 490 1338 524
rect 1456 484 1490 518
rect 1599 501 1633 535
rect 1612 433 1646 467
rect 1714 501 1748 535
rect 1714 433 1748 467
rect 1818 525 1852 559
rect 1946 387 1980 421
rect 2032 469 2066 503
rect 2725 573 2759 607
rect 2142 509 2176 543
rect 2228 509 2262 543
rect 2314 509 2348 543
rect 2418 509 2452 543
rect 2504 509 2538 543
rect 2608 449 2642 483
rect 2608 379 2642 413
rect 2725 473 2759 507
rect 2694 379 2728 413
rect 2811 565 2845 599
rect 2811 471 2845 505
rect 2811 386 2845 420
<< poly >>
rect 606 609 636 635
rect 823 611 853 637
rect 909 611 939 637
rect 1007 615 2119 645
rect 2770 619 2800 645
rect 80 536 110 562
rect 166 536 196 562
rect 238 536 268 562
rect 346 536 376 562
rect 606 436 636 481
rect 80 368 110 408
rect 58 352 124 368
rect 58 318 74 352
rect 108 318 124 352
rect 58 284 124 318
rect 58 250 74 284
rect 108 250 124 284
rect 58 234 124 250
rect 94 212 124 234
rect 166 212 196 408
rect 238 372 268 408
rect 238 356 304 372
rect 238 322 254 356
rect 288 322 304 356
rect 238 306 304 322
rect 346 316 376 408
rect 606 406 683 436
rect 539 342 605 358
rect 539 316 555 342
rect 346 308 555 316
rect 589 308 605 342
rect 252 212 282 306
rect 346 286 605 308
rect 346 264 376 286
rect 324 234 376 264
rect 539 274 605 286
rect 539 240 555 274
rect 589 240 605 274
rect 324 212 354 234
rect 418 212 448 238
rect 539 224 605 240
rect 653 176 683 406
rect 823 365 853 483
rect 909 451 939 483
rect 1007 451 1037 615
rect 1105 547 1135 573
rect 1191 547 1221 615
rect 1263 547 1293 573
rect 1415 547 1445 573
rect 1504 547 1534 573
rect 1673 547 1703 573
rect 559 146 683 176
rect 755 349 853 365
rect 755 315 799 349
rect 833 315 853 349
rect 755 281 853 315
rect 755 247 799 281
rect 833 247 853 281
rect 755 231 853 247
rect 901 435 1037 451
rect 901 401 917 435
rect 951 421 1037 435
rect 951 401 967 421
rect 901 255 967 401
rect 1105 369 1135 463
rect 1191 437 1221 463
rect 1263 441 1293 463
rect 1415 441 1445 463
rect 1263 411 1360 441
rect 1415 411 1462 441
rect 1330 369 1360 411
rect 1060 353 1282 369
rect 1060 319 1076 353
rect 1110 319 1232 353
rect 1266 319 1282 353
rect 1060 303 1282 319
rect 1324 353 1390 369
rect 1324 319 1340 353
rect 1374 319 1390 353
rect 1324 303 1390 319
rect 94 102 124 128
rect 166 54 196 128
rect 252 102 282 128
rect 324 102 354 128
rect 418 54 448 128
rect 559 103 589 146
rect 755 131 785 231
rect 901 225 1135 255
rect 901 183 931 225
rect 841 153 931 183
rect 841 131 871 153
rect 523 87 589 103
rect 523 54 539 87
rect 166 53 539 54
rect 573 53 589 87
rect 166 24 589 53
rect 1105 141 1135 225
rect 1191 141 1221 303
rect 1330 229 1360 303
rect 1432 299 1462 411
rect 1504 377 1534 463
rect 1882 547 1912 573
rect 1991 547 2021 573
rect 1882 419 1912 463
rect 1828 403 1919 419
rect 1504 347 1589 377
rect 1559 341 1589 347
rect 1673 341 1703 379
rect 1828 369 1844 403
rect 1878 369 1919 403
rect 1828 353 1919 369
rect 1559 311 1604 341
rect 1432 283 1502 299
rect 1432 249 1448 283
rect 1482 249 1502 283
rect 1432 233 1502 249
rect 1263 213 1360 229
rect 1263 179 1310 213
rect 1344 179 1360 213
rect 1472 209 1502 233
rect 1574 209 1604 311
rect 1673 325 1739 341
rect 1673 291 1689 325
rect 1723 305 1739 325
rect 1723 291 1847 305
rect 1673 275 1847 291
rect 1817 253 1847 275
rect 1889 253 1919 353
rect 1991 357 2021 379
rect 2089 375 2119 615
rect 2187 567 2217 593
rect 2273 567 2303 593
rect 2463 567 2493 593
rect 2653 495 2683 521
rect 2086 357 2119 375
rect 1991 345 2119 357
rect 1991 327 2116 345
rect 1263 163 1360 179
rect 1263 141 1293 163
rect 2086 209 2116 327
rect 2187 297 2217 483
rect 2273 367 2303 483
rect 2463 451 2493 483
rect 2418 435 2493 451
rect 2418 401 2434 435
rect 2468 401 2493 435
rect 2418 367 2493 401
rect 2266 351 2332 367
rect 2266 317 2282 351
rect 2316 317 2332 351
rect 2418 345 2434 367
rect 2266 301 2332 317
rect 2374 333 2434 345
rect 2468 345 2493 367
rect 2653 345 2683 367
rect 2468 333 2683 345
rect 2374 315 2683 333
rect 2770 325 2800 367
rect 2158 281 2224 297
rect 2158 247 2174 281
rect 2208 247 2224 281
rect 2158 231 2224 247
rect 2194 209 2224 231
rect 2266 231 2302 301
rect 2266 209 2296 231
rect 2374 209 2404 315
rect 2651 237 2681 315
rect 2729 309 2800 325
rect 2729 275 2745 309
rect 2779 275 2800 309
rect 2729 259 2800 275
rect 2753 237 2783 259
rect 2651 127 2681 153
rect 1472 99 1502 125
rect 1574 103 1604 125
rect 1574 87 1640 103
rect 1817 99 1847 125
rect 1889 99 1919 125
rect 2086 99 2116 125
rect 2194 99 2224 125
rect 2266 99 2296 125
rect 2374 99 2404 125
rect 755 21 785 47
rect 841 21 871 47
rect 1105 31 1135 57
rect 1191 31 1221 57
rect 1263 31 1293 57
rect 1574 53 1590 87
rect 1624 53 1640 87
rect 1574 37 1640 53
rect 2753 43 2783 69
<< polycont >>
rect 74 318 108 352
rect 74 250 108 284
rect 254 322 288 356
rect 555 308 589 342
rect 555 240 589 274
rect 799 315 833 349
rect 799 247 833 281
rect 917 401 951 435
rect 1076 319 1110 353
rect 1232 319 1266 353
rect 1340 319 1374 353
rect 539 53 573 87
rect 1844 369 1878 403
rect 1448 249 1482 283
rect 1310 179 1344 213
rect 1689 291 1723 325
rect 2434 401 2468 435
rect 2282 317 2316 351
rect 2434 333 2468 367
rect 2174 247 2208 281
rect 2745 275 2779 309
rect 1590 53 1624 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 19 524 78 540
rect 19 490 35 524
rect 69 490 78 524
rect 19 454 78 490
rect 112 520 171 649
rect 475 598 541 649
rect 475 564 491 598
rect 525 564 541 598
rect 475 562 541 564
rect 577 579 812 613
rect 577 528 611 579
rect 112 486 121 520
rect 155 486 171 520
rect 112 470 171 486
rect 274 511 611 528
rect 274 477 290 511
rect 324 490 611 511
rect 645 529 688 545
rect 645 495 647 529
rect 681 495 688 529
rect 778 533 812 579
rect 848 603 914 649
rect 848 569 864 603
rect 898 569 914 603
rect 948 589 1250 607
rect 948 555 950 589
rect 984 573 1250 589
rect 984 555 1000 573
rect 948 539 1000 555
rect 778 505 914 533
rect 1040 522 1110 538
rect 1040 505 1060 522
rect 778 499 1060 505
rect 324 477 340 490
rect 274 470 340 477
rect 19 420 35 454
rect 69 436 78 454
rect 371 436 387 456
rect 69 422 387 436
rect 421 422 437 456
rect 69 420 437 422
rect 19 402 437 420
rect 31 352 124 368
rect 31 318 74 352
rect 108 318 124 352
rect 31 284 124 318
rect 203 356 451 368
rect 203 322 254 356
rect 288 322 451 356
rect 203 306 451 322
rect 31 250 74 284
rect 108 250 124 284
rect 485 272 519 490
rect 645 358 688 495
rect 880 488 1060 499
rect 1094 488 1110 522
rect 880 471 1110 488
rect 31 234 124 250
rect 191 238 519 272
rect 553 342 688 358
rect 553 308 555 342
rect 589 324 688 342
rect 722 429 755 463
rect 789 437 805 463
rect 1006 459 1110 471
rect 1144 522 1180 538
rect 1144 488 1146 522
rect 789 435 967 437
rect 789 429 917 435
rect 722 401 917 429
rect 951 401 967 435
rect 722 399 967 401
rect 589 308 605 324
rect 553 274 605 308
rect 553 240 555 274
rect 589 240 605 274
rect 33 187 99 200
rect 33 153 49 187
rect 83 153 99 187
rect 33 17 99 153
rect 191 187 257 238
rect 553 204 605 240
rect 191 153 207 187
rect 241 153 257 187
rect 191 137 257 153
rect 349 187 403 203
rect 349 153 365 187
rect 399 153 403 187
rect 443 198 605 204
rect 443 164 459 198
rect 493 164 605 198
rect 443 162 605 164
rect 349 17 403 153
rect 486 87 655 128
rect 722 122 756 399
rect 790 349 857 365
rect 790 315 799 349
rect 833 315 857 349
rect 790 281 857 315
rect 790 247 799 281
rect 833 247 857 281
rect 790 156 857 247
rect 1006 161 1040 459
rect 974 157 1040 161
rect 974 123 990 157
rect 1024 123 1040 157
rect 486 53 539 87
rect 573 53 655 87
rect 694 106 756 122
rect 694 72 710 106
rect 744 72 756 106
rect 694 56 756 72
rect 790 106 840 122
rect 790 72 796 106
rect 830 72 840 106
rect 790 17 840 72
rect 874 106 932 122
rect 974 121 1040 123
rect 1074 353 1110 369
rect 1074 319 1076 353
rect 874 72 882 106
rect 916 87 932 106
rect 1074 87 1110 319
rect 916 72 1110 87
rect 874 53 1110 72
rect 1144 285 1180 488
rect 1216 423 1250 573
rect 1288 524 1344 649
rect 1288 490 1304 524
rect 1338 490 1344 524
rect 1288 474 1344 490
rect 1378 568 1560 602
rect 1378 423 1412 568
rect 1216 389 1412 423
rect 1446 518 1492 534
rect 1446 484 1456 518
rect 1490 484 1492 518
rect 1216 353 1282 389
rect 1446 355 1492 484
rect 1526 397 1560 568
rect 1594 535 1662 649
rect 1802 559 2184 593
rect 1594 501 1599 535
rect 1633 501 1662 535
rect 1594 467 1662 501
rect 1594 433 1612 467
rect 1646 433 1662 467
rect 1594 431 1662 433
rect 1698 535 1764 551
rect 1698 501 1714 535
rect 1748 501 1764 535
rect 1802 525 1818 559
rect 1852 525 1868 559
rect 2126 543 2184 559
rect 1698 491 1764 501
rect 2016 503 2082 525
rect 2016 491 2032 503
rect 1698 469 2032 491
rect 2066 469 2082 503
rect 2126 509 2142 543
rect 2176 509 2184 543
rect 2126 493 2184 509
rect 2218 543 2270 649
rect 2218 509 2228 543
rect 2262 509 2270 543
rect 2218 493 2270 509
rect 2304 543 2352 559
rect 2304 509 2314 543
rect 2348 509 2352 543
rect 1698 467 2082 469
rect 1698 433 1714 467
rect 1748 457 2082 467
rect 1748 433 1764 457
rect 1698 431 1764 433
rect 2304 451 2352 509
rect 2402 543 2468 649
rect 2685 607 2773 649
rect 2685 573 2725 607
rect 2759 573 2773 607
rect 2402 509 2418 543
rect 2452 509 2468 543
rect 2402 493 2468 509
rect 2502 543 2554 559
rect 2502 509 2504 543
rect 2538 509 2554 543
rect 2304 435 2468 451
rect 2304 423 2434 435
rect 1928 421 2434 423
rect 1828 403 1894 421
rect 1828 397 1844 403
rect 1526 369 1844 397
rect 1878 369 1894 403
rect 1526 363 1894 369
rect 1928 387 1946 421
rect 1980 401 2434 421
rect 1980 387 2468 401
rect 1216 319 1232 353
rect 1266 319 1282 353
rect 1324 353 1492 355
rect 1324 319 1340 353
rect 1374 319 1492 353
rect 1673 325 1739 329
rect 1673 291 1689 325
rect 1723 291 1739 325
rect 1673 285 1739 291
rect 1144 283 1739 285
rect 1144 249 1448 283
rect 1482 249 1739 283
rect 1144 145 1180 249
rect 1928 245 2056 387
rect 2418 367 2468 387
rect 1294 213 1463 215
rect 1294 179 1310 213
rect 1344 182 1463 213
rect 1928 211 1930 245
rect 1964 211 2056 245
rect 1344 179 1427 182
rect 1294 167 1427 179
rect 1411 148 1427 167
rect 1461 148 1463 182
rect 1144 115 1184 145
rect 1144 81 1146 115
rect 1180 81 1184 115
rect 1144 65 1184 81
rect 1288 117 1354 133
rect 1411 132 1463 148
rect 1497 198 1771 202
rect 1497 164 1721 198
rect 1755 164 1771 198
rect 1928 201 2056 211
rect 1928 167 2006 201
rect 2040 167 2056 201
rect 1288 83 1304 117
rect 1338 83 1354 117
rect 1288 17 1354 83
rect 1497 17 1531 164
rect 1928 162 2056 167
rect 2090 351 2332 353
rect 2090 317 2282 351
rect 2316 317 2332 351
rect 2418 333 2434 367
rect 2418 317 2468 333
rect 2090 128 2124 317
rect 2502 283 2554 509
rect 2685 507 2773 573
rect 2158 281 2554 283
rect 2158 247 2174 281
rect 2208 247 2554 281
rect 2590 483 2651 499
rect 2590 449 2608 483
rect 2642 449 2651 483
rect 2590 413 2651 449
rect 2590 379 2608 413
rect 2642 379 2651 413
rect 2590 325 2651 379
rect 2685 473 2725 507
rect 2759 473 2773 507
rect 2685 413 2773 473
rect 2685 379 2694 413
rect 2728 379 2773 413
rect 2685 363 2773 379
rect 2807 599 2863 615
rect 2807 565 2811 599
rect 2845 565 2863 599
rect 2807 505 2863 565
rect 2807 471 2811 505
rect 2845 471 2863 505
rect 2807 420 2863 471
rect 2807 386 2811 420
rect 2845 386 2863 420
rect 2807 370 2863 386
rect 2590 309 2779 325
rect 2590 275 2745 309
rect 2590 259 2779 275
rect 1567 87 2124 128
rect 1567 53 1590 87
rect 1624 53 2124 87
rect 2299 183 2365 199
rect 2299 149 2315 183
rect 2349 149 2365 183
rect 2299 17 2365 149
rect 2399 183 2465 247
rect 2399 149 2415 183
rect 2449 149 2465 183
rect 2590 212 2646 259
rect 2813 225 2863 370
rect 2590 178 2606 212
rect 2640 178 2646 212
rect 2590 162 2646 178
rect 2680 191 2696 225
rect 2730 191 2751 225
rect 2399 133 2465 149
rect 2680 115 2751 191
rect 2680 81 2708 115
rect 2742 81 2751 115
rect 2680 17 2751 81
rect 2785 209 2863 225
rect 2785 175 2794 209
rect 2828 175 2863 209
rect 2785 115 2863 175
rect 2785 81 2794 115
rect 2828 81 2863 115
rect 2785 65 2863 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfstp_1
flabel comment s 1174 332 1174 332 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 1342 270 1342 270 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2815 94 2849 128 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2815 168 2849 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2815 242 2849 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2815 316 2849 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2815 390 2849 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2815 464 2849 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2815 538 2849 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 1567 94 1601 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 1663 94 1697 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 1759 94 1793 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 1855 94 1889 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 1951 94 1985 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 2047 94 2081 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2880 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 110164
string GDS_START 89786
<< end >>
