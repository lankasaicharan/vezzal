magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 7 158 293 241
rect 7 49 761 158
rect 0 0 768 49
<< scnmos >>
rect 86 47 116 215
rect 172 47 202 215
rect 289 48 319 132
rect 361 48 391 132
rect 469 48 499 132
rect 541 48 571 132
rect 652 48 682 132
<< scpmoshvt >>
rect 86 367 116 619
rect 172 367 202 619
rect 320 449 350 577
rect 392 449 422 577
rect 478 449 508 577
rect 572 449 602 577
rect 658 449 688 577
<< ndiff >>
rect 33 203 86 215
rect 33 169 41 203
rect 75 169 86 203
rect 33 93 86 169
rect 33 59 41 93
rect 75 59 86 93
rect 33 47 86 59
rect 116 203 172 215
rect 116 169 127 203
rect 161 169 172 203
rect 116 101 172 169
rect 116 67 127 101
rect 161 67 172 101
rect 116 47 172 67
rect 202 132 267 215
rect 202 81 289 132
rect 202 47 225 81
rect 259 48 289 81
rect 319 48 361 132
rect 391 109 469 132
rect 391 75 404 109
rect 438 75 469 109
rect 391 48 469 75
rect 499 48 541 132
rect 571 107 652 132
rect 571 73 597 107
rect 631 73 652 107
rect 571 48 652 73
rect 682 105 735 132
rect 682 71 693 105
rect 727 71 735 105
rect 682 48 735 71
rect 259 47 267 48
rect 217 35 267 47
<< pdiff >>
rect 33 607 86 619
rect 33 573 41 607
rect 75 573 86 607
rect 33 509 86 573
rect 33 475 41 509
rect 75 475 86 509
rect 33 413 86 475
rect 33 379 41 413
rect 75 379 86 413
rect 33 367 86 379
rect 116 599 172 619
rect 116 565 127 599
rect 161 565 172 599
rect 116 505 172 565
rect 116 471 127 505
rect 161 471 172 505
rect 116 420 172 471
rect 116 386 127 420
rect 161 386 172 420
rect 116 367 172 386
rect 202 611 259 619
rect 202 577 213 611
rect 247 577 259 611
rect 202 449 320 577
rect 350 449 392 577
rect 422 553 478 577
rect 422 519 433 553
rect 467 519 478 553
rect 422 449 478 519
rect 508 449 572 577
rect 602 547 658 577
rect 602 513 613 547
rect 647 513 658 547
rect 602 449 658 513
rect 688 563 741 577
rect 688 529 699 563
rect 733 529 741 563
rect 688 495 741 529
rect 688 461 699 495
rect 733 461 741 495
rect 688 449 741 461
rect 202 445 259 449
rect 202 367 252 445
<< ndiffc >>
rect 41 169 75 203
rect 41 59 75 93
rect 127 169 161 203
rect 127 67 161 101
rect 225 47 259 81
rect 404 75 438 109
rect 597 73 631 107
rect 693 71 727 105
<< pdiffc >>
rect 41 573 75 607
rect 41 475 75 509
rect 41 379 75 413
rect 127 565 161 599
rect 127 471 161 505
rect 127 386 161 420
rect 213 577 247 611
rect 433 519 467 553
rect 613 513 647 547
rect 699 529 733 563
rect 699 461 733 495
<< poly >>
rect 86 619 116 645
rect 172 619 202 645
rect 320 577 350 603
rect 392 577 422 603
rect 478 577 508 603
rect 572 577 602 603
rect 658 577 688 603
rect 320 413 350 449
rect 284 397 350 413
rect 86 321 116 367
rect 172 321 202 367
rect 284 363 300 397
rect 334 363 350 397
rect 284 329 350 363
rect 86 305 236 321
rect 86 271 186 305
rect 220 271 236 305
rect 284 295 300 329
rect 334 295 350 329
rect 284 279 350 295
rect 392 309 422 449
rect 478 417 508 449
rect 464 401 530 417
rect 464 367 480 401
rect 514 367 530 401
rect 464 351 530 367
rect 572 370 602 449
rect 658 370 688 449
rect 572 354 688 370
rect 572 340 607 354
rect 580 320 607 340
rect 641 320 688 354
rect 392 292 499 309
rect 392 279 538 292
rect 86 255 236 271
rect 86 215 116 255
rect 172 215 202 255
rect 289 132 319 279
rect 469 276 538 279
rect 469 242 488 276
rect 522 242 538 276
rect 361 221 427 237
rect 361 187 377 221
rect 411 187 427 221
rect 361 171 427 187
rect 469 226 538 242
rect 580 286 688 320
rect 580 252 607 286
rect 641 252 688 286
rect 580 236 688 252
rect 361 132 391 171
rect 469 132 499 226
rect 580 184 610 236
rect 658 188 688 236
rect 541 154 610 184
rect 652 158 688 188
rect 541 132 571 154
rect 652 132 682 158
rect 86 21 116 47
rect 172 21 202 47
rect 289 22 319 48
rect 361 22 391 48
rect 469 22 499 48
rect 541 22 571 48
rect 652 22 682 48
<< polycont >>
rect 300 363 334 397
rect 186 271 220 305
rect 300 295 334 329
rect 480 367 514 401
rect 607 320 641 354
rect 488 242 522 276
rect 377 187 411 221
rect 607 252 641 286
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 25 607 82 649
rect 25 573 41 607
rect 75 573 82 607
rect 25 509 82 573
rect 25 475 41 509
rect 75 475 82 509
rect 25 413 82 475
rect 25 379 41 413
rect 75 379 82 413
rect 25 363 82 379
rect 116 599 161 615
rect 116 565 127 599
rect 197 611 263 649
rect 197 577 213 611
rect 247 577 263 611
rect 197 571 263 577
rect 116 505 161 565
rect 417 553 483 569
rect 417 537 433 553
rect 116 471 127 505
rect 116 420 161 471
rect 116 386 127 420
rect 116 370 161 386
rect 201 519 433 537
rect 467 519 483 553
rect 201 503 483 519
rect 597 547 663 649
rect 597 513 613 547
rect 647 513 663 547
rect 597 503 663 513
rect 697 563 749 579
rect 697 529 699 563
rect 733 529 749 563
rect 116 219 150 370
rect 201 321 235 503
rect 697 495 749 529
rect 697 469 699 495
rect 186 305 235 321
rect 220 271 235 305
rect 284 461 699 469
rect 733 461 749 495
rect 284 435 749 461
rect 284 397 350 435
rect 284 363 300 397
rect 334 363 350 397
rect 284 329 350 363
rect 284 295 300 329
rect 334 295 350 329
rect 284 279 350 295
rect 393 367 480 401
rect 514 367 530 401
rect 393 310 530 367
rect 591 354 655 370
rect 591 320 607 354
rect 641 320 655 354
rect 186 255 235 271
rect 25 203 82 219
rect 25 169 41 203
rect 75 169 82 203
rect 25 93 82 169
rect 25 59 41 93
rect 75 59 82 93
rect 25 17 82 59
rect 116 203 167 219
rect 116 169 127 203
rect 161 169 167 203
rect 116 101 167 169
rect 201 153 235 255
rect 393 237 427 310
rect 591 286 655 320
rect 361 221 427 237
rect 361 187 377 221
rect 411 187 427 221
rect 472 242 488 276
rect 522 242 547 276
rect 201 119 438 153
rect 116 67 127 101
rect 161 67 167 101
rect 386 109 438 119
rect 116 51 167 67
rect 209 81 275 85
rect 209 47 225 81
rect 259 47 275 81
rect 386 75 404 109
rect 472 94 547 242
rect 591 252 607 286
rect 641 252 655 286
rect 591 157 655 252
rect 581 107 647 123
rect 386 51 438 75
rect 581 73 597 107
rect 631 73 647 107
rect 209 17 275 47
rect 581 17 647 73
rect 689 105 749 435
rect 689 71 693 105
rect 727 71 749 105
rect 689 55 749 71
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1670976
string GDS_START 1663624
<< end >>
