magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 1258 241 2008 259
rect 34 49 2008 241
rect 0 0 2016 49
<< scnmos >>
rect 117 47 147 215
rect 203 47 233 215
rect 289 47 319 215
rect 375 47 405 215
rect 461 47 491 215
rect 547 47 577 215
rect 633 47 663 215
rect 719 47 749 215
rect 821 47 851 215
rect 907 47 937 215
rect 993 47 1023 215
rect 1087 47 1117 215
rect 1337 65 1367 233
rect 1455 65 1485 233
rect 1541 65 1571 233
rect 1696 65 1726 233
rect 1782 65 1812 233
rect 1868 65 1898 233
<< scpmoshvt >>
rect 110 367 140 619
rect 196 367 226 619
rect 282 367 312 619
rect 368 367 398 619
rect 454 367 484 619
rect 540 367 570 619
rect 626 367 656 619
rect 712 367 742 619
rect 821 367 851 619
rect 907 367 937 619
rect 1001 367 1031 619
rect 1087 367 1117 619
rect 1337 367 1367 619
rect 1423 367 1453 619
rect 1563 367 1593 619
rect 1649 367 1679 619
rect 1768 367 1798 619
rect 1906 367 1936 619
<< ndiff >>
rect 60 175 117 215
rect 60 141 72 175
rect 106 141 117 175
rect 60 89 117 141
rect 60 55 72 89
rect 106 55 117 89
rect 60 47 117 55
rect 147 203 203 215
rect 147 169 158 203
rect 192 169 203 203
rect 147 101 203 169
rect 147 67 158 101
rect 192 67 203 101
rect 147 47 203 67
rect 233 172 289 215
rect 233 138 244 172
rect 278 138 289 172
rect 233 89 289 138
rect 233 55 244 89
rect 278 55 289 89
rect 233 47 289 55
rect 319 203 375 215
rect 319 169 330 203
rect 364 169 375 203
rect 319 101 375 169
rect 319 67 330 101
rect 364 67 375 101
rect 319 47 375 67
rect 405 127 461 215
rect 405 93 416 127
rect 450 93 461 127
rect 405 47 461 93
rect 491 203 547 215
rect 491 169 502 203
rect 536 169 547 203
rect 491 101 547 169
rect 491 67 502 101
rect 536 67 547 101
rect 491 47 547 67
rect 577 171 633 215
rect 577 137 588 171
rect 622 137 633 171
rect 577 89 633 137
rect 577 55 588 89
rect 622 55 633 89
rect 577 47 633 55
rect 663 203 719 215
rect 663 169 674 203
rect 708 169 719 203
rect 663 101 719 169
rect 663 67 674 101
rect 708 67 719 101
rect 663 47 719 67
rect 749 157 821 215
rect 749 123 762 157
rect 796 123 821 157
rect 749 89 821 123
rect 749 55 762 89
rect 796 55 821 89
rect 749 47 821 55
rect 851 159 907 215
rect 851 125 862 159
rect 896 125 907 159
rect 851 91 907 125
rect 851 57 862 91
rect 896 57 907 91
rect 851 47 907 57
rect 937 171 993 215
rect 937 137 948 171
rect 982 137 993 171
rect 937 47 993 137
rect 1023 161 1087 215
rect 1023 127 1037 161
rect 1071 127 1087 161
rect 1023 93 1087 127
rect 1023 59 1037 93
rect 1071 59 1087 93
rect 1023 47 1087 59
rect 1117 167 1170 215
rect 1117 133 1128 167
rect 1162 133 1170 167
rect 1117 93 1170 133
rect 1117 59 1128 93
rect 1162 59 1170 93
rect 1284 179 1337 233
rect 1284 145 1292 179
rect 1326 145 1337 179
rect 1284 111 1337 145
rect 1284 77 1292 111
rect 1326 77 1337 111
rect 1284 65 1337 77
rect 1367 107 1455 233
rect 1367 73 1394 107
rect 1428 73 1455 107
rect 1367 65 1455 73
rect 1485 181 1541 233
rect 1485 147 1496 181
rect 1530 147 1541 181
rect 1485 107 1541 147
rect 1485 73 1496 107
rect 1530 73 1541 107
rect 1485 65 1541 73
rect 1571 135 1696 233
rect 1571 107 1651 135
rect 1571 73 1582 107
rect 1616 101 1651 107
rect 1685 101 1696 135
rect 1616 73 1696 101
rect 1571 65 1696 73
rect 1726 179 1782 233
rect 1726 145 1737 179
rect 1771 145 1782 179
rect 1726 111 1782 145
rect 1726 77 1737 111
rect 1771 77 1782 111
rect 1726 65 1782 77
rect 1812 225 1868 233
rect 1812 191 1823 225
rect 1857 191 1868 225
rect 1812 157 1868 191
rect 1812 123 1823 157
rect 1857 123 1868 157
rect 1812 65 1868 123
rect 1898 221 1982 233
rect 1898 187 1936 221
rect 1970 187 1982 221
rect 1898 111 1982 187
rect 1898 77 1936 111
rect 1970 77 1982 111
rect 1898 65 1982 77
rect 1117 47 1170 59
<< pdiff >>
rect 1475 630 1533 638
rect 1475 619 1487 630
rect 57 607 110 619
rect 57 573 65 607
rect 99 573 110 607
rect 57 530 110 573
rect 57 496 65 530
rect 99 496 110 530
rect 57 453 110 496
rect 57 419 65 453
rect 99 419 110 453
rect 57 367 110 419
rect 140 599 196 619
rect 140 565 151 599
rect 185 565 196 599
rect 140 508 196 565
rect 140 474 151 508
rect 185 474 196 508
rect 140 413 196 474
rect 140 379 151 413
rect 185 379 196 413
rect 140 367 196 379
rect 226 607 282 619
rect 226 573 237 607
rect 271 573 282 607
rect 226 530 282 573
rect 226 496 237 530
rect 271 496 282 530
rect 226 453 282 496
rect 226 419 237 453
rect 271 419 282 453
rect 226 367 282 419
rect 312 599 368 619
rect 312 565 323 599
rect 357 565 368 599
rect 312 508 368 565
rect 312 474 323 508
rect 357 474 368 508
rect 312 413 368 474
rect 312 379 323 413
rect 357 379 368 413
rect 312 367 368 379
rect 398 607 454 619
rect 398 573 409 607
rect 443 573 454 607
rect 398 504 454 573
rect 398 470 409 504
rect 443 470 454 504
rect 398 412 454 470
rect 398 378 409 412
rect 443 378 454 412
rect 398 367 454 378
rect 484 599 540 619
rect 484 565 495 599
rect 529 565 540 599
rect 484 508 540 565
rect 484 474 495 508
rect 529 474 540 508
rect 484 413 540 474
rect 484 379 495 413
rect 529 379 540 413
rect 484 367 540 379
rect 570 607 626 619
rect 570 573 581 607
rect 615 573 626 607
rect 570 539 626 573
rect 570 505 581 539
rect 615 505 626 539
rect 570 469 626 505
rect 570 435 581 469
rect 615 435 626 469
rect 570 367 626 435
rect 656 599 712 619
rect 656 565 667 599
rect 701 565 712 599
rect 656 508 712 565
rect 656 474 667 508
rect 701 474 712 508
rect 656 413 712 474
rect 656 379 667 413
rect 701 379 712 413
rect 656 367 712 379
rect 742 611 821 619
rect 742 577 753 611
rect 787 577 821 611
rect 742 543 821 577
rect 742 509 753 543
rect 787 509 821 543
rect 742 473 821 509
rect 742 439 753 473
rect 787 439 821 473
rect 742 367 821 439
rect 851 595 907 619
rect 851 561 862 595
rect 896 561 907 595
rect 851 527 907 561
rect 851 493 862 527
rect 896 493 907 527
rect 851 459 907 493
rect 851 425 862 459
rect 896 425 907 459
rect 851 367 907 425
rect 937 607 1001 619
rect 937 573 952 607
rect 986 573 1001 607
rect 937 516 1001 573
rect 937 482 952 516
rect 986 482 1001 516
rect 937 367 1001 482
rect 1031 599 1087 619
rect 1031 565 1042 599
rect 1076 565 1087 599
rect 1031 527 1087 565
rect 1031 493 1042 527
rect 1076 493 1087 527
rect 1031 459 1087 493
rect 1031 425 1042 459
rect 1076 425 1087 459
rect 1031 367 1087 425
rect 1117 607 1170 619
rect 1117 573 1128 607
rect 1162 573 1170 607
rect 1117 516 1170 573
rect 1117 482 1128 516
rect 1162 482 1170 516
rect 1117 367 1170 482
rect 1284 599 1337 619
rect 1284 565 1292 599
rect 1326 565 1337 599
rect 1284 529 1337 565
rect 1284 495 1292 529
rect 1326 495 1337 529
rect 1284 367 1337 495
rect 1367 587 1423 619
rect 1367 553 1378 587
rect 1412 553 1423 587
rect 1367 367 1423 553
rect 1453 596 1487 619
rect 1521 619 1533 630
rect 1521 596 1563 619
rect 1453 367 1563 596
rect 1593 576 1649 619
rect 1593 542 1604 576
rect 1638 542 1649 576
rect 1593 367 1649 542
rect 1679 611 1768 619
rect 1679 577 1706 611
rect 1740 577 1768 611
rect 1679 498 1768 577
rect 1679 464 1706 498
rect 1740 464 1768 498
rect 1679 367 1768 464
rect 1798 607 1906 619
rect 1798 573 1816 607
rect 1850 573 1906 607
rect 1798 539 1906 573
rect 1798 505 1861 539
rect 1895 505 1906 539
rect 1798 471 1906 505
rect 1798 437 1861 471
rect 1895 437 1906 471
rect 1798 367 1906 437
rect 1936 599 1989 619
rect 1936 565 1947 599
rect 1981 565 1989 599
rect 1936 508 1989 565
rect 1936 474 1947 508
rect 1981 474 1989 508
rect 1936 413 1989 474
rect 1936 379 1947 413
rect 1981 379 1989 413
rect 1936 367 1989 379
<< ndiffc >>
rect 72 141 106 175
rect 72 55 106 89
rect 158 169 192 203
rect 158 67 192 101
rect 244 138 278 172
rect 244 55 278 89
rect 330 169 364 203
rect 330 67 364 101
rect 416 93 450 127
rect 502 169 536 203
rect 502 67 536 101
rect 588 137 622 171
rect 588 55 622 89
rect 674 169 708 203
rect 674 67 708 101
rect 762 123 796 157
rect 762 55 796 89
rect 862 125 896 159
rect 862 57 896 91
rect 948 137 982 171
rect 1037 127 1071 161
rect 1037 59 1071 93
rect 1128 133 1162 167
rect 1128 59 1162 93
rect 1292 145 1326 179
rect 1292 77 1326 111
rect 1394 73 1428 107
rect 1496 147 1530 181
rect 1496 73 1530 107
rect 1582 73 1616 107
rect 1651 101 1685 135
rect 1737 145 1771 179
rect 1737 77 1771 111
rect 1823 191 1857 225
rect 1823 123 1857 157
rect 1936 187 1970 221
rect 1936 77 1970 111
<< pdiffc >>
rect 65 573 99 607
rect 65 496 99 530
rect 65 419 99 453
rect 151 565 185 599
rect 151 474 185 508
rect 151 379 185 413
rect 237 573 271 607
rect 237 496 271 530
rect 237 419 271 453
rect 323 565 357 599
rect 323 474 357 508
rect 323 379 357 413
rect 409 573 443 607
rect 409 470 443 504
rect 409 378 443 412
rect 495 565 529 599
rect 495 474 529 508
rect 495 379 529 413
rect 581 573 615 607
rect 581 505 615 539
rect 581 435 615 469
rect 667 565 701 599
rect 667 474 701 508
rect 667 379 701 413
rect 753 577 787 611
rect 753 509 787 543
rect 753 439 787 473
rect 862 561 896 595
rect 862 493 896 527
rect 862 425 896 459
rect 952 573 986 607
rect 952 482 986 516
rect 1042 565 1076 599
rect 1042 493 1076 527
rect 1042 425 1076 459
rect 1128 573 1162 607
rect 1128 482 1162 516
rect 1292 565 1326 599
rect 1292 495 1326 529
rect 1378 553 1412 587
rect 1487 596 1521 630
rect 1604 542 1638 576
rect 1706 577 1740 611
rect 1706 464 1740 498
rect 1816 573 1850 607
rect 1861 505 1895 539
rect 1861 437 1895 471
rect 1947 565 1981 599
rect 1947 474 1981 508
rect 1947 379 1981 413
<< poly >>
rect 110 619 140 645
rect 196 619 226 645
rect 282 619 312 645
rect 368 619 398 645
rect 454 619 484 645
rect 540 619 570 645
rect 626 619 656 645
rect 712 619 742 645
rect 821 619 851 645
rect 907 619 937 645
rect 1001 619 1031 645
rect 1087 619 1117 645
rect 1337 619 1367 645
rect 1423 619 1453 645
rect 1563 619 1593 645
rect 1649 619 1679 645
rect 1768 619 1798 645
rect 1906 619 1936 645
rect 110 329 140 367
rect 196 329 226 367
rect 282 329 312 367
rect 368 329 398 367
rect 110 313 405 329
rect 110 279 151 313
rect 185 279 219 313
rect 253 279 287 313
rect 321 279 355 313
rect 389 279 405 313
rect 110 263 405 279
rect 454 293 484 367
rect 540 329 570 367
rect 626 329 656 367
rect 712 329 742 367
rect 821 335 851 367
rect 540 313 757 329
rect 540 293 571 313
rect 454 279 571 293
rect 605 279 639 313
rect 673 279 707 313
rect 741 279 757 313
rect 454 263 757 279
rect 799 319 865 335
rect 799 285 815 319
rect 849 285 865 319
rect 799 269 865 285
rect 907 283 937 367
rect 1001 319 1031 367
rect 1087 335 1117 367
rect 1087 319 1154 335
rect 979 303 1045 319
rect 979 283 995 303
rect 907 269 995 283
rect 1029 269 1045 303
rect 117 215 147 263
rect 203 215 233 263
rect 289 215 319 263
rect 375 215 405 263
rect 461 215 491 263
rect 547 215 577 263
rect 633 215 663 263
rect 719 215 749 263
rect 821 215 851 269
rect 907 253 1045 269
rect 1087 285 1104 319
rect 1138 285 1154 319
rect 1337 285 1367 367
rect 1423 335 1453 367
rect 1563 335 1593 367
rect 1649 335 1679 367
rect 1087 269 1154 285
rect 1196 269 1367 285
rect 1409 319 1593 335
rect 1409 285 1425 319
rect 1459 305 1593 319
rect 1635 319 1701 335
rect 1459 285 1571 305
rect 1409 269 1571 285
rect 1635 285 1651 319
rect 1685 299 1701 319
rect 1768 331 1798 367
rect 1768 315 1834 331
rect 1685 285 1726 299
rect 1635 269 1726 285
rect 907 215 937 253
rect 993 215 1023 253
rect 1087 215 1117 269
rect 1196 235 1212 269
rect 1246 255 1367 269
rect 1246 235 1262 255
rect 1196 219 1262 235
rect 1337 233 1367 255
rect 1455 233 1485 269
rect 1541 233 1571 269
rect 1696 233 1726 269
rect 1768 281 1784 315
rect 1818 295 1834 315
rect 1906 295 1936 367
rect 1818 281 1936 295
rect 1768 265 1936 281
rect 1782 233 1812 265
rect 1868 233 1898 265
rect 117 21 147 47
rect 203 21 233 47
rect 289 21 319 47
rect 375 21 405 47
rect 461 21 491 47
rect 547 21 577 47
rect 633 21 663 47
rect 719 21 749 47
rect 821 21 851 47
rect 907 21 937 47
rect 993 21 1023 47
rect 1087 21 1117 47
rect 1337 39 1367 65
rect 1455 39 1485 65
rect 1541 39 1571 65
rect 1696 39 1726 65
rect 1782 39 1812 65
rect 1868 39 1898 65
<< polycont >>
rect 151 279 185 313
rect 219 279 253 313
rect 287 279 321 313
rect 355 279 389 313
rect 571 279 605 313
rect 639 279 673 313
rect 707 279 741 313
rect 815 285 849 319
rect 995 269 1029 303
rect 1104 285 1138 319
rect 1425 285 1459 319
rect 1651 285 1685 319
rect 1212 235 1246 269
rect 1784 281 1818 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 49 607 115 649
rect 49 573 65 607
rect 99 573 115 607
rect 49 530 115 573
rect 49 496 65 530
rect 99 496 115 530
rect 49 453 115 496
rect 49 419 65 453
rect 99 419 115 453
rect 149 599 187 615
rect 149 565 151 599
rect 185 565 187 599
rect 149 508 187 565
rect 149 474 151 508
rect 185 474 187 508
rect 149 413 187 474
rect 221 607 287 649
rect 221 573 237 607
rect 271 573 287 607
rect 221 530 287 573
rect 221 496 237 530
rect 271 496 287 530
rect 221 453 287 496
rect 221 419 237 453
rect 271 419 287 453
rect 321 599 366 615
rect 321 565 323 599
rect 357 565 366 599
rect 321 508 366 565
rect 321 474 323 508
rect 357 474 366 508
rect 149 385 151 413
rect 18 379 151 385
rect 185 385 187 413
rect 321 413 366 474
rect 321 385 323 413
rect 185 379 323 385
rect 357 379 366 413
rect 18 351 366 379
rect 400 607 451 649
rect 400 573 409 607
rect 443 573 451 607
rect 400 504 451 573
rect 400 470 409 504
rect 443 470 451 504
rect 400 412 451 470
rect 400 378 409 412
rect 443 378 451 412
rect 400 362 451 378
rect 485 599 545 615
rect 485 565 495 599
rect 529 565 545 599
rect 485 508 545 565
rect 485 474 495 508
rect 529 474 545 508
rect 485 413 545 474
rect 579 607 622 649
rect 579 573 581 607
rect 615 573 622 607
rect 579 539 622 573
rect 579 505 581 539
rect 615 505 622 539
rect 579 469 622 505
rect 579 435 581 469
rect 615 435 622 469
rect 579 419 622 435
rect 656 599 703 615
rect 656 565 667 599
rect 701 565 703 599
rect 656 508 703 565
rect 656 474 667 508
rect 701 474 703 508
rect 485 379 495 413
rect 529 385 545 413
rect 656 413 703 474
rect 737 611 803 649
rect 737 577 753 611
rect 787 577 803 611
rect 737 543 803 577
rect 737 509 753 543
rect 787 509 803 543
rect 737 473 803 509
rect 737 439 753 473
rect 787 439 803 473
rect 839 595 902 611
rect 839 561 862 595
rect 896 561 902 595
rect 839 527 902 561
rect 839 493 862 527
rect 896 493 902 527
rect 839 459 902 493
rect 936 607 1002 649
rect 936 573 952 607
rect 986 573 1002 607
rect 936 516 1002 573
rect 936 482 952 516
rect 986 482 1002 516
rect 936 477 1002 482
rect 1036 599 1078 615
rect 1036 565 1042 599
rect 1076 565 1078 599
rect 1036 527 1078 565
rect 1036 493 1042 527
rect 1076 493 1078 527
rect 656 385 667 413
rect 529 379 667 385
rect 701 379 703 413
rect 839 425 862 459
rect 896 443 902 459
rect 1036 459 1078 493
rect 1112 607 1178 649
rect 1468 630 1537 649
rect 1112 573 1128 607
rect 1162 573 1178 607
rect 1112 516 1178 573
rect 1112 482 1128 516
rect 1162 482 1178 516
rect 1112 477 1178 482
rect 1276 599 1328 615
rect 1276 565 1292 599
rect 1326 565 1328 599
rect 1468 596 1487 630
rect 1521 596 1537 630
rect 1276 529 1328 565
rect 1362 587 1434 591
rect 1468 590 1537 596
rect 1690 611 1756 615
rect 1362 553 1378 587
rect 1412 556 1434 587
rect 1588 576 1654 592
rect 1588 556 1604 576
rect 1412 553 1604 556
rect 1362 549 1604 553
rect 1276 495 1292 529
rect 1326 513 1328 529
rect 1400 542 1604 549
rect 1638 542 1654 576
rect 1400 522 1654 542
rect 1690 577 1706 611
rect 1740 577 1756 611
rect 1326 495 1364 513
rect 1276 488 1364 495
rect 1690 498 1756 577
rect 1790 607 1904 649
rect 1790 573 1816 607
rect 1850 573 1904 607
rect 1790 539 1904 573
rect 1790 526 1861 539
rect 1690 488 1706 498
rect 1276 479 1706 488
rect 1036 443 1042 459
rect 896 425 1042 443
rect 1076 443 1078 459
rect 1330 464 1706 479
rect 1740 490 1756 498
rect 1859 505 1861 526
rect 1895 505 1904 539
rect 1740 464 1825 490
rect 1330 454 1825 464
rect 1076 425 1294 443
rect 839 420 1294 425
rect 839 409 1755 420
rect 839 405 873 409
rect 485 351 703 379
rect 744 371 873 405
rect 1260 386 1755 409
rect 18 243 81 351
rect 135 279 151 313
rect 185 279 219 313
rect 253 279 287 313
rect 321 279 355 313
rect 389 279 449 313
rect 18 209 366 243
rect 156 203 194 209
rect 56 141 72 175
rect 106 141 122 175
rect 56 89 122 141
rect 56 55 72 89
rect 106 55 122 89
rect 56 17 122 55
rect 156 169 158 203
rect 192 169 194 203
rect 328 203 366 209
rect 156 101 194 169
rect 156 67 158 101
rect 192 67 194 101
rect 156 51 194 67
rect 228 172 294 173
rect 228 138 244 172
rect 278 138 294 172
rect 228 89 294 138
rect 228 55 244 89
rect 278 55 294 89
rect 228 17 294 55
rect 328 169 330 203
rect 364 169 366 203
rect 328 101 366 169
rect 415 202 449 279
rect 485 243 519 351
rect 744 313 778 371
rect 909 350 1224 375
rect 909 339 1475 350
rect 909 335 943 339
rect 555 279 571 313
rect 605 279 639 313
rect 673 279 707 313
rect 741 279 778 313
rect 485 209 710 243
rect 500 203 538 209
rect 500 169 502 203
rect 536 169 538 203
rect 672 203 710 209
rect 328 67 330 101
rect 364 67 366 101
rect 328 51 366 67
rect 400 127 466 134
rect 400 93 416 127
rect 450 93 466 127
rect 400 17 466 93
rect 500 101 538 169
rect 500 67 502 101
rect 536 67 538 101
rect 500 51 538 67
rect 572 171 638 173
rect 572 137 588 171
rect 622 137 638 171
rect 572 89 638 137
rect 572 55 588 89
rect 622 55 638 89
rect 572 17 638 55
rect 672 169 674 203
rect 708 169 710 203
rect 744 233 778 279
rect 815 319 943 335
rect 849 285 943 319
rect 1088 319 1475 339
rect 815 269 943 285
rect 979 269 995 303
rect 1029 269 1052 303
rect 1088 285 1104 319
rect 1138 316 1425 319
rect 1138 285 1154 316
rect 1375 285 1425 316
rect 1459 285 1475 319
rect 1567 319 1685 350
rect 1567 303 1651 319
rect 1511 285 1651 303
rect 1511 269 1685 285
rect 1721 315 1755 386
rect 1791 385 1825 454
rect 1859 471 1904 505
rect 1859 437 1861 471
rect 1895 437 1904 471
rect 1859 421 1904 437
rect 1938 599 1997 615
rect 1938 565 1947 599
rect 1981 565 1997 599
rect 1938 508 1997 565
rect 1938 474 1947 508
rect 1981 474 1997 508
rect 1938 413 1997 474
rect 1938 385 1947 413
rect 1791 379 1947 385
rect 1981 379 1997 413
rect 1791 351 1997 379
rect 1721 281 1784 315
rect 1818 281 1834 315
rect 1018 251 1052 269
rect 1196 251 1212 269
rect 1018 235 1212 251
rect 1246 251 1262 269
rect 1511 251 1545 269
rect 1246 235 1545 251
rect 744 199 984 233
rect 1018 217 1545 235
rect 1868 229 1902 351
rect 1807 225 1902 229
rect 672 101 710 169
rect 946 171 984 199
rect 1581 185 1771 219
rect 1581 183 1615 185
rect 672 67 674 101
rect 708 67 710 101
rect 672 51 710 67
rect 744 157 812 161
rect 744 123 762 157
rect 796 123 812 157
rect 744 89 812 123
rect 744 55 762 89
rect 796 55 812 89
rect 744 17 812 55
rect 846 159 912 163
rect 846 125 862 159
rect 896 125 912 159
rect 846 91 912 125
rect 946 137 948 171
rect 982 137 984 171
rect 1121 167 1178 183
rect 946 121 984 137
rect 1021 161 1087 165
rect 1021 127 1037 161
rect 1071 127 1087 161
rect 846 57 862 91
rect 896 87 912 91
rect 1021 93 1087 127
rect 1021 87 1037 93
rect 896 59 1037 87
rect 1071 59 1087 93
rect 896 57 1087 59
rect 846 53 1087 57
rect 1121 133 1128 167
rect 1162 133 1178 167
rect 1121 93 1178 133
rect 1121 59 1128 93
rect 1162 59 1178 93
rect 1276 181 1615 183
rect 1276 179 1496 181
rect 1276 145 1292 179
rect 1326 147 1496 179
rect 1530 147 1615 181
rect 1733 179 1771 185
rect 1326 145 1532 147
rect 1276 111 1342 145
rect 1276 77 1292 111
rect 1326 77 1342 111
rect 1480 107 1532 145
rect 1649 135 1689 151
rect 1649 113 1651 135
rect 1276 73 1342 77
rect 1378 73 1394 107
rect 1428 73 1444 107
rect 1121 17 1178 59
rect 1378 17 1444 73
rect 1480 73 1496 107
rect 1530 73 1532 107
rect 1480 57 1532 73
rect 1566 107 1651 113
rect 1566 73 1582 107
rect 1616 101 1651 107
rect 1685 101 1689 135
rect 1616 73 1689 101
rect 1566 17 1689 73
rect 1733 145 1737 179
rect 1733 111 1771 145
rect 1807 191 1823 225
rect 1857 202 1902 225
rect 1807 168 1855 191
rect 1889 168 1902 202
rect 1807 157 1902 168
rect 1807 123 1823 157
rect 1857 123 1902 157
rect 1936 221 1986 237
rect 1970 187 1986 221
rect 1733 77 1737 111
rect 1936 111 1986 187
rect 1771 77 1936 87
rect 1970 77 1986 111
rect 1733 53 1986 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 415 168 449 202
rect 1855 191 1857 202
rect 1857 191 1889 202
rect 1855 168 1889 191
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 403 202 461 208
rect 403 168 415 202
rect 449 199 461 202
rect 1843 202 1901 208
rect 1843 199 1855 202
rect 449 171 1855 199
rect 449 168 461 171
rect 403 162 461 168
rect 1843 168 1855 171
rect 1889 168 1901 202
rect 1843 162 1901 168
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ha_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6694812
string GDS_START 6678586
<< end >>
