magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 23 49 733 157
rect 0 0 768 49
<< scnmos >>
rect 102 47 132 131
rect 216 47 246 131
rect 288 47 318 131
rect 444 47 474 131
rect 516 47 546 131
rect 624 47 654 131
<< scpmoshvt >>
rect 96 484 126 612
rect 186 484 216 612
rect 272 484 302 612
rect 466 429 496 557
rect 552 429 582 557
rect 652 429 682 557
<< ndiff >>
rect 49 106 102 131
rect 49 72 57 106
rect 91 72 102 106
rect 49 47 102 72
rect 132 95 216 131
rect 132 61 156 95
rect 190 61 216 95
rect 132 47 216 61
rect 246 47 288 131
rect 318 106 444 131
rect 318 72 329 106
rect 363 72 399 106
rect 433 72 444 106
rect 318 47 444 72
rect 474 47 516 131
rect 546 89 624 131
rect 546 55 572 89
rect 606 55 624 89
rect 546 47 624 55
rect 654 106 707 131
rect 654 72 665 106
rect 699 72 707 106
rect 654 47 707 72
<< pdiff >>
rect 43 599 96 612
rect 43 565 51 599
rect 85 565 96 599
rect 43 530 96 565
rect 43 496 51 530
rect 85 496 96 530
rect 43 484 96 496
rect 126 600 186 612
rect 126 566 141 600
rect 175 566 186 600
rect 126 530 186 566
rect 126 496 141 530
rect 175 496 186 530
rect 126 484 186 496
rect 216 599 272 612
rect 216 565 227 599
rect 261 565 272 599
rect 216 526 272 565
rect 216 492 227 526
rect 261 492 272 526
rect 216 484 272 492
rect 302 600 355 612
rect 302 566 313 600
rect 347 566 355 600
rect 302 530 355 566
rect 302 496 313 530
rect 347 496 355 530
rect 302 484 355 496
rect 409 545 466 557
rect 409 511 417 545
rect 451 511 466 545
rect 409 477 466 511
rect 409 443 417 477
rect 451 443 466 477
rect 409 429 466 443
rect 496 545 552 557
rect 496 511 507 545
rect 541 511 552 545
rect 496 471 552 511
rect 496 437 507 471
rect 541 437 552 471
rect 496 429 552 437
rect 582 545 652 557
rect 582 511 607 545
rect 641 511 652 545
rect 582 477 652 511
rect 582 443 607 477
rect 641 443 652 477
rect 582 429 652 443
rect 682 543 735 557
rect 682 509 693 543
rect 727 509 735 543
rect 682 475 735 509
rect 682 441 693 475
rect 727 441 735 475
rect 682 429 735 441
<< ndiffc >>
rect 57 72 91 106
rect 156 61 190 95
rect 329 72 363 106
rect 399 72 433 106
rect 572 55 606 89
rect 665 72 699 106
<< pdiffc >>
rect 51 565 85 599
rect 51 496 85 530
rect 141 566 175 600
rect 141 496 175 530
rect 227 565 261 599
rect 227 492 261 526
rect 313 566 347 600
rect 313 496 347 530
rect 417 511 451 545
rect 417 443 451 477
rect 507 511 541 545
rect 507 437 541 471
rect 607 511 641 545
rect 607 443 641 477
rect 693 509 727 543
rect 693 441 727 475
<< poly >>
rect 96 612 126 638
rect 186 612 216 638
rect 272 612 302 638
rect 466 557 496 583
rect 552 557 582 583
rect 652 557 682 583
rect 96 446 126 484
rect 72 430 138 446
rect 72 396 88 430
rect 122 396 138 430
rect 72 362 138 396
rect 72 328 88 362
rect 122 328 138 362
rect 186 333 216 484
rect 272 411 302 484
rect 272 381 318 411
rect 72 312 138 328
rect 180 317 246 333
rect 102 131 132 312
rect 180 283 196 317
rect 230 283 246 317
rect 180 249 246 283
rect 180 215 196 249
rect 230 215 246 249
rect 180 199 246 215
rect 216 131 246 199
rect 288 321 318 381
rect 466 354 496 429
rect 438 324 496 354
rect 288 305 360 321
rect 288 271 310 305
rect 344 271 360 305
rect 438 302 474 324
rect 288 237 360 271
rect 288 203 310 237
rect 344 203 360 237
rect 288 187 360 203
rect 402 286 474 302
rect 402 252 418 286
rect 452 252 474 286
rect 552 276 582 429
rect 652 333 682 429
rect 402 218 474 252
rect 288 131 318 187
rect 402 184 418 218
rect 452 184 474 218
rect 402 168 474 184
rect 444 131 474 168
rect 516 260 582 276
rect 516 226 532 260
rect 566 226 582 260
rect 516 210 582 226
rect 624 317 722 333
rect 624 283 672 317
rect 706 283 722 317
rect 624 249 722 283
rect 624 215 672 249
rect 706 215 722 249
rect 516 131 546 210
rect 624 199 722 215
rect 624 131 654 199
rect 102 21 132 47
rect 216 21 246 47
rect 288 21 318 47
rect 444 21 474 47
rect 516 21 546 47
rect 624 21 654 47
<< polycont >>
rect 88 396 122 430
rect 88 328 122 362
rect 196 283 230 317
rect 196 215 230 249
rect 310 271 344 305
rect 310 203 344 237
rect 418 252 452 286
rect 418 184 452 218
rect 532 226 566 260
rect 672 283 706 317
rect 672 215 706 249
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 18 599 95 615
rect 18 565 51 599
rect 85 565 95 599
rect 18 530 95 565
rect 18 496 51 530
rect 85 496 95 530
rect 18 480 95 496
rect 129 600 185 649
rect 129 566 141 600
rect 175 566 185 600
rect 129 530 185 566
rect 129 496 141 530
rect 175 496 185 530
rect 129 480 185 496
rect 219 599 270 615
rect 219 565 227 599
rect 261 565 270 599
rect 219 526 270 565
rect 219 492 227 526
rect 261 492 270 526
rect 18 278 54 480
rect 88 430 135 446
rect 122 396 135 430
rect 88 362 135 396
rect 122 328 135 362
rect 219 391 270 492
rect 304 600 363 649
rect 304 566 313 600
rect 347 566 363 600
rect 304 530 363 566
rect 304 496 313 530
rect 347 496 363 530
rect 304 480 363 496
rect 401 581 657 615
rect 401 545 457 581
rect 401 511 417 545
rect 451 511 457 545
rect 401 477 457 511
rect 401 443 417 477
rect 451 443 457 477
rect 401 427 457 443
rect 491 545 557 547
rect 491 511 507 545
rect 541 511 557 545
rect 491 471 557 511
rect 491 437 507 471
rect 541 437 557 471
rect 591 545 657 581
rect 591 511 607 545
rect 641 511 657 545
rect 591 477 657 511
rect 591 443 607 477
rect 641 443 657 477
rect 591 437 657 443
rect 691 543 743 559
rect 691 509 693 543
rect 727 509 743 543
rect 691 475 743 509
rect 691 441 693 475
rect 727 441 743 475
rect 491 391 557 437
rect 691 403 743 441
rect 219 357 557 391
rect 602 369 743 403
rect 88 312 135 328
rect 18 111 67 278
rect 101 179 135 312
rect 180 317 272 323
rect 180 283 196 317
rect 230 283 272 317
rect 180 249 272 283
rect 180 215 196 249
rect 230 215 272 249
rect 180 213 272 215
rect 308 305 369 321
rect 308 271 310 305
rect 344 271 369 305
rect 308 237 369 271
rect 308 203 310 237
rect 344 203 369 237
rect 101 145 274 179
rect 308 168 369 203
rect 403 286 454 302
rect 403 252 418 286
rect 452 252 454 286
rect 403 218 454 252
rect 403 184 418 218
rect 452 184 454 218
rect 499 260 568 317
rect 499 226 532 260
rect 566 226 568 260
rect 499 210 568 226
rect 403 168 454 184
rect 602 163 638 369
rect 672 317 751 333
rect 706 283 751 317
rect 672 249 751 283
rect 706 215 751 249
rect 672 199 751 215
rect 240 122 274 145
rect 488 129 715 163
rect 488 122 522 129
rect 18 106 107 111
rect 18 72 57 106
rect 91 72 107 106
rect 18 56 107 72
rect 143 95 206 111
rect 143 61 156 95
rect 190 61 206 95
rect 143 17 206 61
rect 240 106 522 122
rect 240 72 329 106
rect 363 72 399 106
rect 433 72 522 106
rect 656 106 715 129
rect 240 56 522 72
rect 556 89 622 95
rect 556 55 572 89
rect 606 55 622 89
rect 656 72 665 106
rect 699 72 715 106
rect 656 56 715 72
rect 556 17 622 55
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a221o_0
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6141998
string GDS_START 6134276
<< end >>
