magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3506 1975
<< nwell >>
rect -38 335 2246 704
rect -38 332 622 335
rect 1384 332 2246 335
rect 258 311 622 332
<< pwell >>
rect 279 229 597 248
rect 1072 229 1342 293
rect 2010 230 2207 268
rect 1908 229 2207 230
rect 279 184 2207 229
rect 7 49 2207 184
rect 0 0 2208 49
<< scpmos >>
rect 82 508 118 592
rect 172 508 208 592
rect 365 347 401 547
rect 482 347 518 547
rect 694 457 730 541
rect 784 457 820 541
rect 862 457 898 541
rect 964 457 1000 541
rect 1158 392 1194 592
rect 1344 392 1380 592
rect 1514 508 1550 592
rect 1598 508 1634 592
rect 1706 508 1742 592
rect 1796 508 1832 592
rect 1990 424 2026 592
rect 2091 368 2127 592
<< nmoslvt >>
rect 90 74 120 158
rect 168 74 198 158
rect 371 74 401 222
rect 480 74 510 222
rect 684 119 714 203
rect 820 119 850 203
rect 892 119 922 203
rect 964 119 994 203
rect 1148 119 1178 267
rect 1236 119 1266 267
rect 1520 119 1550 203
rect 1598 119 1628 203
rect 1706 119 1736 203
rect 1784 119 1814 203
rect 1991 94 2021 204
rect 2093 94 2123 242
<< ndiff >>
rect 305 202 371 222
rect 305 168 322 202
rect 356 168 371 202
rect 33 131 90 158
rect 33 97 45 131
rect 79 97 90 131
rect 33 74 90 97
rect 120 74 168 158
rect 198 133 251 158
rect 198 99 209 133
rect 243 99 251 133
rect 198 74 251 99
rect 305 129 371 168
rect 305 95 322 129
rect 356 95 371 129
rect 305 74 371 95
rect 401 124 480 222
rect 401 90 423 124
rect 457 90 480 124
rect 401 74 480 90
rect 510 202 571 222
rect 510 168 529 202
rect 563 168 571 202
rect 510 129 571 168
rect 510 95 529 129
rect 563 95 571 129
rect 510 74 571 95
rect 1098 203 1148 267
rect 631 177 684 203
rect 631 143 639 177
rect 673 143 684 177
rect 631 119 684 143
rect 714 188 820 203
rect 714 154 775 188
rect 809 154 820 188
rect 714 119 820 154
rect 850 119 892 203
rect 922 119 964 203
rect 994 124 1148 203
rect 994 119 1021 124
rect 1009 90 1021 119
rect 1055 119 1148 124
rect 1178 244 1236 267
rect 1178 210 1189 244
rect 1223 210 1236 244
rect 1178 169 1236 210
rect 1178 135 1189 169
rect 1223 135 1236 169
rect 1178 119 1236 135
rect 1266 203 1316 267
rect 2036 210 2093 242
rect 2036 204 2048 210
rect 1266 175 1520 203
rect 1266 141 1341 175
rect 1375 141 1475 175
rect 1509 141 1520 175
rect 1266 119 1520 141
rect 1550 119 1598 203
rect 1628 165 1706 203
rect 1628 131 1650 165
rect 1684 131 1706 165
rect 1628 119 1706 131
rect 1736 119 1784 203
rect 1814 170 1871 203
rect 1814 136 1825 170
rect 1859 136 1871 170
rect 1814 119 1871 136
rect 1934 166 1991 204
rect 1934 132 1946 166
rect 1980 132 1991 166
rect 1055 90 1067 119
rect 1009 78 1067 90
rect 1934 94 1991 132
rect 2021 176 2048 204
rect 2082 176 2093 210
rect 2021 138 2093 176
rect 2021 104 2048 138
rect 2082 104 2093 138
rect 2021 94 2093 104
rect 2123 214 2181 242
rect 2123 180 2134 214
rect 2168 180 2181 214
rect 2123 138 2181 180
rect 2123 104 2134 138
rect 2168 104 2181 138
rect 2123 94 2181 104
<< pdiff >>
rect 27 567 82 592
rect 27 533 38 567
rect 72 533 82 567
rect 27 508 82 533
rect 118 567 172 592
rect 118 533 128 567
rect 162 533 172 567
rect 118 508 172 533
rect 208 567 261 592
rect 208 533 219 567
rect 253 533 261 567
rect 416 547 467 560
rect 208 508 261 533
rect 315 469 365 547
rect 300 400 365 469
rect 300 366 319 400
rect 353 366 365 400
rect 300 347 365 366
rect 401 544 482 547
rect 401 510 425 544
rect 459 510 482 544
rect 401 347 482 510
rect 518 400 571 547
rect 1106 580 1158 592
rect 1106 546 1114 580
rect 1148 546 1158 580
rect 638 516 694 541
rect 638 482 650 516
rect 684 482 694 516
rect 638 457 694 482
rect 730 516 784 541
rect 730 482 740 516
rect 774 482 784 516
rect 730 457 784 482
rect 820 457 862 541
rect 898 516 964 541
rect 898 482 914 516
rect 948 482 964 516
rect 898 457 964 482
rect 1000 516 1052 541
rect 1000 482 1010 516
rect 1044 482 1052 516
rect 1000 457 1052 482
rect 1106 506 1158 546
rect 1106 472 1114 506
rect 1148 472 1158 506
rect 518 366 529 400
rect 563 366 571 400
rect 518 347 571 366
rect 1106 392 1158 472
rect 1194 580 1344 592
rect 1194 546 1205 580
rect 1239 546 1299 580
rect 1333 546 1344 580
rect 1194 512 1344 546
rect 1194 478 1205 512
rect 1239 478 1299 512
rect 1333 478 1344 512
rect 1194 444 1344 478
rect 1194 410 1205 444
rect 1239 410 1299 444
rect 1333 410 1344 444
rect 1194 392 1344 410
rect 1380 557 1514 592
rect 1380 523 1390 557
rect 1424 523 1470 557
rect 1504 523 1514 557
rect 1380 508 1514 523
rect 1550 508 1598 592
rect 1634 567 1706 592
rect 1634 533 1644 567
rect 1678 533 1706 567
rect 1634 508 1706 533
rect 1742 567 1796 592
rect 1742 533 1752 567
rect 1786 533 1796 567
rect 1742 508 1796 533
rect 1832 567 1884 592
rect 1832 533 1842 567
rect 1876 533 1884 567
rect 1832 508 1884 533
rect 1938 580 1990 592
rect 1938 546 1946 580
rect 1980 546 1990 580
rect 1380 392 1430 508
rect 1938 471 1990 546
rect 1938 437 1946 471
rect 1980 437 1990 471
rect 1938 424 1990 437
rect 2026 580 2091 592
rect 2026 546 2046 580
rect 2080 546 2091 580
rect 2026 470 2091 546
rect 2026 436 2046 470
rect 2080 436 2091 470
rect 2026 424 2091 436
rect 2041 368 2091 424
rect 2127 580 2181 592
rect 2127 546 2137 580
rect 2171 546 2181 580
rect 2127 497 2181 546
rect 2127 463 2137 497
rect 2171 463 2181 497
rect 2127 414 2181 463
rect 2127 380 2137 414
rect 2171 380 2181 414
rect 2127 368 2181 380
<< ndiffc >>
rect 322 168 356 202
rect 45 97 79 131
rect 209 99 243 133
rect 322 95 356 129
rect 423 90 457 124
rect 529 168 563 202
rect 529 95 563 129
rect 639 143 673 177
rect 775 154 809 188
rect 1021 90 1055 124
rect 1189 210 1223 244
rect 1189 135 1223 169
rect 1341 141 1375 175
rect 1475 141 1509 175
rect 1650 131 1684 165
rect 1825 136 1859 170
rect 1946 132 1980 166
rect 2048 176 2082 210
rect 2048 104 2082 138
rect 2134 180 2168 214
rect 2134 104 2168 138
<< pdiffc >>
rect 38 533 72 567
rect 128 533 162 567
rect 219 533 253 567
rect 319 366 353 400
rect 425 510 459 544
rect 1114 546 1148 580
rect 650 482 684 516
rect 740 482 774 516
rect 914 482 948 516
rect 1010 482 1044 516
rect 1114 472 1148 506
rect 529 366 563 400
rect 1205 546 1239 580
rect 1299 546 1333 580
rect 1205 478 1239 512
rect 1299 478 1333 512
rect 1205 410 1239 444
rect 1299 410 1333 444
rect 1390 523 1424 557
rect 1470 523 1504 557
rect 1644 533 1678 567
rect 1752 533 1786 567
rect 1842 533 1876 567
rect 1946 546 1980 580
rect 1946 437 1980 471
rect 2046 546 2080 580
rect 2046 436 2080 470
rect 2137 546 2171 580
rect 2137 463 2171 497
rect 2137 380 2171 414
<< poly >>
rect 82 592 118 618
rect 172 615 1000 645
rect 172 592 208 615
rect 365 547 401 573
rect 482 547 518 573
rect 82 414 118 508
rect 57 384 118 414
rect 57 326 87 384
rect 172 336 208 508
rect 694 541 730 567
rect 784 541 820 567
rect 862 541 898 567
rect 964 541 1000 615
rect 1158 592 1194 618
rect 1344 592 1380 618
rect 1514 592 1550 618
rect 1598 592 1634 618
rect 1706 592 1742 618
rect 1796 592 1832 618
rect 1990 592 2026 618
rect 2091 592 2127 618
rect 694 387 730 457
rect 586 357 730 387
rect 784 404 820 457
rect 21 310 87 326
rect 21 276 37 310
rect 71 276 87 310
rect 21 242 87 276
rect 160 320 226 336
rect 365 332 401 347
rect 482 332 518 347
rect 586 332 616 357
rect 160 286 176 320
rect 210 286 226 320
rect 160 270 226 286
rect 270 299 401 332
rect 21 208 37 242
rect 71 222 87 242
rect 71 208 120 222
rect 21 192 120 208
rect 90 158 120 192
rect 168 158 198 270
rect 270 265 305 299
rect 339 265 401 299
rect 270 242 401 265
rect 451 299 616 332
rect 784 315 814 404
rect 862 360 898 457
rect 964 360 1000 457
rect 1514 473 1550 508
rect 1462 457 1544 473
rect 1462 423 1478 457
rect 1512 423 1544 457
rect 1158 360 1194 392
rect 451 265 467 299
rect 501 265 616 299
rect 451 242 616 265
rect 371 222 401 242
rect 480 222 510 242
rect 90 48 120 74
rect 168 48 198 74
rect 371 48 401 74
rect 480 48 510 74
rect 586 51 616 242
rect 684 299 814 315
rect 684 265 707 299
rect 741 279 814 299
rect 856 344 922 360
rect 856 310 872 344
rect 906 310 922 344
rect 856 294 922 310
rect 741 265 757 279
rect 684 249 757 265
rect 684 203 714 249
rect 820 203 850 237
rect 892 203 922 294
rect 964 344 1030 360
rect 964 310 980 344
rect 1014 310 1030 344
rect 964 294 1030 310
rect 1073 344 1194 360
rect 1073 310 1089 344
rect 1123 310 1194 344
rect 1073 294 1194 310
rect 1236 344 1302 360
rect 1236 310 1252 344
rect 1286 310 1302 344
rect 1236 294 1302 310
rect 964 203 994 294
rect 1148 267 1178 294
rect 1236 267 1266 294
rect 1344 291 1380 392
rect 1462 389 1544 423
rect 1462 355 1478 389
rect 1512 355 1544 389
rect 1462 339 1544 355
rect 1598 467 1634 508
rect 1598 451 1664 467
rect 1598 417 1614 451
rect 1648 417 1664 451
rect 1598 401 1664 417
rect 1344 275 1484 291
rect 684 93 714 119
rect 820 51 850 119
rect 892 93 922 119
rect 964 93 994 119
rect 1344 261 1366 275
rect 1350 241 1366 261
rect 1400 241 1434 275
rect 1468 255 1484 275
rect 1468 241 1550 255
rect 1350 225 1550 241
rect 1520 203 1550 225
rect 1598 203 1628 401
rect 1706 359 1742 508
rect 1796 409 1832 508
rect 1990 409 2026 424
rect 1796 379 2026 409
rect 1796 359 1850 379
rect 1676 343 1742 359
rect 1676 309 1692 343
rect 1726 309 1742 343
rect 1676 293 1742 309
rect 1784 343 1850 359
rect 1784 309 1800 343
rect 1834 309 1850 343
rect 2091 330 2127 368
rect 1706 203 1736 293
rect 1784 275 1850 309
rect 1784 241 1800 275
rect 1834 255 1850 275
rect 2063 314 2129 330
rect 2063 280 2079 314
rect 2113 280 2129 314
rect 2063 264 2129 280
rect 1834 241 2021 255
rect 2093 242 2123 264
rect 1784 225 2021 241
rect 1784 203 1814 225
rect 1991 204 2021 225
rect 1148 93 1178 119
rect 1236 51 1266 119
rect 1520 93 1550 119
rect 1598 93 1628 119
rect 1706 93 1736 119
rect 1784 93 1814 119
rect 1991 68 2021 94
rect 2093 68 2123 94
rect 586 21 1266 51
<< polycont >>
rect 37 276 71 310
rect 176 286 210 320
rect 37 208 71 242
rect 305 265 339 299
rect 1478 423 1512 457
rect 467 265 501 299
rect 707 265 741 299
rect 872 310 906 344
rect 980 310 1014 344
rect 1089 310 1123 344
rect 1252 310 1286 344
rect 1478 355 1512 389
rect 1614 417 1648 451
rect 1366 241 1400 275
rect 1434 241 1468 275
rect 1692 309 1726 343
rect 1800 309 1834 343
rect 1800 241 1834 275
rect 2079 280 2113 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 22 567 88 649
rect 22 533 38 567
rect 72 533 88 567
rect 22 504 88 533
rect 128 567 178 596
rect 162 533 178 567
rect 128 476 178 533
rect 212 567 278 649
rect 212 533 219 567
rect 253 533 278 567
rect 212 510 278 533
rect 409 544 475 649
rect 409 510 425 544
rect 459 510 475 544
rect 634 516 688 541
rect 634 482 650 516
rect 684 482 688 516
rect 634 476 688 482
rect 128 470 688 476
rect 108 436 688 470
rect 724 516 811 541
rect 724 482 740 516
rect 774 482 811 516
rect 724 455 811 482
rect 898 516 964 649
rect 1098 580 1164 649
rect 1098 546 1114 580
rect 1148 546 1164 580
rect 898 482 914 516
rect 948 482 964 516
rect 898 472 964 482
rect 998 516 1060 541
rect 998 482 1010 516
rect 1044 482 1060 516
rect 21 310 74 430
rect 21 276 37 310
rect 71 276 74 310
rect 21 242 74 276
rect 21 208 37 242
rect 71 208 74 242
rect 21 192 74 208
rect 108 158 142 436
rect 303 400 479 402
rect 303 366 319 400
rect 353 366 479 400
rect 303 364 479 366
rect 176 350 257 356
rect 176 320 223 350
rect 210 316 223 320
rect 210 286 257 316
rect 429 315 479 364
rect 513 400 588 402
rect 513 366 529 400
rect 563 366 588 400
rect 513 349 588 366
rect 303 310 353 315
rect 176 270 257 286
rect 291 299 353 310
rect 291 265 305 299
rect 339 265 353 299
rect 291 236 353 265
rect 429 299 501 315
rect 429 265 467 299
rect 429 244 501 265
rect 429 202 495 244
rect 535 218 588 349
rect 306 168 322 202
rect 356 168 495 202
rect 306 162 495 168
rect 529 202 588 218
rect 563 168 588 202
rect 29 131 142 158
rect 29 97 45 131
rect 79 97 142 131
rect 29 70 142 97
rect 209 133 249 162
rect 243 99 249 133
rect 209 17 249 99
rect 306 129 373 162
rect 306 95 322 129
rect 356 95 373 129
rect 529 129 588 168
rect 306 79 373 95
rect 407 124 473 128
rect 407 90 423 124
rect 457 90 473 124
rect 407 17 473 90
rect 563 95 588 129
rect 623 368 688 436
rect 775 438 811 455
rect 998 438 1060 482
rect 1098 506 1164 546
rect 1098 472 1114 506
rect 1148 472 1164 506
rect 1198 580 1340 596
rect 1198 546 1205 580
rect 1239 546 1299 580
rect 1333 546 1340 580
rect 1198 512 1340 546
rect 1198 478 1205 512
rect 1239 478 1299 512
rect 1333 478 1340 512
rect 1374 557 1520 573
rect 1374 523 1390 557
rect 1424 523 1470 557
rect 1504 541 1520 557
rect 1628 567 1694 649
rect 1504 523 1580 541
rect 1374 507 1580 523
rect 1198 444 1340 478
rect 775 404 1139 438
rect 1198 428 1205 444
rect 623 177 673 368
rect 623 143 639 177
rect 623 127 673 143
rect 707 299 741 334
rect 529 93 588 95
rect 707 93 741 265
rect 775 215 811 404
rect 856 344 922 360
rect 856 310 872 344
rect 906 310 922 344
rect 856 294 922 310
rect 964 350 1031 360
rect 964 344 991 350
rect 964 310 980 344
rect 1025 316 1031 350
rect 1014 310 1031 316
rect 964 294 1031 310
rect 1073 344 1139 404
rect 1073 310 1089 344
rect 1123 310 1139 344
rect 1073 294 1139 310
rect 1173 410 1205 428
rect 1239 410 1299 444
rect 1333 410 1340 444
rect 1173 394 1340 410
rect 1462 457 1512 473
rect 1462 423 1478 457
rect 888 260 922 294
rect 1173 260 1207 394
rect 1462 389 1512 423
rect 1462 360 1478 389
rect 1241 355 1478 360
rect 1241 344 1512 355
rect 1241 310 1252 344
rect 1286 326 1512 344
rect 1286 310 1302 326
rect 1241 294 1302 310
rect 1350 275 1484 291
rect 888 244 1239 260
rect 1350 259 1366 275
rect 888 226 1189 244
rect 775 188 825 215
rect 1173 210 1189 226
rect 1223 210 1239 244
rect 809 154 825 188
rect 775 127 825 154
rect 859 158 1139 192
rect 859 93 893 158
rect 529 51 893 93
rect 1005 90 1021 124
rect 1055 90 1071 124
rect 1005 17 1071 90
rect 1105 85 1139 158
rect 1173 169 1239 210
rect 1173 135 1189 169
rect 1223 135 1239 169
rect 1173 119 1239 135
rect 1273 241 1366 259
rect 1400 241 1434 275
rect 1468 241 1484 275
rect 1273 225 1484 241
rect 1546 259 1580 507
rect 1628 533 1644 567
rect 1678 533 1694 567
rect 1628 504 1694 533
rect 1736 567 1802 596
rect 1736 533 1752 567
rect 1786 533 1802 567
rect 1736 467 1802 533
rect 1842 567 1892 649
rect 1876 533 1892 567
rect 1842 504 1892 533
rect 1930 580 1996 596
rect 1930 546 1946 580
rect 1980 546 1996 580
rect 1930 471 1996 546
rect 1614 451 1810 467
rect 1930 461 1946 471
rect 1648 427 1810 451
rect 1980 437 1996 471
rect 1648 417 1912 427
rect 1614 393 1912 417
rect 1657 350 1742 359
rect 1657 316 1663 350
rect 1697 343 1742 350
rect 1657 309 1692 316
rect 1726 309 1742 343
rect 1657 293 1742 309
rect 1784 343 1844 359
rect 1784 309 1800 343
rect 1834 309 1844 343
rect 1784 275 1844 309
rect 1784 259 1800 275
rect 1546 241 1800 259
rect 1834 241 1844 275
rect 1546 225 1844 241
rect 1273 85 1307 225
rect 1546 191 1580 225
rect 1878 191 1912 393
rect 1341 175 1580 191
rect 1375 141 1475 175
rect 1509 141 1580 175
rect 1341 125 1580 141
rect 1623 165 1711 181
rect 1623 131 1650 165
rect 1684 131 1711 165
rect 1105 51 1307 85
rect 1623 17 1711 131
rect 1809 170 1912 191
rect 1809 136 1825 170
rect 1859 136 1912 170
rect 1809 115 1912 136
rect 1946 330 1996 437
rect 2030 580 2080 649
rect 2030 546 2046 580
rect 2030 470 2080 546
rect 2030 436 2046 470
rect 2030 420 2080 436
rect 2121 580 2191 596
rect 2121 546 2137 580
rect 2171 546 2191 580
rect 2121 497 2191 546
rect 2121 463 2137 497
rect 2171 463 2191 497
rect 2121 414 2191 463
rect 2121 380 2137 414
rect 2171 380 2191 414
rect 2121 364 2191 380
rect 1946 314 2123 330
rect 1946 280 2079 314
rect 2113 280 2123 314
rect 1946 264 2123 280
rect 1946 166 1996 264
rect 2157 230 2191 364
rect 1980 132 1996 166
rect 1946 106 1996 132
rect 2032 210 2082 226
rect 2032 176 2048 210
rect 2032 138 2082 176
rect 2032 104 2048 138
rect 2032 17 2082 104
rect 2118 214 2191 230
rect 2118 180 2134 214
rect 2168 180 2191 214
rect 2118 138 2191 180
rect 2118 104 2134 138
rect 2168 104 2191 138
rect 2118 88 2191 104
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 223 316 257 350
rect 991 344 1025 350
rect 991 316 1014 344
rect 1014 316 1025 344
rect 1663 343 1697 350
rect 1663 316 1692 343
rect 1692 316 1697 343
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 211 350 269 356
rect 211 316 223 350
rect 257 347 269 350
rect 979 350 1037 356
rect 979 347 991 350
rect 257 319 991 347
rect 257 316 269 319
rect 211 310 269 316
rect 979 316 991 319
rect 1025 347 1037 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1025 319 1663 347
rect 1025 316 1037 319
rect 979 310 1037 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel comment s 892 36 892 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 557 630 557 630 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfrtn_1
flabel comment s 602 297 602 297 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 223 316 257 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 2143 390 2177 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2143 464 2177 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2143 538 2177 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y R90
string GDS_END 3332086
string GDS_START 3315210
<< end >>
