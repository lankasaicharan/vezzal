magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4370 1975
<< nwell >>
rect -38 331 3110 704
<< pwell >>
rect 1 49 543 230
rect 756 229 1034 273
rect 2184 250 2388 276
rect 2184 241 2684 250
rect 2184 232 3069 241
rect 1899 229 3069 232
rect 756 49 1297 229
rect 1475 49 3069 229
rect 0 0 3072 49
<< scnmos >>
rect 80 120 110 204
rect 152 120 182 204
rect 238 120 268 204
rect 332 120 362 204
rect 434 120 464 204
rect 835 119 865 247
rect 1030 119 1060 203
rect 1102 119 1132 203
rect 1188 119 1218 203
rect 1554 119 1584 203
rect 1640 119 1670 203
rect 1978 122 2008 206
rect 2067 122 2097 206
rect 2139 122 2169 206
rect 2279 122 2309 250
rect 2489 56 2519 224
rect 2575 56 2605 224
rect 2680 56 2710 140
rect 2874 47 2904 215
rect 2960 47 2990 215
<< scpmoshvt >>
rect 80 489 110 617
rect 174 489 204 617
rect 246 489 276 617
rect 332 489 362 617
rect 621 481 651 609
rect 858 425 888 593
rect 963 425 993 509
rect 1198 501 1228 585
rect 1284 501 1314 585
rect 1521 395 1551 523
rect 1639 395 1669 523
rect 1984 379 2014 547
rect 2086 463 2116 547
rect 2158 463 2188 547
rect 2273 379 2303 547
rect 2493 367 2523 619
rect 2579 367 2609 619
rect 2684 367 2714 495
rect 2874 367 2904 619
rect 2960 367 2990 619
<< ndiff >>
rect 27 179 80 204
rect 27 145 35 179
rect 69 145 80 179
rect 27 120 80 145
rect 110 120 152 204
rect 182 179 238 204
rect 182 145 193 179
rect 227 145 238 179
rect 182 120 238 145
rect 268 120 332 204
rect 362 167 434 204
rect 362 133 373 167
rect 407 133 434 167
rect 362 120 434 133
rect 464 166 517 204
rect 464 132 475 166
rect 509 132 517 166
rect 464 120 517 132
rect 782 235 835 247
rect 782 201 790 235
rect 824 201 835 235
rect 782 167 835 201
rect 782 133 790 167
rect 824 133 835 167
rect 782 119 835 133
rect 865 229 1008 247
rect 865 195 958 229
rect 992 203 1008 229
rect 2210 236 2279 250
rect 2210 206 2218 236
rect 992 195 1030 203
rect 865 161 1030 195
rect 865 127 958 161
rect 992 127 1030 161
rect 865 119 1030 127
rect 1060 119 1102 203
rect 1132 177 1188 203
rect 1132 143 1143 177
rect 1177 143 1188 177
rect 1132 119 1188 143
rect 1218 179 1271 203
rect 1218 145 1229 179
rect 1263 145 1271 179
rect 1501 178 1554 203
rect 1218 119 1271 145
rect 1501 144 1509 178
rect 1543 144 1554 178
rect 1501 119 1554 144
rect 1584 178 1640 203
rect 1584 144 1595 178
rect 1629 144 1640 178
rect 1584 119 1640 144
rect 1670 178 1723 203
rect 1670 144 1681 178
rect 1715 144 1723 178
rect 1670 119 1723 144
rect 1925 182 1978 206
rect 1925 148 1933 182
rect 1967 148 1978 182
rect 1925 122 1978 148
rect 2008 182 2067 206
rect 2008 148 2022 182
rect 2056 148 2067 182
rect 2008 122 2067 148
rect 2097 122 2139 206
rect 2169 202 2218 206
rect 2252 202 2279 236
rect 2169 168 2279 202
rect 2169 134 2207 168
rect 2241 134 2279 168
rect 2169 122 2279 134
rect 2309 236 2362 250
rect 2309 202 2320 236
rect 2354 202 2362 236
rect 2309 168 2362 202
rect 2309 134 2320 168
rect 2354 134 2362 168
rect 2309 122 2362 134
rect 2436 176 2489 224
rect 2436 142 2444 176
rect 2478 142 2489 176
rect 2436 102 2489 142
rect 2436 68 2444 102
rect 2478 68 2489 102
rect 2436 56 2489 68
rect 2519 216 2575 224
rect 2519 182 2530 216
rect 2564 182 2575 216
rect 2519 102 2575 182
rect 2519 68 2530 102
rect 2564 68 2575 102
rect 2519 56 2575 68
rect 2605 212 2658 224
rect 2605 178 2616 212
rect 2650 178 2658 212
rect 2605 140 2658 178
rect 2817 177 2874 215
rect 2817 143 2825 177
rect 2859 143 2874 177
rect 2605 102 2680 140
rect 2605 68 2635 102
rect 2669 68 2680 102
rect 2605 56 2680 68
rect 2710 115 2763 140
rect 2710 81 2721 115
rect 2755 81 2763 115
rect 2710 56 2763 81
rect 2817 93 2874 143
rect 2817 59 2825 93
rect 2859 59 2874 93
rect 2817 47 2874 59
rect 2904 207 2960 215
rect 2904 173 2915 207
rect 2949 173 2960 207
rect 2904 101 2960 173
rect 2904 67 2915 101
rect 2949 67 2960 101
rect 2904 47 2960 67
rect 2990 202 3043 215
rect 2990 168 3001 202
rect 3035 168 3043 202
rect 2990 93 3043 168
rect 2990 59 3001 93
rect 3035 59 3043 93
rect 2990 47 3043 59
<< pdiff >>
rect 27 603 80 617
rect 27 569 35 603
rect 69 569 80 603
rect 27 535 80 569
rect 27 501 35 535
rect 69 501 80 535
rect 27 489 80 501
rect 110 576 174 617
rect 110 542 125 576
rect 159 542 174 576
rect 110 489 174 542
rect 204 489 246 617
rect 276 576 332 617
rect 276 542 287 576
rect 321 542 332 576
rect 276 489 332 542
rect 362 540 415 617
rect 362 506 373 540
rect 407 506 415 540
rect 362 489 415 506
rect 528 527 621 609
rect 528 493 536 527
rect 570 493 621 527
rect 528 481 621 493
rect 651 593 718 609
rect 651 559 672 593
rect 706 559 718 593
rect 651 481 718 559
rect 778 441 858 593
rect 778 407 790 441
rect 824 425 858 441
rect 888 577 941 593
rect 888 543 899 577
rect 933 543 941 577
rect 888 509 941 543
rect 1015 577 1065 593
rect 1015 543 1023 577
rect 1057 543 1065 577
rect 1015 509 1065 543
rect 888 425 963 509
rect 993 487 1065 509
rect 993 425 1045 487
rect 1125 547 1198 585
rect 1125 513 1137 547
rect 1171 513 1198 547
rect 1125 501 1198 513
rect 1228 547 1284 585
rect 1228 513 1239 547
rect 1273 513 1284 547
rect 1228 501 1284 513
rect 1314 575 1387 585
rect 1314 541 1341 575
rect 1375 541 1387 575
rect 1566 575 1624 585
rect 1314 501 1387 541
rect 1566 541 1578 575
rect 1612 541 1624 575
rect 1566 523 1624 541
rect 824 407 836 425
rect 778 399 836 407
rect 1441 439 1521 523
rect 1441 405 1453 439
rect 1487 405 1521 439
rect 1441 395 1521 405
rect 1551 395 1639 523
rect 1669 439 1726 523
rect 1669 405 1680 439
rect 1714 405 1726 439
rect 1669 395 1726 405
rect 1927 539 1984 547
rect 1927 505 1939 539
rect 1973 505 1984 539
rect 1927 423 1984 505
rect 1927 389 1939 423
rect 1973 389 1984 423
rect 1927 379 1984 389
rect 2014 539 2086 547
rect 2014 505 2025 539
rect 2059 505 2086 539
rect 2014 463 2086 505
rect 2116 463 2158 547
rect 2188 535 2273 547
rect 2188 501 2199 535
rect 2233 501 2273 535
rect 2188 463 2273 501
rect 2014 421 2071 463
rect 2014 387 2025 421
rect 2059 387 2071 421
rect 2014 379 2071 387
rect 2220 429 2228 463
rect 2262 429 2273 463
rect 2220 379 2273 429
rect 2303 535 2356 547
rect 2303 501 2314 535
rect 2348 501 2356 535
rect 2303 425 2356 501
rect 2303 391 2314 425
rect 2348 391 2356 425
rect 2303 379 2356 391
rect 2440 581 2493 619
rect 2440 547 2448 581
rect 2482 547 2493 581
rect 2440 367 2493 547
rect 2523 433 2579 619
rect 2523 399 2534 433
rect 2568 399 2579 433
rect 2523 367 2579 399
rect 2609 581 2662 619
rect 2609 547 2620 581
rect 2654 547 2662 581
rect 2609 495 2662 547
rect 2821 607 2874 619
rect 2821 573 2829 607
rect 2863 573 2874 607
rect 2821 539 2874 573
rect 2821 505 2829 539
rect 2863 505 2874 539
rect 2609 367 2684 495
rect 2714 481 2767 495
rect 2714 447 2725 481
rect 2759 447 2767 481
rect 2714 413 2767 447
rect 2714 379 2725 413
rect 2759 379 2767 413
rect 2714 367 2767 379
rect 2821 471 2874 505
rect 2821 437 2829 471
rect 2863 437 2874 471
rect 2821 367 2874 437
rect 2904 599 2960 619
rect 2904 565 2915 599
rect 2949 565 2960 599
rect 2904 507 2960 565
rect 2904 473 2915 507
rect 2949 473 2960 507
rect 2904 420 2960 473
rect 2904 386 2915 420
rect 2949 386 2960 420
rect 2904 367 2960 386
rect 2990 607 3043 619
rect 2990 573 3001 607
rect 3035 573 3043 607
rect 2990 510 3043 573
rect 2990 476 3001 510
rect 3035 476 3043 510
rect 2990 413 3043 476
rect 2990 379 3001 413
rect 3035 379 3043 413
rect 2990 367 3043 379
<< ndiffc >>
rect 35 145 69 179
rect 193 145 227 179
rect 373 133 407 167
rect 475 132 509 166
rect 790 201 824 235
rect 790 133 824 167
rect 958 195 992 229
rect 958 127 992 161
rect 1143 143 1177 177
rect 1229 145 1263 179
rect 1509 144 1543 178
rect 1595 144 1629 178
rect 1681 144 1715 178
rect 1933 148 1967 182
rect 2022 148 2056 182
rect 2218 202 2252 236
rect 2207 134 2241 168
rect 2320 202 2354 236
rect 2320 134 2354 168
rect 2444 142 2478 176
rect 2444 68 2478 102
rect 2530 182 2564 216
rect 2530 68 2564 102
rect 2616 178 2650 212
rect 2825 143 2859 177
rect 2635 68 2669 102
rect 2721 81 2755 115
rect 2825 59 2859 93
rect 2915 173 2949 207
rect 2915 67 2949 101
rect 3001 168 3035 202
rect 3001 59 3035 93
<< pdiffc >>
rect 35 569 69 603
rect 35 501 69 535
rect 125 542 159 576
rect 287 542 321 576
rect 373 506 407 540
rect 536 493 570 527
rect 672 559 706 593
rect 790 407 824 441
rect 899 543 933 577
rect 1023 543 1057 577
rect 1137 513 1171 547
rect 1239 513 1273 547
rect 1341 541 1375 575
rect 1578 541 1612 575
rect 1453 405 1487 439
rect 1680 405 1714 439
rect 1939 505 1973 539
rect 1939 389 1973 423
rect 2025 505 2059 539
rect 2199 501 2233 535
rect 2025 387 2059 421
rect 2228 429 2262 463
rect 2314 501 2348 535
rect 2314 391 2348 425
rect 2448 547 2482 581
rect 2534 399 2568 433
rect 2620 547 2654 581
rect 2829 573 2863 607
rect 2829 505 2863 539
rect 2725 447 2759 481
rect 2725 379 2759 413
rect 2829 437 2863 471
rect 2915 565 2949 599
rect 2915 473 2949 507
rect 2915 386 2949 420
rect 3001 573 3035 607
rect 3001 476 3035 510
rect 3001 379 3035 413
<< poly >>
rect 80 617 110 643
rect 174 617 204 643
rect 246 617 276 643
rect 332 617 362 643
rect 621 609 651 635
rect 733 615 1110 645
rect 80 360 110 489
rect 174 467 204 489
rect 44 344 110 360
rect 44 310 60 344
rect 94 310 110 344
rect 44 276 110 310
rect 44 242 60 276
rect 94 242 110 276
rect 44 226 110 242
rect 80 204 110 226
rect 152 437 204 467
rect 152 204 182 437
rect 246 395 276 489
rect 224 379 290 395
rect 224 345 240 379
rect 274 345 290 379
rect 224 311 290 345
rect 224 277 240 311
rect 274 277 290 311
rect 224 261 290 277
rect 332 308 362 489
rect 513 396 579 412
rect 513 362 529 396
rect 563 362 579 396
rect 513 328 579 362
rect 513 308 529 328
rect 332 294 529 308
rect 563 294 579 328
rect 332 278 579 294
rect 238 204 268 261
rect 332 204 362 278
rect 434 204 464 230
rect 621 187 651 481
rect 733 299 763 615
rect 858 593 888 615
rect 963 509 993 535
rect 1080 455 1110 615
rect 1198 585 1228 611
rect 1284 607 1771 637
rect 1284 585 1314 607
rect 1521 523 1551 549
rect 1639 523 1669 549
rect 1080 439 1146 455
rect 858 399 888 425
rect 963 385 993 425
rect 1080 405 1096 439
rect 1130 405 1146 439
rect 1080 389 1146 405
rect 963 369 1029 385
rect 963 335 979 369
rect 1013 341 1029 369
rect 1013 335 1060 341
rect 963 311 1060 335
rect 1198 333 1228 501
rect 1284 475 1314 501
rect 1521 363 1551 395
rect 1385 347 1451 363
rect 1385 333 1401 347
rect 733 269 865 299
rect 591 171 657 187
rect 591 137 607 171
rect 641 137 657 171
rect 80 94 110 120
rect 152 52 182 120
rect 238 94 268 120
rect 332 94 362 120
rect 434 52 464 120
rect 591 103 657 137
rect 591 69 607 103
rect 641 69 657 103
rect 591 52 657 69
rect 152 22 657 52
rect 733 51 763 269
rect 835 247 865 269
rect 1030 203 1060 311
rect 1102 313 1401 333
rect 1435 313 1451 347
rect 1102 303 1451 313
rect 1102 203 1132 303
rect 1385 297 1451 303
rect 1518 347 1584 363
rect 1518 313 1534 347
rect 1568 313 1584 347
rect 1518 297 1584 313
rect 1518 255 1548 297
rect 1639 292 1669 395
rect 1741 347 1771 607
rect 2086 615 2407 645
rect 2493 619 2523 645
rect 2579 619 2609 645
rect 2874 619 2904 645
rect 2960 619 2990 645
rect 1984 547 2014 573
rect 2086 547 2116 615
rect 2158 547 2188 573
rect 2273 547 2303 573
rect 2086 437 2116 463
rect 2158 395 2188 463
rect 2122 379 2188 395
rect 1741 331 1811 347
rect 1741 297 1761 331
rect 1795 304 1811 331
rect 1984 304 2014 379
rect 2122 345 2138 379
rect 2172 345 2188 379
rect 2122 329 2188 345
rect 2273 339 2303 379
rect 1795 297 2086 304
rect 1632 276 1698 292
rect 1188 225 1584 255
rect 1632 242 1648 276
rect 1682 242 1698 276
rect 1632 226 1698 242
rect 1741 274 2086 297
rect 1741 263 1811 274
rect 1741 229 1761 263
rect 1795 229 1811 263
rect 2056 262 2086 274
rect 2056 232 2097 262
rect 1188 203 1218 225
rect 1554 203 1584 225
rect 1640 203 1670 226
rect 1741 213 1811 229
rect 1978 206 2008 232
rect 2067 206 2097 232
rect 2139 206 2169 329
rect 2236 323 2309 339
rect 2236 289 2252 323
rect 2286 289 2309 323
rect 2236 273 2309 289
rect 2279 250 2309 273
rect 1299 155 1365 171
rect 1299 121 1315 155
rect 1349 121 1365 155
rect 835 93 865 119
rect 1030 93 1060 119
rect 1102 93 1132 119
rect 1188 93 1218 119
rect 1299 87 1365 121
rect 1299 53 1315 87
rect 1349 53 1365 87
rect 1299 51 1365 53
rect 733 21 1365 51
rect 1413 87 1479 103
rect 1554 93 1584 119
rect 1640 93 1670 119
rect 1413 53 1429 87
rect 1463 53 1479 87
rect 1413 51 1479 53
rect 1978 51 2008 122
rect 2067 96 2097 122
rect 2139 96 2169 122
rect 2279 96 2309 122
rect 2377 51 2407 615
rect 2684 495 2714 521
rect 2493 331 2523 367
rect 2579 331 2609 367
rect 2684 331 2714 367
rect 2489 315 2771 331
rect 2489 281 2517 315
rect 2551 281 2585 315
rect 2619 281 2653 315
rect 2687 281 2721 315
rect 2755 281 2771 315
rect 2874 303 2904 367
rect 2960 303 2990 367
rect 2489 265 2771 281
rect 2825 287 2990 303
rect 2489 224 2519 265
rect 2575 224 2605 265
rect 2680 140 2710 265
rect 2825 253 2841 287
rect 2875 253 2990 287
rect 2825 237 2990 253
rect 2874 215 2904 237
rect 2960 215 2990 237
rect 1413 21 2407 51
rect 2489 30 2519 56
rect 2575 30 2605 56
rect 2680 30 2710 56
rect 2874 21 2904 47
rect 2960 21 2990 47
<< polycont >>
rect 60 310 94 344
rect 60 242 94 276
rect 240 345 274 379
rect 240 277 274 311
rect 529 362 563 396
rect 529 294 563 328
rect 1096 405 1130 439
rect 979 335 1013 369
rect 607 137 641 171
rect 607 69 641 103
rect 1401 313 1435 347
rect 1534 313 1568 347
rect 1761 297 1795 331
rect 2138 345 2172 379
rect 1648 242 1682 276
rect 1761 229 1795 263
rect 2252 289 2286 323
rect 1315 121 1349 155
rect 1315 53 1349 87
rect 1429 53 1463 87
rect 2517 281 2551 315
rect 2585 281 2619 315
rect 2653 281 2687 315
rect 2721 281 2755 315
rect 2841 253 2875 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 19 603 85 615
rect 19 569 35 603
rect 69 569 85 603
rect 19 535 85 569
rect 19 501 35 535
rect 69 501 85 535
rect 119 576 175 649
rect 119 542 125 576
rect 159 542 175 576
rect 119 526 175 542
rect 271 581 638 615
rect 271 576 323 581
rect 271 542 287 576
rect 321 542 323 576
rect 271 526 323 542
rect 357 540 423 547
rect 19 492 85 501
rect 357 506 373 540
rect 407 506 423 540
rect 357 492 423 506
rect 19 458 423 492
rect 17 344 161 424
rect 17 310 60 344
rect 94 310 161 344
rect 17 276 161 310
rect 208 379 370 424
rect 208 345 240 379
rect 274 345 370 379
rect 208 311 370 345
rect 208 277 240 311
rect 274 277 370 311
rect 17 242 60 276
rect 94 242 161 276
rect 459 243 493 581
rect 17 237 161 242
rect 17 229 151 237
rect 195 206 493 243
rect 527 527 570 547
rect 527 493 536 527
rect 527 396 570 493
rect 604 509 638 581
rect 672 593 722 649
rect 706 559 722 593
rect 672 543 722 559
rect 883 577 949 649
rect 883 543 899 577
rect 933 543 949 577
rect 1007 581 1391 615
rect 1007 577 1073 581
rect 1007 543 1023 577
rect 1057 543 1073 577
rect 1325 575 1391 581
rect 1121 513 1137 547
rect 1171 513 1187 547
rect 1121 509 1187 513
rect 604 475 1187 509
rect 1223 513 1239 547
rect 1273 513 1289 547
rect 1325 541 1341 575
rect 1375 541 1391 575
rect 1562 575 1628 649
rect 1562 541 1578 575
rect 1612 541 1628 575
rect 604 407 738 475
rect 1223 441 1289 513
rect 1923 539 1975 555
rect 1923 507 1939 539
rect 527 362 529 396
rect 563 362 570 396
rect 527 328 570 362
rect 527 294 529 328
rect 563 294 570 328
rect 19 179 85 195
rect 19 145 35 179
rect 69 145 85 179
rect 19 17 85 145
rect 177 179 243 206
rect 177 145 193 179
rect 227 145 243 179
rect 527 172 570 294
rect 177 129 243 145
rect 357 167 423 172
rect 357 133 373 167
rect 407 133 423 167
rect 357 17 423 133
rect 459 166 570 172
rect 459 132 475 166
rect 509 132 570 166
rect 459 116 570 132
rect 604 171 657 297
rect 604 137 607 171
rect 641 137 657 171
rect 604 103 657 137
rect 604 69 607 103
rect 641 69 657 103
rect 604 53 657 69
rect 704 93 738 407
rect 774 407 790 441
rect 824 407 1029 441
rect 774 235 840 407
rect 963 369 1029 407
rect 1080 439 1289 441
rect 1080 405 1096 439
rect 1130 405 1289 439
rect 1080 403 1289 405
rect 1325 505 1939 507
rect 1973 505 1975 539
rect 1325 473 1975 505
rect 1325 369 1359 473
rect 963 335 979 369
rect 1013 335 1359 369
rect 1399 405 1453 439
rect 1487 405 1503 439
rect 1399 388 1503 405
rect 1664 405 1680 439
rect 1714 405 1730 439
rect 1399 347 1435 388
rect 1664 354 1730 405
rect 1399 313 1401 347
rect 1518 347 1730 354
rect 1923 423 1975 473
rect 1923 389 1939 423
rect 1973 389 1975 423
rect 1518 313 1534 347
rect 1568 331 1810 347
rect 1568 313 1761 331
rect 774 201 790 235
rect 824 201 840 235
rect 774 167 840 201
rect 774 133 790 167
rect 824 133 840 167
rect 774 127 840 133
rect 874 267 1265 301
rect 874 93 908 267
rect 704 59 908 93
rect 942 229 1008 233
rect 942 195 958 229
rect 992 195 1008 229
rect 942 161 1008 195
rect 942 127 958 161
rect 992 127 1008 161
rect 942 17 1008 127
rect 1127 177 1184 193
rect 1127 143 1143 177
rect 1177 143 1184 177
rect 1127 87 1184 143
rect 1218 179 1265 267
rect 1218 145 1229 179
rect 1263 145 1265 179
rect 1399 194 1435 313
rect 1744 297 1761 313
rect 1795 297 1810 331
rect 1469 276 1710 279
rect 1469 242 1648 276
rect 1682 242 1710 276
rect 1469 228 1710 242
rect 1744 263 1810 297
rect 1744 229 1761 263
rect 1795 229 1810 263
rect 1744 194 1810 229
rect 1399 178 1552 194
rect 1218 129 1265 145
rect 1299 155 1365 171
rect 1299 121 1315 155
rect 1349 121 1365 155
rect 1299 87 1365 121
rect 1127 53 1315 87
rect 1349 53 1365 87
rect 1399 144 1509 178
rect 1543 144 1552 178
rect 1399 128 1552 144
rect 1586 178 1636 194
rect 1586 144 1595 178
rect 1629 144 1636 178
rect 1399 87 1479 128
rect 1399 53 1429 87
rect 1463 53 1479 87
rect 1399 51 1479 53
rect 1586 17 1636 144
rect 1670 178 1810 194
rect 1670 144 1681 178
rect 1715 144 1810 178
rect 1670 128 1810 144
rect 1923 182 1975 389
rect 1923 148 1933 182
rect 1967 148 1975 182
rect 1923 132 1975 148
rect 2009 539 2072 555
rect 2009 505 2025 539
rect 2059 505 2072 539
rect 2009 421 2072 505
rect 2183 535 2278 649
rect 2432 581 2498 649
rect 2183 501 2199 535
rect 2233 501 2278 535
rect 2183 463 2278 501
rect 2183 429 2228 463
rect 2262 429 2278 463
rect 2312 535 2388 551
rect 2432 547 2448 581
rect 2482 547 2498 581
rect 2432 543 2498 547
rect 2604 581 2670 649
rect 2604 547 2620 581
rect 2654 547 2670 581
rect 2604 543 2670 547
rect 2825 607 2867 649
rect 2825 573 2829 607
rect 2863 573 2867 607
rect 2312 501 2314 535
rect 2348 509 2388 535
rect 2825 539 2867 573
rect 2348 501 2664 509
rect 2312 475 2664 501
rect 2825 505 2829 539
rect 2863 505 2867 539
rect 2009 387 2025 421
rect 2059 387 2072 421
rect 2312 425 2388 475
rect 2312 395 2314 425
rect 2009 310 2072 387
rect 2122 391 2314 395
rect 2348 391 2388 425
rect 2122 379 2388 391
rect 2122 345 2138 379
rect 2172 359 2388 379
rect 2172 345 2188 359
rect 2122 344 2188 345
rect 2236 323 2302 325
rect 2236 310 2252 323
rect 2009 289 2252 310
rect 2286 289 2302 323
rect 2009 276 2302 289
rect 2009 182 2072 276
rect 2338 242 2388 359
rect 2009 148 2022 182
rect 2056 148 2072 182
rect 2009 132 2072 148
rect 2202 236 2268 242
rect 2202 202 2218 236
rect 2252 202 2268 236
rect 2202 168 2268 202
rect 2202 134 2207 168
rect 2241 134 2268 168
rect 2202 17 2268 134
rect 2304 236 2388 242
rect 2304 202 2320 236
rect 2354 202 2388 236
rect 2422 433 2584 441
rect 2422 399 2534 433
rect 2568 399 2584 433
rect 2422 375 2584 399
rect 2422 244 2467 375
rect 2630 331 2664 475
rect 2709 481 2775 497
rect 2709 447 2725 481
rect 2759 447 2775 481
rect 2709 413 2775 447
rect 2825 471 2867 505
rect 2825 437 2829 471
rect 2863 437 2867 471
rect 2825 421 2867 437
rect 2911 599 2963 615
rect 2911 565 2915 599
rect 2949 565 2963 599
rect 2911 507 2963 565
rect 2911 473 2915 507
rect 2949 473 2963 507
rect 2709 379 2725 413
rect 2759 385 2775 413
rect 2911 420 2963 473
rect 2911 386 2915 420
rect 2949 386 2963 420
rect 2759 379 2875 385
rect 2709 351 2875 379
rect 2501 317 2664 331
rect 2501 315 2771 317
rect 2501 281 2517 315
rect 2551 281 2585 315
rect 2619 281 2653 315
rect 2687 281 2721 315
rect 2755 281 2771 315
rect 2805 287 2875 351
rect 2805 253 2841 287
rect 2805 245 2875 253
rect 2422 216 2574 244
rect 2422 210 2530 216
rect 2304 168 2388 202
rect 2528 182 2530 210
rect 2564 182 2574 216
rect 2304 134 2320 168
rect 2354 134 2388 168
rect 2304 118 2388 134
rect 2428 142 2444 176
rect 2478 142 2494 176
rect 2428 102 2494 142
rect 2428 68 2444 102
rect 2478 68 2494 102
rect 2428 17 2494 68
rect 2528 102 2574 182
rect 2528 68 2530 102
rect 2564 68 2574 102
rect 2528 52 2574 68
rect 2608 212 2677 228
rect 2608 178 2616 212
rect 2650 178 2677 212
rect 2608 102 2677 178
rect 2608 68 2635 102
rect 2669 68 2677 102
rect 2608 17 2677 68
rect 2711 211 2875 245
rect 2711 115 2771 211
rect 2911 207 2963 386
rect 2997 607 3051 649
rect 2997 573 3001 607
rect 3035 573 3051 607
rect 2997 510 3051 573
rect 2997 476 3001 510
rect 3035 476 3051 510
rect 2997 413 3051 476
rect 2997 379 3001 413
rect 3035 379 3051 413
rect 2997 363 3051 379
rect 2711 81 2721 115
rect 2755 81 2771 115
rect 2711 65 2771 81
rect 2809 143 2825 177
rect 2859 143 2875 177
rect 2809 93 2875 143
rect 2809 59 2825 93
rect 2859 59 2875 93
rect 2809 17 2875 59
rect 2911 173 2915 207
rect 2949 173 2963 207
rect 2911 101 2963 173
rect 2911 67 2915 101
rect 2949 67 2963 101
rect 2911 51 2963 67
rect 2997 202 3051 218
rect 2997 168 3001 202
rect 3035 168 3051 202
rect 2997 93 3051 168
rect 2997 59 3001 93
rect 3035 59 3051 93
rect 2997 17 3051 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 683 3072 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 0 617 3072 649
rect 0 17 3072 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
rect 0 -49 3072 -17
<< labels >>
flabel pwell s 0 0 3072 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 3072 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfxbp_2
flabel comment s 751 325 751 325 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 3072 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 3072 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2911 94 2945 128 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2911 168 2945 202 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2911 242 2945 276 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2911 316 2945 350 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2911 390 2945 424 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2911 464 2945 498 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2911 538 2945 572 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2431 242 2465 276 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3072 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6063138
string GDS_START 6041654
<< end >>
