magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 195 202 671 235
rect 1 49 671 202
rect 0 0 672 49
<< scnmos >>
rect 82 92 112 176
rect 276 125 306 209
rect 394 125 424 209
rect 480 125 510 209
rect 558 125 588 209
<< scpmoshvt >>
rect 124 419 174 619
rect 230 419 280 619
rect 328 419 378 619
rect 434 419 484 619
rect 540 419 590 619
<< ndiff >>
rect 27 151 82 176
rect 27 117 37 151
rect 71 117 82 151
rect 27 92 82 117
rect 112 151 167 176
rect 112 117 123 151
rect 157 117 167 151
rect 221 171 276 209
rect 221 137 231 171
rect 265 137 276 171
rect 221 125 276 137
rect 306 184 394 209
rect 306 150 333 184
rect 367 150 394 184
rect 306 125 394 150
rect 424 184 480 209
rect 424 150 435 184
rect 469 150 480 184
rect 424 125 480 150
rect 510 125 558 209
rect 588 184 645 209
rect 588 150 599 184
rect 633 150 645 184
rect 588 125 645 150
rect 112 92 167 117
<< pdiff >>
rect 67 607 124 619
rect 67 573 79 607
rect 113 573 124 607
rect 67 515 124 573
rect 67 481 79 515
rect 113 481 124 515
rect 67 419 124 481
rect 174 597 230 619
rect 174 563 185 597
rect 219 563 230 597
rect 174 465 230 563
rect 174 431 185 465
rect 219 431 230 465
rect 174 419 230 431
rect 280 419 328 619
rect 378 607 434 619
rect 378 573 389 607
rect 423 573 434 607
rect 378 524 434 573
rect 378 490 389 524
rect 423 490 434 524
rect 378 419 434 490
rect 484 597 540 619
rect 484 563 495 597
rect 529 563 540 597
rect 484 465 540 563
rect 484 431 495 465
rect 529 431 540 465
rect 484 419 540 431
rect 590 607 645 619
rect 590 573 601 607
rect 635 573 645 607
rect 590 524 645 573
rect 590 490 601 524
rect 635 490 645 524
rect 590 419 645 490
<< ndiffc >>
rect 37 117 71 151
rect 123 117 157 151
rect 231 137 265 171
rect 333 150 367 184
rect 435 150 469 184
rect 599 150 633 184
<< pdiffc >>
rect 79 573 113 607
rect 79 481 113 515
rect 185 563 219 597
rect 185 431 219 465
rect 389 573 423 607
rect 389 490 423 524
rect 495 563 529 597
rect 495 431 529 465
rect 601 573 635 607
rect 601 490 635 524
<< poly >>
rect 124 619 174 645
rect 230 619 280 645
rect 328 619 378 645
rect 434 619 484 645
rect 540 619 590 645
rect 124 359 174 419
rect 82 343 174 359
rect 82 309 124 343
rect 158 309 174 343
rect 82 293 174 309
rect 82 176 112 293
rect 230 254 280 419
rect 328 315 378 419
rect 434 315 484 419
rect 540 368 590 419
rect 526 352 592 368
rect 526 318 542 352
rect 576 318 592 352
rect 348 299 469 315
rect 526 302 592 318
rect 348 265 419 299
rect 453 265 469 299
rect 348 254 469 265
rect 230 224 306 254
rect 348 224 510 254
rect 276 209 306 224
rect 394 209 424 224
rect 480 209 510 224
rect 558 209 588 302
rect 82 66 112 92
rect 276 51 306 125
rect 394 99 424 125
rect 480 99 510 125
rect 558 51 588 125
rect 276 21 588 51
<< polycont >>
rect 124 309 158 343
rect 542 318 576 352
rect 419 265 453 299
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 63 607 129 649
rect 63 573 79 607
rect 113 573 129 607
rect 63 515 129 573
rect 63 481 79 515
rect 113 481 129 515
rect 63 465 129 481
rect 169 597 235 613
rect 169 563 185 597
rect 219 563 235 597
rect 169 465 235 563
rect 373 607 439 649
rect 373 573 389 607
rect 423 573 439 607
rect 373 524 439 573
rect 373 490 389 524
rect 423 490 439 524
rect 373 474 439 490
rect 479 597 545 613
rect 479 563 495 597
rect 529 563 545 597
rect 169 431 185 465
rect 219 431 235 465
rect 479 465 545 563
rect 585 607 651 649
rect 585 573 601 607
rect 635 573 651 607
rect 585 524 651 573
rect 585 490 601 524
rect 635 490 651 524
rect 585 474 651 490
rect 479 438 495 465
rect 169 429 235 431
rect 21 395 235 429
rect 271 431 495 438
rect 529 438 545 465
rect 529 431 654 438
rect 271 404 654 431
rect 21 180 71 395
rect 271 359 305 404
rect 108 343 305 359
rect 108 309 124 343
rect 158 309 305 343
rect 108 293 305 309
rect 403 299 469 356
rect 505 352 584 368
rect 505 318 542 352
rect 576 318 584 352
rect 505 302 584 318
rect 403 265 419 299
rect 453 265 469 299
rect 123 223 367 257
rect 403 249 469 265
rect 21 151 87 180
rect 21 117 37 151
rect 71 117 87 151
rect 21 88 87 117
rect 123 151 173 223
rect 157 117 173 151
rect 123 88 173 117
rect 215 171 281 187
rect 215 137 231 171
rect 265 137 281 171
rect 215 17 281 137
rect 317 184 367 223
rect 620 213 654 404
rect 317 150 333 184
rect 317 121 367 150
rect 419 184 469 213
rect 419 150 435 184
rect 419 17 469 150
rect 583 184 654 213
rect 583 150 599 184
rect 633 150 654 184
rect 583 121 654 150
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xnor2_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4270858
string GDS_START 4265224
<< end >>
