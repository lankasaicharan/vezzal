magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 436 157 624 241
rect 8 49 624 157
rect 0 0 672 49
<< scnmos >>
rect 87 47 117 131
rect 173 47 203 131
rect 327 47 357 131
rect 417 47 447 131
rect 515 47 545 215
<< scpmoshvt >>
rect 93 480 123 564
rect 165 480 195 564
rect 237 480 267 564
rect 309 480 339 564
rect 562 367 592 619
<< ndiff >>
rect 462 165 515 215
rect 462 131 470 165
rect 504 131 515 165
rect 34 106 87 131
rect 34 72 42 106
rect 76 72 87 106
rect 34 47 87 72
rect 117 106 173 131
rect 117 72 128 106
rect 162 72 173 106
rect 117 47 173 72
rect 203 93 327 131
rect 203 59 214 93
rect 248 59 282 93
rect 316 59 327 93
rect 203 47 327 59
rect 357 106 417 131
rect 357 72 372 106
rect 406 72 417 106
rect 357 47 417 72
rect 447 93 515 131
rect 447 59 470 93
rect 504 59 515 93
rect 447 47 515 59
rect 545 181 598 215
rect 545 147 556 181
rect 590 147 598 181
rect 545 93 598 147
rect 545 59 556 93
rect 590 59 598 93
rect 545 47 598 59
<< pdiff >>
rect 509 607 562 619
rect 509 573 517 607
rect 551 573 562 607
rect 509 564 562 573
rect 40 539 93 564
rect 40 505 48 539
rect 82 505 93 539
rect 40 480 93 505
rect 123 480 165 564
rect 195 480 237 564
rect 267 480 309 564
rect 339 539 562 564
rect 339 505 350 539
rect 384 505 437 539
rect 471 514 562 539
rect 471 505 517 514
rect 339 480 517 505
rect 551 480 562 514
rect 509 367 562 480
rect 592 599 645 619
rect 592 565 603 599
rect 637 565 645 599
rect 592 504 645 565
rect 592 470 603 504
rect 637 470 645 504
rect 592 413 645 470
rect 592 379 603 413
rect 637 379 645 413
rect 592 367 645 379
<< ndiffc >>
rect 470 131 504 165
rect 42 72 76 106
rect 128 72 162 106
rect 214 59 248 93
rect 282 59 316 93
rect 372 72 406 106
rect 470 59 504 93
rect 556 147 590 181
rect 556 59 590 93
<< pdiffc >>
rect 517 573 551 607
rect 48 505 82 539
rect 350 505 384 539
rect 437 505 471 539
rect 517 480 551 514
rect 603 565 637 599
rect 603 470 637 504
rect 603 379 637 413
<< poly >>
rect 562 619 592 645
rect 93 564 123 590
rect 165 564 195 590
rect 237 564 267 590
rect 309 564 339 590
rect 93 302 123 480
rect 21 286 123 302
rect 21 252 37 286
rect 71 252 123 286
rect 21 218 123 252
rect 21 184 37 218
rect 71 184 123 218
rect 21 168 123 184
rect 165 315 195 480
rect 237 387 267 480
rect 309 459 339 480
rect 309 429 429 459
rect 237 357 303 387
rect 273 335 303 357
rect 399 335 429 429
rect 273 319 357 335
rect 165 299 231 315
rect 165 265 181 299
rect 215 265 231 299
rect 165 231 231 265
rect 165 197 181 231
rect 215 197 231 231
rect 273 285 295 319
rect 329 285 357 319
rect 273 251 357 285
rect 399 319 465 335
rect 399 285 415 319
rect 449 285 465 319
rect 562 303 592 367
rect 399 269 465 285
rect 513 287 592 303
rect 273 217 295 251
rect 329 217 357 251
rect 273 201 357 217
rect 165 181 231 197
rect 87 131 117 168
rect 173 131 203 181
rect 327 131 357 201
rect 417 131 447 269
rect 513 253 529 287
rect 563 253 592 287
rect 513 237 592 253
rect 515 215 545 237
rect 87 21 117 47
rect 173 21 203 47
rect 327 21 357 47
rect 417 21 447 47
rect 515 21 545 47
<< polycont >>
rect 37 252 71 286
rect 37 184 71 218
rect 181 265 215 299
rect 181 197 215 231
rect 295 285 329 319
rect 415 285 449 319
rect 295 217 329 251
rect 529 253 563 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 334 607 567 649
rect 334 573 517 607
rect 551 573 567 607
rect 32 539 98 555
rect 32 505 48 539
rect 82 505 98 539
rect 32 452 98 505
rect 334 539 567 573
rect 334 505 350 539
rect 384 505 437 539
rect 471 514 567 539
rect 471 505 517 514
rect 334 489 517 505
rect 501 480 517 489
rect 551 480 567 514
rect 501 464 567 480
rect 601 599 655 615
rect 601 565 603 599
rect 637 565 655 599
rect 601 504 655 565
rect 601 470 603 504
rect 637 470 655 504
rect 32 430 467 452
rect 32 400 563 430
rect 433 386 563 400
rect 17 286 82 366
rect 17 252 37 286
rect 71 252 82 286
rect 17 218 82 252
rect 17 184 37 218
rect 71 184 82 218
rect 117 299 231 366
rect 117 265 181 299
rect 215 265 231 299
rect 117 231 231 265
rect 117 197 181 231
rect 215 197 231 231
rect 279 319 355 366
rect 279 285 295 319
rect 329 285 355 319
rect 399 319 465 352
rect 399 285 415 319
rect 449 285 465 319
rect 513 287 563 386
rect 279 251 355 285
rect 279 217 295 251
rect 329 217 355 251
rect 513 253 529 287
rect 513 249 563 253
rect 279 201 355 217
rect 389 215 563 249
rect 601 413 655 470
rect 601 379 603 413
rect 637 379 655 413
rect 17 156 82 184
rect 389 163 423 215
rect 601 181 655 379
rect 120 129 423 163
rect 26 106 86 122
rect 26 72 42 106
rect 76 72 86 106
rect 26 17 86 72
rect 120 106 164 129
rect 120 72 128 106
rect 162 72 164 106
rect 366 106 423 129
rect 120 56 164 72
rect 198 93 332 95
rect 198 59 214 93
rect 248 59 282 93
rect 316 59 332 93
rect 198 17 332 59
rect 366 72 372 106
rect 406 72 423 106
rect 366 56 423 72
rect 457 165 506 181
rect 457 131 470 165
rect 504 131 506 165
rect 457 93 506 131
rect 457 59 470 93
rect 504 59 506 93
rect 457 17 506 59
rect 540 147 556 181
rect 590 147 655 181
rect 540 93 655 147
rect 540 59 556 93
rect 590 59 655 93
rect 540 51 655 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or4_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 327160
string GDS_START 319866
<< end >>
