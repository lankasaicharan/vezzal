magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3986 1975
<< nwell >>
rect -38 331 2726 704
rect 2334 315 2561 331
<< pwell >>
rect 1734 281 1844 282
rect 776 237 1186 263
rect 1602 237 1996 281
rect 2499 237 2687 257
rect 776 232 2687 237
rect 4 169 192 173
rect 429 169 539 191
rect 753 169 2687 232
rect 4 49 2687 169
rect 0 0 2688 49
<< scnmos >>
rect 83 63 113 147
rect 331 59 361 143
rect 403 59 433 143
rect 535 59 565 143
rect 619 59 649 143
rect 727 59 757 143
rect 852 69 882 237
rect 1050 47 1080 215
rect 1321 127 1351 211
rect 1407 127 1437 211
rect 1479 127 1509 211
rect 1551 127 1581 211
rect 1708 127 1738 255
rect 1840 127 1870 255
rect 1992 127 2022 211
rect 2064 127 2094 211
rect 2196 127 2226 211
rect 2268 127 2298 211
rect 2473 63 2503 147
rect 2578 63 2608 231
<< scpmoshvt >>
rect 83 367 113 495
rect 282 491 312 619
rect 354 491 384 619
rect 532 491 562 619
rect 604 491 634 619
rect 712 491 742 619
rect 827 367 857 619
rect 1050 367 1080 619
rect 1248 529 1278 613
rect 1334 529 1364 613
rect 1406 529 1436 613
rect 1492 529 1522 613
rect 1801 449 1831 617
rect 1887 449 1917 617
rect 1992 533 2022 617
rect 2064 533 2094 617
rect 2191 533 2221 617
rect 2277 533 2307 617
rect 2423 351 2453 479
rect 2547 367 2577 619
<< ndiff >>
rect 30 122 83 147
rect 30 88 38 122
rect 72 88 83 122
rect 30 63 83 88
rect 113 109 166 147
rect 455 157 513 165
rect 455 143 467 157
rect 113 75 124 109
rect 158 75 166 109
rect 113 63 166 75
rect 278 105 331 143
rect 278 71 286 105
rect 320 71 331 105
rect 278 59 331 71
rect 361 59 403 143
rect 433 123 467 143
rect 501 143 513 157
rect 802 206 852 237
rect 779 143 852 206
rect 501 123 535 143
rect 433 59 535 123
rect 565 59 619 143
rect 649 101 727 143
rect 649 67 660 101
rect 694 67 727 101
rect 649 59 727 67
rect 757 89 852 143
rect 757 59 791 89
rect 779 55 791 59
rect 825 69 852 89
rect 882 229 939 237
rect 882 195 893 229
rect 927 195 939 229
rect 1102 229 1160 237
rect 1102 215 1114 229
rect 882 69 939 195
rect 993 89 1050 215
rect 825 55 837 69
rect 779 47 837 55
rect 993 55 1005 89
rect 1039 55 1050 89
rect 993 47 1050 55
rect 1080 195 1114 215
rect 1148 195 1160 229
rect 1760 255 1818 256
rect 1628 211 1708 255
rect 1080 47 1160 195
rect 1214 175 1321 211
rect 1214 141 1224 175
rect 1258 141 1321 175
rect 1214 127 1321 141
rect 1351 186 1407 211
rect 1351 152 1362 186
rect 1396 152 1407 186
rect 1351 127 1407 152
rect 1437 127 1479 211
rect 1509 127 1551 211
rect 1581 127 1708 211
rect 1738 248 1840 255
rect 1738 214 1772 248
rect 1806 214 1840 248
rect 1738 127 1840 214
rect 1870 243 1970 255
rect 1870 209 1924 243
rect 1958 211 1970 243
rect 1958 209 1992 211
rect 1870 175 1992 209
rect 1870 141 1924 175
rect 1958 141 1992 175
rect 1870 127 1992 141
rect 2022 127 2064 211
rect 2094 169 2196 211
rect 2094 135 2128 169
rect 2162 135 2196 169
rect 2094 127 2196 135
rect 2226 127 2268 211
rect 2298 169 2355 211
rect 2525 215 2578 231
rect 2298 135 2309 169
rect 2343 135 2355 169
rect 2525 181 2533 215
rect 2567 181 2578 215
rect 2525 147 2578 181
rect 2298 127 2355 135
rect 1628 108 1686 127
rect 1628 74 1640 108
rect 1674 74 1686 108
rect 1628 66 1686 74
rect 2420 120 2473 147
rect 2420 86 2428 120
rect 2462 86 2473 120
rect 2420 63 2473 86
rect 2503 109 2578 147
rect 2503 75 2521 109
rect 2555 75 2578 109
rect 2503 63 2578 75
rect 2608 212 2661 231
rect 2608 178 2619 212
rect 2653 178 2661 212
rect 2608 109 2661 178
rect 2608 75 2619 109
rect 2653 75 2661 109
rect 2608 63 2661 75
<< pdiff >>
rect 399 625 517 639
rect 399 619 407 625
rect 229 577 282 619
rect 229 543 237 577
rect 271 543 282 577
rect 30 483 83 495
rect 30 449 38 483
rect 72 449 83 483
rect 30 413 83 449
rect 30 379 38 413
rect 72 379 83 413
rect 30 367 83 379
rect 113 483 166 495
rect 229 491 282 543
rect 312 491 354 619
rect 384 591 407 619
rect 441 591 475 625
rect 509 619 517 625
rect 509 591 532 619
rect 384 491 532 591
rect 562 491 604 619
rect 634 609 712 619
rect 634 575 655 609
rect 689 575 712 609
rect 634 541 712 575
rect 634 507 655 541
rect 689 507 712 541
rect 634 491 712 507
rect 742 593 827 619
rect 742 559 767 593
rect 801 559 827 593
rect 742 491 827 559
rect 113 449 124 483
rect 158 449 166 483
rect 113 413 166 449
rect 113 379 124 413
rect 158 379 166 413
rect 113 367 166 379
rect 774 367 827 491
rect 857 436 910 619
rect 857 402 868 436
rect 902 402 910 436
rect 857 367 910 402
rect 997 593 1050 619
rect 997 559 1005 593
rect 1039 559 1050 593
rect 997 367 1050 559
rect 1080 436 1133 619
rect 1721 631 1779 639
rect 1191 588 1248 613
rect 1191 554 1203 588
rect 1237 554 1248 588
rect 1191 529 1248 554
rect 1278 588 1334 613
rect 1278 554 1289 588
rect 1323 554 1334 588
rect 1278 529 1334 554
rect 1364 529 1406 613
rect 1436 588 1492 613
rect 1436 554 1447 588
rect 1481 554 1492 588
rect 1436 529 1492 554
rect 1522 588 1575 613
rect 1522 554 1533 588
rect 1567 554 1575 588
rect 1522 529 1575 554
rect 1721 597 1733 631
rect 1767 617 1779 631
rect 1767 597 1801 617
rect 1080 402 1091 436
rect 1125 402 1133 436
rect 1080 367 1133 402
rect 1721 449 1801 597
rect 1831 491 1887 617
rect 1831 457 1842 491
rect 1876 457 1887 491
rect 1831 449 1887 457
rect 1917 533 1992 617
rect 2022 533 2064 617
rect 2094 592 2191 617
rect 2094 558 2124 592
rect 2158 558 2191 592
rect 2094 533 2191 558
rect 2221 592 2277 617
rect 2221 558 2232 592
rect 2266 558 2277 592
rect 2221 533 2277 558
rect 2307 592 2360 617
rect 2307 558 2318 592
rect 2352 558 2360 592
rect 2307 533 2360 558
rect 2482 607 2547 619
rect 2482 573 2490 607
rect 2524 573 2547 607
rect 1917 531 1970 533
rect 1917 497 1928 531
rect 1962 497 1970 531
rect 1917 449 1970 497
rect 2482 509 2547 573
rect 2482 479 2490 509
rect 2370 467 2423 479
rect 2370 433 2378 467
rect 2412 433 2423 467
rect 2370 351 2423 433
rect 2453 475 2490 479
rect 2524 475 2547 509
rect 2453 409 2547 475
rect 2453 375 2490 409
rect 2524 375 2547 409
rect 2453 367 2547 375
rect 2577 599 2634 619
rect 2577 565 2592 599
rect 2626 565 2634 599
rect 2577 507 2634 565
rect 2577 473 2592 507
rect 2626 473 2634 507
rect 2577 413 2634 473
rect 2577 379 2592 413
rect 2626 379 2634 413
rect 2577 367 2634 379
rect 2453 351 2525 367
<< ndiffc >>
rect 38 88 72 122
rect 124 75 158 109
rect 286 71 320 105
rect 467 123 501 157
rect 660 67 694 101
rect 791 55 825 89
rect 893 195 927 229
rect 1005 55 1039 89
rect 1114 195 1148 229
rect 1224 141 1258 175
rect 1362 152 1396 186
rect 1772 214 1806 248
rect 1924 209 1958 243
rect 1924 141 1958 175
rect 2128 135 2162 169
rect 2309 135 2343 169
rect 2533 181 2567 215
rect 1640 74 1674 108
rect 2428 86 2462 120
rect 2521 75 2555 109
rect 2619 178 2653 212
rect 2619 75 2653 109
<< pdiffc >>
rect 237 543 271 577
rect 38 449 72 483
rect 38 379 72 413
rect 407 591 441 625
rect 475 591 509 625
rect 655 575 689 609
rect 655 507 689 541
rect 767 559 801 593
rect 124 449 158 483
rect 124 379 158 413
rect 868 402 902 436
rect 1005 559 1039 593
rect 1203 554 1237 588
rect 1289 554 1323 588
rect 1447 554 1481 588
rect 1533 554 1567 588
rect 1733 597 1767 631
rect 1091 402 1125 436
rect 1842 457 1876 491
rect 2124 558 2158 592
rect 2232 558 2266 592
rect 2318 558 2352 592
rect 2490 573 2524 607
rect 1928 497 1962 531
rect 2378 433 2412 467
rect 2490 475 2524 509
rect 2490 375 2524 409
rect 2592 565 2626 599
rect 2592 473 2626 507
rect 2592 379 2626 413
<< poly >>
rect 282 619 312 645
rect 354 619 384 645
rect 83 495 113 521
rect 532 619 562 645
rect 604 619 634 645
rect 712 619 742 645
rect 827 619 857 645
rect 1050 619 1080 645
rect 282 469 312 491
rect 219 443 312 469
rect 219 409 235 443
rect 269 439 312 443
rect 269 409 285 439
rect 219 393 285 409
rect 354 391 384 491
rect 532 437 562 491
rect 441 421 562 437
rect 327 375 393 391
rect 83 277 113 367
rect 327 341 343 375
rect 377 341 393 375
rect 441 387 457 421
rect 491 407 562 421
rect 491 387 532 407
rect 441 371 532 387
rect 327 325 393 341
rect 604 335 634 491
rect 712 439 742 491
rect 580 329 634 335
rect 547 305 634 329
rect 676 423 742 439
rect 676 389 692 423
rect 726 389 742 423
rect 676 355 742 389
rect 1248 613 1278 639
rect 1334 613 1364 639
rect 1406 613 1436 639
rect 1492 613 1522 639
rect 1801 617 1831 643
rect 1887 617 1917 643
rect 1992 617 2022 643
rect 2064 617 2094 643
rect 2191 617 2221 643
rect 2277 617 2307 643
rect 2547 619 2577 645
rect 1248 507 1278 529
rect 1198 477 1278 507
rect 676 321 692 355
rect 726 335 742 355
rect 827 335 857 367
rect 726 321 763 335
rect 676 305 763 321
rect 827 319 945 335
rect 1050 325 1080 367
rect 547 299 610 305
rect 547 280 577 299
rect 83 261 469 277
rect 83 247 419 261
rect 83 147 113 247
rect 403 227 419 247
rect 453 227 469 261
rect 403 211 469 227
rect 511 264 577 280
rect 511 230 527 264
rect 561 230 577 264
rect 511 214 577 230
rect 619 241 685 257
rect 190 195 256 199
rect 190 183 361 195
rect 190 149 206 183
rect 240 165 361 183
rect 240 149 256 165
rect 190 133 256 149
rect 331 143 361 165
rect 403 143 433 211
rect 83 37 113 63
rect 535 143 565 214
rect 619 207 635 241
rect 669 207 685 241
rect 619 191 685 207
rect 619 143 649 191
rect 727 143 757 305
rect 827 285 895 319
rect 929 285 945 319
rect 827 269 945 285
rect 993 315 1080 325
rect 1198 315 1228 477
rect 1334 429 1364 529
rect 1276 413 1364 429
rect 1276 379 1292 413
rect 1326 379 1364 413
rect 1406 429 1436 529
rect 1492 507 1522 529
rect 1623 515 1689 531
rect 1492 477 1581 507
rect 1406 413 1509 429
rect 1406 399 1459 413
rect 1276 363 1364 379
rect 1414 379 1459 399
rect 1493 379 1509 413
rect 1414 363 1509 379
rect 993 309 1437 315
rect 993 275 1009 309
rect 1043 285 1437 309
rect 1043 275 1080 285
rect 852 237 882 269
rect 993 259 1080 275
rect 331 33 361 59
rect 403 33 433 59
rect 535 33 565 59
rect 619 33 649 59
rect 727 33 757 59
rect 1050 215 1080 259
rect 852 43 882 69
rect 1321 211 1351 237
rect 1407 211 1437 285
rect 1479 211 1509 363
rect 1551 349 1581 477
rect 1623 481 1639 515
rect 1673 481 1689 515
rect 1623 447 1689 481
rect 1623 413 1639 447
rect 1673 427 1689 447
rect 1801 427 1831 449
rect 1673 413 1831 427
rect 1887 417 1917 449
rect 1623 397 1831 413
rect 1873 401 1939 417
rect 1551 333 1633 349
rect 1551 299 1583 333
rect 1617 299 1633 333
rect 1551 283 1633 299
rect 1551 211 1581 283
rect 1708 255 1738 397
rect 1873 367 1889 401
rect 1923 367 1939 401
rect 1873 351 1939 367
rect 1992 309 2022 533
rect 1840 279 2022 309
rect 2064 501 2094 533
rect 2064 485 2149 501
rect 2064 451 2099 485
rect 2133 451 2149 485
rect 2064 435 2149 451
rect 1840 255 1870 279
rect 1992 211 2022 237
rect 2064 211 2094 435
rect 2191 393 2221 533
rect 2142 377 2226 393
rect 2142 343 2158 377
rect 2192 343 2226 377
rect 2142 309 2226 343
rect 2142 275 2158 309
rect 2192 275 2226 309
rect 2277 299 2307 533
rect 2423 479 2453 505
rect 2142 259 2226 275
rect 2196 211 2226 259
rect 2268 283 2334 299
rect 2268 249 2284 283
rect 2318 263 2334 283
rect 2423 263 2453 351
rect 2547 319 2577 367
rect 2318 249 2453 263
rect 2533 303 2608 319
rect 2533 269 2549 303
rect 2583 269 2608 303
rect 2533 253 2608 269
rect 2268 233 2453 249
rect 2268 211 2298 233
rect 2423 199 2453 233
rect 2578 231 2608 253
rect 2423 169 2503 199
rect 2473 147 2503 169
rect 1321 105 1351 127
rect 1292 89 1358 105
rect 1292 55 1308 89
rect 1342 55 1358 89
rect 1050 21 1080 47
rect 1292 39 1358 55
rect 1407 51 1437 127
rect 1479 101 1509 127
rect 1551 101 1581 127
rect 1708 101 1738 127
rect 1840 51 1870 127
rect 1992 105 2022 127
rect 1407 21 1870 51
rect 1956 89 2022 105
rect 2064 101 2094 127
rect 2196 101 2226 127
rect 2268 101 2298 127
rect 1956 55 1972 89
rect 2006 55 2022 89
rect 1956 39 2022 55
rect 2473 37 2503 63
rect 2578 37 2608 63
<< polycont >>
rect 235 409 269 443
rect 343 341 377 375
rect 457 387 491 421
rect 692 389 726 423
rect 692 321 726 355
rect 419 227 453 261
rect 527 230 561 264
rect 206 149 240 183
rect 635 207 669 241
rect 895 285 929 319
rect 1292 379 1326 413
rect 1459 379 1493 413
rect 1009 275 1043 309
rect 1639 481 1673 515
rect 1639 413 1673 447
rect 1583 299 1617 333
rect 1889 367 1923 401
rect 2099 451 2133 485
rect 2158 343 2192 377
rect 2158 275 2192 309
rect 2284 249 2318 283
rect 2549 269 2583 303
rect 1308 55 1342 89
rect 1972 55 2006 89
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 22 483 81 649
rect 391 625 525 649
rect 221 577 287 593
rect 391 591 407 625
rect 441 591 475 625
rect 509 591 525 625
rect 639 609 705 613
rect 221 543 237 577
rect 271 557 287 577
rect 639 575 655 609
rect 689 575 705 609
rect 639 557 705 575
rect 271 543 705 557
rect 751 593 817 649
rect 751 559 767 593
rect 801 559 817 593
rect 751 554 817 559
rect 989 593 1055 649
rect 989 559 1005 593
rect 1039 559 1055 593
rect 989 554 1055 559
rect 1183 588 1247 604
rect 1183 554 1203 588
rect 1237 554 1247 588
rect 221 541 705 543
rect 221 523 655 541
rect 639 507 655 523
rect 689 520 705 541
rect 1183 520 1247 554
rect 689 507 1247 520
rect 22 449 38 483
rect 72 449 81 483
rect 22 413 81 449
rect 22 379 38 413
rect 72 379 81 413
rect 22 363 81 379
rect 115 489 162 499
rect 115 483 592 489
rect 115 449 124 483
rect 158 455 592 483
rect 639 486 1247 507
rect 1281 588 1339 604
rect 1281 554 1289 588
rect 1323 554 1339 588
rect 1281 504 1339 554
rect 1431 588 1491 649
rect 1717 631 1783 649
rect 1431 554 1447 588
rect 1481 554 1491 588
rect 1431 538 1491 554
rect 1525 588 1675 604
rect 1717 597 1733 631
rect 1767 597 1783 631
rect 1525 554 1533 588
rect 1567 554 1675 588
rect 1819 581 2063 615
rect 1819 561 1853 581
rect 1525 515 1675 554
rect 1525 504 1639 515
rect 639 473 807 486
rect 158 449 285 455
rect 115 443 285 449
rect 115 413 235 443
rect 115 379 124 413
rect 158 409 235 413
rect 269 409 285 443
rect 558 439 592 455
rect 158 393 285 409
rect 158 379 162 393
rect 115 363 162 379
rect 328 375 377 391
rect 22 122 81 138
rect 22 88 38 122
rect 72 88 81 122
rect 22 17 81 88
rect 115 113 154 363
rect 328 341 343 375
rect 328 219 377 341
rect 190 183 377 219
rect 411 387 457 421
rect 491 387 524 421
rect 558 404 653 439
rect 411 370 524 387
rect 411 315 557 370
rect 411 261 468 315
rect 411 227 419 261
rect 453 227 468 261
rect 411 211 468 227
rect 502 264 577 281
rect 502 230 527 264
rect 561 230 577 264
rect 502 214 577 230
rect 619 241 653 404
rect 692 424 739 439
rect 692 423 703 424
rect 737 390 739 424
rect 726 389 739 390
rect 692 355 739 389
rect 726 321 739 355
rect 692 305 739 321
rect 619 207 635 241
rect 669 207 685 241
rect 190 149 206 183
rect 240 149 377 183
rect 773 171 807 473
rect 1281 481 1639 504
rect 1673 481 1675 515
rect 1281 470 1675 481
rect 1281 464 1400 470
rect 864 436 1043 452
rect 864 402 868 436
rect 902 402 1043 436
rect 864 386 1043 402
rect 895 319 929 350
rect 895 269 929 285
rect 1009 309 1043 386
rect 1009 233 1043 275
rect 877 229 1043 233
rect 877 195 893 229
rect 927 195 1043 229
rect 877 193 1043 195
rect 1079 436 1232 452
rect 1079 402 1091 436
rect 1125 430 1232 436
rect 1125 413 1326 430
rect 1125 402 1292 413
rect 1079 379 1292 402
rect 1079 363 1326 379
rect 1079 259 1164 363
rect 1079 229 1326 259
rect 1079 195 1114 229
rect 1148 225 1326 229
rect 1148 195 1164 225
rect 1079 193 1164 195
rect 451 159 807 171
rect 1208 175 1258 191
rect 1208 159 1224 175
rect 451 157 1224 159
rect 451 123 467 157
rect 501 141 1224 157
rect 501 137 1258 141
rect 501 123 517 137
rect 773 125 1258 137
rect 451 121 517 123
rect 115 109 174 113
rect 115 75 124 109
rect 158 75 174 109
rect 115 59 174 75
rect 270 105 336 109
rect 270 71 286 105
rect 320 87 336 105
rect 644 101 710 103
rect 644 87 660 101
rect 320 71 660 87
rect 270 67 660 71
rect 694 67 710 101
rect 1292 102 1326 225
rect 1360 186 1400 464
rect 1639 447 1675 470
rect 1443 413 1509 429
rect 1443 379 1459 413
rect 1493 379 1509 413
rect 1443 252 1509 379
rect 1551 424 1605 436
rect 1551 390 1567 424
rect 1601 390 1605 424
rect 1673 413 1675 447
rect 1639 397 1675 413
rect 1709 527 1853 561
rect 1926 531 1993 547
rect 1551 349 1605 390
rect 1709 349 1743 527
rect 1926 497 1928 531
rect 1962 497 1993 531
rect 1551 333 1743 349
rect 1551 299 1583 333
rect 1617 299 1743 333
rect 1551 286 1743 299
rect 1788 491 1892 493
rect 1788 457 1842 491
rect 1876 457 1892 491
rect 1926 481 1993 497
rect 1788 453 1892 457
rect 1788 252 1822 453
rect 1443 248 1822 252
rect 1443 214 1772 248
rect 1806 214 1822 248
rect 1443 212 1822 214
rect 1856 401 1925 417
rect 1856 367 1889 401
rect 1923 367 1925 401
rect 1856 351 1925 367
rect 1360 152 1362 186
rect 1396 152 1400 186
rect 1856 178 1890 351
rect 1959 259 1993 481
rect 2029 393 2063 581
rect 2108 592 2174 649
rect 2108 558 2124 592
rect 2158 558 2174 592
rect 2108 542 2174 558
rect 2216 592 2276 615
rect 2216 558 2232 592
rect 2266 558 2276 592
rect 2216 501 2276 558
rect 2310 592 2368 649
rect 2310 558 2318 592
rect 2352 558 2368 592
rect 2310 542 2368 558
rect 2474 607 2542 649
rect 2474 573 2490 607
rect 2524 573 2542 607
rect 2474 517 2542 573
rect 2490 509 2542 517
rect 2099 485 2278 501
rect 2133 451 2278 485
rect 2099 435 2278 451
rect 2244 393 2278 435
rect 2362 467 2456 483
rect 2362 433 2378 467
rect 2412 433 2456 467
rect 2362 427 2456 433
rect 2029 377 2208 393
rect 2029 343 2158 377
rect 2192 343 2208 377
rect 2244 359 2388 393
rect 2029 309 2208 343
rect 2029 275 2158 309
rect 2192 275 2208 309
rect 2268 283 2320 299
rect 1360 136 1400 152
rect 1436 144 1890 178
rect 1436 102 1470 144
rect 270 53 710 67
rect 775 89 841 91
rect 775 55 791 89
rect 825 55 841 89
rect 775 17 841 55
rect 989 89 1055 91
rect 989 55 1005 89
rect 1039 55 1055 89
rect 989 17 1055 55
rect 1292 89 1470 102
rect 1292 55 1308 89
rect 1342 55 1470 89
rect 1292 51 1470 55
rect 1624 108 1690 110
rect 1624 74 1640 108
rect 1674 74 1690 108
rect 1624 17 1690 74
rect 1839 91 1890 144
rect 1924 243 1993 259
rect 1958 241 1993 243
rect 2268 249 2284 283
rect 2318 249 2320 283
rect 2268 241 2320 249
rect 1958 209 2320 241
rect 1924 205 2320 209
rect 1924 175 1993 205
rect 1958 141 1993 175
rect 2354 171 2388 359
rect 1924 125 1993 141
rect 2112 169 2178 171
rect 2112 135 2128 169
rect 2162 135 2178 169
rect 1839 89 2022 91
rect 1839 55 1972 89
rect 2006 55 2022 89
rect 1839 51 2022 55
rect 2112 17 2178 135
rect 2293 169 2388 171
rect 2293 135 2309 169
rect 2343 135 2388 169
rect 2293 119 2388 135
rect 2422 319 2456 427
rect 2524 475 2542 509
rect 2490 409 2542 475
rect 2524 375 2542 409
rect 2490 353 2542 375
rect 2576 599 2669 615
rect 2576 565 2592 599
rect 2626 565 2669 599
rect 2576 507 2669 565
rect 2576 473 2592 507
rect 2626 473 2669 507
rect 2576 413 2669 473
rect 2576 379 2592 413
rect 2626 379 2669 413
rect 2576 363 2669 379
rect 2422 303 2583 319
rect 2422 269 2549 303
rect 2422 253 2583 269
rect 2422 120 2471 253
rect 2422 86 2428 120
rect 2462 86 2471 120
rect 2422 70 2471 86
rect 2505 215 2583 219
rect 2505 181 2533 215
rect 2567 181 2583 215
rect 2505 109 2583 181
rect 2505 75 2521 109
rect 2555 75 2583 109
rect 2505 17 2583 75
rect 2617 212 2669 363
rect 2617 178 2619 212
rect 2653 178 2669 212
rect 2617 109 2669 178
rect 2617 75 2619 109
rect 2653 75 2669 109
rect 2617 59 2669 75
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 703 423 737 424
rect 703 390 726 423
rect 726 390 737 423
rect 1567 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 691 424 749 430
rect 691 390 703 424
rect 737 421 749 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 737 393 1567 421
rect 737 390 749 393
rect 691 384 749 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
flabel pwell s 0 0 2688 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2688 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfrtn_1
flabel metal1 s 0 617 2688 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2688 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 2623 94 2657 128 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 168 2657 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 242 2657 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 316 2657 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 390 2657 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 464 2657 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 2143 316 2177 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 2623 538 2657 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
rlabel metal1 s 1555 421 1613 430 1 RESET_B
port 3 nsew signal input
rlabel metal1 s 1555 384 1613 393 1 RESET_B
port 3 nsew signal input
rlabel metal1 s 691 421 749 430 1 RESET_B
port 3 nsew signal input
rlabel metal1 s 691 393 1613 421 1 RESET_B
port 3 nsew signal input
rlabel metal1 s 691 384 749 393 1 RESET_B
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2688 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4970214
string GDS_START 4950718
<< end >>
