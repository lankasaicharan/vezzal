magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
rect 452 303 1353 331
<< pwell >>
rect 1747 167 2015 202
rect 1 165 433 167
rect 1319 165 2015 167
rect 1 49 2015 165
rect 0 0 2016 49
<< scnmos >>
rect 84 57 114 141
rect 156 57 186 141
rect 248 57 278 141
rect 320 57 350 141
rect 518 55 548 139
rect 590 55 620 139
rect 676 55 706 139
rect 754 55 784 139
rect 856 55 886 139
rect 934 55 964 139
rect 1132 55 1162 139
rect 1204 55 1234 139
rect 1402 57 1432 141
rect 1474 57 1504 141
rect 1560 57 1590 141
rect 1632 57 1662 141
rect 1830 92 1860 176
rect 1902 92 1932 176
<< scpmoshvt >>
rect 90 409 140 609
rect 228 409 278 609
rect 545 339 595 539
rect 667 393 717 593
rect 765 393 815 593
rect 928 393 978 593
rect 1042 393 1092 593
rect 1210 393 1260 593
rect 1506 367 1556 567
rect 1612 367 1662 567
rect 1830 409 1880 609
<< ndiff >>
rect 27 116 84 141
rect 27 82 39 116
rect 73 82 84 116
rect 27 57 84 82
rect 114 57 156 141
rect 186 108 248 141
rect 186 74 197 108
rect 231 74 248 108
rect 186 57 248 74
rect 278 57 320 141
rect 350 116 407 141
rect 1773 151 1830 176
rect 350 82 361 116
rect 395 82 407 116
rect 350 57 407 82
rect 461 115 518 139
rect 461 81 473 115
rect 507 81 518 115
rect 461 55 518 81
rect 548 55 590 139
rect 620 114 676 139
rect 620 80 631 114
rect 665 80 676 114
rect 620 55 676 80
rect 706 55 754 139
rect 784 114 856 139
rect 784 80 811 114
rect 845 80 856 114
rect 784 55 856 80
rect 886 55 934 139
rect 964 114 1132 139
rect 964 80 1023 114
rect 1057 80 1132 114
rect 964 55 1132 80
rect 1162 55 1204 139
rect 1234 115 1291 139
rect 1234 81 1245 115
rect 1279 81 1291 115
rect 1234 55 1291 81
rect 1345 103 1402 141
rect 1345 69 1357 103
rect 1391 69 1402 103
rect 1345 57 1402 69
rect 1432 57 1474 141
rect 1504 116 1560 141
rect 1504 82 1515 116
rect 1549 82 1560 116
rect 1504 57 1560 82
rect 1590 57 1632 141
rect 1662 116 1719 141
rect 1662 82 1673 116
rect 1707 82 1719 116
rect 1773 117 1785 151
rect 1819 117 1830 151
rect 1773 92 1830 117
rect 1860 92 1902 176
rect 1932 151 1989 176
rect 1932 117 1943 151
rect 1977 117 1989 151
rect 1932 92 1989 117
rect 1662 57 1719 82
<< pdiff >>
rect 155 627 213 639
rect 155 609 167 627
rect 33 597 90 609
rect 33 563 45 597
rect 79 563 90 597
rect 33 526 90 563
rect 33 492 45 526
rect 79 492 90 526
rect 33 455 90 492
rect 33 421 45 455
rect 79 421 90 455
rect 33 409 90 421
rect 140 593 167 609
rect 201 609 213 627
rect 201 593 228 609
rect 140 409 228 593
rect 278 455 335 609
rect 1773 597 1830 609
rect 610 569 667 593
rect 610 539 622 569
rect 278 421 289 455
rect 323 421 335 455
rect 278 409 335 421
rect 488 385 545 539
rect 488 351 500 385
rect 534 351 545 385
rect 488 339 545 351
rect 595 535 622 539
rect 656 535 667 569
rect 595 393 667 535
rect 717 393 765 593
rect 815 581 928 593
rect 815 547 842 581
rect 876 547 928 581
rect 815 510 928 547
rect 815 476 842 510
rect 876 476 928 510
rect 815 439 928 476
rect 815 405 842 439
rect 876 405 928 439
rect 815 393 928 405
rect 978 393 1042 593
rect 1092 581 1210 593
rect 1092 547 1114 581
rect 1148 547 1210 581
rect 1092 447 1210 547
rect 1092 413 1114 447
rect 1148 413 1210 447
rect 1092 393 1210 413
rect 1260 581 1317 593
rect 1260 547 1271 581
rect 1305 547 1317 581
rect 1260 510 1317 547
rect 1260 476 1271 510
rect 1305 476 1317 510
rect 1260 439 1317 476
rect 1260 405 1271 439
rect 1305 405 1317 439
rect 1260 393 1317 405
rect 1449 555 1506 567
rect 1449 521 1461 555
rect 1495 521 1506 555
rect 1449 484 1506 521
rect 1449 450 1461 484
rect 1495 450 1506 484
rect 1449 413 1506 450
rect 595 339 645 393
rect 1449 379 1461 413
rect 1495 379 1506 413
rect 1449 367 1506 379
rect 1556 555 1612 567
rect 1556 521 1567 555
rect 1601 521 1612 555
rect 1556 484 1612 521
rect 1556 450 1567 484
rect 1601 450 1612 484
rect 1556 413 1612 450
rect 1556 379 1567 413
rect 1601 379 1612 413
rect 1556 367 1612 379
rect 1662 555 1719 567
rect 1662 521 1673 555
rect 1707 521 1719 555
rect 1662 484 1719 521
rect 1662 450 1673 484
rect 1707 450 1719 484
rect 1662 413 1719 450
rect 1662 379 1673 413
rect 1707 379 1719 413
rect 1773 563 1785 597
rect 1819 563 1830 597
rect 1773 526 1830 563
rect 1773 492 1785 526
rect 1819 492 1830 526
rect 1773 455 1830 492
rect 1773 421 1785 455
rect 1819 421 1830 455
rect 1773 409 1830 421
rect 1880 597 1937 609
rect 1880 563 1891 597
rect 1925 563 1937 597
rect 1880 526 1937 563
rect 1880 492 1891 526
rect 1925 492 1937 526
rect 1880 455 1937 492
rect 1880 421 1891 455
rect 1925 421 1937 455
rect 1880 409 1937 421
rect 1662 367 1719 379
<< ndiffc >>
rect 39 82 73 116
rect 197 74 231 108
rect 361 82 395 116
rect 473 81 507 115
rect 631 80 665 114
rect 811 80 845 114
rect 1023 80 1057 114
rect 1245 81 1279 115
rect 1357 69 1391 103
rect 1515 82 1549 116
rect 1673 82 1707 116
rect 1785 117 1819 151
rect 1943 117 1977 151
<< pdiffc >>
rect 45 563 79 597
rect 45 492 79 526
rect 45 421 79 455
rect 167 593 201 627
rect 289 421 323 455
rect 500 351 534 385
rect 622 535 656 569
rect 842 547 876 581
rect 842 476 876 510
rect 842 405 876 439
rect 1114 547 1148 581
rect 1114 413 1148 447
rect 1271 547 1305 581
rect 1271 476 1305 510
rect 1271 405 1305 439
rect 1461 521 1495 555
rect 1461 450 1495 484
rect 1461 379 1495 413
rect 1567 521 1601 555
rect 1567 450 1601 484
rect 1567 379 1601 413
rect 1673 521 1707 555
rect 1673 450 1707 484
rect 1673 379 1707 413
rect 1785 563 1819 597
rect 1785 492 1819 526
rect 1785 421 1819 455
rect 1891 563 1925 597
rect 1891 492 1925 526
rect 1891 421 1925 455
<< poly >>
rect 90 609 140 635
rect 228 609 278 635
rect 390 613 717 643
rect 390 597 456 613
rect 390 563 406 597
rect 440 563 456 597
rect 667 593 717 613
rect 765 593 815 619
rect 928 593 978 619
rect 1042 593 1092 619
rect 1210 593 1260 619
rect 1830 609 1880 635
rect 390 547 456 563
rect 545 539 595 565
rect 90 356 140 409
rect 228 369 278 409
rect 90 340 186 356
rect 90 306 117 340
rect 151 306 186 340
rect 90 272 186 306
rect 90 252 117 272
rect 84 238 117 252
rect 151 238 186 272
rect 84 222 186 238
rect 228 353 379 369
rect 228 319 329 353
rect 363 319 379 353
rect 1506 567 1556 593
rect 1612 567 1662 593
rect 667 367 717 393
rect 676 362 717 367
rect 228 285 379 319
rect 545 299 595 339
rect 228 251 329 285
rect 363 251 379 285
rect 228 235 379 251
rect 518 283 620 299
rect 518 249 570 283
rect 604 249 620 283
rect 84 141 114 222
rect 156 141 186 222
rect 248 141 278 235
rect 320 141 350 235
rect 518 233 620 249
rect 518 139 548 233
rect 590 139 620 233
rect 676 139 706 362
rect 765 351 815 393
rect 928 361 978 393
rect 1042 361 1092 393
rect 765 335 831 351
rect 765 301 781 335
rect 815 315 831 335
rect 928 345 994 361
rect 815 301 886 315
rect 765 285 886 301
rect 928 311 944 345
rect 978 311 994 345
rect 928 295 994 311
rect 1042 345 1162 361
rect 1042 311 1112 345
rect 1146 311 1162 345
rect 1042 295 1162 311
rect 748 213 814 229
rect 748 179 764 213
rect 798 179 814 213
rect 748 163 814 179
rect 754 139 784 163
rect 856 139 886 285
rect 1042 184 1072 295
rect 1210 291 1260 393
rect 1318 297 1384 313
rect 1204 275 1270 291
rect 1204 241 1220 275
rect 1254 241 1270 275
rect 1204 225 1270 241
rect 1318 263 1334 297
rect 1368 263 1384 297
rect 1318 229 1384 263
rect 1204 184 1234 225
rect 934 154 1072 184
rect 1132 154 1234 184
rect 1318 195 1334 229
rect 1368 209 1384 229
rect 1506 209 1556 367
rect 1612 209 1662 367
rect 1830 352 1880 409
rect 1773 336 1880 352
rect 1773 302 1789 336
rect 1823 302 1880 336
rect 1773 268 1880 302
rect 1773 234 1789 268
rect 1823 248 1880 268
rect 1823 234 1932 248
rect 1773 218 1932 234
rect 1368 195 1662 209
rect 1318 179 1662 195
rect 934 139 964 154
rect 1132 139 1162 154
rect 1204 139 1234 154
rect 1402 141 1432 179
rect 1474 141 1504 179
rect 1560 141 1590 179
rect 1632 141 1662 179
rect 1830 176 1860 218
rect 1902 176 1932 218
rect 84 31 114 57
rect 156 31 186 57
rect 248 31 278 57
rect 320 31 350 57
rect 1830 66 1860 92
rect 1902 66 1932 92
rect 518 29 548 55
rect 590 29 620 55
rect 676 29 706 55
rect 754 29 784 55
rect 856 29 886 55
rect 934 29 964 55
rect 1132 29 1162 55
rect 1204 29 1234 55
rect 1402 31 1432 57
rect 1474 31 1504 57
rect 1560 31 1590 57
rect 1632 31 1662 57
<< polycont >>
rect 406 563 440 597
rect 117 306 151 340
rect 117 238 151 272
rect 329 319 363 353
rect 329 251 363 285
rect 570 249 604 283
rect 781 301 815 335
rect 944 311 978 345
rect 1112 311 1146 345
rect 764 179 798 213
rect 1220 241 1254 275
rect 1334 263 1368 297
rect 1334 195 1368 229
rect 1789 302 1823 336
rect 1789 234 1823 268
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 151 627 217 649
rect 23 597 95 613
rect 23 563 45 597
rect 79 563 95 597
rect 151 593 167 627
rect 201 593 217 627
rect 151 577 217 593
rect 390 597 456 613
rect 23 541 95 563
rect 390 563 406 597
rect 440 563 456 597
rect 390 541 456 563
rect 23 526 456 541
rect 23 492 45 526
rect 79 507 456 526
rect 606 569 672 649
rect 606 535 622 569
rect 656 535 672 569
rect 606 507 672 535
rect 826 581 1062 597
rect 826 547 842 581
rect 876 563 1062 581
rect 876 547 892 563
rect 826 510 892 547
rect 79 492 95 507
rect 23 455 95 492
rect 826 476 842 510
rect 876 476 892 510
rect 23 421 45 455
rect 79 421 95 455
rect 23 405 95 421
rect 243 455 620 471
rect 243 421 289 455
rect 323 437 620 455
rect 323 421 339 437
rect 243 405 339 421
rect 23 145 57 405
rect 101 340 167 356
rect 101 306 117 340
rect 151 306 167 340
rect 101 272 167 306
rect 101 238 117 272
rect 151 238 167 272
rect 101 222 167 238
rect 243 199 277 405
rect 457 385 550 401
rect 313 353 379 369
rect 313 319 329 353
rect 363 319 379 353
rect 313 285 379 319
rect 313 251 329 285
rect 363 251 379 285
rect 313 235 379 251
rect 457 351 500 385
rect 534 351 550 385
rect 457 335 550 351
rect 586 351 620 437
rect 826 439 892 476
rect 826 405 842 439
rect 876 405 892 439
rect 826 389 892 405
rect 586 335 831 351
rect 243 165 411 199
rect 23 116 89 145
rect 23 82 39 116
rect 73 82 89 116
rect 23 53 89 82
rect 181 108 247 129
rect 181 74 197 108
rect 231 74 247 108
rect 181 17 247 74
rect 345 116 411 165
rect 345 82 361 116
rect 395 82 411 116
rect 345 53 411 82
rect 457 197 491 335
rect 586 301 781 335
rect 815 301 831 335
rect 928 345 992 361
rect 928 329 944 345
rect 586 299 831 301
rect 554 285 831 299
rect 867 311 944 329
rect 978 311 992 345
rect 867 295 992 311
rect 554 283 620 285
rect 554 249 570 283
rect 604 249 620 283
rect 554 233 620 249
rect 867 229 901 295
rect 1028 259 1062 563
rect 1098 581 1164 649
rect 1098 547 1114 581
rect 1148 547 1164 581
rect 1098 447 1164 547
rect 1098 413 1114 447
rect 1148 413 1164 447
rect 1098 397 1164 413
rect 1255 581 1321 597
rect 1255 547 1271 581
rect 1305 547 1321 581
rect 1255 510 1321 547
rect 1255 476 1271 510
rect 1305 476 1321 510
rect 1255 439 1321 476
rect 1255 405 1271 439
rect 1305 405 1321 439
rect 1255 361 1321 405
rect 1420 555 1511 578
rect 1420 521 1461 555
rect 1495 521 1511 555
rect 1420 484 1511 521
rect 1420 450 1461 484
rect 1495 450 1511 484
rect 1420 413 1511 450
rect 1420 379 1461 413
rect 1495 379 1511 413
rect 1098 345 1352 361
rect 1098 311 1112 345
rect 1146 327 1352 345
rect 1146 311 1162 327
rect 1098 295 1162 311
rect 1318 313 1352 327
rect 1318 297 1384 313
rect 1204 275 1270 291
rect 1204 259 1220 275
rect 748 213 901 229
rect 748 197 764 213
rect 457 179 764 197
rect 798 179 901 213
rect 457 163 901 179
rect 937 241 1220 259
rect 1254 241 1270 275
rect 937 225 1270 241
rect 1318 263 1334 297
rect 1368 263 1384 297
rect 1318 229 1384 263
rect 457 115 523 163
rect 937 127 971 225
rect 1318 195 1334 229
rect 1368 195 1384 229
rect 1318 189 1384 195
rect 1229 179 1384 189
rect 1420 236 1511 379
rect 1551 555 1617 649
rect 1769 597 1835 649
rect 1551 521 1567 555
rect 1601 521 1617 555
rect 1551 484 1617 521
rect 1551 450 1567 484
rect 1601 450 1617 484
rect 1551 413 1617 450
rect 1551 379 1567 413
rect 1601 379 1617 413
rect 1551 363 1617 379
rect 1657 555 1723 571
rect 1657 521 1673 555
rect 1707 521 1723 555
rect 1657 484 1723 521
rect 1657 450 1673 484
rect 1707 450 1723 484
rect 1657 413 1723 450
rect 1657 379 1673 413
rect 1707 379 1723 413
rect 1769 563 1785 597
rect 1819 563 1835 597
rect 1769 526 1835 563
rect 1769 492 1785 526
rect 1819 492 1835 526
rect 1769 455 1835 492
rect 1769 421 1785 455
rect 1819 421 1835 455
rect 1769 405 1835 421
rect 1875 597 1941 613
rect 1875 563 1891 597
rect 1925 578 1941 597
rect 1925 563 1993 578
rect 1875 526 1993 563
rect 1875 492 1891 526
rect 1925 492 1993 526
rect 1875 455 1993 492
rect 1875 421 1891 455
rect 1925 421 1993 455
rect 1875 405 1993 421
rect 1657 352 1723 379
rect 1657 336 1839 352
rect 1657 318 1789 336
rect 1229 155 1352 179
rect 457 81 473 115
rect 507 81 523 115
rect 457 53 523 81
rect 615 114 681 127
rect 615 80 631 114
rect 665 80 681 114
rect 615 17 681 80
rect 795 114 971 127
rect 795 80 811 114
rect 845 80 971 114
rect 795 67 971 80
rect 1007 114 1073 143
rect 1007 80 1023 114
rect 1057 80 1073 114
rect 1007 17 1073 80
rect 1229 115 1295 155
rect 1420 119 1454 236
rect 1229 81 1245 115
rect 1279 81 1295 115
rect 1229 53 1295 81
rect 1341 103 1454 119
rect 1341 69 1357 103
rect 1391 69 1454 103
rect 1341 53 1454 69
rect 1499 116 1565 145
rect 1499 82 1515 116
rect 1549 82 1565 116
rect 1499 17 1565 82
rect 1657 116 1723 318
rect 1773 302 1789 318
rect 1823 302 1839 336
rect 1773 268 1839 302
rect 1773 234 1789 268
rect 1823 234 1839 268
rect 1773 218 1839 234
rect 1657 82 1673 116
rect 1707 82 1723 116
rect 1657 53 1723 82
rect 1769 151 1835 180
rect 1769 117 1785 151
rect 1819 117 1835 151
rect 1769 17 1835 117
rect 1927 151 1993 405
rect 1927 117 1943 151
rect 1977 117 1993 151
rect 1927 88 1993 117
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlxbp_lp2
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1471 390 1505 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1471 464 1505 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1471 538 1505 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1951 94 1985 128 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 168 1985 202 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 390 1985 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 464 1985 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1951 538 1985 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2280324
string GDS_START 2266002
<< end >>
