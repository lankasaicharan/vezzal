magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 1 49 1123 248
rect 0 0 1152 49
<< scpmos >>
rect 87 368 117 592
rect 186 368 216 592
rect 286 368 316 592
rect 376 368 406 592
rect 476 368 506 592
rect 576 368 606 592
rect 666 368 696 592
rect 758 368 788 592
rect 1036 368 1066 592
<< nmoslvt >>
rect 84 74 114 222
rect 184 74 214 222
rect 289 74 319 222
rect 384 74 414 222
rect 484 74 514 222
rect 598 74 628 222
rect 684 74 714 222
rect 798 74 828 222
rect 996 74 1026 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 182 184 222
rect 114 148 139 182
rect 173 148 184 182
rect 114 74 184 148
rect 214 144 289 222
rect 214 110 239 144
rect 273 110 289 144
rect 214 74 289 110
rect 319 182 384 222
rect 319 148 339 182
rect 373 148 384 182
rect 319 74 384 148
rect 414 210 484 222
rect 414 176 439 210
rect 473 176 484 210
rect 414 120 484 176
rect 414 86 439 120
rect 473 86 484 120
rect 414 74 484 86
rect 514 210 598 222
rect 514 176 539 210
rect 573 176 598 210
rect 514 120 598 176
rect 514 86 539 120
rect 573 86 598 120
rect 514 74 598 86
rect 628 210 684 222
rect 628 176 639 210
rect 673 176 684 210
rect 628 120 684 176
rect 628 86 639 120
rect 673 86 684 120
rect 628 74 684 86
rect 714 210 798 222
rect 714 176 739 210
rect 773 176 798 210
rect 714 120 798 176
rect 714 86 739 120
rect 773 86 798 120
rect 714 74 798 86
rect 828 210 885 222
rect 828 176 839 210
rect 873 176 885 210
rect 828 120 885 176
rect 828 86 839 120
rect 873 86 885 120
rect 828 74 885 86
rect 939 210 996 222
rect 939 176 951 210
rect 985 176 996 210
rect 939 120 996 176
rect 939 86 951 120
rect 985 86 996 120
rect 939 74 996 86
rect 1026 198 1097 222
rect 1026 164 1051 198
rect 1085 164 1097 198
rect 1026 120 1097 164
rect 1026 86 1051 120
rect 1085 86 1097 120
rect 1026 74 1097 86
<< pdiff >>
rect 27 580 87 592
rect 27 546 39 580
rect 73 546 87 580
rect 27 503 87 546
rect 27 469 39 503
rect 73 469 87 503
rect 27 424 87 469
rect 27 390 39 424
rect 73 390 87 424
rect 27 368 87 390
rect 117 540 186 592
rect 117 506 139 540
rect 173 506 186 540
rect 117 424 186 506
rect 117 390 139 424
rect 173 390 186 424
rect 117 368 186 390
rect 216 580 286 592
rect 216 546 239 580
rect 273 546 286 580
rect 216 508 286 546
rect 216 474 239 508
rect 273 474 286 508
rect 216 368 286 474
rect 316 540 376 592
rect 316 506 329 540
rect 363 506 376 540
rect 316 424 376 506
rect 316 390 329 424
rect 363 390 376 424
rect 316 368 376 390
rect 406 580 476 592
rect 406 546 429 580
rect 463 546 476 580
rect 406 497 476 546
rect 406 463 429 497
rect 463 463 476 497
rect 406 414 476 463
rect 406 380 429 414
rect 463 380 476 414
rect 406 368 476 380
rect 506 582 576 592
rect 506 548 529 582
rect 563 548 576 582
rect 506 514 576 548
rect 506 480 529 514
rect 563 480 576 514
rect 506 446 576 480
rect 506 412 529 446
rect 563 412 576 446
rect 506 368 576 412
rect 606 580 666 592
rect 606 546 619 580
rect 653 546 666 580
rect 606 497 666 546
rect 606 463 619 497
rect 653 463 666 497
rect 606 414 666 463
rect 606 380 619 414
rect 653 380 666 414
rect 606 368 666 380
rect 696 582 758 592
rect 696 548 710 582
rect 744 548 758 582
rect 696 514 758 548
rect 696 480 710 514
rect 744 480 758 514
rect 696 446 758 480
rect 696 412 710 446
rect 744 412 758 446
rect 696 368 758 412
rect 788 580 847 592
rect 788 546 801 580
rect 835 546 847 580
rect 788 497 847 546
rect 788 463 801 497
rect 835 463 847 497
rect 788 414 847 463
rect 788 380 801 414
rect 835 380 847 414
rect 788 368 847 380
rect 977 580 1036 592
rect 977 546 989 580
rect 1023 546 1036 580
rect 977 497 1036 546
rect 977 463 989 497
rect 1023 463 1036 497
rect 977 414 1036 463
rect 977 380 989 414
rect 1023 380 1036 414
rect 977 368 1036 380
rect 1066 580 1125 592
rect 1066 546 1079 580
rect 1113 546 1125 580
rect 1066 497 1125 546
rect 1066 463 1079 497
rect 1113 463 1125 497
rect 1066 414 1125 463
rect 1066 380 1079 414
rect 1113 380 1125 414
rect 1066 368 1125 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 148 173 182
rect 239 110 273 144
rect 339 148 373 182
rect 439 176 473 210
rect 439 86 473 120
rect 539 176 573 210
rect 539 86 573 120
rect 639 176 673 210
rect 639 86 673 120
rect 739 176 773 210
rect 739 86 773 120
rect 839 176 873 210
rect 839 86 873 120
rect 951 176 985 210
rect 951 86 985 120
rect 1051 164 1085 198
rect 1051 86 1085 120
<< pdiffc >>
rect 39 546 73 580
rect 39 469 73 503
rect 39 390 73 424
rect 139 506 173 540
rect 139 390 173 424
rect 239 546 273 580
rect 239 474 273 508
rect 329 506 363 540
rect 329 390 363 424
rect 429 546 463 580
rect 429 463 463 497
rect 429 380 463 414
rect 529 548 563 582
rect 529 480 563 514
rect 529 412 563 446
rect 619 546 653 580
rect 619 463 653 497
rect 619 380 653 414
rect 710 548 744 582
rect 710 480 744 514
rect 710 412 744 446
rect 801 546 835 580
rect 801 463 835 497
rect 801 380 835 414
rect 989 546 1023 580
rect 989 463 1023 497
rect 989 380 1023 414
rect 1079 546 1113 580
rect 1079 463 1113 497
rect 1079 380 1113 414
<< poly >>
rect 87 592 117 618
rect 186 592 216 618
rect 286 592 316 618
rect 376 592 406 618
rect 476 592 506 618
rect 576 592 606 618
rect 666 592 696 618
rect 758 592 788 618
rect 879 582 945 598
rect 1036 592 1066 618
rect 879 548 895 582
rect 929 548 945 582
rect 879 514 945 548
rect 879 480 895 514
rect 929 480 945 514
rect 879 446 945 480
rect 879 412 895 446
rect 929 412 945 446
rect 879 378 945 412
rect 87 353 117 368
rect 186 353 216 368
rect 286 353 316 368
rect 376 353 406 368
rect 476 353 506 368
rect 576 353 606 368
rect 666 353 696 368
rect 758 353 788 368
rect 879 353 895 378
rect 84 336 120 353
rect 183 336 219 353
rect 283 336 319 353
rect 84 320 319 336
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 300 319 320
rect 373 300 409 353
rect 473 344 895 353
rect 929 344 945 378
rect 1036 353 1066 368
rect 473 323 945 344
rect 1033 326 1069 353
rect 996 310 1130 326
rect 270 286 414 300
rect 84 270 414 286
rect 996 276 1012 310
rect 1046 276 1080 310
rect 1114 276 1130 310
rect 996 275 1130 276
rect 84 222 114 270
rect 184 222 214 270
rect 289 222 319 270
rect 384 222 414 270
rect 484 245 1130 275
rect 484 222 514 245
rect 598 222 628 245
rect 684 222 714 245
rect 798 222 828 245
rect 996 222 1026 245
rect 84 48 114 74
rect 184 48 214 74
rect 289 48 319 74
rect 384 48 414 74
rect 484 48 514 74
rect 598 48 628 74
rect 684 48 714 74
rect 798 48 828 74
rect 996 48 1026 74
<< polycont >>
rect 895 548 929 582
rect 895 480 929 514
rect 895 412 929 446
rect 100 286 134 320
rect 168 286 202 320
rect 236 286 270 320
rect 895 344 929 378
rect 1012 276 1046 310
rect 1080 276 1114 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 581 479 615
rect 23 580 89 581
rect 23 546 39 580
rect 73 546 89 580
rect 223 580 273 581
rect 23 503 89 546
rect 23 469 39 503
rect 73 469 89 503
rect 23 424 89 469
rect 23 390 39 424
rect 73 390 89 424
rect 123 540 189 547
rect 123 506 139 540
rect 173 506 189 540
rect 123 424 189 506
rect 223 546 239 580
rect 413 580 479 581
rect 223 508 273 546
rect 223 474 239 508
rect 223 458 273 474
rect 313 540 379 547
rect 313 506 329 540
rect 363 506 379 540
rect 313 424 379 506
rect 123 390 139 424
rect 173 390 329 424
rect 363 390 379 424
rect 25 320 286 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 286 320
rect 25 270 286 286
rect 323 236 379 390
rect 413 546 429 580
rect 463 546 479 580
rect 413 497 479 546
rect 413 463 429 497
rect 463 463 479 497
rect 413 414 479 463
rect 413 380 429 414
rect 463 380 479 414
rect 513 582 563 649
rect 513 548 529 582
rect 513 514 563 548
rect 513 480 529 514
rect 513 446 563 480
rect 513 412 529 446
rect 513 396 563 412
rect 603 580 653 596
rect 603 546 619 580
rect 603 497 653 546
rect 603 463 619 497
rect 603 414 653 463
rect 413 362 479 380
rect 603 380 619 414
rect 693 582 745 649
rect 879 596 957 598
rect 693 548 710 582
rect 744 548 745 582
rect 693 514 745 548
rect 693 480 710 514
rect 744 480 745 514
rect 693 446 745 480
rect 693 412 710 446
rect 744 412 745 446
rect 693 396 745 412
rect 785 580 835 596
rect 785 546 801 580
rect 785 497 835 546
rect 785 463 801 497
rect 785 414 835 463
rect 603 362 653 380
rect 785 380 801 414
rect 785 362 835 380
rect 413 328 835 362
rect 879 582 1039 596
rect 879 548 895 582
rect 929 580 1039 582
rect 929 548 989 580
rect 879 546 989 548
rect 1023 546 1039 580
rect 879 514 1039 546
rect 879 480 895 514
rect 929 497 1039 514
rect 929 480 989 497
rect 879 463 989 480
rect 1023 463 1039 497
rect 879 446 1039 463
rect 879 412 895 446
rect 929 414 1039 446
rect 929 412 989 414
rect 879 380 989 412
rect 1023 380 1039 414
rect 879 378 1039 380
rect 879 344 895 378
rect 929 364 1039 378
rect 1079 580 1129 649
rect 1113 546 1129 580
rect 1079 497 1129 546
rect 1113 463 1129 497
rect 1079 414 1129 463
rect 1113 380 1129 414
rect 1079 364 1129 380
rect 929 344 957 364
rect 879 328 957 344
rect 423 260 889 294
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 123 202 389 236
rect 123 182 189 202
rect 123 148 139 182
rect 173 148 189 182
rect 323 182 389 202
rect 123 132 189 148
rect 223 144 289 160
rect 23 86 39 120
rect 73 86 89 120
rect 23 85 89 86
rect 223 110 239 144
rect 273 110 289 144
rect 323 148 339 182
rect 373 148 389 182
rect 323 132 389 148
rect 423 210 489 260
rect 423 176 439 210
rect 473 176 489 210
rect 223 85 289 110
rect 423 120 489 176
rect 423 86 439 120
rect 473 86 489 120
rect 423 85 489 86
rect 23 51 489 85
rect 523 210 589 226
rect 523 176 539 210
rect 573 176 589 210
rect 523 120 589 176
rect 523 86 539 120
rect 573 86 589 120
rect 523 17 589 86
rect 623 210 689 260
rect 623 176 639 210
rect 673 176 689 210
rect 623 120 689 176
rect 623 86 639 120
rect 673 86 689 120
rect 623 70 689 86
rect 723 210 789 226
rect 723 176 739 210
rect 773 176 789 210
rect 723 120 789 176
rect 723 86 739 120
rect 773 86 789 120
rect 723 17 789 86
rect 823 210 889 260
rect 823 176 839 210
rect 873 176 889 210
rect 823 120 889 176
rect 823 86 839 120
rect 873 86 889 120
rect 823 70 889 86
rect 923 226 957 328
rect 996 310 1130 326
rect 996 276 1012 310
rect 1046 276 1080 310
rect 1114 276 1130 310
rect 996 260 1130 276
rect 1081 236 1130 260
rect 923 210 1001 226
rect 923 176 951 210
rect 985 176 1001 210
rect 923 120 1001 176
rect 923 86 951 120
rect 985 86 1001 120
rect 923 70 1001 86
rect 1035 198 1101 202
rect 1035 164 1051 198
rect 1085 164 1101 198
rect 1035 120 1101 164
rect 1035 86 1051 120
rect 1085 86 1101 120
rect 1035 17 1101 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 einvp_4
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 2064652
string GDS_START 2055208
<< end >>
