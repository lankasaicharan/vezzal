magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 332 1478 704
<< pwell >>
rect 806 274 1401 277
rect 177 49 1401 274
rect 0 0 1440 49
<< scpmos >>
rect 98 368 128 592
rect 188 368 218 592
rect 278 368 308 592
rect 368 368 398 592
rect 610 392 640 592
rect 700 392 730 592
rect 790 392 820 592
rect 880 392 910 592
rect 976 392 1006 592
rect 1109 392 1139 592
rect 1199 392 1229 592
rect 1289 392 1319 592
<< nmoslvt >>
rect 256 100 286 248
rect 342 100 372 248
rect 428 100 458 248
rect 514 100 544 248
rect 615 120 645 248
rect 701 120 731 248
rect 787 120 817 248
rect 882 123 912 251
rect 1034 123 1064 251
rect 1120 123 1150 251
rect 1206 123 1236 251
rect 1292 123 1322 251
<< ndiff >>
rect 832 248 882 251
rect 203 178 256 248
rect 203 144 211 178
rect 245 144 256 178
rect 203 100 256 144
rect 286 236 342 248
rect 286 202 297 236
rect 331 202 342 236
rect 286 146 342 202
rect 286 112 297 146
rect 331 112 342 146
rect 286 100 342 112
rect 372 149 428 248
rect 372 115 383 149
rect 417 115 428 149
rect 372 100 428 115
rect 458 220 514 248
rect 458 186 469 220
rect 503 186 514 220
rect 458 146 514 186
rect 458 112 469 146
rect 503 112 514 146
rect 458 100 514 112
rect 544 167 615 248
rect 544 133 555 167
rect 589 133 615 167
rect 544 120 615 133
rect 645 166 701 248
rect 645 132 656 166
rect 690 132 701 166
rect 645 120 701 132
rect 731 235 787 248
rect 731 201 742 235
rect 776 201 787 235
rect 731 120 787 201
rect 817 167 882 248
rect 817 133 832 167
rect 866 133 882 167
rect 817 123 882 133
rect 912 169 1034 251
rect 912 135 923 169
rect 957 135 1034 169
rect 912 123 1034 135
rect 1064 169 1120 251
rect 1064 135 1075 169
rect 1109 135 1120 169
rect 1064 123 1120 135
rect 1150 238 1206 251
rect 1150 204 1161 238
rect 1195 204 1206 238
rect 1150 123 1206 204
rect 1236 239 1292 251
rect 1236 205 1247 239
rect 1281 205 1292 239
rect 1236 169 1292 205
rect 1236 135 1247 169
rect 1281 135 1292 169
rect 1236 123 1292 135
rect 1322 239 1375 251
rect 1322 205 1333 239
rect 1367 205 1375 239
rect 1322 169 1375 205
rect 1322 135 1333 169
rect 1367 135 1375 169
rect 1322 123 1375 135
rect 817 120 867 123
rect 544 100 597 120
<< pdiff >>
rect 43 580 98 592
rect 43 546 51 580
rect 85 546 98 580
rect 43 497 98 546
rect 43 463 51 497
rect 85 463 98 497
rect 43 414 98 463
rect 43 380 51 414
rect 85 380 98 414
rect 43 368 98 380
rect 128 580 188 592
rect 128 546 141 580
rect 175 546 188 580
rect 128 497 188 546
rect 128 463 141 497
rect 175 463 188 497
rect 128 414 188 463
rect 128 380 141 414
rect 175 380 188 414
rect 128 368 188 380
rect 218 580 278 592
rect 218 546 231 580
rect 265 546 278 580
rect 218 497 278 546
rect 218 463 231 497
rect 265 463 278 497
rect 218 414 278 463
rect 218 380 231 414
rect 265 380 278 414
rect 218 368 278 380
rect 308 580 368 592
rect 308 546 321 580
rect 355 546 368 580
rect 308 497 368 546
rect 308 463 321 497
rect 355 463 368 497
rect 308 414 368 463
rect 308 380 321 414
rect 355 380 368 414
rect 308 368 368 380
rect 398 580 453 592
rect 398 546 411 580
rect 445 546 453 580
rect 398 500 453 546
rect 398 466 411 500
rect 445 466 453 500
rect 398 420 453 466
rect 398 386 411 420
rect 445 386 453 420
rect 555 531 610 592
rect 555 497 563 531
rect 597 497 610 531
rect 555 438 610 497
rect 555 404 563 438
rect 597 404 610 438
rect 555 392 610 404
rect 640 573 700 592
rect 640 539 653 573
rect 687 539 700 573
rect 640 392 700 539
rect 730 498 790 592
rect 730 464 743 498
rect 777 464 790 498
rect 730 392 790 464
rect 820 573 880 592
rect 820 539 833 573
rect 867 539 880 573
rect 820 392 880 539
rect 910 580 976 592
rect 910 546 923 580
rect 957 546 976 580
rect 910 509 976 546
rect 910 475 923 509
rect 957 475 976 509
rect 910 438 976 475
rect 910 404 923 438
rect 957 404 976 438
rect 910 392 976 404
rect 1006 580 1109 592
rect 1006 546 1037 580
rect 1071 546 1109 580
rect 1006 492 1109 546
rect 1006 458 1037 492
rect 1071 458 1109 492
rect 1006 392 1109 458
rect 1139 580 1199 592
rect 1139 546 1152 580
rect 1186 546 1199 580
rect 1139 510 1199 546
rect 1139 476 1152 510
rect 1186 476 1199 510
rect 1139 440 1199 476
rect 1139 406 1152 440
rect 1186 406 1199 440
rect 1139 392 1199 406
rect 1229 580 1289 592
rect 1229 546 1242 580
rect 1276 546 1289 580
rect 1229 492 1289 546
rect 1229 458 1242 492
rect 1276 458 1289 492
rect 1229 392 1289 458
rect 1319 580 1374 592
rect 1319 546 1332 580
rect 1366 546 1374 580
rect 1319 509 1374 546
rect 1319 475 1332 509
rect 1366 475 1374 509
rect 1319 438 1374 475
rect 1319 404 1332 438
rect 1366 404 1374 438
rect 1319 392 1374 404
rect 398 368 453 386
<< ndiffc >>
rect 211 144 245 178
rect 297 202 331 236
rect 297 112 331 146
rect 383 115 417 149
rect 469 186 503 220
rect 469 112 503 146
rect 555 133 589 167
rect 656 132 690 166
rect 742 201 776 235
rect 832 133 866 167
rect 923 135 957 169
rect 1075 135 1109 169
rect 1161 204 1195 238
rect 1247 205 1281 239
rect 1247 135 1281 169
rect 1333 205 1367 239
rect 1333 135 1367 169
<< pdiffc >>
rect 51 546 85 580
rect 51 463 85 497
rect 51 380 85 414
rect 141 546 175 580
rect 141 463 175 497
rect 141 380 175 414
rect 231 546 265 580
rect 231 463 265 497
rect 231 380 265 414
rect 321 546 355 580
rect 321 463 355 497
rect 321 380 355 414
rect 411 546 445 580
rect 411 466 445 500
rect 411 386 445 420
rect 563 497 597 531
rect 563 404 597 438
rect 653 539 687 573
rect 743 464 777 498
rect 833 539 867 573
rect 923 546 957 580
rect 923 475 957 509
rect 923 404 957 438
rect 1037 546 1071 580
rect 1037 458 1071 492
rect 1152 546 1186 580
rect 1152 476 1186 510
rect 1152 406 1186 440
rect 1242 546 1276 580
rect 1242 458 1276 492
rect 1332 546 1366 580
rect 1332 475 1366 509
rect 1332 404 1366 438
<< poly >>
rect 98 592 128 618
rect 188 592 218 618
rect 278 592 308 618
rect 368 592 398 618
rect 610 592 640 618
rect 700 592 730 618
rect 790 592 820 618
rect 880 592 910 618
rect 976 592 1006 618
rect 1109 592 1139 618
rect 1199 592 1229 618
rect 1289 592 1319 618
rect 610 377 640 392
rect 700 377 730 392
rect 790 377 820 392
rect 880 377 910 392
rect 976 377 1006 392
rect 1109 377 1139 392
rect 1199 377 1229 392
rect 1289 377 1319 392
rect 98 353 128 368
rect 188 353 218 368
rect 278 353 308 368
rect 368 353 398 368
rect 607 353 643 377
rect 697 353 733 377
rect 787 353 823 377
rect 877 354 913 377
rect 95 336 131 353
rect 185 336 221 353
rect 275 336 311 353
rect 365 336 401 353
rect 589 337 655 353
rect 95 320 544 336
rect 95 306 407 320
rect 256 248 286 306
rect 342 286 407 306
rect 441 286 494 320
rect 528 286 544 320
rect 589 303 605 337
rect 639 303 655 337
rect 589 287 655 303
rect 697 337 823 353
rect 697 303 715 337
rect 749 303 823 337
rect 697 287 823 303
rect 865 338 931 354
rect 865 304 881 338
rect 915 304 931 338
rect 865 288 931 304
rect 973 296 1009 377
rect 1106 356 1142 377
rect 1196 356 1232 377
rect 1106 340 1236 356
rect 1106 306 1122 340
rect 1156 306 1236 340
rect 342 270 544 286
rect 342 248 372 270
rect 428 248 458 270
rect 514 248 544 270
rect 615 248 645 287
rect 701 248 731 287
rect 787 248 817 287
rect 882 251 912 288
rect 973 266 1064 296
rect 1106 290 1236 306
rect 1034 251 1064 266
rect 1120 251 1150 290
rect 1206 251 1236 290
rect 1286 266 1322 377
rect 1292 251 1322 266
rect 256 74 286 100
rect 342 74 372 100
rect 428 74 458 100
rect 514 74 544 100
rect 615 94 645 120
rect 701 94 731 120
rect 787 94 817 120
rect 882 97 912 123
rect 1034 101 1064 123
rect 998 85 1064 101
rect 1120 97 1150 123
rect 1206 97 1236 123
rect 998 51 1014 85
rect 1048 55 1064 85
rect 1292 55 1322 123
rect 1048 51 1322 55
rect 998 25 1322 51
<< polycont >>
rect 407 286 441 320
rect 494 286 528 320
rect 605 303 639 337
rect 715 303 749 337
rect 881 304 915 338
rect 1122 306 1156 340
rect 1014 51 1048 85
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 35 580 101 649
rect 35 546 51 580
rect 85 546 101 580
rect 35 497 101 546
rect 35 463 51 497
rect 85 463 101 497
rect 35 414 101 463
rect 35 380 51 414
rect 85 380 101 414
rect 141 580 175 596
rect 141 497 175 546
rect 141 414 175 463
rect 141 330 175 380
rect 215 580 265 649
rect 215 546 231 580
rect 215 497 265 546
rect 215 463 231 497
rect 215 414 265 463
rect 215 380 231 414
rect 215 364 265 380
rect 305 580 371 596
rect 305 546 321 580
rect 355 546 371 580
rect 305 497 371 546
rect 305 463 321 497
rect 355 463 371 497
rect 305 414 371 463
rect 305 380 321 414
rect 355 380 371 414
rect 305 330 371 380
rect 411 580 461 649
rect 445 546 461 580
rect 411 500 461 546
rect 445 466 461 500
rect 411 420 461 466
rect 445 386 461 420
rect 411 370 461 386
rect 495 596 703 615
rect 495 581 883 596
rect 495 336 529 581
rect 637 573 883 581
rect 563 531 597 547
rect 637 539 653 573
rect 687 539 833 573
rect 867 539 883 573
rect 637 532 883 539
rect 923 580 973 596
rect 957 546 973 580
rect 923 509 973 546
rect 597 497 743 498
rect 563 464 743 497
rect 777 475 923 498
rect 957 475 973 509
rect 777 464 973 475
rect 563 438 597 464
rect 923 438 973 464
rect 1007 580 1102 649
rect 1007 546 1037 580
rect 1071 546 1102 580
rect 1007 492 1102 546
rect 1007 458 1037 492
rect 1071 458 1102 492
rect 1136 580 1186 596
rect 1136 546 1152 580
rect 1136 510 1186 546
rect 1136 476 1152 510
rect 563 388 597 404
rect 631 387 839 430
rect 957 424 973 438
rect 1136 440 1186 476
rect 1226 580 1292 649
rect 1226 546 1242 580
rect 1276 546 1292 580
rect 1226 492 1292 546
rect 1226 458 1242 492
rect 1276 458 1292 492
rect 1332 580 1382 596
rect 1366 546 1382 580
rect 1332 509 1382 546
rect 1366 475 1382 509
rect 1136 424 1152 440
rect 957 406 1152 424
rect 1332 438 1382 475
rect 1186 406 1332 424
rect 957 404 1332 406
rect 1366 404 1382 438
rect 923 390 1382 404
rect 923 388 973 390
rect 1332 388 1382 390
rect 631 353 665 387
rect 805 354 839 387
rect 605 337 665 353
rect 141 282 371 330
rect 25 236 371 282
rect 405 320 571 336
rect 405 286 407 320
rect 441 286 494 320
rect 528 286 571 320
rect 639 303 665 337
rect 605 287 665 303
rect 699 337 765 353
rect 699 303 715 337
rect 749 303 765 337
rect 699 287 765 303
rect 805 338 931 354
rect 805 304 881 338
rect 915 304 931 338
rect 805 288 931 304
rect 1081 340 1223 356
rect 1081 306 1122 340
rect 1156 306 1223 340
rect 1081 290 1223 306
rect 405 270 571 286
rect 537 253 571 270
rect 1145 253 1211 255
rect 537 238 1211 253
rect 25 228 297 236
rect 281 202 297 228
rect 331 220 503 236
rect 331 202 469 220
rect 195 178 245 194
rect 195 144 211 178
rect 195 17 245 144
rect 281 146 331 202
rect 453 186 469 202
rect 537 235 1161 238
rect 537 219 742 235
rect 726 201 742 219
rect 776 219 1161 235
rect 776 201 792 219
rect 1145 204 1161 219
rect 1195 204 1211 238
rect 1145 203 1211 204
rect 1247 239 1281 255
rect 726 200 792 201
rect 281 112 297 146
rect 281 96 331 112
rect 367 149 417 168
rect 367 115 383 149
rect 367 17 417 115
rect 453 146 503 186
rect 453 112 469 146
rect 453 96 503 112
rect 539 167 605 185
rect 539 133 555 167
rect 589 133 605 167
rect 828 167 871 185
rect 828 166 832 167
rect 539 17 605 133
rect 640 132 656 166
rect 690 133 832 166
rect 866 133 871 167
rect 690 132 871 133
rect 640 116 871 132
rect 907 169 957 185
rect 1247 169 1281 205
rect 907 135 923 169
rect 1059 135 1075 169
rect 1109 135 1247 169
rect 907 17 957 135
rect 991 101 1025 134
rect 1247 119 1281 135
rect 1317 239 1383 255
rect 1317 205 1333 239
rect 1367 205 1383 239
rect 1317 169 1383 205
rect 1317 135 1333 169
rect 1367 135 1383 169
rect 991 85 1064 101
rect 991 51 1014 85
rect 1048 51 1064 85
rect 1317 17 1383 135
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a22o_4
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 991 94 1025 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 1183298
string GDS_START 1171942
<< end >>
