magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 23 157 351 180
rect 974 157 1608 267
rect 23 49 1608 157
rect 0 0 1632 49
<< scnmos >>
rect 102 70 132 154
rect 242 70 272 154
rect 467 47 497 131
rect 569 47 599 131
rect 641 47 671 131
rect 749 47 779 131
rect 857 47 887 131
rect 1053 73 1083 241
rect 1155 73 1185 241
rect 1241 73 1271 241
rect 1327 73 1357 241
rect 1413 73 1443 241
rect 1499 73 1529 241
<< scpmoshvt >>
rect 102 464 132 592
rect 237 464 267 592
rect 467 469 497 597
rect 621 469 651 597
rect 693 469 723 597
rect 798 469 828 553
rect 873 469 903 553
rect 1053 367 1083 619
rect 1139 367 1169 619
rect 1240 367 1270 619
rect 1326 367 1356 619
rect 1412 367 1442 619
rect 1498 367 1528 619
<< ndiff >>
rect 49 129 102 154
rect 49 95 57 129
rect 91 95 102 129
rect 49 70 102 95
rect 132 118 242 154
rect 132 84 197 118
rect 231 84 242 118
rect 132 70 242 84
rect 272 129 325 154
rect 272 95 283 129
rect 317 95 325 129
rect 272 70 325 95
rect 414 95 467 131
rect 414 61 422 95
rect 456 61 467 95
rect 414 47 467 61
rect 497 92 569 131
rect 497 58 524 92
rect 558 58 569 92
rect 497 47 569 58
rect 599 47 641 131
rect 671 91 749 131
rect 671 57 704 91
rect 738 57 749 91
rect 671 47 749 57
rect 779 47 857 131
rect 887 95 940 131
rect 887 61 898 95
rect 932 61 940 95
rect 887 47 940 61
rect 1000 190 1053 241
rect 1000 156 1008 190
rect 1042 156 1053 190
rect 1000 122 1053 156
rect 1000 88 1008 122
rect 1042 88 1053 122
rect 1000 73 1053 88
rect 1083 73 1155 241
rect 1185 133 1241 241
rect 1185 99 1196 133
rect 1230 99 1241 133
rect 1185 73 1241 99
rect 1271 231 1327 241
rect 1271 197 1282 231
rect 1316 197 1327 231
rect 1271 121 1327 197
rect 1271 87 1282 121
rect 1316 87 1327 121
rect 1271 73 1327 87
rect 1357 163 1413 241
rect 1357 129 1368 163
rect 1402 129 1413 163
rect 1357 73 1413 129
rect 1443 229 1499 241
rect 1443 195 1454 229
rect 1488 195 1499 229
rect 1443 119 1499 195
rect 1443 85 1454 119
rect 1488 85 1499 119
rect 1443 73 1499 85
rect 1529 187 1582 241
rect 1529 153 1540 187
rect 1574 153 1582 187
rect 1529 119 1582 153
rect 1529 85 1540 119
rect 1574 85 1582 119
rect 1529 73 1582 85
<< pdiff >>
rect 49 578 102 592
rect 49 544 57 578
rect 91 544 102 578
rect 49 510 102 544
rect 49 476 57 510
rect 91 476 102 510
rect 49 464 102 476
rect 132 580 237 592
rect 132 546 145 580
rect 179 546 237 580
rect 132 464 237 546
rect 267 517 325 592
rect 267 483 283 517
rect 317 483 325 517
rect 267 464 325 483
rect 414 531 467 597
rect 414 497 422 531
rect 456 497 467 531
rect 414 469 467 497
rect 497 585 621 597
rect 497 551 569 585
rect 603 551 621 585
rect 497 517 621 551
rect 497 483 569 517
rect 603 483 621 517
rect 497 469 621 483
rect 651 469 693 597
rect 723 553 776 597
rect 1000 568 1053 619
rect 1000 553 1008 568
rect 723 527 798 553
rect 723 493 734 527
rect 768 493 798 527
rect 723 469 798 493
rect 828 469 873 553
rect 903 534 1008 553
rect 1042 534 1053 568
rect 903 469 1053 534
rect 1000 367 1053 469
rect 1083 599 1139 619
rect 1083 565 1094 599
rect 1128 565 1139 599
rect 1083 510 1139 565
rect 1083 476 1094 510
rect 1128 476 1139 510
rect 1083 367 1139 476
rect 1169 568 1240 619
rect 1169 534 1186 568
rect 1220 534 1240 568
rect 1169 367 1240 534
rect 1270 599 1326 619
rect 1270 565 1281 599
rect 1315 565 1326 599
rect 1270 503 1326 565
rect 1270 469 1281 503
rect 1315 469 1326 503
rect 1270 413 1326 469
rect 1270 379 1281 413
rect 1315 379 1326 413
rect 1270 367 1326 379
rect 1356 607 1412 619
rect 1356 573 1367 607
rect 1401 573 1412 607
rect 1356 526 1412 573
rect 1356 492 1367 526
rect 1401 492 1412 526
rect 1356 451 1412 492
rect 1356 417 1367 451
rect 1401 417 1412 451
rect 1356 367 1412 417
rect 1442 599 1498 619
rect 1442 565 1453 599
rect 1487 565 1498 599
rect 1442 503 1498 565
rect 1442 469 1453 503
rect 1487 469 1498 503
rect 1442 413 1498 469
rect 1442 379 1453 413
rect 1487 379 1498 413
rect 1442 367 1498 379
rect 1528 607 1581 619
rect 1528 573 1539 607
rect 1573 573 1581 607
rect 1528 526 1581 573
rect 1528 492 1539 526
rect 1573 492 1581 526
rect 1528 451 1581 492
rect 1528 417 1539 451
rect 1573 417 1581 451
rect 1528 367 1581 417
<< ndiffc >>
rect 57 95 91 129
rect 197 84 231 118
rect 283 95 317 129
rect 422 61 456 95
rect 524 58 558 92
rect 704 57 738 91
rect 898 61 932 95
rect 1008 156 1042 190
rect 1008 88 1042 122
rect 1196 99 1230 133
rect 1282 197 1316 231
rect 1282 87 1316 121
rect 1368 129 1402 163
rect 1454 195 1488 229
rect 1454 85 1488 119
rect 1540 153 1574 187
rect 1540 85 1574 119
<< pdiffc >>
rect 57 544 91 578
rect 57 476 91 510
rect 145 546 179 580
rect 283 483 317 517
rect 422 497 456 531
rect 569 551 603 585
rect 569 483 603 517
rect 734 493 768 527
rect 1008 534 1042 568
rect 1094 565 1128 599
rect 1094 476 1128 510
rect 1186 534 1220 568
rect 1281 565 1315 599
rect 1281 469 1315 503
rect 1281 379 1315 413
rect 1367 573 1401 607
rect 1367 492 1401 526
rect 1367 417 1401 451
rect 1453 565 1487 599
rect 1453 469 1487 503
rect 1453 379 1487 413
rect 1539 573 1573 607
rect 1539 492 1573 526
rect 1539 417 1573 451
<< poly >>
rect 102 592 132 618
rect 237 592 267 618
rect 467 597 497 623
rect 621 597 651 623
rect 693 597 723 623
rect 1053 619 1083 645
rect 1139 619 1169 645
rect 1240 619 1270 645
rect 1326 619 1356 645
rect 1412 619 1442 645
rect 1498 619 1528 645
rect 798 553 828 579
rect 873 553 903 579
rect 102 310 132 464
rect 237 310 267 464
rect 327 416 393 432
rect 327 382 343 416
rect 377 382 393 416
rect 327 348 393 382
rect 327 314 343 348
rect 377 328 393 348
rect 467 328 497 469
rect 621 433 651 469
rect 377 314 497 328
rect 102 294 177 310
rect 102 260 127 294
rect 161 260 177 294
rect 102 226 177 260
rect 102 192 127 226
rect 161 192 177 226
rect 102 176 177 192
rect 219 294 285 310
rect 327 298 497 314
rect 539 417 651 433
rect 539 383 555 417
rect 589 383 651 417
rect 539 349 651 383
rect 539 315 555 349
rect 589 315 651 349
rect 539 299 651 315
rect 693 323 723 469
rect 798 437 828 469
rect 873 437 903 469
rect 765 421 831 437
rect 765 387 781 421
rect 815 387 831 421
rect 765 371 831 387
rect 873 421 939 437
rect 873 387 889 421
rect 923 387 939 421
rect 873 371 939 387
rect 219 260 235 294
rect 269 260 285 294
rect 219 226 285 260
rect 219 192 235 226
rect 269 192 285 226
rect 467 219 497 298
rect 563 245 599 299
rect 693 293 779 323
rect 749 265 779 293
rect 219 176 285 192
rect 449 203 515 219
rect 102 154 132 176
rect 242 154 272 176
rect 449 169 465 203
rect 499 169 515 203
rect 449 153 515 169
rect 467 131 497 153
rect 569 131 599 245
rect 641 235 707 251
rect 641 201 657 235
rect 691 201 707 235
rect 641 185 707 201
rect 749 249 815 265
rect 749 215 765 249
rect 799 215 815 249
rect 749 199 815 215
rect 641 131 671 185
rect 749 131 779 199
rect 873 183 903 371
rect 1053 345 1083 367
rect 981 329 1083 345
rect 1139 329 1169 367
rect 1240 345 1270 367
rect 1326 345 1356 367
rect 1412 345 1442 367
rect 1498 345 1528 367
rect 1240 331 1528 345
rect 945 315 1083 329
rect 945 313 1011 315
rect 945 279 961 313
rect 995 279 1011 313
rect 945 263 1011 279
rect 1125 313 1191 329
rect 1125 279 1141 313
rect 1175 279 1191 313
rect 857 153 903 183
rect 857 131 887 153
rect 102 44 132 70
rect 242 44 272 70
rect 955 51 985 263
rect 1053 241 1083 267
rect 1125 263 1191 279
rect 1233 315 1528 331
rect 1233 281 1249 315
rect 1283 281 1317 315
rect 1351 281 1385 315
rect 1419 295 1528 315
rect 1419 281 1529 295
rect 1233 265 1529 281
rect 1155 241 1185 263
rect 1241 241 1271 265
rect 1327 241 1357 265
rect 1413 241 1443 265
rect 1499 241 1529 265
rect 1053 51 1083 73
rect 467 21 497 47
rect 569 21 599 47
rect 641 21 671 47
rect 749 21 779 47
rect 857 21 887 47
rect 955 21 1083 51
rect 1155 47 1185 73
rect 1241 47 1271 73
rect 1327 47 1357 73
rect 1413 47 1443 73
rect 1499 47 1529 73
<< polycont >>
rect 343 382 377 416
rect 343 314 377 348
rect 127 260 161 294
rect 127 192 161 226
rect 555 383 589 417
rect 555 315 589 349
rect 781 387 815 421
rect 889 387 923 421
rect 235 260 269 294
rect 235 192 269 226
rect 465 169 499 203
rect 657 201 691 235
rect 765 215 799 249
rect 961 279 995 313
rect 1141 279 1175 313
rect 1249 281 1283 315
rect 1317 281 1351 315
rect 1385 281 1419 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 41 578 95 594
rect 41 544 57 578
rect 91 544 95 578
rect 41 510 95 544
rect 129 580 179 649
rect 129 546 145 580
rect 129 528 179 546
rect 213 581 533 615
rect 41 476 57 510
rect 91 494 95 510
rect 213 494 247 581
rect 91 476 247 494
rect 41 460 247 476
rect 281 517 343 533
rect 281 483 283 517
rect 317 483 343 517
rect 281 460 343 483
rect 406 531 465 547
rect 406 497 422 531
rect 456 497 465 531
rect 406 481 465 497
rect 41 129 91 460
rect 309 431 343 460
rect 41 95 57 129
rect 41 79 91 95
rect 125 294 175 426
rect 125 260 127 294
rect 161 260 175 294
rect 125 226 175 260
rect 125 192 127 226
rect 161 192 175 226
rect 125 168 175 192
rect 209 294 275 426
rect 209 260 235 294
rect 269 260 275 294
rect 209 226 275 260
rect 209 192 235 226
rect 269 192 275 226
rect 209 168 275 192
rect 309 416 393 431
rect 309 382 343 416
rect 377 382 393 416
rect 309 348 393 382
rect 309 314 343 348
rect 377 314 393 348
rect 309 307 393 314
rect 125 94 161 168
rect 309 134 343 307
rect 429 273 465 481
rect 499 433 533 581
rect 567 585 607 649
rect 567 551 569 585
rect 603 551 607 585
rect 567 517 607 551
rect 567 483 569 517
rect 603 483 607 517
rect 567 467 607 483
rect 641 577 842 615
rect 499 417 605 433
rect 499 383 555 417
rect 589 383 605 417
rect 499 349 605 383
rect 499 315 555 349
rect 589 315 605 349
rect 499 307 605 315
rect 641 273 675 577
rect 711 527 774 543
rect 711 493 734 527
rect 768 493 774 527
rect 711 477 774 493
rect 711 329 745 477
rect 808 437 842 577
rect 992 568 1058 649
rect 992 534 1008 568
rect 1042 534 1058 568
rect 992 526 1058 534
rect 1092 599 1132 615
rect 1092 565 1094 599
rect 1128 565 1132 599
rect 1092 510 1132 565
rect 1170 568 1236 649
rect 1170 534 1186 568
rect 1220 534 1236 568
rect 1170 526 1236 534
rect 1279 599 1317 615
rect 1279 565 1281 599
rect 1315 565 1317 599
rect 1092 492 1094 510
rect 779 421 842 437
rect 779 387 781 421
rect 815 387 842 421
rect 779 371 842 387
rect 876 476 1094 492
rect 1128 492 1132 510
rect 1279 503 1317 565
rect 1128 476 1245 492
rect 876 458 1245 476
rect 876 421 939 458
rect 876 387 889 421
rect 923 387 939 421
rect 876 371 939 387
rect 711 313 1011 329
rect 711 295 961 313
rect 195 118 233 134
rect 195 84 197 118
rect 231 84 233 118
rect 195 17 233 84
rect 267 129 343 134
rect 267 95 283 129
rect 317 95 343 129
rect 267 79 343 95
rect 379 251 675 273
rect 851 279 961 295
rect 995 279 1011 313
rect 851 263 1011 279
rect 1063 313 1177 424
rect 1063 279 1141 313
rect 1175 279 1177 313
rect 379 239 707 251
rect 379 97 413 239
rect 641 235 707 239
rect 449 203 515 205
rect 449 169 465 203
rect 499 169 515 203
rect 641 201 657 235
rect 691 201 707 235
rect 641 199 707 201
rect 749 249 815 261
rect 749 215 765 249
rect 799 215 815 249
rect 749 213 815 215
rect 449 165 515 169
rect 749 165 783 213
rect 851 179 885 263
rect 1063 242 1177 279
rect 1211 315 1245 458
rect 1279 469 1281 503
rect 1315 469 1317 503
rect 1279 413 1317 469
rect 1351 607 1417 649
rect 1351 573 1367 607
rect 1401 573 1417 607
rect 1351 526 1417 573
rect 1351 492 1367 526
rect 1401 492 1417 526
rect 1351 451 1417 492
rect 1351 417 1367 451
rect 1401 417 1417 451
rect 1451 599 1489 615
rect 1451 565 1453 599
rect 1487 565 1489 599
rect 1451 503 1489 565
rect 1451 469 1453 503
rect 1487 469 1489 503
rect 1279 379 1281 413
rect 1315 383 1317 413
rect 1451 413 1489 469
rect 1523 607 1589 649
rect 1523 573 1539 607
rect 1573 573 1589 607
rect 1523 526 1589 573
rect 1523 492 1539 526
rect 1573 492 1589 526
rect 1523 451 1589 492
rect 1523 417 1539 451
rect 1573 417 1589 451
rect 1451 383 1453 413
rect 1315 379 1453 383
rect 1487 383 1489 413
rect 1487 379 1615 383
rect 1279 349 1615 379
rect 1211 281 1249 315
rect 1283 281 1317 315
rect 1351 281 1385 315
rect 1419 281 1435 315
rect 1211 208 1246 281
rect 1469 247 1615 349
rect 449 131 783 165
rect 817 145 885 179
rect 1004 190 1246 208
rect 1004 156 1008 190
rect 1042 174 1246 190
rect 1280 231 1615 247
rect 1280 197 1282 231
rect 1316 229 1615 231
rect 1316 213 1454 229
rect 1316 197 1325 213
rect 1042 156 1046 174
rect 817 97 853 145
rect 1004 122 1046 156
rect 379 95 472 97
rect 379 61 422 95
rect 456 61 472 95
rect 379 57 472 61
rect 508 92 574 97
rect 508 58 524 92
rect 558 58 574 92
rect 508 17 574 58
rect 688 91 853 97
rect 688 57 704 91
rect 738 57 853 91
rect 688 53 853 57
rect 887 95 948 111
rect 887 61 898 95
rect 932 61 948 95
rect 1004 88 1008 122
rect 1042 88 1046 122
rect 1004 72 1046 88
rect 1180 133 1246 140
rect 1180 99 1196 133
rect 1230 99 1246 133
rect 887 17 948 61
rect 1180 17 1246 99
rect 1280 121 1325 197
rect 1445 195 1454 213
rect 1488 221 1615 229
rect 1488 211 1499 221
rect 1488 195 1490 211
rect 1280 87 1282 121
rect 1316 87 1325 121
rect 1280 71 1325 87
rect 1359 163 1411 179
rect 1359 129 1368 163
rect 1402 129 1411 163
rect 1359 17 1411 129
rect 1445 119 1490 195
rect 1445 85 1454 119
rect 1488 85 1490 119
rect 1445 69 1490 85
rect 1524 153 1540 187
rect 1574 153 1590 187
rect 1524 119 1590 153
rect 1524 85 1540 119
rect 1574 85 1590 119
rect 1524 17 1590 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrtp_4
flabel comment s 442 315 442 315 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1087 390 1121 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1922682
string GDS_START 1909410
<< end >>
