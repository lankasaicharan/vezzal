magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 4274 1975
<< nwell >>
rect -38 356 3014 704
rect -38 332 797 356
rect 1167 332 3014 356
rect 1625 311 1929 332
<< pwell >>
rect 830 248 1125 293
rect 830 228 1726 248
rect 830 206 1821 228
rect 811 191 1821 206
rect 199 184 1821 191
rect 2313 184 2975 248
rect 1 49 2975 184
rect 0 0 2976 49
<< scnmos >>
rect 84 74 114 158
rect 282 81 312 165
rect 385 81 415 165
rect 542 81 572 165
rect 614 81 644 165
rect 700 81 730 165
rect 906 119 936 267
rect 1016 119 1046 267
rect 1206 138 1236 222
rect 1292 138 1322 222
rect 1367 138 1397 222
rect 1445 138 1475 222
rect 1620 74 1650 222
rect 1715 74 1745 202
rect 1925 74 1955 158
rect 2003 74 2033 158
rect 2111 74 2141 158
rect 2183 74 2213 158
rect 2396 74 2426 222
rect 2482 74 2512 222
rect 2568 74 2598 222
rect 2776 74 2806 222
rect 2862 74 2892 222
<< scpmoshvt >>
rect 86 464 116 592
rect 310 464 340 592
rect 394 464 424 592
rect 484 464 514 592
rect 592 464 622 592
rect 706 464 736 592
rect 914 392 944 592
rect 1004 392 1034 592
rect 1212 463 1242 547
rect 1312 463 1342 547
rect 1390 463 1420 547
rect 1518 463 1548 547
rect 1720 347 1750 547
rect 1810 347 1840 547
rect 1952 508 1982 592
rect 2036 508 2066 592
rect 2173 508 2203 592
rect 2280 508 2310 592
rect 2393 368 2423 536
rect 2483 368 2513 536
rect 2590 368 2620 592
rect 2680 368 2710 592
rect 2770 368 2800 592
rect 2860 368 2890 592
<< ndiff >>
rect 856 180 906 267
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 128 171 158
rect 114 94 125 128
rect 159 94 171 128
rect 114 74 171 94
rect 225 127 282 165
rect 225 93 237 127
rect 271 93 282 127
rect 225 81 282 93
rect 312 81 385 165
rect 415 153 542 165
rect 415 119 483 153
rect 517 119 542 153
rect 415 81 542 119
rect 572 81 614 165
rect 644 134 700 165
rect 644 100 655 134
rect 689 100 700 134
rect 644 81 700 100
rect 730 134 783 165
rect 730 100 741 134
rect 775 100 783 134
rect 730 81 783 100
rect 837 150 906 180
rect 837 116 849 150
rect 883 119 906 150
rect 936 150 1016 267
rect 936 119 959 150
rect 883 116 891 119
rect 837 98 891 116
rect 951 116 959 119
rect 993 119 1016 150
rect 1046 234 1099 267
rect 1046 200 1057 234
rect 1091 200 1099 234
rect 1046 166 1099 200
rect 1046 132 1057 166
rect 1091 132 1099 166
rect 1153 197 1206 222
rect 1153 163 1161 197
rect 1195 163 1206 197
rect 1153 138 1206 163
rect 1236 191 1292 222
rect 1236 157 1247 191
rect 1281 157 1292 191
rect 1236 138 1292 157
rect 1322 138 1367 222
rect 1397 138 1445 222
rect 1475 138 1620 222
rect 1046 119 1099 132
rect 993 116 1001 119
rect 951 98 1001 116
rect 1490 82 1620 138
rect 1490 48 1502 82
rect 1536 74 1620 82
rect 1650 202 1700 222
rect 1650 179 1715 202
rect 1650 145 1670 179
rect 1704 145 1715 179
rect 1650 74 1715 145
rect 1745 158 1795 202
rect 2339 210 2396 222
rect 2339 176 2351 210
rect 2385 176 2396 210
rect 1745 131 1925 158
rect 1745 97 1864 131
rect 1898 97 1925 131
rect 1745 74 1925 97
rect 1955 74 2003 158
rect 2033 120 2111 158
rect 2033 86 2055 120
rect 2089 86 2111 120
rect 2033 74 2111 86
rect 2141 74 2183 158
rect 2213 127 2285 158
rect 2213 93 2231 127
rect 2265 93 2285 127
rect 2213 74 2285 93
rect 2339 120 2396 176
rect 2339 86 2351 120
rect 2385 86 2396 120
rect 2339 74 2396 86
rect 2426 204 2482 222
rect 2426 170 2437 204
rect 2471 170 2482 204
rect 2426 120 2482 170
rect 2426 86 2437 120
rect 2471 86 2482 120
rect 2426 74 2482 86
rect 2512 204 2568 222
rect 2512 170 2523 204
rect 2557 170 2568 204
rect 2512 120 2568 170
rect 2512 86 2523 120
rect 2557 86 2568 120
rect 2512 74 2568 86
rect 2598 136 2776 222
rect 2598 102 2609 136
rect 2643 102 2731 136
rect 2765 102 2776 136
rect 2598 74 2776 102
rect 2806 210 2862 222
rect 2806 176 2817 210
rect 2851 176 2862 210
rect 2806 120 2862 176
rect 2806 86 2817 120
rect 2851 86 2862 120
rect 2806 74 2862 86
rect 2892 210 2949 222
rect 2892 176 2903 210
rect 2937 176 2949 210
rect 2892 120 2949 176
rect 2892 86 2903 120
rect 2937 86 2949 120
rect 2892 74 2949 86
rect 1536 48 1548 74
rect 1490 36 1548 48
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 464 86 476
rect 116 580 310 592
rect 116 546 139 580
rect 173 546 263 580
rect 297 546 310 580
rect 116 510 310 546
rect 116 476 139 510
rect 173 476 263 510
rect 297 476 310 510
rect 116 464 310 476
rect 340 464 394 592
rect 424 580 484 592
rect 424 546 437 580
rect 471 546 484 580
rect 424 510 484 546
rect 424 476 437 510
rect 471 476 484 510
rect 424 464 484 476
rect 514 464 592 592
rect 622 575 706 592
rect 622 541 635 575
rect 669 541 706 575
rect 622 464 706 541
rect 736 580 795 592
rect 736 546 749 580
rect 783 546 795 580
rect 736 510 795 546
rect 736 476 749 510
rect 783 476 795 510
rect 736 464 795 476
rect 855 434 914 592
rect 855 400 867 434
rect 901 400 914 434
rect 855 392 914 400
rect 944 584 1004 592
rect 944 550 957 584
rect 991 550 1004 584
rect 944 392 1004 550
rect 1034 434 1093 592
rect 1034 400 1047 434
rect 1081 400 1093 434
rect 1034 392 1093 400
rect 1438 582 1500 594
rect 1438 548 1452 582
rect 1486 548 1500 582
rect 1438 547 1500 548
rect 1858 560 1952 592
rect 1858 547 1887 560
rect 1153 522 1212 547
rect 1153 488 1165 522
rect 1199 488 1212 522
rect 1153 463 1212 488
rect 1242 535 1312 547
rect 1242 501 1265 535
rect 1299 501 1312 535
rect 1242 463 1312 501
rect 1342 463 1390 547
rect 1420 463 1518 547
rect 1548 524 1607 547
rect 1548 490 1561 524
rect 1595 490 1607 524
rect 1548 463 1607 490
rect 1661 535 1720 547
rect 1661 501 1673 535
rect 1707 501 1720 535
rect 1661 467 1720 501
rect 1661 433 1673 467
rect 1707 433 1720 467
rect 1661 399 1720 433
rect 1661 365 1673 399
rect 1707 365 1720 399
rect 1661 347 1720 365
rect 1750 535 1810 547
rect 1750 501 1763 535
rect 1797 501 1810 535
rect 1750 464 1810 501
rect 1750 430 1763 464
rect 1797 430 1810 464
rect 1750 393 1810 430
rect 1750 359 1763 393
rect 1797 359 1810 393
rect 1750 347 1810 359
rect 1840 526 1887 547
rect 1921 526 1952 560
rect 1840 508 1952 526
rect 1982 508 2036 592
rect 2066 567 2173 592
rect 2066 533 2109 567
rect 2143 533 2173 567
rect 2066 508 2173 533
rect 2203 567 2280 592
rect 2203 533 2216 567
rect 2250 533 2280 567
rect 2203 508 2280 533
rect 2310 536 2375 592
rect 2531 580 2590 592
rect 2531 546 2543 580
rect 2577 546 2590 580
rect 2531 536 2590 546
rect 2310 524 2393 536
rect 2310 508 2346 524
rect 1840 347 1893 508
rect 2333 490 2346 508
rect 2380 490 2393 524
rect 2333 414 2393 490
rect 2333 380 2346 414
rect 2380 380 2393 414
rect 2333 368 2393 380
rect 2423 524 2483 536
rect 2423 490 2436 524
rect 2470 490 2483 524
rect 2423 414 2483 490
rect 2423 380 2436 414
rect 2470 380 2483 414
rect 2423 368 2483 380
rect 2513 497 2590 536
rect 2513 463 2543 497
rect 2577 463 2590 497
rect 2513 414 2590 463
rect 2513 380 2543 414
rect 2577 380 2590 414
rect 2513 368 2590 380
rect 2620 580 2680 592
rect 2620 546 2633 580
rect 2667 546 2680 580
rect 2620 497 2680 546
rect 2620 463 2633 497
rect 2667 463 2680 497
rect 2620 414 2680 463
rect 2620 380 2633 414
rect 2667 380 2680 414
rect 2620 368 2680 380
rect 2710 580 2770 592
rect 2710 546 2723 580
rect 2757 546 2770 580
rect 2710 472 2770 546
rect 2710 438 2723 472
rect 2757 438 2770 472
rect 2710 368 2770 438
rect 2800 580 2860 592
rect 2800 546 2813 580
rect 2847 546 2860 580
rect 2800 497 2860 546
rect 2800 463 2813 497
rect 2847 463 2860 497
rect 2800 414 2860 463
rect 2800 380 2813 414
rect 2847 380 2860 414
rect 2800 368 2860 380
rect 2890 580 2949 592
rect 2890 546 2903 580
rect 2937 546 2949 580
rect 2890 472 2949 546
rect 2890 438 2903 472
rect 2937 438 2949 472
rect 2890 368 2949 438
<< ndiffc >>
rect 39 99 73 133
rect 125 94 159 128
rect 237 93 271 127
rect 483 119 517 153
rect 655 100 689 134
rect 741 100 775 134
rect 849 116 883 150
rect 959 116 993 150
rect 1057 200 1091 234
rect 1057 132 1091 166
rect 1161 163 1195 197
rect 1247 157 1281 191
rect 1502 48 1536 82
rect 1670 145 1704 179
rect 2351 176 2385 210
rect 1864 97 1898 131
rect 2055 86 2089 120
rect 2231 93 2265 127
rect 2351 86 2385 120
rect 2437 170 2471 204
rect 2437 86 2471 120
rect 2523 170 2557 204
rect 2523 86 2557 120
rect 2609 102 2643 136
rect 2731 102 2765 136
rect 2817 176 2851 210
rect 2817 86 2851 120
rect 2903 176 2937 210
rect 2903 86 2937 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 139 546 173 580
rect 263 546 297 580
rect 139 476 173 510
rect 263 476 297 510
rect 437 546 471 580
rect 437 476 471 510
rect 635 541 669 575
rect 749 546 783 580
rect 749 476 783 510
rect 867 400 901 434
rect 957 550 991 584
rect 1047 400 1081 434
rect 1452 548 1486 582
rect 1165 488 1199 522
rect 1265 501 1299 535
rect 1561 490 1595 524
rect 1673 501 1707 535
rect 1673 433 1707 467
rect 1673 365 1707 399
rect 1763 501 1797 535
rect 1763 430 1797 464
rect 1763 359 1797 393
rect 1887 526 1921 560
rect 2109 533 2143 567
rect 2216 533 2250 567
rect 2543 546 2577 580
rect 2346 490 2380 524
rect 2346 380 2380 414
rect 2436 490 2470 524
rect 2436 380 2470 414
rect 2543 463 2577 497
rect 2543 380 2577 414
rect 2633 546 2667 580
rect 2633 463 2667 497
rect 2633 380 2667 414
rect 2723 546 2757 580
rect 2723 438 2757 472
rect 2813 546 2847 580
rect 2813 463 2847 497
rect 2813 380 2847 414
rect 2903 546 2937 580
rect 2903 438 2937 472
<< poly >>
rect 86 592 116 618
rect 310 592 340 618
rect 394 592 424 618
rect 484 592 514 618
rect 592 592 622 618
rect 706 592 736 618
rect 914 592 944 618
rect 1004 592 1034 618
rect 1108 615 1843 645
rect 86 449 116 464
rect 310 449 340 464
rect 394 449 424 464
rect 484 449 514 464
rect 592 449 622 464
rect 706 449 736 464
rect 83 367 119 449
rect 307 367 343 449
rect 83 351 343 367
rect 83 317 137 351
rect 171 317 205 351
rect 239 317 273 351
rect 307 317 343 351
rect 83 301 343 317
rect 84 158 114 301
rect 391 253 427 449
rect 481 432 517 449
rect 474 416 540 432
rect 474 382 490 416
rect 524 382 540 416
rect 474 366 540 382
rect 588 422 625 449
rect 696 432 739 449
rect 588 406 654 422
rect 588 372 604 406
rect 638 372 654 406
rect 588 338 654 372
rect 162 237 228 253
rect 162 203 178 237
rect 212 217 228 237
rect 354 237 427 253
rect 480 302 546 318
rect 480 268 496 302
rect 530 268 546 302
rect 588 304 604 338
rect 638 304 654 338
rect 588 288 654 304
rect 696 416 823 432
rect 696 382 773 416
rect 807 382 823 416
rect 696 366 823 382
rect 480 252 546 268
rect 212 203 312 217
rect 162 187 312 203
rect 354 203 370 237
rect 404 203 427 237
rect 516 240 546 252
rect 516 210 572 240
rect 354 187 427 203
rect 282 165 312 187
rect 385 165 415 187
rect 542 165 572 210
rect 614 165 644 288
rect 696 212 726 366
rect 914 360 944 392
rect 1004 360 1034 392
rect 865 324 944 360
rect 768 308 944 324
rect 768 274 784 308
rect 818 282 944 308
rect 990 339 1056 360
rect 990 305 1006 339
rect 1040 312 1056 339
rect 1108 312 1138 615
rect 1212 547 1242 573
rect 1309 562 1345 615
rect 1312 547 1342 562
rect 1390 547 1420 573
rect 1518 547 1548 573
rect 1720 547 1750 573
rect 1807 562 1843 615
rect 1952 592 1982 618
rect 2036 592 2066 618
rect 2173 592 2203 618
rect 2280 592 2310 618
rect 2590 592 2620 618
rect 2680 592 2710 618
rect 2770 592 2800 618
rect 2860 592 2890 618
rect 1810 547 1840 562
rect 1212 448 1242 463
rect 1209 383 1245 448
rect 1312 437 1342 463
rect 1390 448 1420 463
rect 1518 448 1548 463
rect 1387 389 1423 448
rect 1515 430 1551 448
rect 1515 414 1629 430
rect 1180 367 1246 383
rect 1180 333 1196 367
rect 1230 347 1246 367
rect 1367 373 1471 389
rect 1230 333 1322 347
rect 1180 317 1322 333
rect 1040 305 1138 312
rect 990 300 1138 305
rect 990 295 1141 300
rect 990 282 1144 295
rect 818 274 834 282
rect 768 258 834 274
rect 906 267 936 282
rect 1016 267 1046 282
rect 1110 278 1144 282
rect 1114 267 1144 278
rect 696 193 730 212
rect 700 165 730 193
rect 906 93 936 119
rect 1114 237 1236 267
rect 1206 222 1236 237
rect 1292 222 1322 317
rect 1367 339 1421 373
rect 1455 339 1471 373
rect 1515 380 1579 414
rect 1613 380 1629 414
rect 1515 364 1629 380
rect 1367 323 1471 339
rect 1367 222 1397 323
rect 1519 267 1549 364
rect 2393 536 2423 562
rect 2483 536 2513 562
rect 1952 493 1982 508
rect 2036 493 2066 508
rect 2173 493 2203 508
rect 2280 493 2310 508
rect 1949 476 1985 493
rect 1925 460 1991 476
rect 1925 426 1941 460
rect 1975 426 1991 460
rect 1925 410 1991 426
rect 1720 332 1750 347
rect 1810 332 1840 347
rect 1717 319 1753 332
rect 1445 237 1549 267
rect 1597 299 1753 319
rect 1807 302 1955 332
rect 2033 311 2069 493
rect 2170 430 2206 493
rect 1597 265 1613 299
rect 1647 289 1753 299
rect 1647 265 1663 289
rect 1597 249 1663 265
rect 1445 222 1475 237
rect 1620 222 1650 249
rect 1715 231 1883 247
rect 1016 93 1046 119
rect 1206 112 1236 138
rect 1292 112 1322 138
rect 1367 112 1397 138
rect 84 48 114 74
rect 282 55 312 81
rect 385 55 415 81
rect 542 55 572 81
rect 614 55 644 81
rect 700 51 730 81
rect 1445 51 1475 138
rect 700 21 1475 51
rect 1715 217 1833 231
rect 1715 202 1745 217
rect 1817 197 1833 217
rect 1867 197 1883 231
rect 1817 181 1883 197
rect 1925 158 1955 302
rect 2003 295 2069 311
rect 2003 261 2019 295
rect 2053 261 2069 295
rect 2003 245 2069 261
rect 2111 414 2206 430
rect 2111 380 2133 414
rect 2167 380 2206 414
rect 2111 364 2206 380
rect 2003 158 2033 245
rect 2111 158 2141 364
rect 2277 315 2313 493
rect 2393 353 2423 368
rect 2483 353 2513 368
rect 2590 353 2620 368
rect 2680 353 2710 368
rect 2770 353 2800 368
rect 2860 353 2890 368
rect 2390 323 2516 353
rect 2277 267 2307 315
rect 2396 267 2426 323
rect 2587 320 2623 353
rect 2677 320 2713 353
rect 2767 320 2803 353
rect 2857 320 2893 353
rect 2568 304 2893 320
rect 2568 275 2584 304
rect 2183 237 2426 267
rect 2183 230 2307 237
rect 2183 196 2199 230
rect 2233 196 2307 230
rect 2396 222 2426 237
rect 2482 270 2584 275
rect 2618 270 2652 304
rect 2686 270 2720 304
rect 2754 290 2893 304
rect 2754 270 2892 290
rect 2482 245 2892 270
rect 2482 222 2512 245
rect 2568 222 2598 245
rect 2776 222 2806 245
rect 2862 222 2892 245
rect 2183 180 2307 196
rect 2183 158 2213 180
rect 1620 48 1650 74
rect 1715 48 1745 74
rect 1925 48 1955 74
rect 2003 48 2033 74
rect 2111 48 2141 74
rect 2183 48 2213 74
rect 2396 48 2426 74
rect 2482 48 2512 74
rect 2568 48 2598 74
rect 2776 48 2806 74
rect 2862 48 2892 74
<< polycont >>
rect 137 317 171 351
rect 205 317 239 351
rect 273 317 307 351
rect 490 382 524 416
rect 604 372 638 406
rect 178 203 212 237
rect 496 268 530 302
rect 604 304 638 338
rect 773 382 807 416
rect 370 203 404 237
rect 784 274 818 308
rect 1006 305 1040 339
rect 1196 333 1230 367
rect 1421 339 1455 373
rect 1579 380 1613 414
rect 1941 426 1975 460
rect 1613 265 1647 299
rect 1833 197 1867 231
rect 2019 261 2053 295
rect 2133 380 2167 414
rect 2199 196 2233 230
rect 2584 270 2618 304
rect 2652 270 2686 304
rect 2720 270 2754 304
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 435 89 476
rect 123 580 313 649
rect 123 546 139 580
rect 173 546 263 580
rect 297 546 313 580
rect 123 510 313 546
rect 123 476 139 510
rect 173 476 263 510
rect 297 476 313 510
rect 123 469 313 476
rect 421 580 487 596
rect 421 546 437 580
rect 471 546 487 580
rect 421 510 487 546
rect 619 575 685 649
rect 619 541 635 575
rect 669 541 685 575
rect 619 537 685 541
rect 723 580 799 596
rect 723 546 749 580
rect 783 546 799 580
rect 941 584 1007 649
rect 941 550 957 584
rect 991 550 1007 584
rect 1434 582 1504 649
rect 421 476 437 510
rect 471 503 487 510
rect 723 518 799 546
rect 1149 522 1215 551
rect 723 516 929 518
rect 1149 516 1165 522
rect 723 510 1165 516
rect 723 503 749 510
rect 471 476 749 503
rect 783 488 1165 510
rect 1199 488 1215 522
rect 783 484 1215 488
rect 1249 535 1377 551
rect 1249 501 1265 535
rect 1299 501 1377 535
rect 1434 548 1452 582
rect 1486 548 1504 582
rect 1434 532 1504 548
rect 1249 498 1377 501
rect 1545 524 1611 551
rect 1545 498 1561 524
rect 1249 490 1561 498
rect 1595 490 1611 524
rect 1249 485 1611 490
rect 783 476 799 484
rect 916 482 1215 484
rect 421 469 799 476
rect 689 466 799 469
rect 23 416 541 435
rect 23 401 490 416
rect 23 253 57 401
rect 475 382 490 401
rect 524 382 541 416
rect 121 351 359 367
rect 475 366 541 382
rect 589 406 655 430
rect 589 372 604 406
rect 638 372 655 406
rect 121 317 137 351
rect 171 317 205 351
rect 239 317 273 351
rect 307 332 359 351
rect 589 338 655 372
rect 307 317 547 332
rect 121 302 547 317
rect 121 298 496 302
rect 481 268 496 298
rect 530 268 547 302
rect 589 304 604 338
rect 638 304 655 338
rect 589 288 655 304
rect 23 237 228 253
rect 23 203 178 237
rect 212 203 228 237
rect 23 187 228 203
rect 313 237 420 253
rect 481 252 547 268
rect 313 203 370 237
rect 404 203 420 237
rect 689 218 723 466
rect 1165 451 1215 482
rect 1343 464 1611 485
rect 1673 535 1707 649
rect 1854 560 2059 576
rect 1673 467 1707 501
rect 867 434 903 450
rect 757 424 833 432
rect 757 416 799 424
rect 757 382 773 416
rect 807 382 833 390
rect 757 366 833 382
rect 901 400 903 434
rect 867 398 903 400
rect 1031 434 1131 448
rect 1031 400 1047 434
rect 1081 400 1131 434
rect 1165 417 1309 451
rect 867 364 995 398
rect 1031 383 1131 400
rect 1031 382 1241 383
rect 961 348 995 364
rect 1090 367 1241 382
rect 961 339 1056 348
rect 768 308 927 318
rect 768 274 784 308
rect 818 274 927 308
rect 768 252 927 274
rect 961 305 1006 339
rect 1040 305 1056 339
rect 961 282 1056 305
rect 1090 333 1196 367
rect 1230 333 1241 367
rect 1090 317 1241 333
rect 768 236 839 252
rect 961 218 995 282
rect 1090 248 1124 317
rect 1275 283 1309 417
rect 23 133 73 187
rect 313 162 420 203
rect 513 184 723 218
rect 873 184 995 218
rect 1039 234 1124 248
rect 1039 200 1057 234
rect 1091 200 1124 234
rect 1039 184 1124 200
rect 513 169 547 184
rect 454 153 547 169
rect 23 99 39 133
rect 23 70 73 99
rect 109 128 175 153
rect 109 94 125 128
rect 159 94 175 128
rect 109 17 175 94
rect 221 127 287 128
rect 221 93 237 127
rect 271 93 287 127
rect 454 119 483 153
rect 517 119 547 153
rect 873 150 907 184
rect 1043 166 1124 184
rect 645 134 700 150
rect 221 85 287 93
rect 645 100 655 134
rect 689 100 700 134
rect 645 85 700 100
rect 221 51 700 85
rect 734 134 799 150
rect 734 100 741 134
rect 775 100 799 134
rect 833 116 849 150
rect 883 116 907 150
rect 833 110 907 116
rect 943 116 959 150
rect 993 116 1009 150
rect 734 17 799 100
rect 943 17 1009 116
rect 1043 132 1057 166
rect 1091 132 1124 166
rect 1158 249 1309 283
rect 1158 197 1198 249
rect 1343 215 1377 464
rect 1158 163 1161 197
rect 1195 163 1198 197
rect 1158 134 1198 163
rect 1232 191 1377 215
rect 1232 157 1247 191
rect 1281 181 1377 191
rect 1411 373 1465 389
rect 1411 339 1421 373
rect 1455 339 1465 373
rect 1411 218 1465 339
rect 1499 315 1533 464
rect 1567 424 1629 430
rect 1601 414 1629 424
rect 1567 380 1579 390
rect 1613 380 1629 414
rect 1567 364 1629 380
rect 1673 399 1707 433
rect 1673 349 1707 365
rect 1747 535 1813 551
rect 1747 501 1763 535
rect 1797 501 1813 535
rect 1854 526 1887 560
rect 1921 526 2059 560
rect 1854 510 2059 526
rect 1747 464 1813 501
rect 1747 430 1763 464
rect 1797 430 1813 464
rect 1747 393 1813 430
rect 1747 359 1763 393
rect 1797 359 1813 393
rect 1747 315 1813 359
rect 1499 299 1663 315
rect 1499 265 1613 299
rect 1647 265 1663 299
rect 1499 252 1663 265
rect 1697 281 1813 315
rect 1849 460 1991 476
rect 1849 426 1941 460
rect 1975 426 1991 460
rect 1849 413 1991 426
rect 1697 218 1731 281
rect 1849 247 1883 413
rect 2025 379 2059 510
rect 2093 567 2159 649
rect 2093 533 2109 567
rect 2143 533 2159 567
rect 2093 504 2159 533
rect 2200 567 2266 596
rect 2200 533 2216 567
rect 2250 533 2266 567
rect 2200 504 2266 533
rect 1411 184 1731 218
rect 1281 157 1294 181
rect 1232 134 1294 157
rect 1654 179 1731 184
rect 1043 100 1124 132
rect 1411 116 1620 150
rect 1654 145 1670 179
rect 1704 145 1731 179
rect 1654 119 1731 145
rect 1765 231 1883 247
rect 1765 197 1833 231
rect 1867 197 1883 231
rect 1765 181 1883 197
rect 1917 345 2059 379
rect 2117 424 2183 430
rect 2117 414 2143 424
rect 2117 380 2133 414
rect 2177 390 2183 424
rect 2167 380 2183 390
rect 2117 364 2183 380
rect 1917 211 1951 345
rect 2232 311 2266 504
rect 2330 524 2380 649
rect 2527 580 2577 649
rect 2527 546 2543 580
rect 2330 490 2346 524
rect 2330 414 2380 490
rect 2330 380 2346 414
rect 2330 364 2380 380
rect 2420 524 2486 540
rect 2420 490 2436 524
rect 2470 490 2486 524
rect 2420 414 2486 490
rect 2420 380 2436 414
rect 2470 380 2486 414
rect 2420 320 2486 380
rect 2527 497 2577 546
rect 2527 463 2543 497
rect 2527 414 2577 463
rect 2527 380 2543 414
rect 2527 364 2577 380
rect 2617 580 2683 596
rect 2617 546 2633 580
rect 2667 546 2683 580
rect 2617 497 2683 546
rect 2617 463 2633 497
rect 2667 463 2683 497
rect 2617 414 2683 463
rect 2723 580 2773 649
rect 2757 546 2773 580
rect 2723 472 2773 546
rect 2757 438 2773 472
rect 2723 422 2773 438
rect 2813 580 2856 596
rect 2847 546 2856 580
rect 2813 497 2856 546
rect 2847 463 2856 497
rect 2617 380 2633 414
rect 2667 388 2683 414
rect 2813 414 2856 463
rect 2894 580 2953 649
rect 2894 546 2903 580
rect 2937 546 2953 580
rect 2894 472 2953 546
rect 2894 438 2903 472
rect 2937 438 2953 472
rect 2894 422 2953 438
rect 2667 380 2813 388
rect 2847 388 2856 414
rect 2847 380 2951 388
rect 2617 354 2951 380
rect 2003 295 2317 311
rect 2003 261 2019 295
rect 2053 277 2317 295
rect 2053 261 2069 277
rect 2003 245 2069 261
rect 2183 230 2249 243
rect 2183 211 2199 230
rect 1917 196 2199 211
rect 2233 196 2249 230
rect 1411 100 1445 116
rect 1043 66 1445 100
rect 1586 85 1620 116
rect 1765 85 1799 181
rect 1917 177 2249 196
rect 1917 147 1951 177
rect 1486 48 1502 82
rect 1536 48 1552 82
rect 1586 51 1799 85
rect 1833 131 1951 147
rect 2283 143 2317 277
rect 1833 97 1864 131
rect 1898 97 1951 131
rect 1833 81 1951 97
rect 2028 120 2116 136
rect 2028 86 2055 120
rect 2089 86 2116 120
rect 1486 17 1552 48
rect 2028 17 2116 86
rect 2208 127 2317 143
rect 2208 93 2231 127
rect 2265 93 2317 127
rect 2208 77 2317 93
rect 2351 304 2770 320
rect 2351 270 2584 304
rect 2618 270 2652 304
rect 2686 270 2720 304
rect 2754 270 2770 304
rect 2351 254 2770 270
rect 2817 260 2951 354
rect 2351 210 2385 254
rect 2817 220 2851 260
rect 2351 120 2385 176
rect 2351 70 2385 86
rect 2421 204 2473 220
rect 2421 170 2437 204
rect 2471 170 2473 204
rect 2421 120 2473 170
rect 2421 86 2437 120
rect 2471 86 2473 120
rect 2421 17 2473 86
rect 2507 210 2851 220
rect 2507 204 2817 210
rect 2507 170 2523 204
rect 2557 186 2817 204
rect 2557 170 2573 186
rect 2507 120 2573 170
rect 2507 86 2523 120
rect 2557 86 2573 120
rect 2507 70 2573 86
rect 2607 136 2781 152
rect 2607 102 2609 136
rect 2643 102 2731 136
rect 2765 102 2781 136
rect 2607 17 2781 102
rect 2817 120 2851 176
rect 2817 70 2851 86
rect 2887 210 2953 226
rect 2887 176 2903 210
rect 2937 176 2953 210
rect 2887 120 2953 176
rect 2887 86 2903 120
rect 2937 86 2953 120
rect 2887 17 2953 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 799 416 833 424
rect 799 390 807 416
rect 807 390 833 416
rect 1567 414 1601 424
rect 1567 390 1579 414
rect 1579 390 1601 414
rect 2143 414 2177 424
rect 2143 390 2167 414
rect 2167 390 2177 414
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< metal1 >>
rect 0 683 2976 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 0 617 2976 649
rect 787 424 845 430
rect 787 390 799 424
rect 833 421 845 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 833 393 1567 421
rect 833 390 845 393
rect 787 384 845 390
rect 1555 390 1567 393
rect 1601 421 1613 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1601 393 2143 421
rect 1601 390 1613 393
rect 1555 384 1613 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 2976 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
rect 0 -49 2976 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfrtp_4
flabel comment s 1507 630 1507 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 1119 36 1119 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel pwell s 0 0 2976 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2976 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 2143 390 2177 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 0 2976 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 0 617 2976 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2911 316 2945 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2976 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y R90
string GDS_END 1721550
string GDS_START 1699480
<< end >>
