magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
<< pwell >>
rect 1 49 2111 241
rect 0 0 2112 49
<< scnmos >>
rect 84 47 114 215
rect 170 47 200 215
rect 270 47 300 215
rect 356 47 386 215
rect 442 47 472 215
rect 528 47 558 215
rect 614 47 644 215
rect 700 47 730 215
rect 786 47 816 215
rect 872 47 902 215
rect 982 47 1012 215
rect 1068 47 1098 215
rect 1154 47 1184 215
rect 1240 47 1270 215
rect 1326 47 1356 215
rect 1412 47 1442 215
rect 1498 47 1528 215
rect 1598 47 1628 215
rect 1698 47 1728 215
rect 1798 47 1828 215
rect 1898 47 1928 215
rect 1994 47 2024 215
<< scpmoshvt >>
rect 84 367 114 619
rect 170 367 200 619
rect 256 367 286 619
rect 342 367 372 619
rect 428 367 458 619
rect 514 367 544 619
rect 606 367 636 619
rect 692 367 722 619
rect 778 367 808 619
rect 864 367 894 619
rect 950 367 980 619
rect 1036 367 1066 619
rect 1122 367 1152 619
rect 1208 367 1238 619
rect 1308 367 1338 619
rect 1408 367 1438 619
rect 1508 367 1538 619
rect 1608 367 1638 619
rect 1708 367 1738 619
rect 1808 367 1838 619
rect 1908 367 1938 619
rect 1994 367 2024 619
<< ndiff >>
rect 27 203 84 215
rect 27 169 39 203
rect 73 169 84 203
rect 27 101 84 169
rect 27 67 39 101
rect 73 67 84 101
rect 27 47 84 67
rect 114 114 170 215
rect 114 80 125 114
rect 159 80 170 114
rect 114 47 170 80
rect 200 170 270 215
rect 200 136 225 170
rect 259 136 270 170
rect 200 47 270 136
rect 300 186 356 215
rect 300 152 311 186
rect 345 152 356 186
rect 300 101 356 152
rect 300 67 311 101
rect 345 67 356 101
rect 300 47 356 67
rect 386 105 442 215
rect 386 71 397 105
rect 431 71 442 105
rect 386 47 442 71
rect 472 187 528 215
rect 472 153 483 187
rect 517 153 528 187
rect 472 101 528 153
rect 472 67 483 101
rect 517 67 528 101
rect 472 47 528 67
rect 558 203 614 215
rect 558 169 569 203
rect 603 169 614 203
rect 558 93 614 169
rect 558 59 569 93
rect 603 59 614 93
rect 558 47 614 59
rect 644 203 700 215
rect 644 169 655 203
rect 689 169 700 203
rect 644 101 700 169
rect 644 67 655 101
rect 689 67 700 101
rect 644 47 700 67
rect 730 114 786 215
rect 730 80 741 114
rect 775 80 786 114
rect 730 47 786 80
rect 816 203 872 215
rect 816 169 827 203
rect 861 169 872 203
rect 816 101 872 169
rect 816 67 827 101
rect 861 67 872 101
rect 816 47 872 67
rect 902 114 982 215
rect 902 80 913 114
rect 947 80 982 114
rect 902 47 982 80
rect 1012 203 1068 215
rect 1012 169 1023 203
rect 1057 169 1068 203
rect 1012 101 1068 169
rect 1012 67 1023 101
rect 1057 67 1068 101
rect 1012 47 1068 67
rect 1098 114 1154 215
rect 1098 80 1109 114
rect 1143 80 1154 114
rect 1098 47 1154 80
rect 1184 203 1240 215
rect 1184 169 1195 203
rect 1229 169 1240 203
rect 1184 101 1240 169
rect 1184 67 1195 101
rect 1229 67 1240 101
rect 1184 47 1240 67
rect 1270 186 1326 215
rect 1270 152 1281 186
rect 1315 152 1326 186
rect 1270 47 1326 152
rect 1356 118 1412 215
rect 1356 84 1367 118
rect 1401 84 1412 118
rect 1356 47 1412 84
rect 1442 186 1498 215
rect 1442 152 1453 186
rect 1487 152 1498 186
rect 1442 47 1498 152
rect 1528 122 1598 215
rect 1528 88 1553 122
rect 1587 88 1598 122
rect 1528 47 1598 88
rect 1628 178 1698 215
rect 1628 144 1653 178
rect 1687 144 1698 178
rect 1628 47 1698 144
rect 1728 122 1798 215
rect 1728 88 1753 122
rect 1787 88 1798 122
rect 1728 47 1798 88
rect 1828 186 1898 215
rect 1828 152 1853 186
rect 1887 152 1898 186
rect 1828 47 1898 152
rect 1928 118 1994 215
rect 1928 84 1939 118
rect 1973 84 1994 118
rect 1928 47 1994 84
rect 2024 114 2085 215
rect 2024 80 2039 114
rect 2073 80 2085 114
rect 2024 47 2085 80
<< pdiff >>
rect 27 599 84 619
rect 27 565 39 599
rect 73 565 84 599
rect 27 506 84 565
rect 27 472 39 506
rect 73 472 84 506
rect 27 413 84 472
rect 27 379 39 413
rect 73 379 84 413
rect 27 367 84 379
rect 114 599 170 619
rect 114 565 125 599
rect 159 565 170 599
rect 114 519 170 565
rect 114 485 125 519
rect 159 485 170 519
rect 114 439 170 485
rect 114 405 125 439
rect 159 405 170 439
rect 114 367 170 405
rect 200 531 256 619
rect 200 497 211 531
rect 245 497 256 531
rect 200 413 256 497
rect 200 379 211 413
rect 245 379 256 413
rect 200 367 256 379
rect 286 599 342 619
rect 286 565 297 599
rect 331 565 342 599
rect 286 527 342 565
rect 286 493 297 527
rect 331 493 342 527
rect 286 455 342 493
rect 286 421 297 455
rect 331 421 342 455
rect 286 367 342 421
rect 372 607 428 619
rect 372 573 383 607
rect 417 573 428 607
rect 372 523 428 573
rect 372 489 383 523
rect 417 489 428 523
rect 372 367 428 489
rect 458 599 514 619
rect 458 565 469 599
rect 503 565 514 599
rect 458 527 514 565
rect 458 493 469 527
rect 503 493 514 527
rect 458 455 514 493
rect 458 421 469 455
rect 503 421 514 455
rect 458 367 514 421
rect 544 607 606 619
rect 544 573 555 607
rect 589 573 606 607
rect 544 531 606 573
rect 544 497 555 531
rect 589 497 606 531
rect 544 455 606 497
rect 544 421 555 455
rect 589 421 606 455
rect 544 367 606 421
rect 636 599 692 619
rect 636 565 647 599
rect 681 565 692 599
rect 636 506 692 565
rect 636 472 647 506
rect 681 472 692 506
rect 636 413 692 472
rect 636 379 647 413
rect 681 379 692 413
rect 636 367 692 379
rect 722 607 778 619
rect 722 573 733 607
rect 767 573 778 607
rect 722 539 778 573
rect 722 505 733 539
rect 767 505 778 539
rect 722 471 778 505
rect 722 437 733 471
rect 767 437 778 471
rect 722 367 778 437
rect 808 599 864 619
rect 808 565 819 599
rect 853 565 864 599
rect 808 506 864 565
rect 808 472 819 506
rect 853 472 864 506
rect 808 413 864 472
rect 808 379 819 413
rect 853 379 864 413
rect 808 367 864 379
rect 894 607 950 619
rect 894 573 905 607
rect 939 573 950 607
rect 894 539 950 573
rect 894 505 905 539
rect 939 505 950 539
rect 894 471 950 505
rect 894 437 905 471
rect 939 437 950 471
rect 894 367 950 437
rect 980 599 1036 619
rect 980 565 991 599
rect 1025 565 1036 599
rect 980 506 1036 565
rect 980 472 991 506
rect 1025 472 1036 506
rect 980 413 1036 472
rect 980 379 991 413
rect 1025 379 1036 413
rect 980 367 1036 379
rect 1066 607 1122 619
rect 1066 573 1077 607
rect 1111 573 1122 607
rect 1066 539 1122 573
rect 1066 505 1077 539
rect 1111 505 1122 539
rect 1066 471 1122 505
rect 1066 437 1077 471
rect 1111 437 1122 471
rect 1066 367 1122 437
rect 1152 599 1208 619
rect 1152 565 1163 599
rect 1197 565 1208 599
rect 1152 506 1208 565
rect 1152 472 1163 506
rect 1197 472 1208 506
rect 1152 413 1208 472
rect 1152 379 1163 413
rect 1197 379 1208 413
rect 1152 367 1208 379
rect 1238 531 1308 619
rect 1238 497 1263 531
rect 1297 497 1308 531
rect 1238 413 1308 497
rect 1238 379 1263 413
rect 1297 379 1308 413
rect 1238 367 1308 379
rect 1338 599 1408 619
rect 1338 565 1363 599
rect 1397 565 1408 599
rect 1338 471 1408 565
rect 1338 437 1363 471
rect 1397 437 1408 471
rect 1338 367 1408 437
rect 1438 531 1508 619
rect 1438 497 1463 531
rect 1497 497 1508 531
rect 1438 413 1508 497
rect 1438 379 1463 413
rect 1497 379 1508 413
rect 1438 367 1508 379
rect 1538 599 1608 619
rect 1538 565 1563 599
rect 1597 565 1608 599
rect 1538 471 1608 565
rect 1538 437 1563 471
rect 1597 437 1608 471
rect 1538 367 1608 437
rect 1638 531 1708 619
rect 1638 497 1663 531
rect 1697 497 1708 531
rect 1638 413 1708 497
rect 1638 379 1663 413
rect 1697 379 1708 413
rect 1638 367 1708 379
rect 1738 599 1808 619
rect 1738 565 1763 599
rect 1797 565 1808 599
rect 1738 471 1808 565
rect 1738 437 1763 471
rect 1797 437 1808 471
rect 1738 367 1808 437
rect 1838 531 1908 619
rect 1838 497 1863 531
rect 1897 497 1908 531
rect 1838 413 1908 497
rect 1838 379 1863 413
rect 1897 379 1908 413
rect 1838 367 1908 379
rect 1938 599 1994 619
rect 1938 565 1949 599
rect 1983 565 1994 599
rect 1938 471 1994 565
rect 1938 437 1949 471
rect 1983 437 1994 471
rect 1938 367 1994 437
rect 2024 607 2081 619
rect 2024 573 2035 607
rect 2069 573 2081 607
rect 2024 539 2081 573
rect 2024 505 2035 539
rect 2069 505 2081 539
rect 2024 471 2081 505
rect 2024 437 2035 471
rect 2069 437 2081 471
rect 2024 367 2081 437
<< ndiffc >>
rect 39 169 73 203
rect 39 67 73 101
rect 125 80 159 114
rect 225 136 259 170
rect 311 152 345 186
rect 311 67 345 101
rect 397 71 431 105
rect 483 153 517 187
rect 483 67 517 101
rect 569 169 603 203
rect 569 59 603 93
rect 655 169 689 203
rect 655 67 689 101
rect 741 80 775 114
rect 827 169 861 203
rect 827 67 861 101
rect 913 80 947 114
rect 1023 169 1057 203
rect 1023 67 1057 101
rect 1109 80 1143 114
rect 1195 169 1229 203
rect 1195 67 1229 101
rect 1281 152 1315 186
rect 1367 84 1401 118
rect 1453 152 1487 186
rect 1553 88 1587 122
rect 1653 144 1687 178
rect 1753 88 1787 122
rect 1853 152 1887 186
rect 1939 84 1973 118
rect 2039 80 2073 114
<< pdiffc >>
rect 39 565 73 599
rect 39 472 73 506
rect 39 379 73 413
rect 125 565 159 599
rect 125 485 159 519
rect 125 405 159 439
rect 211 497 245 531
rect 211 379 245 413
rect 297 565 331 599
rect 297 493 331 527
rect 297 421 331 455
rect 383 573 417 607
rect 383 489 417 523
rect 469 565 503 599
rect 469 493 503 527
rect 469 421 503 455
rect 555 573 589 607
rect 555 497 589 531
rect 555 421 589 455
rect 647 565 681 599
rect 647 472 681 506
rect 647 379 681 413
rect 733 573 767 607
rect 733 505 767 539
rect 733 437 767 471
rect 819 565 853 599
rect 819 472 853 506
rect 819 379 853 413
rect 905 573 939 607
rect 905 505 939 539
rect 905 437 939 471
rect 991 565 1025 599
rect 991 472 1025 506
rect 991 379 1025 413
rect 1077 573 1111 607
rect 1077 505 1111 539
rect 1077 437 1111 471
rect 1163 565 1197 599
rect 1163 472 1197 506
rect 1163 379 1197 413
rect 1263 497 1297 531
rect 1263 379 1297 413
rect 1363 565 1397 599
rect 1363 437 1397 471
rect 1463 497 1497 531
rect 1463 379 1497 413
rect 1563 565 1597 599
rect 1563 437 1597 471
rect 1663 497 1697 531
rect 1663 379 1697 413
rect 1763 565 1797 599
rect 1763 437 1797 471
rect 1863 497 1897 531
rect 1863 379 1897 413
rect 1949 565 1983 599
rect 1949 437 1983 471
rect 2035 573 2069 607
rect 2035 505 2069 539
rect 2035 437 2069 471
<< poly >>
rect 84 619 114 645
rect 170 619 200 645
rect 256 619 286 645
rect 342 619 372 645
rect 428 619 458 645
rect 514 619 544 645
rect 606 619 636 645
rect 692 619 722 645
rect 778 619 808 645
rect 864 619 894 645
rect 950 619 980 645
rect 1036 619 1066 645
rect 1122 619 1152 645
rect 1208 619 1238 645
rect 1308 619 1338 645
rect 1408 619 1438 645
rect 1508 619 1538 645
rect 1608 619 1638 645
rect 1708 619 1738 645
rect 1808 619 1838 645
rect 1908 619 1938 645
rect 1994 619 2024 645
rect 84 303 114 367
rect 170 303 200 367
rect 256 303 286 367
rect 342 303 372 367
rect 428 303 458 367
rect 514 303 544 367
rect 606 319 636 367
rect 692 319 722 367
rect 778 319 808 367
rect 864 319 894 367
rect 950 319 980 367
rect 1036 319 1066 367
rect 1122 319 1152 367
rect 1208 319 1238 367
rect 1308 319 1338 367
rect 1408 319 1438 367
rect 1508 319 1538 367
rect 1608 319 1638 367
rect 1708 319 1738 367
rect 1808 319 1838 367
rect 1908 319 1938 367
rect 1994 319 2024 367
rect 606 303 2024 319
rect 84 287 558 303
rect 84 253 123 287
rect 157 253 191 287
rect 225 253 259 287
rect 293 253 327 287
rect 361 253 395 287
rect 429 253 463 287
rect 497 253 558 287
rect 606 269 622 303
rect 656 269 690 303
rect 724 269 758 303
rect 792 269 826 303
rect 860 269 894 303
rect 928 269 962 303
rect 996 269 1030 303
rect 1064 269 1098 303
rect 1132 269 1166 303
rect 1200 269 1234 303
rect 1268 269 1302 303
rect 1336 269 1370 303
rect 1404 269 1438 303
rect 1472 269 1506 303
rect 1540 269 1574 303
rect 1608 269 1642 303
rect 1676 269 1710 303
rect 1744 269 1778 303
rect 1812 269 1846 303
rect 1880 269 1914 303
rect 1948 269 2024 303
rect 606 253 2024 269
rect 84 237 558 253
rect 84 215 114 237
rect 170 215 200 237
rect 270 215 300 237
rect 356 215 386 237
rect 442 215 472 237
rect 528 215 558 237
rect 614 215 644 253
rect 700 215 730 253
rect 786 215 816 253
rect 872 215 902 253
rect 982 215 1012 253
rect 1068 215 1098 253
rect 1154 215 1184 253
rect 1240 215 1270 253
rect 1326 215 1356 253
rect 1412 215 1442 253
rect 1498 215 1528 253
rect 1598 215 1628 253
rect 1698 215 1728 253
rect 1798 215 1828 253
rect 1898 215 1928 253
rect 1994 215 2024 253
rect 84 21 114 47
rect 170 21 200 47
rect 270 21 300 47
rect 356 21 386 47
rect 442 21 472 47
rect 528 21 558 47
rect 614 21 644 47
rect 700 21 730 47
rect 786 21 816 47
rect 872 21 902 47
rect 982 21 1012 47
rect 1068 21 1098 47
rect 1154 21 1184 47
rect 1240 21 1270 47
rect 1326 21 1356 47
rect 1412 21 1442 47
rect 1498 21 1528 47
rect 1598 21 1628 47
rect 1698 21 1728 47
rect 1798 21 1828 47
rect 1898 21 1928 47
rect 1994 21 2024 47
<< polycont >>
rect 123 253 157 287
rect 191 253 225 287
rect 259 253 293 287
rect 327 253 361 287
rect 395 253 429 287
rect 463 253 497 287
rect 622 269 656 303
rect 690 269 724 303
rect 758 269 792 303
rect 826 269 860 303
rect 894 269 928 303
rect 962 269 996 303
rect 1030 269 1064 303
rect 1098 269 1132 303
rect 1166 269 1200 303
rect 1234 269 1268 303
rect 1302 269 1336 303
rect 1370 269 1404 303
rect 1438 269 1472 303
rect 1506 269 1540 303
rect 1574 269 1608 303
rect 1642 269 1676 303
rect 1710 269 1744 303
rect 1778 269 1812 303
rect 1846 269 1880 303
rect 1914 269 1948 303
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 23 599 73 615
rect 23 565 39 599
rect 23 506 73 565
rect 23 472 39 506
rect 23 413 73 472
rect 23 379 39 413
rect 109 599 347 615
rect 109 565 125 599
rect 159 581 297 599
rect 159 565 175 581
rect 109 519 175 565
rect 281 565 297 581
rect 331 565 347 599
rect 109 485 125 519
rect 159 485 175 519
rect 109 439 175 485
rect 109 405 125 439
rect 159 405 175 439
rect 211 531 245 547
rect 211 413 245 497
rect 23 371 73 379
rect 281 527 347 565
rect 281 493 297 527
rect 331 493 347 527
rect 281 455 347 493
rect 383 607 417 649
rect 383 523 417 573
rect 383 473 417 489
rect 453 599 519 615
rect 453 565 469 599
rect 503 565 519 599
rect 453 527 519 565
rect 453 493 469 527
rect 503 493 519 527
rect 281 421 297 455
rect 331 439 347 455
rect 453 455 519 493
rect 453 439 469 455
rect 331 421 469 439
rect 503 421 519 455
rect 281 405 519 421
rect 555 607 589 649
rect 555 531 589 573
rect 555 455 589 497
rect 555 405 589 421
rect 631 599 697 615
rect 631 565 647 599
rect 681 565 697 599
rect 631 506 697 565
rect 631 472 647 506
rect 681 472 697 506
rect 631 413 697 472
rect 733 607 767 649
rect 733 539 767 573
rect 733 471 767 505
rect 733 421 767 437
rect 803 599 869 615
rect 803 565 819 599
rect 853 565 869 599
rect 803 506 869 565
rect 803 472 819 506
rect 853 472 869 506
rect 211 371 245 379
rect 631 379 647 413
rect 681 387 697 413
rect 803 413 869 472
rect 905 607 939 649
rect 905 539 939 573
rect 905 471 939 505
rect 905 421 939 437
rect 975 599 1041 615
rect 975 565 991 599
rect 1025 565 1041 599
rect 975 506 1041 565
rect 975 472 991 506
rect 1025 472 1041 506
rect 803 387 819 413
rect 681 379 819 387
rect 853 387 869 413
rect 975 413 1041 472
rect 1077 607 1111 649
rect 1077 539 1111 573
rect 1077 471 1111 505
rect 1077 421 1111 437
rect 1147 599 1983 615
rect 1147 565 1163 599
rect 1197 581 1363 599
rect 1197 565 1213 581
rect 1147 506 1213 565
rect 1347 565 1363 581
rect 1397 581 1563 599
rect 1397 565 1413 581
rect 1147 472 1163 506
rect 1197 472 1213 506
rect 975 387 991 413
rect 853 379 991 387
rect 1025 387 1041 413
rect 1147 413 1213 472
rect 1147 387 1163 413
rect 1025 379 1163 387
rect 1197 379 1213 413
rect 23 337 597 371
rect 631 353 1213 379
rect 1247 531 1313 547
rect 1247 497 1263 531
rect 1297 497 1313 531
rect 1247 413 1313 497
rect 1347 471 1413 565
rect 1547 565 1563 581
rect 1597 581 1763 599
rect 1597 565 1613 581
rect 1347 437 1363 471
rect 1397 437 1413 471
rect 1347 421 1413 437
rect 1447 531 1513 547
rect 1447 497 1463 531
rect 1497 497 1513 531
rect 1247 379 1263 413
rect 1297 387 1313 413
rect 1447 413 1513 497
rect 1547 471 1613 565
rect 1747 565 1763 581
rect 1797 581 1949 599
rect 1797 565 1813 581
rect 1547 437 1563 471
rect 1597 437 1613 471
rect 1547 421 1613 437
rect 1647 531 1713 547
rect 1647 497 1663 531
rect 1697 497 1713 531
rect 1447 387 1463 413
rect 1297 379 1463 387
rect 1497 387 1513 413
rect 1647 413 1713 497
rect 1747 471 1813 565
rect 1747 437 1763 471
rect 1797 437 1813 471
rect 1747 421 1813 437
rect 1847 531 1913 547
rect 1847 497 1863 531
rect 1897 497 1913 531
rect 1647 387 1663 413
rect 1497 379 1663 387
rect 1697 387 1713 413
rect 1847 413 1913 497
rect 1949 471 1983 565
rect 1949 421 1983 437
rect 2019 607 2085 649
rect 2019 573 2035 607
rect 2069 573 2085 607
rect 2019 539 2085 573
rect 2019 505 2035 539
rect 2069 505 2085 539
rect 2019 471 2085 505
rect 2019 437 2035 471
rect 2069 437 2085 471
rect 2019 421 2085 437
rect 1847 387 1863 413
rect 1697 379 1863 387
rect 1897 387 1913 413
rect 1897 379 2087 387
rect 1247 353 2087 379
rect 39 219 73 337
rect 563 319 597 337
rect 563 303 1964 319
rect 107 287 513 303
rect 107 253 123 287
rect 157 253 191 287
rect 225 253 259 287
rect 293 253 327 287
rect 361 253 395 287
rect 429 253 463 287
rect 497 253 513 287
rect 563 269 622 303
rect 656 269 690 303
rect 724 269 758 303
rect 792 269 826 303
rect 860 269 894 303
rect 928 269 962 303
rect 996 269 1030 303
rect 1064 269 1098 303
rect 1132 269 1166 303
rect 1200 269 1234 303
rect 1268 269 1302 303
rect 1336 269 1370 303
rect 1404 269 1438 303
rect 1472 269 1506 303
rect 1540 269 1574 303
rect 1608 269 1642 303
rect 1676 269 1710 303
rect 1744 269 1778 303
rect 1812 269 1846 303
rect 1880 269 1914 303
rect 1948 269 1964 303
rect 563 253 1964 269
rect 107 237 513 253
rect 107 236 451 237
rect 1999 219 2087 353
rect 23 203 73 219
rect 569 203 603 219
rect 23 169 39 203
rect 467 202 533 203
rect 73 170 275 202
rect 73 169 225 170
rect 23 168 225 169
rect 23 101 73 168
rect 209 136 225 168
rect 259 136 275 170
rect 23 67 39 101
rect 23 51 73 67
rect 109 114 175 134
rect 209 119 275 136
rect 311 187 533 202
rect 311 186 483 187
rect 345 155 483 186
rect 109 80 125 114
rect 159 85 175 114
rect 311 101 345 152
rect 467 153 483 155
rect 517 153 533 187
rect 159 80 311 85
rect 109 67 311 80
rect 109 51 345 67
rect 381 105 431 121
rect 381 71 397 105
rect 381 17 431 71
rect 467 101 533 153
rect 467 67 483 101
rect 517 67 533 101
rect 467 51 533 67
rect 569 93 603 169
rect 569 17 603 59
rect 639 203 1245 219
rect 639 169 655 203
rect 689 185 827 203
rect 639 101 689 169
rect 811 169 827 185
rect 861 185 1023 203
rect 639 67 655 101
rect 639 51 689 67
rect 725 114 775 151
rect 725 80 741 114
rect 725 17 775 80
rect 811 101 861 169
rect 1007 169 1023 185
rect 1057 185 1195 203
rect 811 67 827 101
rect 811 51 861 67
rect 897 114 963 151
rect 897 80 913 114
rect 947 80 963 114
rect 897 17 963 80
rect 1007 101 1057 169
rect 1179 169 1195 185
rect 1229 169 1245 203
rect 1007 67 1023 101
rect 1007 51 1057 67
rect 1093 114 1143 151
rect 1093 80 1109 114
rect 1093 17 1143 80
rect 1179 101 1245 169
rect 1281 186 2087 219
rect 1315 185 1453 186
rect 1281 119 1315 152
rect 1487 185 1853 186
rect 1487 152 1503 185
rect 1179 67 1195 101
rect 1229 85 1245 101
rect 1351 118 1417 151
rect 1453 119 1503 152
rect 1637 178 1703 185
rect 1537 122 1603 151
rect 1351 85 1367 118
rect 1229 84 1367 85
rect 1401 85 1417 118
rect 1537 88 1553 122
rect 1587 88 1603 122
rect 1637 144 1653 178
rect 1687 144 1703 178
rect 1837 152 1853 185
rect 1887 185 2087 186
rect 1887 152 1903 185
rect 1637 119 1703 144
rect 1737 122 1803 151
rect 1537 85 1603 88
rect 1737 88 1753 122
rect 1787 88 1803 122
rect 1837 119 1903 152
rect 1737 85 1803 88
rect 1939 118 1989 151
rect 1401 84 1939 85
rect 1973 84 1989 118
rect 1229 67 1989 84
rect 1179 51 1989 67
rect 2023 114 2089 151
rect 2023 80 2039 114
rect 2073 80 2089 114
rect 2023 17 2089 80
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 buflp_8
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6962294
string GDS_START 6946532
<< end >>
