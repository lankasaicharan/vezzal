magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1304 -1309 2065 1975
<< nwell >>
rect -44 331 805 704
<< pwell >>
rect 1 49 753 203
rect 0 0 768 49
<< scnmos >>
rect 80 93 110 177
rect 152 93 182 177
rect 238 93 268 177
rect 310 93 340 177
rect 408 93 438 177
rect 480 93 510 177
rect 572 93 602 177
rect 644 93 674 177
<< scpmoshvt >>
rect 124 489 154 573
rect 202 489 232 573
rect 310 489 340 573
rect 382 489 412 573
rect 572 367 602 619
rect 644 367 674 619
<< ndiff >>
rect 27 161 80 177
rect 27 127 35 161
rect 69 127 80 161
rect 27 93 80 127
rect 110 93 152 177
rect 182 159 238 177
rect 182 125 193 159
rect 227 125 238 159
rect 182 93 238 125
rect 268 93 310 177
rect 340 160 408 177
rect 340 126 363 160
rect 397 126 408 160
rect 340 93 408 126
rect 438 93 480 177
rect 510 161 572 177
rect 510 127 521 161
rect 555 127 572 161
rect 510 93 572 127
rect 602 93 644 177
rect 674 161 727 177
rect 674 127 685 161
rect 719 127 727 161
rect 674 93 727 127
<< pdiff >>
rect 519 607 572 619
rect 519 573 527 607
rect 561 573 572 607
rect 71 548 124 573
rect 71 514 79 548
rect 113 514 124 548
rect 71 489 124 514
rect 154 489 202 573
rect 232 548 310 573
rect 232 514 254 548
rect 288 514 310 548
rect 232 489 310 514
rect 340 489 382 573
rect 412 556 465 573
rect 412 522 423 556
rect 457 522 465 556
rect 412 489 465 522
rect 519 493 572 573
rect 519 459 527 493
rect 561 459 572 493
rect 519 367 572 459
rect 602 367 644 619
rect 674 599 727 619
rect 674 565 685 599
rect 719 565 727 599
rect 674 507 727 565
rect 674 473 685 507
rect 719 473 727 507
rect 674 413 727 473
rect 674 379 685 413
rect 719 379 727 413
rect 674 367 727 379
<< ndiffc >>
rect 35 127 69 161
rect 193 125 227 159
rect 363 126 397 160
rect 521 127 555 161
rect 685 127 719 161
<< pdiffc >>
rect 527 573 561 607
rect 79 514 113 548
rect 254 514 288 548
rect 423 522 457 556
rect 527 459 561 493
rect 685 565 719 599
rect 685 473 719 507
rect 685 379 719 413
<< poly >>
rect 572 619 602 645
rect 644 619 674 645
rect 124 573 154 599
rect 202 573 232 599
rect 310 573 340 599
rect 382 573 412 599
rect 124 398 154 489
rect 202 398 232 489
rect 98 382 232 398
rect 310 397 340 489
rect 98 294 114 382
rect 80 280 114 294
rect 216 280 232 382
rect 80 264 232 280
rect 274 381 340 397
rect 274 347 290 381
rect 324 347 340 381
rect 274 313 340 347
rect 274 279 290 313
rect 324 279 340 313
rect 80 177 110 264
rect 152 177 182 264
rect 274 222 340 279
rect 382 329 412 489
rect 572 338 602 367
rect 644 338 674 367
rect 382 313 516 329
rect 382 279 398 313
rect 432 279 466 313
rect 500 279 516 313
rect 382 263 516 279
rect 572 319 674 338
rect 572 285 595 319
rect 629 285 674 319
rect 238 192 340 222
rect 238 177 268 192
rect 310 177 340 192
rect 408 177 438 263
rect 480 177 510 263
rect 572 251 674 285
rect 572 217 595 251
rect 629 217 674 251
rect 572 201 674 217
rect 572 177 602 201
rect 644 177 674 201
rect 80 67 110 93
rect 152 67 182 93
rect 238 67 268 93
rect 310 67 340 93
rect 408 67 438 93
rect 480 67 510 93
rect 572 67 602 93
rect 644 67 674 93
<< polycont >>
rect 114 280 216 382
rect 290 347 324 381
rect 290 279 324 313
rect 398 279 432 313
rect 466 279 500 313
rect 595 285 629 319
rect 595 217 629 251
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 69 548 118 564
rect 69 514 79 548
rect 113 514 118 548
rect 69 466 118 514
rect 238 548 304 649
rect 505 607 582 649
rect 238 514 254 548
rect 288 514 304 548
rect 238 500 304 514
rect 419 556 461 576
rect 419 522 423 556
rect 457 522 461 556
rect 25 432 340 466
rect 25 177 74 432
rect 108 382 232 398
rect 108 280 114 382
rect 216 280 232 382
rect 108 232 232 280
rect 274 381 340 432
rect 419 425 461 522
rect 505 573 527 607
rect 561 573 582 607
rect 505 493 582 573
rect 505 459 527 493
rect 561 459 582 493
rect 679 599 751 615
rect 679 565 685 599
rect 719 565 751 599
rect 679 507 751 565
rect 679 473 685 507
rect 719 473 751 507
rect 419 391 645 425
rect 274 347 290 381
rect 324 347 340 381
rect 274 313 340 347
rect 274 279 290 313
rect 324 279 340 313
rect 382 313 516 350
rect 382 279 398 313
rect 432 279 466 313
rect 500 279 516 313
rect 579 319 645 391
rect 579 285 595 319
rect 629 285 645 319
rect 274 263 340 279
rect 579 251 645 285
rect 579 245 595 251
rect 374 217 595 245
rect 629 217 645 251
rect 374 211 645 217
rect 679 413 751 473
rect 679 379 685 413
rect 719 379 751 413
rect 374 177 413 211
rect 24 161 73 177
rect 24 127 35 161
rect 69 127 73 161
rect 24 86 73 127
rect 177 159 303 177
rect 177 128 193 159
rect 227 128 303 159
rect 177 94 187 128
rect 227 125 259 128
rect 221 94 259 125
rect 293 94 303 128
rect 177 86 303 94
rect 347 160 413 177
rect 347 126 363 160
rect 397 126 413 160
rect 347 86 413 126
rect 505 161 631 177
rect 505 128 521 161
rect 555 128 631 161
rect 505 94 515 128
rect 555 127 587 128
rect 549 94 587 127
rect 621 94 631 128
rect 505 86 631 94
rect 679 161 751 379
rect 679 127 685 161
rect 719 127 751 161
rect 679 93 751 127
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 187 125 193 128
rect 193 125 221 128
rect 187 94 221 125
rect 259 94 293 128
rect 515 127 521 128
rect 521 127 549 128
rect 515 94 549 127
rect 587 94 621 128
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 14 128 754 134
rect 14 94 187 128
rect 221 94 259 128
rect 293 94 515 128
rect 549 94 587 128
rect 621 94 754 128
rect 14 88 754 94
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel locali s 703 168 737 202 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 200 0 0 0 SLEEP_B
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 200 0 0 0 SLEEP_B
port 3 nsew signal input
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 iso1n_lp
flabel metal1 s 14 88 754 134 0 FreeSans 340 0 0 0 KAGND
port 2 nsew ground input
flabel metal1 s 0 617 768 666 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2855482
string GDS_START 2848718
<< end >>
