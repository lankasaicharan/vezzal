magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 1 49 1151 248
rect 0 0 1152 49
<< scnmos >>
rect 84 74 114 222
rect 179 74 209 222
rect 265 74 295 222
rect 351 74 381 222
rect 437 74 467 222
rect 537 74 567 222
rect 623 74 653 222
rect 737 74 767 222
rect 823 74 853 222
rect 937 74 967 222
rect 1024 74 1054 222
<< scpmoshvt >>
rect 87 368 117 592
rect 177 368 207 592
rect 267 368 297 592
rect 357 368 387 592
rect 457 368 487 592
rect 557 368 587 592
rect 647 368 677 592
rect 747 368 777 592
rect 837 368 867 592
rect 934 368 964 592
rect 1027 368 1057 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 152 179 222
rect 114 118 125 152
rect 159 118 179 152
rect 114 74 179 118
rect 209 210 265 222
rect 209 176 220 210
rect 254 176 265 210
rect 209 120 265 176
rect 209 86 220 120
rect 254 86 265 120
rect 209 74 265 86
rect 295 152 351 222
rect 295 118 306 152
rect 340 118 351 152
rect 295 74 351 118
rect 381 210 437 222
rect 381 176 392 210
rect 426 176 437 210
rect 381 120 437 176
rect 381 86 392 120
rect 426 86 437 120
rect 381 74 437 86
rect 467 142 537 222
rect 467 108 478 142
rect 512 108 537 142
rect 467 74 537 108
rect 567 210 623 222
rect 567 176 578 210
rect 612 176 623 210
rect 567 120 623 176
rect 567 86 578 120
rect 612 86 623 120
rect 567 74 623 86
rect 653 142 737 222
rect 653 108 678 142
rect 712 108 737 142
rect 653 74 737 108
rect 767 210 823 222
rect 767 176 778 210
rect 812 176 823 210
rect 767 120 823 176
rect 767 86 778 120
rect 812 86 823 120
rect 767 74 823 86
rect 853 142 937 222
rect 853 108 878 142
rect 912 108 937 142
rect 853 74 937 108
rect 967 210 1024 222
rect 967 176 978 210
rect 1012 176 1024 210
rect 967 120 1024 176
rect 967 86 978 120
rect 1012 86 1024 120
rect 967 74 1024 86
rect 1054 210 1125 222
rect 1054 176 1079 210
rect 1113 176 1125 210
rect 1054 120 1125 176
rect 1054 86 1079 120
rect 1113 86 1125 120
rect 1054 74 1125 86
<< pdiff >>
rect 28 580 87 592
rect 28 546 40 580
rect 74 546 87 580
rect 28 510 87 546
rect 28 476 40 510
rect 74 476 87 510
rect 28 440 87 476
rect 28 406 40 440
rect 74 406 87 440
rect 28 368 87 406
rect 117 580 177 592
rect 117 546 130 580
rect 164 546 177 580
rect 117 508 177 546
rect 117 474 130 508
rect 164 474 177 508
rect 117 368 177 474
rect 207 580 267 592
rect 207 546 220 580
rect 254 546 267 580
rect 207 510 267 546
rect 207 476 220 510
rect 254 476 267 510
rect 207 440 267 476
rect 207 406 220 440
rect 254 406 267 440
rect 207 368 267 406
rect 297 580 357 592
rect 297 546 310 580
rect 344 546 357 580
rect 297 508 357 546
rect 297 474 310 508
rect 344 474 357 508
rect 297 368 357 474
rect 387 580 457 592
rect 387 546 410 580
rect 444 546 457 580
rect 387 497 457 546
rect 387 463 410 497
rect 444 463 457 497
rect 387 414 457 463
rect 387 380 410 414
rect 444 380 457 414
rect 387 368 457 380
rect 487 580 557 592
rect 487 546 500 580
rect 534 546 557 580
rect 487 478 557 546
rect 487 444 500 478
rect 534 444 557 478
rect 487 368 557 444
rect 587 580 647 592
rect 587 546 600 580
rect 634 546 647 580
rect 587 497 647 546
rect 587 463 600 497
rect 634 463 647 497
rect 587 414 647 463
rect 587 380 600 414
rect 634 380 647 414
rect 587 368 647 380
rect 677 580 747 592
rect 677 546 690 580
rect 724 546 747 580
rect 677 478 747 546
rect 677 444 690 478
rect 724 444 747 478
rect 677 368 747 444
rect 777 580 837 592
rect 777 546 790 580
rect 824 546 837 580
rect 777 497 837 546
rect 777 463 790 497
rect 824 463 837 497
rect 777 414 837 463
rect 777 380 790 414
rect 824 380 837 414
rect 777 368 837 380
rect 867 580 934 592
rect 867 546 880 580
rect 914 546 934 580
rect 867 478 934 546
rect 867 444 880 478
rect 914 444 934 478
rect 867 368 934 444
rect 964 580 1027 592
rect 964 546 980 580
rect 1014 546 1027 580
rect 964 497 1027 546
rect 964 463 980 497
rect 1014 463 1027 497
rect 964 414 1027 463
rect 964 380 980 414
rect 1014 380 1027 414
rect 964 368 1027 380
rect 1057 580 1116 592
rect 1057 546 1070 580
rect 1104 546 1116 580
rect 1057 497 1116 546
rect 1057 463 1070 497
rect 1104 463 1116 497
rect 1057 414 1116 463
rect 1057 380 1070 414
rect 1104 380 1116 414
rect 1057 368 1116 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 118 159 152
rect 220 176 254 210
rect 220 86 254 120
rect 306 118 340 152
rect 392 176 426 210
rect 392 86 426 120
rect 478 108 512 142
rect 578 176 612 210
rect 578 86 612 120
rect 678 108 712 142
rect 778 176 812 210
rect 778 86 812 120
rect 878 108 912 142
rect 978 176 1012 210
rect 978 86 1012 120
rect 1079 176 1113 210
rect 1079 86 1113 120
<< pdiffc >>
rect 40 546 74 580
rect 40 476 74 510
rect 40 406 74 440
rect 130 546 164 580
rect 130 474 164 508
rect 220 546 254 580
rect 220 476 254 510
rect 220 406 254 440
rect 310 546 344 580
rect 310 474 344 508
rect 410 546 444 580
rect 410 463 444 497
rect 410 380 444 414
rect 500 546 534 580
rect 500 444 534 478
rect 600 546 634 580
rect 600 463 634 497
rect 600 380 634 414
rect 690 546 724 580
rect 690 444 724 478
rect 790 546 824 580
rect 790 463 824 497
rect 790 380 824 414
rect 880 546 914 580
rect 880 444 914 478
rect 980 546 1014 580
rect 980 463 1014 497
rect 980 380 1014 414
rect 1070 546 1104 580
rect 1070 463 1104 497
rect 1070 380 1104 414
<< poly >>
rect 87 592 117 618
rect 177 592 207 618
rect 267 592 297 618
rect 357 592 387 618
rect 457 592 487 618
rect 557 592 587 618
rect 647 592 677 618
rect 747 592 777 618
rect 837 592 867 618
rect 934 592 964 618
rect 1027 592 1057 618
rect 87 353 117 368
rect 177 353 207 368
rect 267 353 297 368
rect 357 353 387 368
rect 457 353 487 368
rect 557 353 587 368
rect 647 353 677 368
rect 747 353 777 368
rect 837 353 867 368
rect 934 353 964 368
rect 1027 353 1057 368
rect 84 336 120 353
rect 174 336 210 353
rect 264 336 300 353
rect 84 320 300 336
rect 354 326 390 353
rect 454 326 490 353
rect 554 326 590 353
rect 644 326 680 353
rect 744 326 780 353
rect 834 326 870 353
rect 931 326 967 353
rect 1024 326 1060 353
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 300 320
rect 84 270 300 286
rect 351 310 1060 326
rect 351 276 367 310
rect 401 276 435 310
rect 469 276 503 310
rect 537 276 571 310
rect 605 276 639 310
rect 673 276 707 310
rect 741 276 775 310
rect 809 276 843 310
rect 877 276 911 310
rect 945 276 1060 310
rect 84 222 114 270
rect 179 222 209 270
rect 265 222 295 270
rect 351 260 1060 276
rect 351 222 381 260
rect 437 222 467 260
rect 537 222 567 260
rect 623 222 653 260
rect 737 222 767 260
rect 823 222 853 260
rect 937 222 967 260
rect 1024 222 1054 260
rect 84 48 114 74
rect 179 48 209 74
rect 265 48 295 74
rect 351 48 381 74
rect 437 48 467 74
rect 537 48 567 74
rect 623 48 653 74
rect 737 48 767 74
rect 823 48 853 74
rect 937 48 967 74
rect 1024 48 1054 74
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 236 286 270 320
rect 367 276 401 310
rect 435 276 469 310
rect 503 276 537 310
rect 571 276 605 310
rect 639 276 673 310
rect 707 276 741 310
rect 775 276 809 310
rect 843 276 877 310
rect 911 276 945 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 24 580 90 596
rect 24 546 40 580
rect 74 546 90 580
rect 24 510 90 546
rect 24 476 40 510
rect 74 476 90 510
rect 24 440 90 476
rect 130 580 164 649
rect 130 508 164 546
rect 130 458 164 474
rect 204 580 270 596
rect 204 546 220 580
rect 254 546 270 580
rect 204 510 270 546
rect 204 476 220 510
rect 254 476 270 510
rect 24 406 40 440
rect 74 424 90 440
rect 204 440 270 476
rect 310 580 360 649
rect 344 546 360 580
rect 310 508 360 546
rect 344 474 360 508
rect 310 458 360 474
rect 394 580 460 596
rect 394 546 410 580
rect 444 546 460 580
rect 394 497 460 546
rect 394 463 410 497
rect 444 463 460 497
rect 204 424 220 440
rect 74 406 220 424
rect 254 424 270 440
rect 254 406 354 424
rect 24 390 354 406
rect 25 320 286 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 286 320
rect 25 270 286 286
rect 320 326 354 390
rect 394 414 460 463
rect 500 580 550 649
rect 534 546 550 580
rect 500 478 550 546
rect 534 444 550 478
rect 500 428 550 444
rect 584 580 650 596
rect 584 546 600 580
rect 634 546 650 580
rect 584 497 650 546
rect 584 463 600 497
rect 634 463 650 497
rect 394 380 410 414
rect 444 394 460 414
rect 584 414 650 463
rect 690 580 740 649
rect 724 546 740 580
rect 690 478 740 546
rect 724 444 740 478
rect 690 428 740 444
rect 774 580 840 596
rect 774 546 790 580
rect 824 546 840 580
rect 774 497 840 546
rect 774 463 790 497
rect 824 463 840 497
rect 584 394 600 414
rect 444 380 600 394
rect 634 394 650 414
rect 774 414 840 463
rect 880 580 930 649
rect 914 546 930 580
rect 880 478 930 546
rect 914 444 930 478
rect 880 428 930 444
rect 964 580 1031 596
rect 964 546 980 580
rect 1014 546 1031 580
rect 964 497 1031 546
rect 964 463 980 497
rect 1014 463 1031 497
rect 774 394 790 414
rect 634 380 790 394
rect 824 394 840 414
rect 964 414 1031 463
rect 964 394 980 414
rect 824 380 980 394
rect 1014 380 1031 414
rect 394 360 1031 380
rect 1070 580 1120 649
rect 1104 546 1120 580
rect 1070 497 1120 546
rect 1104 463 1120 497
rect 1070 414 1120 463
rect 1104 380 1120 414
rect 1070 364 1120 380
rect 320 310 961 326
rect 320 276 367 310
rect 401 276 435 310
rect 469 276 503 310
rect 537 276 571 310
rect 605 276 639 310
rect 673 276 707 310
rect 741 276 775 310
rect 809 276 843 310
rect 877 276 911 310
rect 945 276 961 310
rect 320 260 961 276
rect 320 236 354 260
rect 23 210 354 236
rect 995 226 1029 360
rect 23 176 39 210
rect 73 202 220 210
rect 23 120 73 176
rect 254 202 354 210
rect 392 210 1029 226
rect 23 86 39 120
rect 23 70 73 86
rect 109 152 175 168
rect 109 118 125 152
rect 159 118 175 152
rect 109 17 175 118
rect 220 120 254 176
rect 426 192 578 210
rect 220 70 254 86
rect 290 152 356 168
rect 290 118 306 152
rect 340 118 356 152
rect 290 17 356 118
rect 392 120 426 176
rect 562 176 578 192
rect 612 192 778 210
rect 612 176 628 192
rect 392 70 426 86
rect 462 142 528 158
rect 462 108 478 142
rect 512 108 528 142
rect 462 17 528 108
rect 562 120 628 176
rect 762 176 778 192
rect 812 192 978 210
rect 812 176 828 192
rect 562 86 578 120
rect 612 86 628 120
rect 562 70 628 86
rect 662 142 728 158
rect 662 108 678 142
rect 712 108 728 142
rect 662 17 728 108
rect 762 120 828 176
rect 962 176 978 192
rect 1012 176 1029 210
rect 762 86 778 120
rect 812 86 828 120
rect 762 70 828 86
rect 862 142 928 158
rect 862 108 878 142
rect 912 108 928 142
rect 862 17 928 108
rect 962 120 1029 176
rect 962 86 978 120
rect 1012 86 1029 120
rect 962 70 1029 86
rect 1063 210 1129 226
rect 1063 176 1079 210
rect 1113 176 1129 210
rect 1063 120 1129 176
rect 1063 86 1079 120
rect 1113 86 1129 120
rect 1063 17 1129 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buf_8
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 464 1025 498 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 538 1025 572 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 2994842
string GDS_START 2985050
<< end >>
