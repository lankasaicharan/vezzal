magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2065 1975
<< nwell >>
rect -38 331 805 704
<< pwell >>
rect 1 49 753 203
rect 0 0 768 49
<< scnmos >>
rect 82 93 112 177
rect 154 93 184 177
rect 310 93 340 177
rect 382 93 412 177
rect 572 93 602 177
rect 644 93 674 177
<< scpmoshvt >>
rect 82 417 132 617
rect 292 417 342 617
rect 402 417 452 617
rect 624 417 674 617
<< ndiff >>
rect 27 161 82 177
rect 27 127 37 161
rect 71 127 82 161
rect 27 93 82 127
rect 112 93 154 177
rect 184 152 310 177
rect 184 118 195 152
rect 229 118 265 152
rect 299 118 310 152
rect 184 93 310 118
rect 340 93 382 177
rect 412 161 465 177
rect 412 127 423 161
rect 457 127 465 161
rect 412 93 465 127
rect 519 161 572 177
rect 519 127 527 161
rect 561 127 572 161
rect 519 93 572 127
rect 602 93 644 177
rect 674 161 727 177
rect 674 127 685 161
rect 719 127 727 161
rect 674 93 727 127
<< pdiff >>
rect 27 599 82 617
rect 27 565 37 599
rect 71 565 82 599
rect 27 531 82 565
rect 27 497 37 531
rect 71 497 82 531
rect 27 463 82 497
rect 27 429 37 463
rect 71 429 82 463
rect 27 417 82 429
rect 132 609 292 617
rect 132 575 143 609
rect 177 575 247 609
rect 281 575 292 609
rect 132 496 292 575
rect 132 462 143 496
rect 177 462 247 496
rect 281 462 292 496
rect 132 417 292 462
rect 342 599 402 617
rect 342 565 357 599
rect 391 565 402 599
rect 342 531 402 565
rect 342 497 357 531
rect 391 497 402 531
rect 342 463 402 497
rect 342 429 357 463
rect 391 429 402 463
rect 342 417 402 429
rect 452 609 624 617
rect 452 575 463 609
rect 497 575 579 609
rect 613 575 624 609
rect 452 496 624 575
rect 452 462 463 496
rect 497 462 579 496
rect 613 462 624 496
rect 452 417 624 462
rect 674 599 727 617
rect 674 565 685 599
rect 719 565 727 599
rect 674 531 727 565
rect 674 497 685 531
rect 719 497 727 531
rect 674 463 727 497
rect 674 429 685 463
rect 719 429 727 463
rect 674 417 727 429
<< ndiffc >>
rect 37 127 71 161
rect 195 118 229 152
rect 265 118 299 152
rect 423 127 457 161
rect 527 127 561 161
rect 685 127 719 161
<< pdiffc >>
rect 37 565 71 599
rect 37 497 71 531
rect 37 429 71 463
rect 143 575 177 609
rect 247 575 281 609
rect 143 462 177 496
rect 247 462 281 496
rect 357 565 391 599
rect 357 497 391 531
rect 357 429 391 463
rect 463 575 497 609
rect 579 575 613 609
rect 463 462 497 496
rect 579 462 613 496
rect 685 565 719 599
rect 685 497 719 531
rect 685 429 719 463
<< poly >>
rect 82 617 132 645
rect 292 617 342 645
rect 402 617 452 645
rect 624 617 674 645
rect 82 337 132 417
rect 82 320 184 337
rect 292 336 342 417
rect 82 286 125 320
rect 159 286 184 320
rect 82 252 184 286
rect 82 218 125 252
rect 159 218 184 252
rect 82 202 184 218
rect 240 320 342 336
rect 402 329 452 417
rect 624 337 674 417
rect 240 286 269 320
rect 303 286 342 320
rect 240 265 342 286
rect 396 313 530 329
rect 396 279 412 313
rect 446 279 480 313
rect 514 279 530 313
rect 240 252 340 265
rect 240 218 269 252
rect 303 218 340 252
rect 396 263 530 279
rect 572 319 674 337
rect 572 285 595 319
rect 629 285 674 319
rect 396 229 426 263
rect 240 202 340 218
rect 82 177 112 202
rect 154 177 184 202
rect 310 177 340 202
rect 382 199 426 229
rect 572 251 674 285
rect 572 217 595 251
rect 629 217 674 251
rect 572 201 674 217
rect 382 177 412 199
rect 572 177 602 201
rect 644 177 674 201
rect 82 67 112 93
rect 154 67 184 93
rect 310 67 340 93
rect 382 67 412 93
rect 572 67 602 93
rect 644 67 674 93
<< polycont >>
rect 125 286 159 320
rect 125 218 159 252
rect 269 286 303 320
rect 412 279 446 313
rect 480 279 514 313
rect 269 218 303 252
rect 595 285 629 319
rect 595 217 629 251
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 31 599 75 615
rect 31 565 37 599
rect 71 565 75 599
rect 31 531 75 565
rect 31 497 37 531
rect 71 497 75 531
rect 31 463 75 497
rect 31 429 37 463
rect 71 429 75 463
rect 127 609 297 615
rect 127 575 143 609
rect 177 575 247 609
rect 281 575 297 609
rect 127 572 297 575
rect 127 538 143 572
rect 177 538 247 572
rect 281 538 297 572
rect 127 496 297 538
rect 127 462 143 496
rect 177 462 247 496
rect 281 462 297 496
rect 127 458 297 462
rect 353 599 395 615
rect 353 565 357 599
rect 391 565 395 599
rect 353 531 395 565
rect 353 497 357 531
rect 391 497 395 531
rect 353 463 395 497
rect 31 424 75 429
rect 353 429 357 463
rect 391 429 395 463
rect 447 609 629 615
rect 447 575 463 609
rect 497 575 579 609
rect 613 575 629 609
rect 447 572 629 575
rect 447 538 463 572
rect 497 538 579 572
rect 613 538 629 572
rect 447 496 629 538
rect 447 462 463 496
rect 497 462 579 496
rect 613 462 629 496
rect 447 459 629 462
rect 680 599 751 615
rect 680 565 685 599
rect 719 565 751 599
rect 680 531 751 565
rect 680 497 685 531
rect 719 497 751 531
rect 680 463 751 497
rect 353 425 395 429
rect 680 429 685 463
rect 719 429 751 463
rect 31 390 319 424
rect 353 391 646 425
rect 31 161 75 390
rect 109 320 184 356
rect 109 286 125 320
rect 159 286 184 320
rect 109 252 184 286
rect 109 218 125 252
rect 159 218 184 252
rect 109 202 184 218
rect 240 320 319 390
rect 240 286 269 320
rect 303 286 319 320
rect 240 252 319 286
rect 396 313 551 350
rect 396 279 412 313
rect 446 279 480 313
rect 514 279 551 313
rect 585 319 646 391
rect 585 285 595 319
rect 629 285 646 319
rect 240 218 269 252
rect 303 218 319 252
rect 585 251 646 285
rect 585 245 595 251
rect 240 202 319 218
rect 419 217 595 245
rect 629 217 646 251
rect 419 201 646 217
rect 31 127 37 161
rect 71 127 75 161
rect 31 86 75 127
rect 179 152 315 168
rect 179 118 195 152
rect 229 118 265 152
rect 299 118 315 152
rect 179 17 315 118
rect 419 161 461 201
rect 419 127 423 161
rect 457 127 461 161
rect 419 86 461 127
rect 510 161 577 167
rect 510 127 527 161
rect 561 127 577 161
rect 510 17 577 127
rect 680 161 751 429
rect 680 127 685 161
rect 719 127 751 161
rect 680 93 751 127
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 143 538 177 572
rect 247 538 281 572
rect 463 538 497 572
rect 579 538 613 572
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 14 572 754 578
rect 14 538 143 572
rect 177 538 247 572
rect 281 538 463 572
rect 497 538 579 572
rect 613 538 754 572
rect 14 532 754 538
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel locali s 511 316 545 350 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 200 0 0 0 SLEEP
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 200 0 0 0 SLEEP
port 2 nsew signal input
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 iso0p_lp2
flabel metal1 s 14 532 754 578 0 FreeSans 340 0 0 0 KAPWR
port 3 nsew power bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5919108
string GDS_START 5911916
<< end >>
