magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 5 246 451 259
rect 5 49 907 246
rect 0 0 960 49
<< scnmos >>
rect 84 65 114 233
rect 170 65 200 233
rect 256 65 286 233
rect 342 65 372 233
rect 540 52 570 220
rect 626 52 656 220
rect 712 52 742 220
rect 798 52 828 220
<< scpmoshvt >>
rect 84 367 114 619
rect 170 367 200 619
rect 256 367 286 619
rect 342 367 372 619
rect 540 367 570 619
rect 626 367 656 619
rect 712 367 742 619
rect 798 367 828 619
<< ndiff >>
rect 31 192 84 233
rect 31 158 39 192
rect 73 158 84 192
rect 31 111 84 158
rect 31 77 39 111
rect 73 77 84 111
rect 31 65 84 77
rect 114 225 170 233
rect 114 191 125 225
rect 159 191 170 225
rect 114 153 170 191
rect 114 119 125 153
rect 159 119 170 153
rect 114 65 170 119
rect 200 192 256 233
rect 200 158 211 192
rect 245 158 256 192
rect 200 111 256 158
rect 200 77 211 111
rect 245 77 256 111
rect 200 65 256 77
rect 286 201 342 233
rect 286 167 297 201
rect 331 167 342 201
rect 286 65 342 167
rect 372 113 425 233
rect 372 79 383 113
rect 417 79 425 113
rect 372 65 425 79
rect 487 121 540 220
rect 487 87 495 121
rect 529 87 540 121
rect 487 52 540 87
rect 570 208 626 220
rect 570 174 581 208
rect 615 174 626 208
rect 570 101 626 174
rect 570 67 581 101
rect 615 67 626 101
rect 570 52 626 67
rect 656 182 712 220
rect 656 148 667 182
rect 701 148 712 182
rect 656 98 712 148
rect 656 64 667 98
rect 701 64 712 98
rect 656 52 712 64
rect 742 208 798 220
rect 742 174 753 208
rect 787 174 798 208
rect 742 101 798 174
rect 742 67 753 101
rect 787 67 798 101
rect 742 52 798 67
rect 828 208 881 220
rect 828 174 839 208
rect 873 174 881 208
rect 828 98 881 174
rect 828 64 839 98
rect 873 64 881 98
rect 828 52 881 64
<< pdiff >>
rect 31 607 84 619
rect 31 573 39 607
rect 73 573 84 607
rect 31 510 84 573
rect 31 476 39 510
rect 73 476 84 510
rect 31 418 84 476
rect 31 384 39 418
rect 73 384 84 418
rect 31 367 84 384
rect 114 599 170 619
rect 114 565 125 599
rect 159 565 170 599
rect 114 503 170 565
rect 114 469 125 503
rect 159 469 170 503
rect 114 420 170 469
rect 114 386 125 420
rect 159 386 170 420
rect 114 367 170 386
rect 200 607 256 619
rect 200 573 211 607
rect 245 573 256 607
rect 200 528 256 573
rect 200 494 211 528
rect 245 494 256 528
rect 200 454 256 494
rect 200 420 211 454
rect 245 420 256 454
rect 200 367 256 420
rect 286 599 342 619
rect 286 565 297 599
rect 331 565 342 599
rect 286 508 342 565
rect 286 474 297 508
rect 331 474 342 508
rect 286 413 342 474
rect 286 379 297 413
rect 331 379 342 413
rect 286 367 342 379
rect 372 607 425 619
rect 372 573 383 607
rect 417 573 425 607
rect 372 539 425 573
rect 372 505 383 539
rect 417 505 425 539
rect 372 454 425 505
rect 372 420 383 454
rect 417 420 425 454
rect 372 367 425 420
rect 487 599 540 619
rect 487 565 495 599
rect 529 565 540 599
rect 487 470 540 565
rect 487 436 495 470
rect 529 436 540 470
rect 487 367 540 436
rect 570 547 626 619
rect 570 513 581 547
rect 615 513 626 547
rect 570 479 626 513
rect 570 445 581 479
rect 615 445 626 479
rect 570 411 626 445
rect 570 377 581 411
rect 615 377 626 411
rect 570 367 626 377
rect 656 599 712 619
rect 656 565 667 599
rect 701 565 712 599
rect 656 504 712 565
rect 656 470 667 504
rect 701 470 712 504
rect 656 413 712 470
rect 656 379 667 413
rect 701 379 712 413
rect 656 367 712 379
rect 742 607 798 619
rect 742 573 753 607
rect 787 573 798 607
rect 742 529 798 573
rect 742 495 753 529
rect 787 495 798 529
rect 742 454 798 495
rect 742 420 753 454
rect 787 420 798 454
rect 742 367 798 420
rect 828 599 881 619
rect 828 565 839 599
rect 873 565 881 599
rect 828 504 881 565
rect 828 470 839 504
rect 873 470 881 504
rect 828 413 881 470
rect 828 379 839 413
rect 873 379 881 413
rect 828 367 881 379
<< ndiffc >>
rect 39 158 73 192
rect 39 77 73 111
rect 125 191 159 225
rect 125 119 159 153
rect 211 158 245 192
rect 211 77 245 111
rect 297 167 331 201
rect 383 79 417 113
rect 495 87 529 121
rect 581 174 615 208
rect 581 67 615 101
rect 667 148 701 182
rect 667 64 701 98
rect 753 174 787 208
rect 753 67 787 101
rect 839 174 873 208
rect 839 64 873 98
<< pdiffc >>
rect 39 573 73 607
rect 39 476 73 510
rect 39 384 73 418
rect 125 565 159 599
rect 125 469 159 503
rect 125 386 159 420
rect 211 573 245 607
rect 211 494 245 528
rect 211 420 245 454
rect 297 565 331 599
rect 297 474 331 508
rect 297 379 331 413
rect 383 573 417 607
rect 383 505 417 539
rect 383 420 417 454
rect 495 565 529 599
rect 495 436 529 470
rect 581 513 615 547
rect 581 445 615 479
rect 581 377 615 411
rect 667 565 701 599
rect 667 470 701 504
rect 667 379 701 413
rect 753 573 787 607
rect 753 495 787 529
rect 753 420 787 454
rect 839 565 873 599
rect 839 470 873 504
rect 839 379 873 413
<< poly >>
rect 84 619 114 645
rect 170 619 200 645
rect 256 619 286 645
rect 342 619 372 645
rect 540 619 570 645
rect 626 619 656 645
rect 712 619 742 645
rect 798 619 828 645
rect 84 321 114 367
rect 170 321 200 367
rect 256 321 286 367
rect 342 321 372 367
rect 540 334 570 367
rect 626 334 656 367
rect 23 305 200 321
rect 23 271 39 305
rect 73 271 200 305
rect 23 255 200 271
rect 247 305 381 321
rect 540 318 656 334
rect 540 308 606 318
rect 247 271 263 305
rect 297 271 331 305
rect 365 271 381 305
rect 247 255 381 271
rect 495 292 606 308
rect 495 258 511 292
rect 545 284 606 292
rect 640 284 656 318
rect 545 258 656 284
rect 84 233 114 255
rect 170 233 200 255
rect 256 233 286 255
rect 342 233 372 255
rect 495 242 656 258
rect 540 220 570 242
rect 626 220 656 242
rect 712 334 742 367
rect 798 334 828 367
rect 712 318 828 334
rect 712 284 728 318
rect 762 308 828 318
rect 762 292 873 308
rect 762 284 823 292
rect 712 258 823 284
rect 857 258 873 292
rect 712 242 873 258
rect 712 220 742 242
rect 798 220 828 242
rect 84 39 114 65
rect 170 39 200 65
rect 256 39 286 65
rect 342 39 372 65
rect 540 26 570 52
rect 626 26 656 52
rect 712 26 742 52
rect 798 26 828 52
<< polycont >>
rect 39 271 73 305
rect 263 271 297 305
rect 331 271 365 305
rect 511 258 545 292
rect 606 284 640 318
rect 728 284 762 318
rect 823 258 857 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 607 89 649
rect 23 573 39 607
rect 73 573 89 607
rect 23 510 89 573
rect 23 476 39 510
rect 73 476 89 510
rect 23 418 89 476
rect 23 384 39 418
rect 73 384 89 418
rect 123 599 161 615
rect 123 565 125 599
rect 159 565 161 599
rect 123 503 161 565
rect 123 469 125 503
rect 159 469 161 503
rect 123 420 161 469
rect 195 607 261 649
rect 195 573 211 607
rect 245 573 261 607
rect 195 528 261 573
rect 195 494 211 528
rect 245 494 261 528
rect 195 454 261 494
rect 195 420 211 454
rect 245 420 261 454
rect 295 599 333 615
rect 295 565 297 599
rect 331 565 333 599
rect 295 508 333 565
rect 295 474 297 508
rect 331 474 333 508
rect 123 386 125 420
rect 159 386 161 420
rect 295 413 333 474
rect 367 607 433 649
rect 367 573 383 607
rect 417 573 433 607
rect 367 539 433 573
rect 367 505 383 539
rect 417 505 433 539
rect 367 454 433 505
rect 367 420 383 454
rect 417 420 433 454
rect 479 599 703 615
rect 479 565 495 599
rect 529 581 667 599
rect 529 565 531 581
rect 479 470 531 565
rect 665 565 667 581
rect 701 565 703 599
rect 479 436 495 470
rect 529 436 531 470
rect 479 420 531 436
rect 565 513 581 547
rect 615 513 631 547
rect 565 479 631 513
rect 565 445 581 479
rect 615 445 631 479
rect 295 386 297 413
rect 123 379 297 386
rect 331 386 333 413
rect 565 411 631 445
rect 565 386 581 411
rect 331 379 581 386
rect 123 377 581 379
rect 615 377 631 411
rect 123 352 631 377
rect 665 504 703 565
rect 665 470 667 504
rect 701 470 703 504
rect 665 413 703 470
rect 737 607 803 649
rect 737 573 753 607
rect 787 573 803 607
rect 737 529 803 573
rect 737 495 753 529
rect 787 495 803 529
rect 737 454 803 495
rect 737 420 753 454
rect 787 420 803 454
rect 837 599 889 615
rect 837 565 839 599
rect 873 565 889 599
rect 837 504 889 565
rect 837 470 839 504
rect 873 470 889 504
rect 665 379 667 413
rect 701 386 703 413
rect 837 413 889 470
rect 837 386 839 413
rect 701 379 839 386
rect 873 379 889 413
rect 665 352 889 379
rect 17 305 89 350
rect 17 271 39 305
rect 73 271 89 305
rect 17 257 89 271
rect 17 242 77 257
rect 123 229 175 352
rect 209 271 263 305
rect 297 271 331 305
rect 365 271 381 305
rect 209 242 381 271
rect 415 292 606 318
rect 415 258 511 292
rect 545 284 606 292
rect 640 284 656 318
rect 712 284 728 318
rect 762 292 943 318
rect 762 284 823 292
rect 545 258 547 284
rect 415 239 547 258
rect 857 258 943 292
rect 109 225 175 229
rect 19 192 75 208
rect 19 158 39 192
rect 73 158 75 192
rect 19 111 75 158
rect 109 191 125 225
rect 159 191 175 225
rect 581 216 789 250
rect 823 242 943 258
rect 581 208 617 216
rect 109 153 175 191
rect 109 119 125 153
rect 159 119 175 153
rect 209 192 247 208
rect 209 158 211 192
rect 245 158 247 192
rect 281 201 581 205
rect 281 167 297 201
rect 331 174 581 201
rect 615 174 617 208
rect 751 208 789 216
rect 331 167 617 174
rect 281 163 617 167
rect 209 129 247 158
rect 19 77 39 111
rect 73 85 75 111
rect 209 113 433 129
rect 209 111 383 113
rect 209 85 211 111
rect 73 77 211 85
rect 245 79 383 111
rect 417 79 433 113
rect 245 77 433 79
rect 19 51 433 77
rect 479 121 545 129
rect 479 87 495 121
rect 529 87 545 121
rect 479 17 545 87
rect 579 101 617 163
rect 579 67 581 101
rect 615 67 617 101
rect 579 51 617 67
rect 651 148 667 182
rect 701 148 717 182
rect 651 98 717 148
rect 651 64 667 98
rect 701 64 717 98
rect 651 17 717 64
rect 751 174 753 208
rect 787 174 789 208
rect 751 101 789 174
rect 751 67 753 101
rect 787 67 789 101
rect 751 51 789 67
rect 823 174 839 208
rect 873 174 889 208
rect 823 98 889 174
rect 823 64 839 98
rect 873 64 889 98
rect 823 17 889 64
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o211ai_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6903808
string GDS_START 6894108
<< end >>
