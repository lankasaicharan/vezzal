magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 5 49 2015 259
rect 0 0 2016 49
<< scnmos >>
rect 88 65 118 233
rect 190 65 220 233
rect 276 65 306 233
rect 362 65 392 233
rect 448 65 478 233
rect 534 65 564 233
rect 620 65 650 233
rect 722 65 752 233
rect 808 65 838 233
rect 894 65 924 233
rect 982 65 1012 233
rect 1082 65 1112 233
rect 1288 65 1318 233
rect 1390 65 1420 233
rect 1476 65 1506 233
rect 1562 65 1592 233
rect 1648 65 1678 233
rect 1734 65 1764 233
rect 1820 65 1850 233
rect 1906 65 1936 233
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 284 367 314 619
rect 370 367 400 619
rect 456 367 486 619
rect 542 367 572 619
rect 628 367 658 619
rect 714 367 744 619
rect 808 367 838 619
rect 894 367 924 619
rect 1125 367 1155 619
rect 1211 367 1241 619
rect 1297 367 1327 619
rect 1383 367 1413 619
rect 1469 367 1499 619
rect 1555 367 1585 619
rect 1641 367 1671 619
rect 1727 367 1757 619
rect 1813 367 1843 619
rect 1899 367 1929 619
<< ndiff >>
rect 31 181 88 233
rect 31 147 43 181
rect 77 147 88 181
rect 31 109 88 147
rect 31 75 43 109
rect 77 75 88 109
rect 31 65 88 75
rect 118 107 190 233
rect 118 73 143 107
rect 177 73 190 107
rect 118 65 190 73
rect 220 181 276 233
rect 220 147 231 181
rect 265 147 276 181
rect 220 113 276 147
rect 220 79 231 113
rect 265 79 276 113
rect 220 65 276 79
rect 306 107 362 233
rect 306 73 317 107
rect 351 73 362 107
rect 306 65 362 73
rect 392 181 448 233
rect 392 147 403 181
rect 437 147 448 181
rect 392 113 448 147
rect 392 79 403 113
rect 437 79 448 113
rect 392 65 448 79
rect 478 107 534 233
rect 478 73 489 107
rect 523 73 534 107
rect 478 65 534 73
rect 564 181 620 233
rect 564 147 575 181
rect 609 147 620 181
rect 564 107 620 147
rect 564 73 575 107
rect 609 73 620 107
rect 564 65 620 73
rect 650 107 722 233
rect 650 73 661 107
rect 695 73 722 107
rect 650 65 722 73
rect 752 181 808 233
rect 752 147 763 181
rect 797 147 808 181
rect 752 107 808 147
rect 752 73 763 107
rect 797 73 808 107
rect 752 65 808 73
rect 838 171 894 233
rect 838 137 849 171
rect 883 137 894 171
rect 838 65 894 137
rect 924 181 982 233
rect 924 147 937 181
rect 971 147 982 181
rect 924 107 982 147
rect 924 73 937 107
rect 971 73 982 107
rect 924 65 982 73
rect 1012 225 1082 233
rect 1012 191 1037 225
rect 1071 191 1082 225
rect 1012 153 1082 191
rect 1012 119 1037 153
rect 1071 119 1082 153
rect 1012 65 1082 119
rect 1112 183 1181 233
rect 1112 149 1137 183
rect 1171 149 1181 183
rect 1112 111 1181 149
rect 1112 77 1137 111
rect 1171 77 1181 111
rect 1112 65 1181 77
rect 1235 183 1288 233
rect 1235 149 1243 183
rect 1277 149 1288 183
rect 1235 111 1288 149
rect 1235 77 1243 111
rect 1277 77 1288 111
rect 1235 65 1288 77
rect 1318 107 1390 233
rect 1318 73 1343 107
rect 1377 73 1390 107
rect 1318 65 1390 73
rect 1420 183 1476 233
rect 1420 149 1431 183
rect 1465 149 1476 183
rect 1420 107 1476 149
rect 1420 73 1431 107
rect 1465 73 1476 107
rect 1420 65 1476 73
rect 1506 107 1562 233
rect 1506 73 1517 107
rect 1551 73 1562 107
rect 1506 65 1562 73
rect 1592 167 1648 233
rect 1592 133 1603 167
rect 1637 133 1648 167
rect 1592 65 1648 133
rect 1678 225 1734 233
rect 1678 191 1689 225
rect 1723 191 1734 225
rect 1678 157 1734 191
rect 1678 123 1689 157
rect 1723 123 1734 157
rect 1678 65 1734 123
rect 1764 163 1820 233
rect 1764 129 1775 163
rect 1809 129 1820 163
rect 1764 65 1820 129
rect 1850 225 1906 233
rect 1850 191 1861 225
rect 1895 191 1906 225
rect 1850 157 1906 191
rect 1850 123 1861 157
rect 1895 123 1906 157
rect 1850 65 1906 123
rect 1936 163 1989 233
rect 1936 129 1947 163
rect 1981 129 1989 163
rect 1936 65 1989 129
<< pdiff >>
rect 211 630 269 638
rect 211 619 223 630
rect 27 607 80 619
rect 27 573 35 607
rect 69 573 80 607
rect 27 490 80 573
rect 27 456 35 490
rect 69 456 80 490
rect 27 367 80 456
rect 110 574 166 619
rect 110 540 121 574
rect 155 540 166 574
rect 110 367 166 540
rect 196 596 223 619
rect 257 619 269 630
rect 257 596 284 619
rect 196 367 284 596
rect 314 576 370 619
rect 314 542 325 576
rect 359 542 370 576
rect 314 367 370 542
rect 400 490 456 619
rect 400 456 411 490
rect 445 456 456 490
rect 400 367 456 456
rect 486 576 542 619
rect 486 542 497 576
rect 531 542 542 576
rect 486 367 542 542
rect 572 490 628 619
rect 572 456 583 490
rect 617 456 628 490
rect 572 367 628 456
rect 658 576 714 619
rect 658 542 669 576
rect 703 542 714 576
rect 658 367 714 542
rect 744 566 808 619
rect 744 532 759 566
rect 793 532 808 566
rect 744 367 808 532
rect 838 599 894 619
rect 838 565 849 599
rect 883 565 894 599
rect 838 529 894 565
rect 838 495 849 529
rect 883 495 894 529
rect 838 461 894 495
rect 838 427 849 461
rect 883 427 894 461
rect 838 367 894 427
rect 924 611 1125 619
rect 924 577 963 611
rect 997 577 1080 611
rect 1114 577 1125 611
rect 924 543 1125 577
rect 924 509 963 543
rect 997 523 1125 543
rect 997 509 1080 523
rect 924 489 1080 509
rect 1114 489 1125 523
rect 924 367 1125 489
rect 1155 599 1211 619
rect 1155 565 1166 599
rect 1200 565 1211 599
rect 1155 527 1211 565
rect 1155 493 1166 527
rect 1200 493 1211 527
rect 1155 455 1211 493
rect 1155 421 1166 455
rect 1200 421 1211 455
rect 1155 367 1211 421
rect 1241 611 1297 619
rect 1241 577 1252 611
rect 1286 577 1297 611
rect 1241 543 1297 577
rect 1241 509 1252 543
rect 1286 509 1297 543
rect 1241 475 1297 509
rect 1241 441 1252 475
rect 1286 441 1297 475
rect 1241 367 1297 441
rect 1327 599 1383 619
rect 1327 565 1338 599
rect 1372 565 1383 599
rect 1327 507 1383 565
rect 1327 473 1338 507
rect 1372 473 1383 507
rect 1327 409 1383 473
rect 1327 375 1338 409
rect 1372 375 1383 409
rect 1327 367 1383 375
rect 1413 611 1469 619
rect 1413 577 1424 611
rect 1458 577 1469 611
rect 1413 536 1469 577
rect 1413 502 1424 536
rect 1458 502 1469 536
rect 1413 459 1469 502
rect 1413 425 1424 459
rect 1458 425 1469 459
rect 1413 367 1469 425
rect 1499 599 1555 619
rect 1499 565 1510 599
rect 1544 565 1555 599
rect 1499 507 1555 565
rect 1499 473 1510 507
rect 1544 473 1555 507
rect 1499 409 1555 473
rect 1499 375 1510 409
rect 1544 375 1555 409
rect 1499 367 1555 375
rect 1585 611 1641 619
rect 1585 577 1596 611
rect 1630 577 1641 611
rect 1585 490 1641 577
rect 1585 456 1596 490
rect 1630 456 1641 490
rect 1585 367 1641 456
rect 1671 599 1727 619
rect 1671 565 1682 599
rect 1716 565 1727 599
rect 1671 507 1727 565
rect 1671 473 1682 507
rect 1716 473 1727 507
rect 1671 418 1727 473
rect 1671 384 1682 418
rect 1716 384 1727 418
rect 1671 367 1727 384
rect 1757 611 1813 619
rect 1757 577 1768 611
rect 1802 577 1813 611
rect 1757 490 1813 577
rect 1757 456 1768 490
rect 1802 456 1813 490
rect 1757 367 1813 456
rect 1843 599 1899 619
rect 1843 565 1854 599
rect 1888 565 1899 599
rect 1843 507 1899 565
rect 1843 473 1854 507
rect 1888 473 1899 507
rect 1843 418 1899 473
rect 1843 384 1854 418
rect 1888 384 1899 418
rect 1843 367 1899 384
rect 1929 607 1982 619
rect 1929 573 1940 607
rect 1974 573 1982 607
rect 1929 490 1982 573
rect 1929 456 1940 490
rect 1974 456 1982 490
rect 1929 367 1982 456
<< ndiffc >>
rect 43 147 77 181
rect 43 75 77 109
rect 143 73 177 107
rect 231 147 265 181
rect 231 79 265 113
rect 317 73 351 107
rect 403 147 437 181
rect 403 79 437 113
rect 489 73 523 107
rect 575 147 609 181
rect 575 73 609 107
rect 661 73 695 107
rect 763 147 797 181
rect 763 73 797 107
rect 849 137 883 171
rect 937 147 971 181
rect 937 73 971 107
rect 1037 191 1071 225
rect 1037 119 1071 153
rect 1137 149 1171 183
rect 1137 77 1171 111
rect 1243 149 1277 183
rect 1243 77 1277 111
rect 1343 73 1377 107
rect 1431 149 1465 183
rect 1431 73 1465 107
rect 1517 73 1551 107
rect 1603 133 1637 167
rect 1689 191 1723 225
rect 1689 123 1723 157
rect 1775 129 1809 163
rect 1861 191 1895 225
rect 1861 123 1895 157
rect 1947 129 1981 163
<< pdiffc >>
rect 35 573 69 607
rect 35 456 69 490
rect 121 540 155 574
rect 223 596 257 630
rect 325 542 359 576
rect 411 456 445 490
rect 497 542 531 576
rect 583 456 617 490
rect 669 542 703 576
rect 759 532 793 566
rect 849 565 883 599
rect 849 495 883 529
rect 849 427 883 461
rect 963 577 997 611
rect 1080 577 1114 611
rect 963 509 997 543
rect 1080 489 1114 523
rect 1166 565 1200 599
rect 1166 493 1200 527
rect 1166 421 1200 455
rect 1252 577 1286 611
rect 1252 509 1286 543
rect 1252 441 1286 475
rect 1338 565 1372 599
rect 1338 473 1372 507
rect 1338 375 1372 409
rect 1424 577 1458 611
rect 1424 502 1458 536
rect 1424 425 1458 459
rect 1510 565 1544 599
rect 1510 473 1544 507
rect 1510 375 1544 409
rect 1596 577 1630 611
rect 1596 456 1630 490
rect 1682 565 1716 599
rect 1682 473 1716 507
rect 1682 384 1716 418
rect 1768 577 1802 611
rect 1768 456 1802 490
rect 1854 565 1888 599
rect 1854 473 1888 507
rect 1854 384 1888 418
rect 1940 573 1974 607
rect 1940 456 1974 490
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 284 619 314 645
rect 370 619 400 645
rect 456 619 486 645
rect 542 619 572 645
rect 628 619 658 645
rect 714 619 744 645
rect 808 619 838 645
rect 894 619 924 645
rect 1125 619 1155 645
rect 1211 619 1241 645
rect 1297 619 1327 645
rect 1383 619 1413 645
rect 1469 619 1499 645
rect 1555 619 1585 645
rect 1641 619 1671 645
rect 1727 619 1757 645
rect 1813 619 1843 645
rect 1899 619 1929 645
rect 80 335 110 367
rect 166 335 196 367
rect 284 335 314 367
rect 370 335 400 367
rect 456 335 486 367
rect 542 335 572 367
rect 628 335 658 367
rect 714 335 744 367
rect 80 319 314 335
rect 80 285 105 319
rect 139 285 173 319
rect 207 285 241 319
rect 275 285 314 319
rect 80 269 314 285
rect 362 319 658 335
rect 362 285 378 319
rect 412 285 446 319
rect 480 285 514 319
rect 548 285 582 319
rect 616 305 658 319
rect 700 319 766 335
rect 616 285 650 305
rect 362 269 650 285
rect 700 285 716 319
rect 750 285 766 319
rect 700 269 766 285
rect 808 333 838 367
rect 894 333 924 367
rect 1125 333 1155 367
rect 1211 333 1241 367
rect 1297 335 1327 367
rect 1383 335 1413 367
rect 1469 335 1499 367
rect 1555 335 1585 367
rect 1641 345 1671 367
rect 1727 345 1757 367
rect 1813 345 1843 367
rect 1899 345 1929 367
rect 1641 335 1929 345
rect 808 317 1246 333
rect 808 283 824 317
rect 858 283 892 317
rect 926 283 960 317
rect 994 283 1028 317
rect 1062 283 1096 317
rect 1130 283 1164 317
rect 1198 283 1246 317
rect 88 233 118 269
rect 190 233 220 269
rect 276 233 306 269
rect 362 233 392 269
rect 448 233 478 269
rect 534 233 564 269
rect 620 233 650 269
rect 722 233 752 269
rect 808 267 1246 283
rect 1288 319 1592 335
rect 1288 285 1320 319
rect 1354 285 1388 319
rect 1422 285 1456 319
rect 1490 285 1524 319
rect 1558 285 1592 319
rect 1641 319 1936 335
rect 1641 315 1664 319
rect 1288 269 1592 285
rect 808 233 838 267
rect 894 233 924 267
rect 982 233 1012 267
rect 1082 233 1112 267
rect 1288 233 1318 269
rect 1390 233 1420 269
rect 1476 233 1506 269
rect 1562 233 1592 269
rect 1648 285 1664 315
rect 1698 285 1732 319
rect 1766 285 1800 319
rect 1834 285 1868 319
rect 1902 285 1936 319
rect 1648 269 1936 285
rect 1648 233 1678 269
rect 1734 233 1764 269
rect 1820 233 1850 269
rect 1906 233 1936 269
rect 88 39 118 65
rect 190 39 220 65
rect 276 39 306 65
rect 362 39 392 65
rect 448 39 478 65
rect 534 39 564 65
rect 620 39 650 65
rect 722 39 752 65
rect 808 39 838 65
rect 894 39 924 65
rect 982 39 1012 65
rect 1082 39 1112 65
rect 1288 39 1318 65
rect 1390 39 1420 65
rect 1476 39 1506 65
rect 1562 39 1592 65
rect 1648 39 1678 65
rect 1734 39 1764 65
rect 1820 39 1850 65
rect 1906 39 1936 65
<< polycont >>
rect 105 285 139 319
rect 173 285 207 319
rect 241 285 275 319
rect 378 285 412 319
rect 446 285 480 319
rect 514 285 548 319
rect 582 285 616 319
rect 716 285 750 319
rect 824 283 858 317
rect 892 283 926 317
rect 960 283 994 317
rect 1028 283 1062 317
rect 1096 283 1130 317
rect 1164 283 1198 317
rect 1320 285 1354 319
rect 1388 285 1422 319
rect 1456 285 1490 319
rect 1524 285 1558 319
rect 1664 285 1698 319
rect 1732 285 1766 319
rect 1800 285 1834 319
rect 1868 285 1902 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 19 607 85 649
rect 19 573 35 607
rect 69 573 85 607
rect 207 630 273 649
rect 207 596 223 630
rect 257 596 273 630
rect 207 592 273 596
rect 19 490 85 573
rect 119 574 173 590
rect 119 540 121 574
rect 155 558 173 574
rect 307 576 709 592
rect 307 558 325 576
rect 155 542 325 558
rect 359 542 497 576
rect 531 542 669 576
rect 703 542 709 576
rect 155 540 709 542
rect 119 524 709 540
rect 743 566 809 649
rect 743 532 759 566
rect 793 532 809 566
rect 743 524 809 532
rect 843 599 929 615
rect 843 565 849 599
rect 883 565 929 599
rect 843 529 929 565
rect 843 495 849 529
rect 883 495 929 529
rect 843 490 929 495
rect 19 456 35 490
rect 69 456 85 490
rect 19 452 85 456
rect 189 456 411 490
rect 445 456 583 490
rect 617 461 929 490
rect 963 611 1130 649
rect 997 577 1080 611
rect 1114 577 1130 611
rect 963 543 1130 577
rect 997 523 1130 543
rect 997 509 1080 523
rect 963 489 1080 509
rect 1114 489 1130 523
rect 1164 599 1216 615
rect 1164 565 1166 599
rect 1200 565 1216 599
rect 1164 527 1216 565
rect 1164 493 1166 527
rect 1200 493 1216 527
rect 617 456 849 461
rect 189 454 849 456
rect 189 418 223 454
rect 833 427 849 454
rect 883 455 929 461
rect 1164 455 1216 493
rect 883 427 1166 455
rect 833 421 1166 427
rect 1200 421 1216 455
rect 1250 611 1294 649
rect 1250 577 1252 611
rect 1286 577 1294 611
rect 1250 543 1294 577
rect 1250 509 1252 543
rect 1286 509 1294 543
rect 1250 475 1294 509
rect 1250 441 1252 475
rect 1286 441 1294 475
rect 1250 425 1294 441
rect 1329 599 1374 615
rect 1329 565 1338 599
rect 1372 565 1374 599
rect 1329 507 1374 565
rect 1329 473 1338 507
rect 1372 473 1374 507
rect 19 384 223 418
rect 257 387 734 420
rect 1329 409 1374 473
rect 1408 611 1474 649
rect 1408 577 1424 611
rect 1458 577 1474 611
rect 1408 536 1474 577
rect 1408 502 1424 536
rect 1458 502 1474 536
rect 1408 459 1474 502
rect 1408 425 1424 459
rect 1458 425 1474 459
rect 1508 599 1546 615
rect 1508 565 1510 599
rect 1544 565 1546 599
rect 1508 507 1546 565
rect 1508 473 1510 507
rect 1544 473 1546 507
rect 257 386 1295 387
rect 19 249 55 384
rect 257 350 314 386
rect 700 353 1295 386
rect 1329 375 1338 409
rect 1372 389 1374 409
rect 1508 418 1546 473
rect 1580 611 1646 649
rect 1580 577 1596 611
rect 1630 577 1646 611
rect 1580 490 1646 577
rect 1580 456 1596 490
rect 1630 456 1646 490
rect 1580 452 1646 456
rect 1680 599 1718 615
rect 1680 565 1682 599
rect 1716 565 1718 599
rect 1680 507 1718 565
rect 1680 473 1682 507
rect 1716 473 1718 507
rect 1680 418 1718 473
rect 1752 611 1818 649
rect 1752 577 1768 611
rect 1802 577 1818 611
rect 1752 490 1818 577
rect 1752 456 1768 490
rect 1802 456 1818 490
rect 1752 452 1818 456
rect 1852 599 1890 615
rect 1852 565 1854 599
rect 1888 565 1890 599
rect 1852 507 1890 565
rect 1852 473 1854 507
rect 1888 473 1890 507
rect 1852 418 1890 473
rect 1924 607 1990 649
rect 1924 573 1940 607
rect 1974 573 1990 607
rect 1924 490 1990 573
rect 1924 456 1940 490
rect 1974 456 1990 490
rect 1924 452 1990 456
rect 1508 409 1682 418
rect 1508 389 1510 409
rect 1372 375 1510 389
rect 1544 384 1682 409
rect 1716 384 1854 418
rect 1888 384 1998 418
rect 1544 375 1560 384
rect 1329 355 1560 375
rect 89 319 314 350
rect 449 319 632 350
rect 89 285 105 319
rect 139 285 173 319
rect 207 285 241 319
rect 275 285 314 319
rect 89 283 314 285
rect 362 285 378 319
rect 412 316 415 319
rect 412 285 446 316
rect 480 285 514 319
rect 548 285 582 319
rect 616 285 632 319
rect 362 283 632 285
rect 700 319 766 353
rect 700 285 716 319
rect 750 285 766 319
rect 1261 319 1295 353
rect 700 283 766 285
rect 808 283 824 317
rect 858 283 892 317
rect 926 283 960 317
rect 994 283 1028 317
rect 1062 283 1096 317
rect 1130 283 1164 317
rect 1198 283 1227 317
rect 1261 285 1320 319
rect 1354 285 1388 319
rect 1422 285 1456 319
rect 1490 285 1524 319
rect 1558 285 1592 319
rect 1648 316 1663 350
rect 1697 319 1918 350
rect 1648 285 1664 316
rect 1698 285 1732 319
rect 1766 285 1800 319
rect 1834 285 1868 319
rect 1902 285 1918 319
rect 1125 251 1227 283
rect 1954 251 1998 384
rect 19 225 1087 249
rect 19 215 1037 225
rect 27 147 43 181
rect 77 147 231 181
rect 265 147 403 181
rect 437 147 575 181
rect 609 147 763 181
rect 797 147 813 181
rect 27 109 93 147
rect 231 113 267 147
rect 401 113 439 147
rect 27 75 43 109
rect 77 75 93 109
rect 27 59 93 75
rect 127 107 193 113
rect 127 73 143 107
rect 177 73 193 107
rect 127 17 193 73
rect 265 79 267 113
rect 231 57 267 79
rect 301 107 367 113
rect 301 73 317 107
rect 351 73 367 107
rect 301 17 367 73
rect 401 79 403 113
rect 437 79 439 113
rect 401 57 439 79
rect 473 107 539 113
rect 473 73 489 107
rect 523 73 539 107
rect 473 17 539 73
rect 573 107 611 147
rect 573 73 575 107
rect 609 73 611 107
rect 573 57 611 73
rect 645 107 711 113
rect 645 73 661 107
rect 695 73 711 107
rect 645 17 711 73
rect 747 107 813 147
rect 847 171 887 215
rect 1021 191 1037 215
rect 1071 191 1087 225
rect 1125 225 1998 251
rect 1125 217 1689 225
rect 847 137 849 171
rect 883 137 887 171
rect 847 121 887 137
rect 921 147 937 181
rect 971 147 987 181
rect 747 73 763 107
rect 797 87 813 107
rect 921 107 987 147
rect 1021 153 1087 191
rect 1673 191 1689 217
rect 1723 213 1861 225
rect 1723 191 1739 213
rect 1021 119 1037 153
rect 1071 119 1087 153
rect 1121 149 1137 183
rect 1171 149 1187 183
rect 921 87 937 107
rect 797 73 937 87
rect 971 85 987 107
rect 1121 111 1187 149
rect 1121 85 1137 111
rect 971 77 1137 85
rect 1171 77 1187 111
rect 971 73 1187 77
rect 747 51 1187 73
rect 1227 149 1243 183
rect 1277 149 1431 183
rect 1465 167 1639 183
rect 1465 149 1603 167
rect 1227 111 1293 149
rect 1227 77 1243 111
rect 1277 77 1293 111
rect 1227 61 1293 77
rect 1327 107 1393 115
rect 1327 73 1343 107
rect 1377 73 1393 107
rect 1327 17 1393 73
rect 1427 107 1467 149
rect 1601 133 1603 149
rect 1637 133 1639 167
rect 1427 73 1431 107
rect 1465 73 1467 107
rect 1427 57 1467 73
rect 1501 107 1567 115
rect 1501 73 1517 107
rect 1551 73 1567 107
rect 1501 17 1567 73
rect 1601 87 1639 133
rect 1673 157 1739 191
rect 1845 191 1861 213
rect 1895 213 1998 225
rect 1895 191 1911 213
rect 1673 123 1689 157
rect 1723 123 1739 157
rect 1773 163 1811 179
rect 1773 129 1775 163
rect 1809 129 1811 163
rect 1773 87 1811 129
rect 1845 157 1911 191
rect 1845 123 1861 157
rect 1895 123 1911 157
rect 1945 163 1997 179
rect 1945 129 1947 163
rect 1981 129 1997 163
rect 1601 85 1811 87
rect 1945 85 1997 129
rect 1601 51 1997 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 415 319 449 350
rect 415 316 446 319
rect 446 316 449 319
rect 1663 319 1697 350
rect 1663 316 1664 319
rect 1664 316 1697 319
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 403 350 461 356
rect 403 316 415 350
rect 449 347 461 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 449 319 1663 347
rect 449 316 461 319
rect 403 310 461 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xnor2_4
flabel metal1 s 1663 316 1697 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 464 929 498 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 895 538 929 572 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4285878
string GDS_START 4270914
<< end >>
