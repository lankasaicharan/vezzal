magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 1 49 863 157
rect 0 0 864 49
<< scnmos >>
rect 84 47 114 131
rect 156 47 186 131
rect 354 47 384 131
rect 426 47 456 131
rect 504 47 534 131
rect 582 47 612 131
rect 678 47 708 131
rect 750 47 780 131
<< scpmoshvt >>
rect 120 419 170 619
rect 226 419 276 619
rect 332 419 382 619
rect 500 419 550 619
rect 606 419 656 619
rect 720 419 770 619
<< ndiff >>
rect 27 111 84 131
rect 27 77 39 111
rect 73 77 84 111
rect 27 47 84 77
rect 114 47 156 131
rect 186 106 243 131
rect 186 72 197 106
rect 231 72 243 106
rect 186 47 243 72
rect 297 111 354 131
rect 297 77 309 111
rect 343 77 354 111
rect 297 47 354 77
rect 384 47 426 131
rect 456 47 504 131
rect 534 47 582 131
rect 612 97 678 131
rect 612 63 623 97
rect 657 63 678 97
rect 612 47 678 63
rect 708 47 750 131
rect 780 97 837 131
rect 780 63 791 97
rect 825 63 837 97
rect 780 47 837 63
<< pdiff >>
rect 63 597 120 619
rect 63 563 75 597
rect 109 563 120 597
rect 63 465 120 563
rect 63 431 75 465
rect 109 431 120 465
rect 63 419 120 431
rect 170 607 226 619
rect 170 573 181 607
rect 215 573 226 607
rect 170 536 226 573
rect 170 502 181 536
rect 215 502 226 536
rect 170 465 226 502
rect 170 431 181 465
rect 215 431 226 465
rect 170 419 226 431
rect 276 597 332 619
rect 276 563 287 597
rect 321 563 332 597
rect 276 508 332 563
rect 276 474 287 508
rect 321 474 332 508
rect 276 419 332 474
rect 382 598 500 619
rect 382 564 393 598
rect 427 564 500 598
rect 382 419 500 564
rect 550 597 606 619
rect 550 563 561 597
rect 595 563 606 597
rect 550 516 606 563
rect 550 482 561 516
rect 595 482 606 516
rect 550 419 606 482
rect 656 607 720 619
rect 656 573 667 607
rect 701 573 720 607
rect 656 516 720 573
rect 656 482 667 516
rect 701 482 720 516
rect 656 419 720 482
rect 770 597 827 619
rect 770 563 781 597
rect 815 563 827 597
rect 770 465 827 563
rect 770 431 781 465
rect 815 431 827 465
rect 770 419 827 431
<< ndiffc >>
rect 39 77 73 111
rect 197 72 231 106
rect 309 77 343 111
rect 623 63 657 97
rect 791 63 825 97
<< pdiffc >>
rect 75 563 109 597
rect 75 431 109 465
rect 181 573 215 607
rect 181 502 215 536
rect 181 431 215 465
rect 287 563 321 597
rect 287 474 321 508
rect 393 564 427 598
rect 561 563 595 597
rect 561 482 595 516
rect 667 573 701 607
rect 667 482 701 516
rect 781 563 815 597
rect 781 431 815 465
<< poly >>
rect 120 619 170 645
rect 226 619 276 645
rect 332 619 382 645
rect 500 619 550 645
rect 606 619 656 645
rect 720 619 770 645
rect 120 305 170 419
rect 226 379 276 419
rect 218 363 284 379
rect 218 329 234 363
rect 268 329 284 363
rect 332 352 382 419
rect 500 387 550 419
rect 606 387 656 419
rect 498 371 564 387
rect 84 289 159 305
rect 84 255 109 289
rect 143 255 159 289
rect 84 221 159 255
rect 218 295 284 329
rect 218 261 234 295
rect 268 261 284 295
rect 218 245 284 261
rect 84 187 109 221
rect 143 197 159 221
rect 143 187 186 197
rect 84 167 186 187
rect 84 131 114 167
rect 156 131 186 167
rect 254 176 284 245
rect 352 336 456 352
rect 352 302 406 336
rect 440 302 456 336
rect 498 337 514 371
rect 548 337 564 371
rect 498 321 564 337
rect 606 371 672 387
rect 606 337 622 371
rect 656 337 672 371
rect 606 321 672 337
rect 352 268 456 302
rect 352 234 406 268
rect 440 234 456 268
rect 352 218 456 234
rect 254 146 384 176
rect 354 131 384 146
rect 426 131 456 218
rect 504 131 534 321
rect 606 176 636 321
rect 720 219 770 419
rect 582 146 636 176
rect 678 203 780 219
rect 678 169 694 203
rect 728 169 780 203
rect 678 153 780 169
rect 582 131 612 146
rect 678 131 708 153
rect 750 131 780 153
rect 84 21 114 47
rect 156 21 186 47
rect 354 21 384 47
rect 426 21 456 47
rect 504 21 534 47
rect 582 21 612 47
rect 678 21 708 47
rect 750 21 780 47
<< polycont >>
rect 234 329 268 363
rect 109 255 143 289
rect 234 261 268 295
rect 109 187 143 221
rect 406 302 440 336
rect 514 337 548 371
rect 622 337 656 371
rect 406 234 440 268
rect 694 169 728 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 597 125 613
rect 23 563 75 597
rect 109 563 125 597
rect 23 465 125 563
rect 23 431 75 465
rect 109 431 125 465
rect 23 379 125 431
rect 165 607 231 649
rect 165 573 181 607
rect 215 573 231 607
rect 165 536 231 573
rect 165 502 181 536
rect 215 502 231 536
rect 165 465 231 502
rect 165 431 181 465
rect 215 431 231 465
rect 271 597 337 613
rect 271 563 287 597
rect 321 563 337 597
rect 271 508 337 563
rect 377 598 443 649
rect 377 564 393 598
rect 427 564 443 598
rect 377 540 443 564
rect 545 597 611 613
rect 545 563 561 597
rect 595 563 611 597
rect 271 474 287 508
rect 321 504 337 508
rect 545 516 611 563
rect 545 504 561 516
rect 321 482 561 504
rect 595 482 611 516
rect 321 474 611 482
rect 271 466 611 474
rect 651 607 717 649
rect 651 573 667 607
rect 701 573 717 607
rect 651 516 717 573
rect 651 482 667 516
rect 701 482 717 516
rect 651 466 717 482
rect 765 597 841 613
rect 765 563 781 597
rect 815 563 841 597
rect 271 458 337 466
rect 165 415 231 431
rect 409 422 455 466
rect 765 465 841 563
rect 765 431 781 465
rect 815 431 841 465
rect 320 388 455 422
rect 23 363 284 379
rect 23 345 234 363
rect 23 135 57 345
rect 218 329 234 345
rect 268 329 284 363
rect 93 289 167 305
rect 93 255 109 289
rect 143 255 167 289
rect 93 221 167 255
rect 218 295 284 329
rect 218 261 234 295
rect 268 261 284 295
rect 218 245 284 261
rect 93 187 109 221
rect 143 187 167 221
rect 93 171 167 187
rect 320 135 354 388
rect 498 371 564 430
rect 390 336 456 352
rect 390 302 406 336
rect 440 302 456 336
rect 498 337 514 371
rect 548 337 564 371
rect 498 323 564 337
rect 601 371 672 430
rect 601 337 622 371
rect 656 337 672 371
rect 601 323 672 337
rect 390 287 456 302
rect 765 287 841 431
rect 390 268 841 287
rect 390 234 406 268
rect 440 253 841 268
rect 440 234 456 253
rect 390 218 456 234
rect 505 203 744 217
rect 505 169 694 203
rect 728 169 744 203
rect 505 153 744 169
rect 23 111 89 135
rect 23 77 39 111
rect 73 77 89 111
rect 23 53 89 77
rect 181 106 247 135
rect 181 72 197 106
rect 231 72 247 106
rect 181 17 247 72
rect 293 111 359 135
rect 807 117 841 253
rect 293 77 309 111
rect 343 77 359 111
rect 293 53 359 77
rect 607 97 673 117
rect 607 63 623 97
rect 657 63 673 97
rect 607 17 673 63
rect 775 97 841 117
rect 775 63 791 97
rect 825 63 841 97
rect 775 59 841 63
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4bb_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5690218
string GDS_START 5682912
<< end >>
