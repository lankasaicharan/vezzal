magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 16 49 1110 263
rect 0 0 1152 49
<< scnmos >>
rect 95 69 125 237
rect 181 69 211 237
rect 267 69 297 237
rect 353 69 383 237
rect 555 69 585 237
rect 641 69 671 237
rect 743 69 773 237
rect 829 69 859 237
rect 915 69 945 237
rect 1001 69 1031 237
<< scpmoshvt >>
rect 95 367 125 619
rect 181 367 211 619
rect 267 367 297 619
rect 353 367 383 619
rect 555 367 585 619
rect 641 367 671 619
rect 735 367 765 619
rect 821 367 851 619
rect 915 367 945 619
rect 1001 367 1031 619
<< ndiff >>
rect 42 225 95 237
rect 42 191 50 225
rect 84 191 95 225
rect 42 115 95 191
rect 42 81 50 115
rect 84 81 95 115
rect 42 69 95 81
rect 125 202 181 237
rect 125 168 136 202
rect 170 168 181 202
rect 125 111 181 168
rect 125 77 136 111
rect 170 77 181 111
rect 125 69 181 77
rect 211 204 267 237
rect 211 170 222 204
rect 256 170 267 204
rect 211 69 267 170
rect 297 116 353 237
rect 297 82 308 116
rect 342 82 353 116
rect 297 69 353 82
rect 383 124 436 237
rect 383 90 394 124
rect 428 90 436 124
rect 383 69 436 90
rect 502 225 555 237
rect 502 191 510 225
rect 544 191 555 225
rect 502 115 555 191
rect 502 81 510 115
rect 544 81 555 115
rect 502 69 555 81
rect 585 229 641 237
rect 585 195 596 229
rect 630 195 641 229
rect 585 153 641 195
rect 585 119 596 153
rect 630 119 641 153
rect 585 69 641 119
rect 671 192 743 237
rect 671 158 690 192
rect 724 158 743 192
rect 671 111 743 158
rect 671 77 690 111
rect 724 77 743 111
rect 671 69 743 77
rect 773 132 829 237
rect 773 98 784 132
rect 818 98 829 132
rect 773 69 829 98
rect 859 208 915 237
rect 859 174 870 208
rect 904 174 915 208
rect 859 115 915 174
rect 859 81 870 115
rect 904 81 915 115
rect 859 69 915 81
rect 945 132 1001 237
rect 945 98 956 132
rect 990 98 1001 132
rect 945 69 1001 98
rect 1031 192 1084 237
rect 1031 158 1042 192
rect 1076 158 1084 192
rect 1031 115 1084 158
rect 1031 81 1042 115
rect 1076 81 1084 115
rect 1031 69 1084 81
<< pdiff >>
rect 42 607 95 619
rect 42 573 50 607
rect 84 573 95 607
rect 42 492 95 573
rect 42 458 50 492
rect 84 458 95 492
rect 42 367 95 458
rect 125 599 181 619
rect 125 565 136 599
rect 170 565 181 599
rect 125 502 181 565
rect 125 468 136 502
rect 170 468 181 502
rect 125 367 181 468
rect 211 562 267 619
rect 211 528 222 562
rect 256 528 267 562
rect 211 367 267 528
rect 297 599 353 619
rect 297 565 308 599
rect 342 565 353 599
rect 297 486 353 565
rect 297 452 308 486
rect 342 452 353 486
rect 297 367 353 452
rect 383 611 555 619
rect 383 577 510 611
rect 544 577 555 611
rect 383 574 555 577
rect 383 540 394 574
rect 428 540 555 574
rect 383 516 555 540
rect 383 482 510 516
rect 544 482 555 516
rect 383 413 555 482
rect 383 379 510 413
rect 544 379 555 413
rect 383 367 555 379
rect 585 599 641 619
rect 585 565 596 599
rect 630 565 641 599
rect 585 504 641 565
rect 585 470 596 504
rect 630 470 641 504
rect 585 409 641 470
rect 585 375 596 409
rect 630 375 641 409
rect 585 367 641 375
rect 671 602 735 619
rect 671 568 686 602
rect 720 568 735 602
rect 671 367 735 568
rect 765 596 821 619
rect 765 562 776 596
rect 810 562 821 596
rect 765 367 821 562
rect 851 502 915 619
rect 851 468 866 502
rect 900 468 915 502
rect 851 367 915 468
rect 945 599 1001 619
rect 945 565 956 599
rect 990 565 1001 599
rect 945 502 1001 565
rect 945 468 956 502
rect 990 468 1001 502
rect 945 367 1001 468
rect 1031 607 1084 619
rect 1031 573 1042 607
rect 1076 573 1084 607
rect 1031 490 1084 573
rect 1031 456 1042 490
rect 1076 456 1084 490
rect 1031 367 1084 456
<< ndiffc >>
rect 50 191 84 225
rect 50 81 84 115
rect 136 168 170 202
rect 136 77 170 111
rect 222 170 256 204
rect 308 82 342 116
rect 394 90 428 124
rect 510 191 544 225
rect 510 81 544 115
rect 596 195 630 229
rect 596 119 630 153
rect 690 158 724 192
rect 690 77 724 111
rect 784 98 818 132
rect 870 174 904 208
rect 870 81 904 115
rect 956 98 990 132
rect 1042 158 1076 192
rect 1042 81 1076 115
<< pdiffc >>
rect 50 573 84 607
rect 50 458 84 492
rect 136 565 170 599
rect 136 468 170 502
rect 222 528 256 562
rect 308 565 342 599
rect 308 452 342 486
rect 510 577 544 611
rect 394 540 428 574
rect 510 482 544 516
rect 510 379 544 413
rect 596 565 630 599
rect 596 470 630 504
rect 596 375 630 409
rect 686 568 720 602
rect 776 562 810 596
rect 866 468 900 502
rect 956 565 990 599
rect 956 468 990 502
rect 1042 573 1076 607
rect 1042 456 1076 490
<< poly >>
rect 95 619 125 645
rect 181 619 211 645
rect 267 619 297 645
rect 353 619 383 645
rect 555 619 585 645
rect 641 619 671 645
rect 735 619 765 645
rect 821 619 851 645
rect 915 619 945 645
rect 1001 619 1031 645
rect 95 335 125 367
rect 59 319 125 335
rect 59 285 75 319
rect 109 285 125 319
rect 59 269 125 285
rect 95 237 125 269
rect 181 325 211 367
rect 267 325 297 367
rect 353 325 383 367
rect 181 309 297 325
rect 181 275 213 309
rect 247 275 297 309
rect 181 259 297 275
rect 339 309 405 325
rect 339 275 355 309
rect 389 275 405 309
rect 339 259 405 275
rect 447 309 513 325
rect 447 275 463 309
rect 497 289 513 309
rect 555 289 585 367
rect 641 289 671 367
rect 735 335 765 367
rect 497 275 671 289
rect 447 259 671 275
rect 713 319 779 335
rect 713 285 729 319
rect 763 285 779 319
rect 713 269 779 285
rect 821 325 851 367
rect 915 325 945 367
rect 1001 325 1031 367
rect 821 309 955 325
rect 821 275 837 309
rect 871 275 905 309
rect 939 275 955 309
rect 181 237 211 259
rect 267 237 297 259
rect 353 237 383 259
rect 555 237 585 259
rect 641 237 671 259
rect 743 237 773 269
rect 821 259 955 275
rect 1001 309 1131 325
rect 1001 275 1081 309
rect 1115 275 1131 309
rect 1001 259 1131 275
rect 829 237 859 259
rect 915 237 945 259
rect 1001 237 1031 259
rect 95 43 125 69
rect 181 43 211 69
rect 267 43 297 69
rect 353 43 383 69
rect 555 43 585 69
rect 641 43 671 69
rect 743 43 773 69
rect 829 43 859 69
rect 915 43 945 69
rect 1001 43 1031 69
<< polycont >>
rect 75 285 109 319
rect 213 275 247 309
rect 355 275 389 309
rect 463 275 497 309
rect 729 285 763 319
rect 837 275 871 309
rect 905 275 939 309
rect 1081 275 1115 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 34 607 100 649
rect 34 573 50 607
rect 84 573 100 607
rect 34 492 100 573
rect 34 458 50 492
rect 84 458 100 492
rect 34 454 100 458
rect 134 599 172 615
rect 134 565 136 599
rect 170 565 172 599
rect 134 502 172 565
rect 206 562 272 649
rect 206 528 222 562
rect 256 528 272 562
rect 206 520 272 528
rect 306 599 351 615
rect 306 565 308 599
rect 342 565 351 599
rect 134 468 136 502
rect 170 486 172 502
rect 306 490 351 565
rect 385 611 546 649
rect 385 577 510 611
rect 544 577 546 611
rect 385 574 546 577
rect 385 540 394 574
rect 428 540 546 574
rect 385 524 546 540
rect 504 516 546 524
rect 306 486 470 490
rect 170 468 308 486
rect 134 452 308 468
rect 342 452 470 486
rect 17 384 402 418
rect 17 319 161 384
rect 17 285 75 319
rect 109 285 161 319
rect 17 275 161 285
rect 197 309 291 350
rect 197 275 213 309
rect 247 275 291 309
rect 197 242 291 275
rect 339 309 402 384
rect 339 275 355 309
rect 389 275 402 309
rect 339 259 402 275
rect 436 325 470 452
rect 504 482 510 516
rect 544 482 546 516
rect 504 413 546 482
rect 504 379 510 413
rect 544 379 546 413
rect 504 363 546 379
rect 580 599 646 615
rect 580 565 596 599
rect 630 565 646 599
rect 580 518 646 565
rect 680 602 726 649
rect 680 568 686 602
rect 720 568 726 602
rect 680 552 726 568
rect 760 599 990 615
rect 760 596 956 599
rect 760 562 776 596
rect 810 565 956 596
rect 810 562 990 565
rect 760 552 990 562
rect 580 504 910 518
rect 580 470 596 504
rect 630 502 910 504
rect 630 470 866 502
rect 580 468 866 470
rect 900 468 910 502
rect 580 452 910 468
rect 944 502 990 552
rect 944 468 956 502
rect 944 452 990 468
rect 1026 607 1092 649
rect 1026 573 1042 607
rect 1076 573 1092 607
rect 1026 490 1092 573
rect 1026 456 1042 490
rect 1076 456 1092 490
rect 1026 452 1092 456
rect 580 409 646 452
rect 580 375 596 409
rect 630 375 646 409
rect 436 309 513 325
rect 436 275 463 309
rect 497 275 513 309
rect 34 225 95 241
rect 34 191 50 225
rect 84 191 95 225
rect 34 115 95 191
rect 34 81 50 115
rect 84 81 95 115
rect 34 17 95 81
rect 129 202 172 218
rect 436 208 470 275
rect 129 168 136 202
rect 170 168 172 202
rect 129 132 172 168
rect 206 204 470 208
rect 206 170 222 204
rect 256 170 470 204
rect 206 166 470 170
rect 504 225 546 241
rect 504 191 510 225
rect 544 191 546 225
rect 129 116 342 132
rect 129 111 308 116
rect 129 77 136 111
rect 170 82 308 111
rect 170 77 342 82
rect 129 61 342 77
rect 378 124 444 132
rect 378 90 394 124
rect 428 90 444 124
rect 378 17 444 90
rect 504 115 546 191
rect 580 229 646 375
rect 713 384 1135 418
rect 713 319 763 384
rect 713 285 729 319
rect 713 269 763 285
rect 799 309 1031 350
rect 799 275 837 309
rect 871 275 905 309
rect 939 275 1031 309
rect 799 242 1031 275
rect 1065 309 1135 384
rect 1065 275 1081 309
rect 1115 275 1135 309
rect 1065 259 1135 275
rect 580 195 596 229
rect 630 195 646 229
rect 580 153 646 195
rect 580 119 596 153
rect 630 119 646 153
rect 682 192 870 208
rect 682 158 690 192
rect 724 174 870 192
rect 904 192 1092 208
rect 904 174 1042 192
rect 724 158 734 174
rect 504 81 510 115
rect 544 85 546 115
rect 682 111 734 158
rect 682 85 690 111
rect 544 81 690 85
rect 504 77 690 81
rect 724 77 734 111
rect 504 51 734 77
rect 768 132 834 140
rect 768 98 784 132
rect 818 98 834 132
rect 768 17 834 98
rect 868 115 906 174
rect 1040 158 1042 174
rect 1076 158 1092 192
rect 868 81 870 115
rect 904 81 906 115
rect 868 65 906 81
rect 940 132 1006 140
rect 940 98 956 132
rect 990 98 1006 132
rect 940 17 1006 98
rect 1040 115 1092 158
rect 1040 81 1042 115
rect 1076 81 1092 115
rect 1040 65 1092 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2bb2ai_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4090354
string GDS_START 4079916
<< end >>
