magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 331 1478 704
rect 737 285 905 331
<< pwell >>
rect 741 241 1153 243
rect 7 230 196 241
rect 7 191 199 230
rect 741 191 1429 241
rect 7 49 1429 191
rect 0 0 1440 49
<< scnmos >>
rect 90 47 120 215
rect 228 81 258 165
rect 300 81 330 165
rect 386 81 416 165
rect 480 81 510 165
rect 589 81 619 165
rect 847 133 877 217
rect 972 133 1002 217
rect 1044 133 1074 217
rect 1234 47 1264 215
rect 1320 47 1350 215
<< scpmoshvt >>
rect 87 367 117 619
rect 212 465 242 593
rect 284 465 314 593
rect 392 465 422 549
rect 464 465 494 549
rect 589 391 619 519
rect 891 367 921 495
rect 1009 367 1039 495
rect 1114 367 1144 495
rect 1234 367 1264 619
rect 1320 367 1350 619
<< ndiff >>
rect 33 203 90 215
rect 33 169 41 203
rect 75 169 90 203
rect 33 101 90 169
rect 33 67 41 101
rect 75 67 90 101
rect 33 47 90 67
rect 120 204 170 215
rect 120 165 173 204
rect 767 209 847 217
rect 767 175 779 209
rect 813 175 847 209
rect 120 95 228 165
rect 120 61 131 95
rect 165 81 228 95
rect 258 81 300 165
rect 330 155 386 165
rect 330 121 341 155
rect 375 121 386 155
rect 330 81 386 121
rect 416 81 480 165
rect 510 137 589 165
rect 510 103 540 137
rect 574 103 589 137
rect 510 81 589 103
rect 619 135 672 165
rect 619 101 630 135
rect 664 101 672 135
rect 767 133 847 175
rect 877 133 972 217
rect 1002 133 1044 217
rect 1074 192 1127 217
rect 1074 158 1085 192
rect 1119 158 1127 192
rect 1074 133 1127 158
rect 1181 167 1234 215
rect 1181 133 1189 167
rect 1223 133 1234 167
rect 619 81 672 101
rect 165 61 173 81
rect 120 47 173 61
rect 892 69 950 133
rect 892 35 904 69
rect 938 35 950 69
rect 1181 93 1234 133
rect 1181 59 1189 93
rect 1223 59 1234 93
rect 1181 47 1234 59
rect 1264 203 1320 215
rect 1264 169 1275 203
rect 1309 169 1320 203
rect 1264 101 1320 169
rect 1264 67 1275 101
rect 1309 67 1320 101
rect 1264 47 1320 67
rect 1350 203 1403 215
rect 1350 169 1361 203
rect 1395 169 1403 203
rect 1350 93 1403 169
rect 1350 59 1361 93
rect 1395 59 1403 93
rect 1350 47 1403 59
rect 892 27 950 35
<< pdiff >>
rect 132 630 190 638
rect 132 619 144 630
rect 34 556 87 619
rect 34 522 42 556
rect 76 522 87 556
rect 34 488 87 522
rect 34 454 42 488
rect 76 454 87 488
rect 34 420 87 454
rect 34 386 42 420
rect 76 386 87 420
rect 34 367 87 386
rect 117 596 144 619
rect 178 596 190 630
rect 117 593 190 596
rect 117 465 212 593
rect 242 465 284 593
rect 314 549 367 593
rect 516 573 574 581
rect 516 549 528 573
rect 314 531 392 549
rect 314 497 325 531
rect 359 497 392 531
rect 314 465 392 497
rect 422 465 464 549
rect 494 539 528 549
rect 562 539 574 573
rect 1181 607 1234 619
rect 936 573 994 581
rect 494 519 574 539
rect 936 539 948 573
rect 982 539 994 573
rect 494 465 589 519
rect 117 367 190 465
rect 516 393 589 465
rect 539 391 589 393
rect 619 433 676 519
rect 936 495 994 539
rect 1181 573 1189 607
rect 1223 573 1234 607
rect 1181 525 1234 573
rect 1181 495 1189 525
rect 619 399 630 433
rect 664 399 676 433
rect 619 391 676 399
rect 811 367 891 495
rect 921 367 1009 495
rect 1039 483 1114 495
rect 1039 449 1060 483
rect 1094 449 1114 483
rect 1039 413 1114 449
rect 1039 379 1060 413
rect 1094 379 1114 413
rect 1039 367 1114 379
rect 1144 491 1189 495
rect 1223 491 1234 525
rect 1144 443 1234 491
rect 1144 409 1171 443
rect 1205 409 1234 443
rect 1144 367 1234 409
rect 1264 599 1320 619
rect 1264 565 1275 599
rect 1309 565 1320 599
rect 1264 507 1320 565
rect 1264 473 1275 507
rect 1309 473 1320 507
rect 1264 413 1320 473
rect 1264 379 1275 413
rect 1309 379 1320 413
rect 1264 367 1320 379
rect 1350 607 1403 619
rect 1350 573 1361 607
rect 1395 573 1403 607
rect 1350 507 1403 573
rect 1350 473 1361 507
rect 1395 473 1403 507
rect 1350 413 1403 473
rect 1350 379 1361 413
rect 1395 379 1403 413
rect 1350 367 1403 379
rect 811 363 869 367
rect 811 329 823 363
rect 857 329 869 363
rect 811 321 869 329
<< ndiffc >>
rect 41 169 75 203
rect 41 67 75 101
rect 779 175 813 209
rect 131 61 165 95
rect 341 121 375 155
rect 540 103 574 137
rect 630 101 664 135
rect 1085 158 1119 192
rect 1189 133 1223 167
rect 904 35 938 69
rect 1189 59 1223 93
rect 1275 169 1309 203
rect 1275 67 1309 101
rect 1361 169 1395 203
rect 1361 59 1395 93
<< pdiffc >>
rect 42 522 76 556
rect 42 454 76 488
rect 42 386 76 420
rect 144 596 178 630
rect 325 497 359 531
rect 528 539 562 573
rect 948 539 982 573
rect 1189 573 1223 607
rect 630 399 664 433
rect 1060 449 1094 483
rect 1060 379 1094 413
rect 1189 491 1223 525
rect 1171 409 1205 443
rect 1275 565 1309 599
rect 1275 473 1309 507
rect 1275 379 1309 413
rect 1361 573 1395 607
rect 1361 473 1395 507
rect 1361 379 1395 413
rect 823 329 857 363
<< poly >>
rect 87 619 117 645
rect 212 593 242 619
rect 284 593 314 619
rect 464 605 733 626
rect 1234 619 1264 645
rect 1320 619 1350 645
rect 464 596 683 605
rect 392 549 422 575
rect 464 549 494 596
rect 667 571 683 596
rect 717 571 733 605
rect 667 555 733 571
rect 589 519 619 545
rect 87 335 117 367
rect 78 319 144 335
rect 78 285 94 319
rect 128 285 144 319
rect 212 292 242 465
rect 284 433 314 465
rect 284 417 350 433
rect 284 383 300 417
rect 334 383 350 417
rect 284 367 350 383
rect 392 361 422 465
rect 464 439 494 465
rect 891 495 921 521
rect 1009 495 1039 521
rect 1114 495 1144 521
rect 392 345 507 361
rect 392 325 457 345
rect 300 311 457 325
rect 491 311 507 345
rect 300 295 507 311
rect 589 321 619 391
rect 703 326 769 342
rect 589 305 655 321
rect 78 269 144 285
rect 192 276 258 292
rect 90 215 120 269
rect 192 242 208 276
rect 242 242 258 276
rect 192 217 258 242
rect 228 165 258 217
rect 300 165 330 295
rect 589 271 605 305
rect 639 271 655 305
rect 703 292 719 326
rect 753 306 769 326
rect 891 345 921 367
rect 1009 345 1039 367
rect 891 315 1039 345
rect 1114 321 1144 367
rect 1234 335 1264 367
rect 891 306 1002 315
rect 753 292 1002 306
rect 703 276 1002 292
rect 372 237 438 253
rect 372 203 388 237
rect 422 203 438 237
rect 372 187 438 203
rect 480 237 546 253
rect 480 203 496 237
rect 530 203 546 237
rect 480 187 546 203
rect 589 237 655 271
rect 589 203 605 237
rect 639 203 655 237
rect 847 217 877 276
rect 972 217 1002 276
rect 1081 305 1147 321
rect 1081 273 1097 305
rect 1044 271 1097 273
rect 1131 271 1147 305
rect 1044 243 1147 271
rect 1189 319 1264 335
rect 1189 285 1205 319
rect 1239 299 1264 319
rect 1320 299 1350 367
rect 1239 285 1350 299
rect 1189 269 1350 285
rect 1044 217 1074 243
rect 589 187 655 203
rect 386 165 416 187
rect 480 165 510 187
rect 589 165 619 187
rect 1234 215 1264 269
rect 1320 215 1350 269
rect 847 107 877 133
rect 228 55 258 81
rect 300 55 330 81
rect 386 55 416 81
rect 480 55 510 81
rect 589 55 619 81
rect 972 107 1002 133
rect 1044 107 1074 133
rect 90 21 120 47
rect 1234 21 1264 47
rect 1320 21 1350 47
<< polycont >>
rect 683 571 717 605
rect 94 285 128 319
rect 300 383 334 417
rect 457 311 491 345
rect 208 242 242 276
rect 605 271 639 305
rect 719 292 753 326
rect 388 203 422 237
rect 496 203 530 237
rect 605 203 639 237
rect 1097 271 1131 305
rect 1205 285 1239 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 128 630 194 649
rect 128 596 144 630
rect 178 596 194 630
rect 128 594 194 596
rect 230 581 433 615
rect 230 560 264 581
rect 24 556 264 560
rect 24 522 42 556
rect 76 526 264 556
rect 309 531 365 547
rect 76 522 92 526
rect 24 488 92 522
rect 309 497 325 531
rect 359 497 365 531
rect 309 490 365 497
rect 24 454 42 488
rect 76 454 92 488
rect 24 420 92 454
rect 24 386 42 420
rect 76 386 92 420
rect 24 382 92 386
rect 214 456 365 490
rect 399 503 433 581
rect 512 573 578 649
rect 512 539 528 573
rect 562 539 578 573
rect 512 537 578 539
rect 667 605 733 615
rect 667 571 683 605
rect 717 571 733 605
rect 667 503 733 571
rect 932 573 998 649
rect 932 539 948 573
rect 982 539 998 573
rect 932 537 998 539
rect 1155 607 1239 649
rect 1155 573 1189 607
rect 1223 573 1239 607
rect 1155 525 1239 573
rect 399 469 1009 503
rect 24 219 58 382
rect 214 346 248 456
rect 614 433 941 435
rect 614 422 630 433
rect 284 417 630 422
rect 284 383 300 417
rect 334 399 630 417
rect 664 399 941 433
rect 334 397 941 399
rect 334 386 680 397
rect 334 383 405 386
rect 284 380 405 383
rect 92 319 335 346
rect 92 285 94 319
rect 128 312 335 319
rect 128 285 144 312
rect 92 269 144 285
rect 192 276 267 278
rect 192 242 208 276
rect 242 242 267 276
rect 192 226 267 242
rect 24 203 91 219
rect 24 169 41 203
rect 75 169 91 203
rect 24 167 91 169
rect 301 169 335 312
rect 371 253 405 380
rect 441 345 647 352
rect 441 311 457 345
rect 491 311 647 345
rect 441 305 647 311
rect 441 295 605 305
rect 639 271 647 305
rect 687 326 769 352
rect 687 292 719 326
rect 753 292 769 326
rect 807 329 823 363
rect 857 329 873 363
rect 371 237 438 253
rect 371 203 388 237
rect 422 203 438 237
rect 472 237 546 253
rect 472 203 496 237
rect 530 203 546 237
rect 472 187 546 203
rect 605 237 647 271
rect 639 213 647 237
rect 807 213 873 329
rect 639 209 873 213
rect 639 203 779 209
rect 24 133 251 167
rect 24 101 81 133
rect 24 67 41 101
rect 75 67 81 101
rect 24 51 81 67
rect 115 95 181 99
rect 115 61 131 95
rect 165 61 181 95
rect 115 17 181 61
rect 215 87 251 133
rect 301 155 391 169
rect 301 121 341 155
rect 375 121 391 155
rect 472 87 506 187
rect 605 175 779 203
rect 813 175 873 209
rect 215 53 506 87
rect 540 137 578 153
rect 907 139 941 397
rect 975 307 1009 469
rect 1043 483 1110 499
rect 1043 449 1060 483
rect 1094 449 1110 483
rect 1043 413 1110 449
rect 1043 379 1060 413
rect 1094 379 1110 413
rect 1155 491 1189 525
rect 1223 491 1239 525
rect 1155 443 1239 491
rect 1155 409 1171 443
rect 1205 409 1239 443
rect 1273 599 1318 615
rect 1273 565 1275 599
rect 1309 565 1318 599
rect 1273 507 1318 565
rect 1273 473 1275 507
rect 1309 473 1318 507
rect 1273 413 1318 473
rect 1043 375 1110 379
rect 1273 379 1275 413
rect 1309 379 1318 413
rect 1043 341 1239 375
rect 1189 319 1239 341
rect 975 305 1147 307
rect 975 271 1097 305
rect 1131 271 1147 305
rect 975 269 1147 271
rect 1189 285 1205 319
rect 1189 235 1239 285
rect 1069 201 1239 235
rect 1273 203 1318 379
rect 1357 607 1411 649
rect 1357 573 1361 607
rect 1395 573 1411 607
rect 1357 507 1411 573
rect 1357 473 1361 507
rect 1395 473 1411 507
rect 1357 413 1411 473
rect 1357 379 1361 413
rect 1395 379 1411 413
rect 1357 363 1411 379
rect 1069 192 1135 201
rect 1069 158 1085 192
rect 1119 158 1135 192
rect 1273 169 1275 203
rect 1309 169 1318 203
rect 1069 142 1135 158
rect 574 103 578 137
rect 540 17 578 103
rect 614 135 941 139
rect 614 101 630 135
rect 664 105 941 135
rect 1173 133 1189 167
rect 1223 133 1239 167
rect 664 101 680 105
rect 614 97 680 101
rect 1173 93 1239 133
rect 888 35 904 69
rect 938 35 954 69
rect 888 17 954 35
rect 1173 59 1189 93
rect 1223 59 1239 93
rect 1173 17 1239 59
rect 1273 101 1318 169
rect 1273 67 1275 101
rect 1309 67 1318 101
rect 1273 51 1318 67
rect 1352 203 1411 219
rect 1352 169 1361 203
rect 1395 169 1411 203
rect 1352 93 1411 169
rect 1352 59 1361 93
rect 1395 59 1411 93
rect 1352 17 1411 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlclkp_2
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 1279 94 1313 128 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1279 168 1313 202 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1279 464 1313 498 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1279 538 1313 572 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3513240
string GDS_START 3501994
<< end >>
