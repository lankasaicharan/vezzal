magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 7 49 671 241
rect 0 0 672 49
<< scnmos >>
rect 86 47 116 215
rect 165 47 195 215
rect 355 47 385 215
rect 463 47 493 215
rect 562 47 592 215
<< scpmoshvt >>
rect 86 367 116 619
rect 172 367 202 619
rect 355 367 385 619
rect 463 367 493 619
rect 562 367 592 619
<< ndiff >>
rect 33 187 86 215
rect 33 153 41 187
rect 75 153 86 187
rect 33 93 86 153
rect 33 59 41 93
rect 75 59 86 93
rect 33 47 86 59
rect 116 47 165 215
rect 195 183 248 215
rect 195 149 206 183
rect 240 149 248 183
rect 195 93 248 149
rect 195 59 206 93
rect 240 59 248 93
rect 195 47 248 59
rect 302 183 355 215
rect 302 149 310 183
rect 344 149 355 183
rect 302 93 355 149
rect 302 59 310 93
rect 344 59 355 93
rect 302 47 355 59
rect 385 108 463 215
rect 385 74 410 108
rect 444 74 463 108
rect 385 47 463 74
rect 493 183 562 215
rect 493 149 517 183
rect 551 149 562 183
rect 493 93 562 149
rect 493 59 517 93
rect 551 59 562 93
rect 493 47 562 59
rect 592 203 645 215
rect 592 169 603 203
rect 637 169 645 203
rect 592 101 645 169
rect 592 67 603 101
rect 637 67 645 101
rect 592 47 645 67
<< pdiff >>
rect 33 607 86 619
rect 33 573 41 607
rect 75 573 86 607
rect 33 502 86 573
rect 33 468 41 502
rect 75 468 86 502
rect 33 367 86 468
rect 116 599 172 619
rect 116 565 127 599
rect 161 565 172 599
rect 116 486 172 565
rect 116 452 127 486
rect 161 452 172 486
rect 116 367 172 452
rect 202 562 355 619
rect 202 528 213 562
rect 247 528 310 562
rect 344 528 355 562
rect 202 367 355 528
rect 385 367 463 619
rect 493 599 562 619
rect 493 565 517 599
rect 551 565 562 599
rect 493 511 562 565
rect 493 477 517 511
rect 551 477 562 511
rect 493 367 562 477
rect 592 587 645 619
rect 592 553 603 587
rect 637 553 645 587
rect 592 367 645 553
<< ndiffc >>
rect 41 153 75 187
rect 41 59 75 93
rect 206 149 240 183
rect 206 59 240 93
rect 310 149 344 183
rect 310 59 344 93
rect 410 74 444 108
rect 517 149 551 183
rect 517 59 551 93
rect 603 169 637 203
rect 603 67 637 101
<< pdiffc >>
rect 41 573 75 607
rect 41 468 75 502
rect 127 565 161 599
rect 127 452 161 486
rect 213 528 247 562
rect 310 528 344 562
rect 517 565 551 599
rect 517 477 551 511
rect 603 553 637 587
<< poly >>
rect 86 619 116 645
rect 172 619 202 645
rect 355 619 385 645
rect 463 619 493 645
rect 562 619 592 645
rect 86 303 116 367
rect 172 335 202 367
rect 355 335 385 367
rect 463 335 493 367
rect 562 335 592 367
rect 38 287 116 303
rect 38 253 54 287
rect 88 253 116 287
rect 38 237 116 253
rect 158 319 385 335
rect 158 285 174 319
rect 208 285 281 319
rect 315 285 385 319
rect 158 237 385 285
rect 427 319 493 335
rect 427 285 443 319
rect 477 285 493 319
rect 427 269 493 285
rect 535 319 601 335
rect 535 285 551 319
rect 585 285 601 319
rect 535 269 601 285
rect 86 215 116 237
rect 165 215 195 237
rect 355 215 385 237
rect 463 215 493 269
rect 562 215 592 269
rect 86 21 116 47
rect 165 21 195 47
rect 355 21 385 47
rect 463 21 493 47
rect 562 21 592 47
<< polycont >>
rect 54 253 88 287
rect 174 285 208 319
rect 281 285 315 319
rect 443 285 477 319
rect 551 285 585 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 25 607 77 649
rect 25 573 41 607
rect 75 573 77 607
rect 25 502 77 573
rect 25 468 41 502
rect 75 468 77 502
rect 25 452 77 468
rect 111 599 163 615
rect 111 565 127 599
rect 161 565 163 599
rect 111 486 163 565
rect 197 562 365 649
rect 197 528 213 562
rect 247 528 310 562
rect 344 528 365 562
rect 197 520 365 528
rect 501 599 553 615
rect 501 565 517 599
rect 551 565 553 599
rect 501 511 553 565
rect 587 587 653 649
rect 587 553 603 587
rect 637 553 653 587
rect 587 545 653 553
rect 111 452 127 486
rect 161 452 467 486
rect 501 477 517 511
rect 551 477 655 511
rect 501 471 655 477
rect 433 437 467 452
rect 17 384 399 418
rect 433 403 569 437
rect 17 287 88 384
rect 365 369 399 384
rect 17 253 54 287
rect 127 319 331 350
rect 127 285 174 319
rect 208 285 281 319
rect 315 285 331 319
rect 365 319 493 369
rect 365 285 443 319
rect 477 285 493 319
rect 535 335 569 403
rect 603 369 655 471
rect 535 319 585 335
rect 535 285 551 319
rect 17 237 88 253
rect 535 269 585 285
rect 535 251 569 269
rect 122 217 569 251
rect 619 235 655 369
rect 122 203 156 217
rect 25 187 156 203
rect 25 153 41 187
rect 75 169 156 187
rect 603 203 655 235
rect 75 153 91 169
rect 25 93 91 153
rect 25 59 41 93
rect 75 59 91 93
rect 25 53 91 59
rect 190 149 206 183
rect 240 149 256 183
rect 190 93 256 149
rect 190 59 206 93
rect 240 59 256 93
rect 190 17 256 59
rect 294 149 310 183
rect 344 149 517 183
rect 551 149 567 183
rect 294 93 360 149
rect 294 59 310 93
rect 344 59 360 93
rect 294 51 360 59
rect 394 108 460 115
rect 394 74 410 108
rect 444 74 460 108
rect 394 17 460 74
rect 501 93 567 149
rect 501 59 517 93
rect 551 59 567 93
rect 501 51 567 59
rect 637 169 655 203
rect 603 101 655 169
rect 637 67 655 101
rect 603 51 655 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xnor2_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4292220
string GDS_START 4285934
<< end >>
