magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 1361 241 1629 247
rect 1 157 433 212
rect 1092 157 1629 241
rect 1 49 1629 157
rect 0 0 1632 49
<< scnmos >>
rect 84 102 114 186
rect 156 102 186 186
rect 248 102 278 186
rect 320 102 350 186
rect 554 47 584 131
rect 632 47 662 131
rect 760 47 790 131
rect 838 47 868 131
rect 952 47 982 131
rect 1030 47 1060 131
rect 1168 47 1198 215
rect 1246 47 1276 215
rect 1444 53 1474 221
rect 1516 53 1546 221
<< scpmoshvt >>
rect 84 470 114 598
rect 162 470 192 598
rect 248 470 278 598
rect 320 470 350 598
rect 520 491 550 619
rect 598 491 628 619
rect 716 491 746 619
rect 794 491 824 619
rect 903 535 933 619
rect 1027 535 1057 619
rect 1174 367 1204 619
rect 1246 367 1276 619
rect 1444 367 1474 619
rect 1516 367 1546 619
<< ndiff >>
rect 27 161 84 186
rect 27 127 39 161
rect 73 127 84 161
rect 27 102 84 127
rect 114 102 156 186
rect 186 161 248 186
rect 186 127 197 161
rect 231 127 248 161
rect 186 102 248 127
rect 278 102 320 186
rect 350 161 407 186
rect 350 127 361 161
rect 395 127 407 161
rect 1118 131 1168 215
rect 350 102 407 127
rect 497 111 554 131
rect 497 77 509 111
rect 543 77 554 111
rect 497 47 554 77
rect 584 47 632 131
rect 662 93 760 131
rect 662 59 673 93
rect 707 59 760 93
rect 662 47 760 59
rect 790 47 838 131
rect 868 111 952 131
rect 868 77 907 111
rect 941 77 952 111
rect 868 47 952 77
rect 982 47 1030 131
rect 1060 106 1168 131
rect 1060 72 1072 106
rect 1106 72 1168 106
rect 1060 47 1168 72
rect 1198 47 1246 215
rect 1276 203 1333 215
rect 1276 169 1287 203
rect 1321 169 1333 203
rect 1276 103 1333 169
rect 1276 69 1287 103
rect 1321 69 1333 103
rect 1276 47 1333 69
rect 1387 209 1444 221
rect 1387 175 1399 209
rect 1433 175 1444 209
rect 1387 99 1444 175
rect 1387 65 1399 99
rect 1433 65 1444 99
rect 1387 53 1444 65
rect 1474 53 1516 221
rect 1546 209 1603 221
rect 1546 175 1557 209
rect 1591 175 1603 209
rect 1546 103 1603 175
rect 1546 69 1557 103
rect 1591 69 1603 103
rect 1546 53 1603 69
<< pdiff >>
rect 643 619 701 627
rect 27 586 84 598
rect 27 552 39 586
rect 73 552 84 586
rect 27 516 84 552
rect 27 482 39 516
rect 73 482 84 516
rect 27 470 84 482
rect 114 470 162 598
rect 192 586 248 598
rect 192 552 203 586
rect 237 552 248 586
rect 192 516 248 552
rect 192 482 203 516
rect 237 482 248 516
rect 192 470 248 482
rect 278 470 320 598
rect 350 586 407 598
rect 350 552 361 586
rect 395 552 407 586
rect 350 516 407 552
rect 350 482 361 516
rect 395 482 407 516
rect 463 567 520 619
rect 463 533 475 567
rect 509 533 520 567
rect 463 491 520 533
rect 550 491 598 619
rect 628 615 716 619
rect 628 581 655 615
rect 689 581 716 615
rect 628 491 716 581
rect 746 491 794 619
rect 824 603 903 619
rect 824 569 835 603
rect 869 569 903 603
rect 824 535 903 569
rect 933 535 1027 619
rect 1057 607 1174 619
rect 1057 573 1129 607
rect 1163 573 1174 607
rect 1057 535 1174 573
rect 824 491 881 535
rect 350 470 407 482
rect 1117 510 1174 535
rect 1117 476 1129 510
rect 1163 476 1174 510
rect 1117 413 1174 476
rect 1117 379 1129 413
rect 1163 379 1174 413
rect 1117 367 1174 379
rect 1204 367 1246 619
rect 1276 597 1333 619
rect 1276 563 1287 597
rect 1321 563 1333 597
rect 1276 505 1333 563
rect 1276 471 1287 505
rect 1321 471 1333 505
rect 1276 413 1333 471
rect 1276 379 1287 413
rect 1321 379 1333 413
rect 1276 367 1333 379
rect 1387 607 1444 619
rect 1387 573 1399 607
rect 1433 573 1444 607
rect 1387 510 1444 573
rect 1387 476 1399 510
rect 1433 476 1444 510
rect 1387 413 1444 476
rect 1387 379 1399 413
rect 1433 379 1444 413
rect 1387 367 1444 379
rect 1474 367 1516 619
rect 1546 597 1603 619
rect 1546 563 1557 597
rect 1591 563 1603 597
rect 1546 505 1603 563
rect 1546 471 1557 505
rect 1591 471 1603 505
rect 1546 413 1603 471
rect 1546 379 1557 413
rect 1591 379 1603 413
rect 1546 367 1603 379
<< ndiffc >>
rect 39 127 73 161
rect 197 127 231 161
rect 361 127 395 161
rect 509 77 543 111
rect 673 59 707 93
rect 907 77 941 111
rect 1072 72 1106 106
rect 1287 169 1321 203
rect 1287 69 1321 103
rect 1399 175 1433 209
rect 1399 65 1433 99
rect 1557 175 1591 209
rect 1557 69 1591 103
<< pdiffc >>
rect 39 552 73 586
rect 39 482 73 516
rect 203 552 237 586
rect 203 482 237 516
rect 361 552 395 586
rect 361 482 395 516
rect 475 533 509 567
rect 655 581 689 615
rect 835 569 869 603
rect 1129 573 1163 607
rect 1129 476 1163 510
rect 1129 379 1163 413
rect 1287 563 1321 597
rect 1287 471 1321 505
rect 1287 379 1321 413
rect 1399 573 1433 607
rect 1399 476 1433 510
rect 1399 379 1433 413
rect 1557 563 1591 597
rect 1557 471 1591 505
rect 1557 379 1591 413
<< poly >>
rect 84 598 114 624
rect 162 598 192 624
rect 248 598 278 624
rect 320 598 350 624
rect 520 619 550 645
rect 598 619 628 645
rect 716 619 746 645
rect 794 619 824 645
rect 903 619 933 645
rect 1027 619 1057 645
rect 1174 619 1204 645
rect 1246 619 1276 645
rect 1444 619 1474 645
rect 1516 619 1546 645
rect 903 503 933 535
rect 84 430 114 470
rect 162 430 192 470
rect 84 414 192 430
rect 84 380 131 414
rect 165 380 192 414
rect 84 346 192 380
rect 84 312 131 346
rect 165 312 192 346
rect 84 296 192 312
rect 248 430 278 470
rect 320 430 350 470
rect 248 414 350 430
rect 248 380 270 414
rect 304 380 350 414
rect 248 364 350 380
rect 84 186 114 296
rect 156 186 186 296
rect 248 186 278 364
rect 320 186 350 364
rect 520 315 550 491
rect 598 351 628 491
rect 716 459 746 491
rect 680 443 746 459
rect 680 409 696 443
rect 730 409 746 443
rect 680 393 746 409
rect 794 395 824 491
rect 903 487 979 503
rect 903 453 929 487
rect 963 453 979 487
rect 903 437 979 453
rect 1027 437 1057 535
rect 1027 407 1060 437
rect 596 335 662 351
rect 596 315 612 335
rect 520 301 612 315
rect 646 301 662 335
rect 520 285 662 301
rect 520 237 550 285
rect 520 207 584 237
rect 554 131 584 207
rect 632 131 662 285
rect 710 281 740 393
rect 788 379 854 395
rect 788 345 804 379
rect 838 359 854 379
rect 838 345 982 359
rect 788 329 982 345
rect 710 265 790 281
rect 710 231 726 265
rect 760 231 790 265
rect 710 215 790 231
rect 760 131 790 215
rect 838 221 904 237
rect 838 187 854 221
rect 888 187 904 221
rect 838 171 904 187
rect 838 131 868 171
rect 952 131 982 329
rect 1030 251 1060 407
rect 1174 321 1204 367
rect 1246 321 1276 367
rect 1444 327 1474 367
rect 1516 327 1546 367
rect 1168 305 1276 321
rect 1168 271 1184 305
rect 1218 271 1276 305
rect 1168 255 1276 271
rect 1439 311 1546 327
rect 1439 277 1455 311
rect 1489 277 1546 311
rect 1439 261 1546 277
rect 1030 235 1096 251
rect 1030 201 1046 235
rect 1080 201 1096 235
rect 1168 215 1198 255
rect 1246 215 1276 255
rect 1444 221 1474 261
rect 1516 221 1546 261
rect 1030 185 1096 201
rect 1030 131 1060 185
rect 84 76 114 102
rect 156 76 186 102
rect 248 76 278 102
rect 320 76 350 102
rect 554 21 584 47
rect 632 21 662 47
rect 760 21 790 47
rect 838 21 868 47
rect 952 21 982 47
rect 1030 21 1060 47
rect 1168 21 1198 47
rect 1246 21 1276 47
rect 1444 27 1474 53
rect 1516 27 1546 53
<< polycont >>
rect 131 380 165 414
rect 131 312 165 346
rect 270 380 304 414
rect 696 409 730 443
rect 929 453 963 487
rect 612 301 646 335
rect 804 345 838 379
rect 726 231 760 265
rect 854 187 888 221
rect 1184 271 1218 305
rect 1455 277 1489 311
rect 1046 201 1080 235
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 586 73 602
rect 23 552 39 586
rect 23 516 73 552
rect 23 482 39 516
rect 23 260 73 482
rect 187 586 253 649
rect 639 615 705 649
rect 187 552 203 586
rect 237 552 253 586
rect 187 516 253 552
rect 187 482 203 516
rect 237 482 253 516
rect 187 466 253 482
rect 345 586 411 602
rect 345 552 361 586
rect 395 552 411 586
rect 345 516 411 552
rect 345 482 361 516
rect 395 482 411 516
rect 459 567 525 613
rect 459 533 475 567
rect 509 533 525 567
rect 639 581 655 615
rect 689 581 705 615
rect 1113 607 1179 649
rect 639 565 705 581
rect 819 603 1049 607
rect 819 569 835 603
rect 869 569 1049 603
rect 819 565 1049 569
rect 459 529 525 533
rect 459 495 979 529
rect 459 487 525 495
rect 890 487 979 495
rect 345 466 411 482
rect 115 414 181 430
rect 115 380 131 414
rect 165 380 181 414
rect 115 346 181 380
rect 217 414 320 430
rect 217 380 270 414
rect 304 380 320 414
rect 377 427 411 466
rect 680 443 746 459
rect 680 427 696 443
rect 377 409 696 427
rect 730 409 746 443
rect 377 393 746 409
rect 890 453 929 487
rect 963 453 979 487
rect 890 437 979 453
rect 217 364 320 380
rect 788 379 854 395
rect 788 351 804 379
rect 115 312 131 346
rect 165 312 181 346
rect 596 345 804 351
rect 838 345 854 379
rect 596 335 854 345
rect 596 319 612 335
rect 115 296 181 312
rect 275 301 612 319
rect 646 317 854 335
rect 646 301 662 317
rect 275 285 662 301
rect 275 260 309 285
rect 23 226 309 260
rect 710 265 776 281
rect 710 249 726 265
rect 345 231 726 249
rect 760 231 776 265
rect 890 237 924 437
rect 1015 321 1049 565
rect 1113 573 1129 607
rect 1163 573 1179 607
rect 1113 510 1179 573
rect 1113 476 1129 510
rect 1163 476 1179 510
rect 1113 413 1179 476
rect 1113 379 1129 413
rect 1163 379 1179 413
rect 1113 363 1179 379
rect 1271 597 1337 613
rect 1271 563 1287 597
rect 1321 563 1337 597
rect 1271 505 1337 563
rect 1271 471 1287 505
rect 1321 471 1337 505
rect 1271 413 1337 471
rect 1271 379 1287 413
rect 1321 379 1337 413
rect 1271 327 1337 379
rect 1383 607 1449 649
rect 1383 573 1399 607
rect 1433 573 1449 607
rect 1383 510 1449 573
rect 1383 476 1399 510
rect 1433 476 1449 510
rect 1383 413 1449 476
rect 1383 379 1399 413
rect 1433 379 1449 413
rect 1383 363 1449 379
rect 1541 597 1607 613
rect 1541 563 1557 597
rect 1591 563 1607 597
rect 1541 505 1607 563
rect 1541 471 1557 505
rect 1591 471 1607 505
rect 1541 413 1607 471
rect 1541 379 1557 413
rect 1591 379 1607 413
rect 23 161 89 226
rect 345 215 776 231
rect 821 221 924 237
rect 23 127 39 161
rect 73 127 89 161
rect 23 98 89 127
rect 181 161 247 190
rect 181 127 197 161
rect 231 127 247 161
rect 181 17 247 127
rect 345 161 411 215
rect 821 187 854 221
rect 888 187 924 221
rect 821 179 924 187
rect 345 127 361 161
rect 395 127 411 161
rect 345 98 411 127
rect 493 171 924 179
rect 960 305 1234 321
rect 960 287 1184 305
rect 493 145 855 171
rect 493 111 559 145
rect 960 135 994 287
rect 1168 271 1184 287
rect 1218 271 1234 305
rect 1168 255 1234 271
rect 1271 311 1505 327
rect 1271 277 1455 311
rect 1489 277 1505 311
rect 1271 261 1505 277
rect 1030 235 1096 251
rect 1030 201 1046 235
rect 1080 219 1096 235
rect 1271 219 1337 261
rect 1080 203 1337 219
rect 1080 201 1287 203
rect 1030 185 1287 201
rect 1271 169 1287 185
rect 1321 169 1337 203
rect 493 77 509 111
rect 543 77 559 111
rect 891 111 994 135
rect 493 53 559 77
rect 657 93 723 109
rect 657 59 673 93
rect 707 59 723 93
rect 657 17 723 59
rect 891 77 907 111
rect 941 101 994 111
rect 1056 106 1122 135
rect 941 77 957 101
rect 891 53 957 77
rect 1056 72 1072 106
rect 1106 72 1122 106
rect 1056 17 1122 72
rect 1271 103 1337 169
rect 1271 69 1287 103
rect 1321 69 1337 103
rect 1271 53 1337 69
rect 1383 209 1449 225
rect 1383 175 1399 209
rect 1433 175 1449 209
rect 1383 99 1449 175
rect 1383 65 1399 99
rect 1433 65 1449 99
rect 1383 17 1449 65
rect 1541 209 1607 379
rect 1541 175 1557 209
rect 1591 175 1607 209
rect 1541 103 1607 175
rect 1541 69 1557 103
rect 1591 69 1607 103
rect 1541 53 1607 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlxtp_lp
flabel comment s 722 344 722 344 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 27054
string GDS_START 15672
<< end >>
