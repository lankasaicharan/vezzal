magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 23 49 1097 241
rect 0 0 1152 49
<< scnmos >>
rect 102 47 132 215
rect 188 47 218 215
rect 354 47 384 215
rect 440 47 470 215
rect 526 47 556 215
rect 612 47 642 215
rect 730 47 760 215
rect 816 47 846 215
rect 902 47 932 215
rect 988 47 1018 215
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 356 367 386 619
rect 442 367 472 619
rect 528 367 558 619
rect 614 367 644 619
rect 708 367 738 619
rect 816 367 846 619
rect 902 367 932 619
rect 988 367 1018 619
<< ndiff >>
rect 49 192 102 215
rect 49 158 57 192
rect 91 158 102 192
rect 49 93 102 158
rect 49 59 57 93
rect 91 59 102 93
rect 49 47 102 59
rect 132 183 188 215
rect 132 149 143 183
rect 177 149 188 183
rect 132 115 188 149
rect 132 81 143 115
rect 177 81 188 115
rect 132 47 188 81
rect 218 115 354 215
rect 218 81 229 115
rect 263 81 305 115
rect 339 81 354 115
rect 218 47 354 81
rect 384 107 440 215
rect 384 73 395 107
rect 429 73 440 107
rect 384 47 440 73
rect 470 195 526 215
rect 470 161 481 195
rect 515 161 526 195
rect 470 47 526 161
rect 556 107 612 215
rect 556 73 567 107
rect 601 73 612 107
rect 556 47 612 73
rect 642 113 730 215
rect 642 79 668 113
rect 702 79 730 113
rect 642 47 730 79
rect 760 93 816 215
rect 760 59 771 93
rect 805 59 816 93
rect 760 47 816 59
rect 846 183 902 215
rect 846 149 857 183
rect 891 149 902 183
rect 846 47 902 149
rect 932 203 988 215
rect 932 169 943 203
rect 977 169 988 203
rect 932 93 988 169
rect 932 59 943 93
rect 977 59 988 93
rect 932 47 988 59
rect 1018 192 1071 215
rect 1018 158 1029 192
rect 1063 158 1071 192
rect 1018 93 1071 158
rect 1018 59 1029 93
rect 1063 59 1071 93
rect 1018 47 1071 59
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 511 80 565
rect 27 477 35 511
rect 69 477 80 511
rect 27 435 80 477
rect 27 401 35 435
rect 69 401 80 435
rect 27 367 80 401
rect 110 543 166 619
rect 110 509 121 543
rect 155 509 166 543
rect 110 422 166 509
rect 110 388 121 422
rect 155 388 166 422
rect 110 367 166 388
rect 196 599 249 619
rect 196 565 207 599
rect 241 565 249 599
rect 196 515 249 565
rect 196 481 207 515
rect 241 481 249 515
rect 196 441 249 481
rect 196 407 207 441
rect 241 407 249 441
rect 196 367 249 407
rect 303 599 356 619
rect 303 565 311 599
rect 345 565 356 599
rect 303 509 356 565
rect 303 475 311 509
rect 345 475 356 509
rect 303 367 356 475
rect 386 543 442 619
rect 386 509 397 543
rect 431 509 442 543
rect 386 425 442 509
rect 386 391 397 425
rect 431 391 442 425
rect 386 367 442 391
rect 472 599 528 619
rect 472 565 483 599
rect 517 565 528 599
rect 472 509 528 565
rect 472 475 483 509
rect 517 475 528 509
rect 472 367 528 475
rect 558 543 614 619
rect 558 509 569 543
rect 603 509 614 543
rect 558 425 614 509
rect 558 391 569 425
rect 603 391 614 425
rect 558 367 614 391
rect 644 599 708 619
rect 644 565 655 599
rect 689 565 708 599
rect 644 513 708 565
rect 644 479 655 513
rect 689 479 708 513
rect 644 441 708 479
rect 644 407 655 441
rect 689 407 708 441
rect 644 367 708 407
rect 738 607 816 619
rect 738 573 760 607
rect 794 573 816 607
rect 738 497 816 573
rect 738 463 760 497
rect 794 463 816 497
rect 738 367 816 463
rect 846 599 902 619
rect 846 565 857 599
rect 891 565 902 599
rect 846 513 902 565
rect 846 479 857 513
rect 891 479 902 513
rect 846 425 902 479
rect 846 391 857 425
rect 891 391 902 425
rect 846 367 902 391
rect 932 607 988 619
rect 932 573 943 607
rect 977 573 988 607
rect 932 497 988 573
rect 932 463 943 497
rect 977 463 988 497
rect 932 367 988 463
rect 1018 599 1071 619
rect 1018 565 1029 599
rect 1063 565 1071 599
rect 1018 513 1071 565
rect 1018 479 1029 513
rect 1063 479 1071 513
rect 1018 425 1071 479
rect 1018 391 1029 425
rect 1063 391 1071 425
rect 1018 367 1071 391
<< ndiffc >>
rect 57 158 91 192
rect 57 59 91 93
rect 143 149 177 183
rect 143 81 177 115
rect 229 81 263 115
rect 305 81 339 115
rect 395 73 429 107
rect 481 161 515 195
rect 567 73 601 107
rect 668 79 702 113
rect 771 59 805 93
rect 857 149 891 183
rect 943 169 977 203
rect 943 59 977 93
rect 1029 158 1063 192
rect 1029 59 1063 93
<< pdiffc >>
rect 35 565 69 599
rect 35 477 69 511
rect 35 401 69 435
rect 121 509 155 543
rect 121 388 155 422
rect 207 565 241 599
rect 207 481 241 515
rect 207 407 241 441
rect 311 565 345 599
rect 311 475 345 509
rect 397 509 431 543
rect 397 391 431 425
rect 483 565 517 599
rect 483 475 517 509
rect 569 509 603 543
rect 569 391 603 425
rect 655 565 689 599
rect 655 479 689 513
rect 655 407 689 441
rect 760 573 794 607
rect 760 463 794 497
rect 857 565 891 599
rect 857 479 891 513
rect 857 391 891 425
rect 943 573 977 607
rect 943 463 977 497
rect 1029 565 1063 599
rect 1029 479 1063 513
rect 1029 391 1063 425
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 356 619 386 645
rect 442 619 472 645
rect 528 619 558 645
rect 614 619 644 645
rect 708 619 738 645
rect 816 619 846 645
rect 902 619 932 645
rect 988 619 1018 645
rect 80 308 110 367
rect 166 308 196 367
rect 356 335 386 367
rect 41 292 196 308
rect 41 258 57 292
rect 91 272 196 292
rect 332 319 398 335
rect 332 285 348 319
rect 382 285 398 319
rect 442 303 472 367
rect 528 303 558 367
rect 614 325 644 367
rect 708 335 738 367
rect 91 258 218 272
rect 332 269 398 285
rect 440 287 558 303
rect 41 242 218 258
rect 102 215 132 242
rect 188 215 218 242
rect 354 215 384 269
rect 440 253 501 287
rect 535 273 558 287
rect 600 309 666 325
rect 600 275 616 309
rect 650 275 666 309
rect 535 253 556 273
rect 600 259 666 275
rect 708 319 774 335
rect 708 285 724 319
rect 758 285 774 319
rect 708 269 774 285
rect 816 303 846 367
rect 902 303 932 367
rect 816 287 932 303
rect 440 237 556 253
rect 440 215 470 237
rect 526 215 556 237
rect 612 215 642 259
rect 730 215 760 269
rect 816 253 832 287
rect 866 253 932 287
rect 816 237 932 253
rect 816 215 846 237
rect 902 215 932 237
rect 988 308 1018 367
rect 988 292 1131 308
rect 988 258 1081 292
rect 1115 258 1131 292
rect 988 242 1131 258
rect 988 215 1018 242
rect 102 21 132 47
rect 188 21 218 47
rect 354 21 384 47
rect 440 21 470 47
rect 526 21 556 47
rect 612 21 642 47
rect 730 21 760 47
rect 816 21 846 47
rect 902 21 932 47
rect 988 21 1018 47
<< polycont >>
rect 57 258 91 292
rect 348 285 382 319
rect 501 253 535 287
rect 616 275 650 309
rect 724 285 758 319
rect 832 253 866 287
rect 1081 258 1115 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 19 599 257 615
rect 19 565 35 599
rect 69 581 207 599
rect 69 565 71 581
rect 19 511 71 565
rect 205 565 207 581
rect 241 565 257 599
rect 19 477 35 511
rect 69 477 71 511
rect 19 435 71 477
rect 19 401 35 435
rect 69 401 71 435
rect 19 385 71 401
rect 105 543 171 547
rect 105 509 121 543
rect 155 509 171 543
rect 105 422 171 509
rect 105 388 121 422
rect 155 388 171 422
rect 205 515 257 565
rect 205 481 207 515
rect 241 481 257 515
rect 205 441 257 481
rect 295 599 710 615
rect 295 565 311 599
rect 345 581 483 599
rect 345 565 347 581
rect 295 509 347 565
rect 481 565 483 581
rect 517 581 655 599
rect 517 565 519 581
rect 295 475 311 509
rect 345 475 347 509
rect 295 459 347 475
rect 381 543 447 547
rect 381 509 397 543
rect 431 509 447 543
rect 205 407 207 441
rect 241 425 257 441
rect 381 425 447 509
rect 481 509 519 565
rect 653 565 655 581
rect 689 565 710 599
rect 481 475 483 509
rect 517 475 519 509
rect 481 459 519 475
rect 553 543 619 547
rect 553 509 569 543
rect 603 509 619 543
rect 553 425 619 509
rect 241 407 397 425
rect 205 391 397 407
rect 431 391 569 425
rect 603 391 619 425
rect 653 513 710 565
rect 653 479 655 513
rect 689 479 710 513
rect 653 441 710 479
rect 744 607 810 649
rect 744 573 760 607
rect 794 573 810 607
rect 744 497 810 573
rect 744 463 760 497
rect 794 463 810 497
rect 744 459 810 463
rect 844 599 891 615
rect 844 565 857 599
rect 844 513 891 565
rect 844 479 857 513
rect 653 407 655 441
rect 689 425 710 441
rect 844 425 891 479
rect 927 607 993 649
rect 927 573 943 607
rect 977 573 993 607
rect 927 497 993 573
rect 927 463 943 497
rect 977 463 993 497
rect 927 459 993 463
rect 1029 599 1079 615
rect 1063 565 1079 599
rect 1029 513 1079 565
rect 1063 479 1079 513
rect 1029 425 1079 479
rect 689 407 857 425
rect 653 391 857 407
rect 891 391 1029 425
rect 1063 391 1079 425
rect 105 384 171 388
rect 17 292 93 350
rect 17 258 57 292
rect 91 258 93 292
rect 17 242 93 258
rect 127 208 171 384
rect 205 323 666 357
rect 205 319 451 323
rect 205 285 348 319
rect 382 285 451 319
rect 600 309 666 323
rect 485 287 563 289
rect 485 253 501 287
rect 535 253 563 287
rect 600 275 616 309
rect 650 275 666 309
rect 708 323 1135 357
rect 708 319 758 323
rect 708 285 724 319
rect 1067 292 1135 323
rect 708 269 758 285
rect 792 287 1033 289
rect 485 242 563 253
rect 792 253 832 287
rect 866 253 1033 287
rect 792 242 1033 253
rect 1067 258 1081 292
rect 1115 258 1135 292
rect 1067 242 1135 258
rect 41 192 93 208
rect 41 158 57 192
rect 91 158 93 192
rect 41 93 93 158
rect 41 59 57 93
rect 91 59 93 93
rect 41 17 93 59
rect 127 195 893 208
rect 127 183 481 195
rect 127 149 143 183
rect 177 161 481 183
rect 515 183 893 195
rect 515 161 857 183
rect 177 157 857 161
rect 177 149 179 157
rect 127 115 179 149
rect 841 149 857 157
rect 891 149 893 183
rect 841 133 893 149
rect 927 203 993 208
rect 927 169 943 203
rect 977 169 993 203
rect 127 81 143 115
rect 177 81 179 115
rect 127 51 179 81
rect 213 115 355 123
rect 213 81 229 115
rect 263 81 305 115
rect 339 81 355 115
rect 213 17 355 81
rect 391 107 617 123
rect 391 73 395 107
rect 429 73 567 107
rect 601 73 617 107
rect 391 57 617 73
rect 652 113 718 123
rect 652 79 668 113
rect 702 79 718 113
rect 927 97 993 169
rect 652 17 718 79
rect 755 93 993 97
rect 755 59 771 93
rect 805 59 943 93
rect 977 59 993 93
rect 755 51 993 59
rect 1027 192 1079 208
rect 1027 158 1029 192
rect 1063 158 1079 192
rect 1027 93 1079 158
rect 1027 59 1029 93
rect 1063 59 1079 93
rect 1027 17 1079 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a221oi_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3946100
string GDS_START 3935320
<< end >>
