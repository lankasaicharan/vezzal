magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 2 49 1144 241
rect 0 0 1152 49
<< scnmos >>
rect 81 47 111 215
rect 167 47 197 215
rect 253 47 283 215
rect 339 47 369 215
rect 425 47 455 215
rect 511 47 541 215
rect 597 47 627 215
rect 683 47 713 215
rect 777 47 807 215
rect 863 47 893 215
rect 949 47 979 215
rect 1035 47 1065 215
<< scpmoshvt >>
rect 81 367 111 619
rect 167 367 197 619
rect 253 367 283 619
rect 339 367 369 619
rect 425 367 455 619
rect 511 367 541 619
rect 597 367 627 619
rect 691 367 721 619
rect 777 367 807 619
rect 863 367 893 619
rect 949 367 979 619
rect 1035 367 1065 619
<< ndiff >>
rect 28 203 81 215
rect 28 169 36 203
rect 70 169 81 203
rect 28 93 81 169
rect 28 59 36 93
rect 70 59 81 93
rect 28 47 81 59
rect 111 203 167 215
rect 111 169 122 203
rect 156 169 167 203
rect 111 101 167 169
rect 111 67 122 101
rect 156 67 167 101
rect 111 47 167 67
rect 197 173 253 215
rect 197 139 208 173
rect 242 139 253 173
rect 197 93 253 139
rect 197 59 208 93
rect 242 59 253 93
rect 197 47 253 59
rect 283 203 339 215
rect 283 169 294 203
rect 328 169 339 203
rect 283 101 339 169
rect 283 67 294 101
rect 328 67 339 101
rect 283 47 339 67
rect 369 202 425 215
rect 369 168 380 202
rect 414 168 425 202
rect 369 47 425 168
rect 455 112 511 215
rect 455 78 466 112
rect 500 78 511 112
rect 455 47 511 78
rect 541 202 597 215
rect 541 168 552 202
rect 586 168 597 202
rect 541 47 597 168
rect 627 112 683 215
rect 627 78 638 112
rect 672 78 683 112
rect 627 47 683 78
rect 713 122 777 215
rect 713 88 728 122
rect 762 88 777 122
rect 713 47 777 88
rect 807 203 863 215
rect 807 169 818 203
rect 852 169 863 203
rect 807 101 863 169
rect 807 67 818 101
rect 852 67 863 101
rect 807 47 863 67
rect 893 183 949 215
rect 893 149 904 183
rect 938 149 949 183
rect 893 93 949 149
rect 893 59 904 93
rect 938 59 949 93
rect 893 47 949 59
rect 979 203 1035 215
rect 979 169 990 203
rect 1024 169 1035 203
rect 979 101 1035 169
rect 979 67 990 101
rect 1024 67 1035 101
rect 979 47 1035 67
rect 1065 183 1118 215
rect 1065 149 1076 183
rect 1110 149 1118 183
rect 1065 93 1118 149
rect 1065 59 1076 93
rect 1110 59 1118 93
rect 1065 47 1118 59
<< pdiff >>
rect 28 599 81 619
rect 28 565 36 599
rect 70 565 81 599
rect 28 523 81 565
rect 28 489 36 523
rect 70 489 81 523
rect 28 441 81 489
rect 28 407 36 441
rect 70 407 81 441
rect 28 367 81 407
rect 111 607 167 619
rect 111 573 122 607
rect 156 573 167 607
rect 111 499 167 573
rect 111 465 122 499
rect 156 465 167 499
rect 111 367 167 465
rect 197 599 253 619
rect 197 565 208 599
rect 242 565 253 599
rect 197 523 253 565
rect 197 489 208 523
rect 242 489 253 523
rect 197 441 253 489
rect 197 407 208 441
rect 242 407 253 441
rect 197 367 253 407
rect 283 607 339 619
rect 283 573 294 607
rect 328 573 339 607
rect 283 499 339 573
rect 283 465 294 499
rect 328 465 339 499
rect 283 367 339 465
rect 369 599 425 619
rect 369 565 380 599
rect 414 565 425 599
rect 369 523 425 565
rect 369 489 380 523
rect 414 489 425 523
rect 369 441 425 489
rect 369 407 380 441
rect 414 407 425 441
rect 369 367 425 407
rect 455 607 511 619
rect 455 573 466 607
rect 500 573 511 607
rect 455 499 511 573
rect 455 465 466 499
rect 500 465 511 499
rect 455 367 511 465
rect 541 599 597 619
rect 541 565 552 599
rect 586 565 597 599
rect 541 523 597 565
rect 541 489 552 523
rect 586 489 597 523
rect 541 441 597 489
rect 541 407 552 441
rect 586 407 597 441
rect 541 367 597 407
rect 627 607 691 619
rect 627 573 638 607
rect 672 573 691 607
rect 627 499 691 573
rect 627 465 638 499
rect 672 465 691 499
rect 627 367 691 465
rect 721 599 777 619
rect 721 565 732 599
rect 766 565 777 599
rect 721 523 777 565
rect 721 489 732 523
rect 766 489 777 523
rect 721 441 777 489
rect 721 407 732 441
rect 766 407 777 441
rect 721 367 777 407
rect 807 531 863 619
rect 807 497 818 531
rect 852 497 863 531
rect 807 436 863 497
rect 807 402 818 436
rect 852 402 863 436
rect 807 367 863 402
rect 893 599 949 619
rect 893 565 904 599
rect 938 565 949 599
rect 893 511 949 565
rect 893 477 904 511
rect 938 477 949 511
rect 893 367 949 477
rect 979 531 1035 619
rect 979 497 990 531
rect 1024 497 1035 531
rect 979 436 1035 497
rect 979 402 990 436
rect 1024 402 1035 436
rect 979 367 1035 402
rect 1065 599 1118 619
rect 1065 565 1076 599
rect 1110 565 1118 599
rect 1065 511 1118 565
rect 1065 477 1076 511
rect 1110 477 1118 511
rect 1065 367 1118 477
<< ndiffc >>
rect 36 169 70 203
rect 36 59 70 93
rect 122 169 156 203
rect 122 67 156 101
rect 208 139 242 173
rect 208 59 242 93
rect 294 169 328 203
rect 294 67 328 101
rect 380 168 414 202
rect 466 78 500 112
rect 552 168 586 202
rect 638 78 672 112
rect 728 88 762 122
rect 818 169 852 203
rect 818 67 852 101
rect 904 149 938 183
rect 904 59 938 93
rect 990 169 1024 203
rect 990 67 1024 101
rect 1076 149 1110 183
rect 1076 59 1110 93
<< pdiffc >>
rect 36 565 70 599
rect 36 489 70 523
rect 36 407 70 441
rect 122 573 156 607
rect 122 465 156 499
rect 208 565 242 599
rect 208 489 242 523
rect 208 407 242 441
rect 294 573 328 607
rect 294 465 328 499
rect 380 565 414 599
rect 380 489 414 523
rect 380 407 414 441
rect 466 573 500 607
rect 466 465 500 499
rect 552 565 586 599
rect 552 489 586 523
rect 552 407 586 441
rect 638 573 672 607
rect 638 465 672 499
rect 732 565 766 599
rect 732 489 766 523
rect 732 407 766 441
rect 818 497 852 531
rect 818 402 852 436
rect 904 565 938 599
rect 904 477 938 511
rect 990 497 1024 531
rect 990 402 1024 436
rect 1076 565 1110 599
rect 1076 477 1110 511
<< poly >>
rect 81 619 111 645
rect 167 619 197 645
rect 253 619 283 645
rect 339 619 369 645
rect 425 619 455 645
rect 511 619 541 645
rect 597 619 627 645
rect 691 619 721 645
rect 777 619 807 645
rect 863 619 893 645
rect 949 619 979 645
rect 1035 619 1065 645
rect 81 325 111 367
rect 167 325 197 367
rect 253 325 283 367
rect 21 309 291 325
rect 21 275 37 309
rect 71 275 105 309
rect 139 275 173 309
rect 207 275 241 309
rect 275 275 291 309
rect 21 259 291 275
rect 339 303 369 367
rect 425 303 455 367
rect 511 303 541 367
rect 597 303 627 367
rect 691 335 721 367
rect 777 335 807 367
rect 863 335 893 367
rect 949 335 979 367
rect 1035 335 1065 367
rect 339 287 627 303
rect 81 215 111 259
rect 167 215 197 259
rect 253 215 283 259
rect 339 253 411 287
rect 445 253 479 287
rect 513 253 547 287
rect 581 253 627 287
rect 669 319 735 335
rect 669 285 685 319
rect 719 285 735 319
rect 669 269 735 285
rect 777 319 1065 335
rect 777 285 793 319
rect 827 285 861 319
rect 895 285 929 319
rect 963 285 997 319
rect 1031 285 1065 319
rect 777 269 1065 285
rect 339 237 627 253
rect 339 215 369 237
rect 425 215 455 237
rect 511 215 541 237
rect 597 215 627 237
rect 683 215 713 269
rect 777 215 807 269
rect 863 215 893 269
rect 949 215 979 269
rect 1035 215 1065 269
rect 81 21 111 47
rect 167 21 197 47
rect 253 21 283 47
rect 339 21 369 47
rect 425 21 455 47
rect 511 21 541 47
rect 597 21 627 47
rect 683 21 713 47
rect 777 21 807 47
rect 863 21 893 47
rect 949 21 979 47
rect 1035 21 1065 47
<< polycont >>
rect 37 275 71 309
rect 105 275 139 309
rect 173 275 207 309
rect 241 275 275 309
rect 411 253 445 287
rect 479 253 513 287
rect 547 253 581 287
rect 685 285 719 319
rect 793 285 827 319
rect 861 285 895 319
rect 929 285 963 319
rect 997 285 1031 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 20 599 72 615
rect 20 565 36 599
rect 70 565 72 599
rect 20 523 72 565
rect 20 489 36 523
rect 70 489 72 523
rect 20 441 72 489
rect 106 607 172 649
rect 106 573 122 607
rect 156 573 172 607
rect 106 499 172 573
rect 106 465 122 499
rect 156 465 172 499
rect 106 459 172 465
rect 206 599 244 615
rect 206 565 208 599
rect 242 565 244 599
rect 206 523 244 565
rect 206 489 208 523
rect 242 489 244 523
rect 20 407 36 441
rect 70 425 72 441
rect 206 441 244 489
rect 278 607 344 649
rect 278 573 294 607
rect 328 573 344 607
rect 278 499 344 573
rect 278 465 294 499
rect 328 465 344 499
rect 278 459 344 465
rect 380 599 416 615
rect 414 565 416 599
rect 380 523 416 565
rect 414 489 416 523
rect 206 425 208 441
rect 70 407 208 425
rect 242 425 244 441
rect 380 441 416 489
rect 450 607 516 649
rect 450 573 466 607
rect 500 573 516 607
rect 450 499 516 573
rect 450 465 466 499
rect 500 465 516 499
rect 450 459 516 465
rect 550 599 588 615
rect 550 565 552 599
rect 586 565 588 599
rect 550 523 588 565
rect 550 489 552 523
rect 586 489 588 523
rect 242 407 380 425
rect 414 425 416 441
rect 550 441 588 489
rect 622 607 688 649
rect 622 573 638 607
rect 672 573 688 607
rect 622 499 688 573
rect 622 465 638 499
rect 672 465 688 499
rect 622 459 688 465
rect 722 599 1126 615
rect 722 565 732 599
rect 766 581 904 599
rect 766 565 777 581
rect 722 523 777 565
rect 893 565 904 581
rect 938 581 1076 599
rect 938 565 948 581
rect 722 489 732 523
rect 766 489 777 523
rect 550 425 552 441
rect 414 407 552 425
rect 586 425 588 441
rect 722 441 777 489
rect 722 425 732 441
rect 586 407 732 425
rect 766 407 777 441
rect 20 391 777 407
rect 811 531 859 547
rect 811 497 818 531
rect 852 497 859 531
rect 811 436 859 497
rect 893 511 948 565
rect 1065 565 1076 581
rect 1110 565 1126 599
rect 893 477 904 511
rect 938 477 948 511
rect 893 454 948 477
rect 982 531 1031 547
rect 982 497 990 531
rect 1024 497 1031 531
rect 811 402 818 436
rect 852 420 859 436
rect 982 436 1031 497
rect 1065 511 1126 565
rect 1065 477 1076 511
rect 1110 477 1126 511
rect 1065 454 1126 477
rect 982 420 990 436
rect 852 402 990 420
rect 1024 420 1031 436
rect 1024 402 1117 420
rect 811 386 1117 402
rect 21 323 735 357
rect 21 309 353 323
rect 21 275 37 309
rect 71 275 105 309
rect 139 275 173 309
rect 207 275 241 309
rect 275 275 353 309
rect 680 319 735 323
rect 395 253 411 287
rect 445 253 479 287
rect 513 253 547 287
rect 581 253 646 287
rect 680 285 685 319
rect 719 285 735 319
rect 777 319 1047 352
rect 777 285 793 319
rect 827 285 861 319
rect 895 285 929 319
rect 963 285 997 319
rect 1031 285 1047 319
rect 680 269 735 285
rect 20 203 78 219
rect 20 169 36 203
rect 70 169 78 203
rect 20 93 78 169
rect 20 59 36 93
rect 70 59 78 93
rect 20 17 78 59
rect 112 207 330 241
rect 395 240 646 253
rect 1083 251 1117 386
rect 112 203 158 207
rect 112 169 122 203
rect 156 169 158 203
rect 292 203 330 207
rect 814 217 1117 251
rect 814 206 852 217
rect 112 101 158 169
rect 112 67 122 101
rect 156 67 158 101
rect 112 51 158 67
rect 192 139 208 173
rect 242 139 258 173
rect 192 93 258 139
rect 192 59 208 93
rect 242 59 258 93
rect 192 17 258 59
rect 292 169 294 203
rect 328 169 330 203
rect 292 128 330 169
rect 364 203 852 206
rect 364 202 818 203
rect 364 168 380 202
rect 414 168 552 202
rect 586 169 818 202
rect 988 203 1026 217
rect 586 168 852 169
rect 364 164 852 168
rect 292 112 676 128
rect 292 101 466 112
rect 292 67 294 101
rect 328 78 466 101
rect 500 78 638 112
rect 672 78 676 112
rect 328 67 676 78
rect 292 51 676 67
rect 712 122 778 130
rect 712 88 728 122
rect 762 88 778 122
rect 712 17 778 88
rect 812 101 852 164
rect 812 67 818 101
rect 812 51 852 67
rect 888 149 904 183
rect 938 149 954 183
rect 888 93 954 149
rect 888 59 904 93
rect 938 59 954 93
rect 888 17 954 59
rect 988 169 990 203
rect 1024 169 1026 203
rect 988 101 1026 169
rect 988 67 990 101
rect 1024 67 1026 101
rect 988 51 1026 67
rect 1060 149 1076 183
rect 1110 149 1126 183
rect 1060 93 1126 149
rect 1060 59 1076 93
rect 1110 59 1126 93
rect 1060 17 1126 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21oi_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3677928
string GDS_START 3666920
<< end >>
