magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 7 241 453 243
rect 7 49 1319 241
rect 0 0 1344 49
<< scnmos >>
rect 86 49 116 217
rect 172 49 202 217
rect 258 49 288 217
rect 344 49 374 217
rect 578 47 608 215
rect 664 47 694 215
rect 750 47 780 215
rect 836 47 866 215
rect 938 47 968 215
rect 1038 47 1068 215
rect 1124 47 1154 215
rect 1210 47 1240 215
<< scpmoshvt >>
rect 219 367 249 619
rect 305 367 335 619
rect 391 367 421 619
rect 477 367 507 619
rect 578 367 608 619
rect 664 367 694 619
rect 750 367 780 619
rect 836 367 866 619
rect 952 367 982 619
rect 1038 367 1068 619
rect 1124 367 1154 619
rect 1210 367 1240 619
<< ndiff >>
rect 33 173 86 217
rect 33 139 41 173
rect 75 139 86 173
rect 33 95 86 139
rect 33 61 41 95
rect 75 61 86 95
rect 33 49 86 61
rect 116 205 172 217
rect 116 171 127 205
rect 161 171 172 205
rect 116 101 172 171
rect 116 67 127 101
rect 161 67 172 101
rect 116 49 172 67
rect 202 173 258 217
rect 202 139 213 173
rect 247 139 258 173
rect 202 91 258 139
rect 202 57 213 91
rect 247 57 258 91
rect 202 49 258 57
rect 288 205 344 217
rect 288 171 299 205
rect 333 171 344 205
rect 288 101 344 171
rect 288 67 299 101
rect 333 67 344 101
rect 288 49 344 67
rect 374 205 427 217
rect 374 171 385 205
rect 419 171 427 205
rect 374 95 427 171
rect 374 61 385 95
rect 419 61 427 95
rect 374 49 427 61
rect 525 187 578 215
rect 525 153 533 187
rect 567 153 578 187
rect 525 47 578 153
rect 608 97 664 215
rect 608 63 619 97
rect 653 63 664 97
rect 608 47 664 63
rect 694 175 750 215
rect 694 141 705 175
rect 739 141 750 175
rect 694 47 750 141
rect 780 97 836 215
rect 780 63 791 97
rect 825 63 836 97
rect 780 47 836 63
rect 866 181 938 215
rect 866 147 893 181
rect 927 147 938 181
rect 866 101 938 147
rect 866 67 893 101
rect 927 67 938 101
rect 866 47 938 67
rect 968 105 1038 215
rect 968 71 985 105
rect 1019 71 1038 105
rect 968 47 1038 71
rect 1068 181 1124 215
rect 1068 147 1079 181
rect 1113 147 1124 181
rect 1068 101 1124 147
rect 1068 67 1079 101
rect 1113 67 1124 101
rect 1068 47 1124 67
rect 1154 105 1210 215
rect 1154 71 1165 105
rect 1199 71 1210 105
rect 1154 47 1210 71
rect 1240 187 1293 215
rect 1240 153 1251 187
rect 1285 153 1293 187
rect 1240 101 1293 153
rect 1240 67 1251 101
rect 1285 67 1293 101
rect 1240 47 1293 67
<< pdiff >>
rect 166 607 219 619
rect 166 573 174 607
rect 208 573 219 607
rect 166 531 219 573
rect 166 497 174 531
rect 208 497 219 531
rect 166 453 219 497
rect 166 419 174 453
rect 208 419 219 453
rect 166 367 219 419
rect 249 599 305 619
rect 249 565 260 599
rect 294 565 305 599
rect 249 506 305 565
rect 249 472 260 506
rect 294 472 305 506
rect 249 413 305 472
rect 249 379 260 413
rect 294 379 305 413
rect 249 367 305 379
rect 335 607 391 619
rect 335 573 346 607
rect 380 573 391 607
rect 335 531 391 573
rect 335 497 346 531
rect 380 497 391 531
rect 335 455 391 497
rect 335 421 346 455
rect 380 421 391 455
rect 335 367 391 421
rect 421 599 477 619
rect 421 565 432 599
rect 466 565 477 599
rect 421 506 477 565
rect 421 472 432 506
rect 466 472 477 506
rect 421 413 477 472
rect 421 379 432 413
rect 466 379 477 413
rect 421 367 477 379
rect 507 607 578 619
rect 507 573 525 607
rect 559 573 578 607
rect 507 498 578 573
rect 507 464 525 498
rect 559 464 578 498
rect 507 367 578 464
rect 608 599 664 619
rect 608 565 619 599
rect 653 565 664 599
rect 608 504 664 565
rect 608 470 619 504
rect 653 470 664 504
rect 608 367 664 470
rect 694 540 750 619
rect 694 506 705 540
rect 739 506 750 540
rect 694 436 750 506
rect 694 402 705 436
rect 739 402 750 436
rect 694 367 750 402
rect 780 599 836 619
rect 780 565 791 599
rect 825 565 836 599
rect 780 504 836 565
rect 780 470 791 504
rect 825 470 836 504
rect 780 367 836 470
rect 866 607 952 619
rect 866 573 892 607
rect 926 573 952 607
rect 866 493 952 573
rect 866 459 892 493
rect 926 459 952 493
rect 866 367 952 459
rect 982 599 1038 619
rect 982 565 993 599
rect 1027 565 1038 599
rect 982 504 1038 565
rect 982 470 993 504
rect 1027 470 1038 504
rect 982 367 1038 470
rect 1068 541 1124 619
rect 1068 507 1079 541
rect 1113 507 1124 541
rect 1068 436 1124 507
rect 1068 402 1079 436
rect 1113 402 1124 436
rect 1068 367 1124 402
rect 1154 599 1210 619
rect 1154 565 1165 599
rect 1199 565 1210 599
rect 1154 514 1210 565
rect 1154 480 1165 514
rect 1199 480 1210 514
rect 1154 438 1210 480
rect 1154 404 1165 438
rect 1199 404 1210 438
rect 1154 367 1210 404
rect 1240 607 1293 619
rect 1240 573 1251 607
rect 1285 573 1293 607
rect 1240 510 1293 573
rect 1240 476 1251 510
rect 1285 476 1293 510
rect 1240 422 1293 476
rect 1240 388 1251 422
rect 1285 388 1293 422
rect 1240 367 1293 388
<< ndiffc >>
rect 41 139 75 173
rect 41 61 75 95
rect 127 171 161 205
rect 127 67 161 101
rect 213 139 247 173
rect 213 57 247 91
rect 299 171 333 205
rect 299 67 333 101
rect 385 171 419 205
rect 385 61 419 95
rect 533 153 567 187
rect 619 63 653 97
rect 705 141 739 175
rect 791 63 825 97
rect 893 147 927 181
rect 893 67 927 101
rect 985 71 1019 105
rect 1079 147 1113 181
rect 1079 67 1113 101
rect 1165 71 1199 105
rect 1251 153 1285 187
rect 1251 67 1285 101
<< pdiffc >>
rect 174 573 208 607
rect 174 497 208 531
rect 174 419 208 453
rect 260 565 294 599
rect 260 472 294 506
rect 260 379 294 413
rect 346 573 380 607
rect 346 497 380 531
rect 346 421 380 455
rect 432 565 466 599
rect 432 472 466 506
rect 432 379 466 413
rect 525 573 559 607
rect 525 464 559 498
rect 619 565 653 599
rect 619 470 653 504
rect 705 506 739 540
rect 705 402 739 436
rect 791 565 825 599
rect 791 470 825 504
rect 892 573 926 607
rect 892 459 926 493
rect 993 565 1027 599
rect 993 470 1027 504
rect 1079 507 1113 541
rect 1079 402 1113 436
rect 1165 565 1199 599
rect 1165 480 1199 514
rect 1165 404 1199 438
rect 1251 573 1285 607
rect 1251 476 1285 510
rect 1251 388 1285 422
<< poly >>
rect 219 619 249 645
rect 305 619 335 645
rect 391 619 421 645
rect 477 619 507 645
rect 578 619 608 645
rect 664 619 694 645
rect 750 619 780 645
rect 836 619 866 645
rect 952 619 982 645
rect 1038 619 1068 645
rect 1124 619 1154 645
rect 1210 619 1240 645
rect 219 331 249 367
rect 305 331 335 367
rect 391 331 421 367
rect 477 331 507 367
rect 86 315 507 331
rect 86 281 171 315
rect 205 281 239 315
rect 273 281 307 315
rect 341 281 375 315
rect 409 281 443 315
rect 477 281 507 315
rect 578 305 608 367
rect 664 335 694 367
rect 750 335 780 367
rect 664 319 780 335
rect 86 265 507 281
rect 556 289 622 305
rect 86 217 116 265
rect 172 217 202 265
rect 258 217 288 265
rect 344 217 374 265
rect 556 255 572 289
rect 606 255 622 289
rect 556 239 622 255
rect 664 285 730 319
rect 764 285 780 319
rect 836 303 866 367
rect 952 303 982 367
rect 1038 335 1068 367
rect 1124 335 1154 367
rect 1038 319 1154 335
rect 664 269 780 285
rect 578 215 608 239
rect 664 215 694 269
rect 750 215 780 269
rect 822 287 888 303
rect 822 253 838 287
rect 872 253 888 287
rect 822 237 888 253
rect 930 287 996 303
rect 930 253 946 287
rect 980 253 996 287
rect 930 237 996 253
rect 1038 285 1054 319
rect 1088 285 1154 319
rect 1038 269 1154 285
rect 836 215 866 237
rect 938 215 968 237
rect 1038 215 1068 269
rect 1124 215 1154 269
rect 1210 303 1240 367
rect 1210 287 1276 303
rect 1210 253 1226 287
rect 1260 253 1276 287
rect 1210 237 1276 253
rect 1210 215 1240 237
rect 86 23 116 49
rect 172 23 202 49
rect 258 23 288 49
rect 344 23 374 49
rect 578 21 608 47
rect 664 21 694 47
rect 750 21 780 47
rect 836 21 866 47
rect 938 21 968 47
rect 1038 21 1068 47
rect 1124 21 1154 47
rect 1210 21 1240 47
<< polycont >>
rect 171 281 205 315
rect 239 281 273 315
rect 307 281 341 315
rect 375 281 409 315
rect 443 281 477 315
rect 572 255 606 289
rect 730 285 764 319
rect 838 253 872 287
rect 946 253 980 287
rect 1054 285 1088 319
rect 1226 253 1260 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 158 607 224 649
rect 158 573 174 607
rect 208 573 224 607
rect 158 531 224 573
rect 158 497 174 531
rect 208 497 224 531
rect 158 453 224 497
rect 158 419 174 453
rect 208 419 224 453
rect 258 599 296 615
rect 258 565 260 599
rect 294 565 296 599
rect 258 506 296 565
rect 258 472 260 506
rect 294 472 296 506
rect 258 413 296 472
rect 330 607 396 649
rect 330 573 346 607
rect 380 573 396 607
rect 330 531 396 573
rect 330 497 346 531
rect 380 497 396 531
rect 330 455 396 497
rect 330 421 346 455
rect 380 421 396 455
rect 430 599 468 615
rect 430 565 432 599
rect 466 565 468 599
rect 430 506 468 565
rect 430 472 432 506
rect 466 472 468 506
rect 258 385 260 413
rect 17 379 260 385
rect 294 385 296 413
rect 430 413 468 472
rect 509 607 575 649
rect 509 573 525 607
rect 559 573 575 607
rect 509 498 575 573
rect 509 464 525 498
rect 559 464 575 498
rect 509 454 575 464
rect 609 599 841 615
rect 609 565 619 599
rect 653 581 791 599
rect 653 565 655 581
rect 609 504 655 565
rect 789 565 791 581
rect 825 565 841 599
rect 609 470 619 504
rect 653 470 655 504
rect 609 454 655 470
rect 689 540 755 547
rect 689 506 705 540
rect 739 506 755 540
rect 689 436 755 506
rect 789 504 841 565
rect 789 470 791 504
rect 825 470 841 504
rect 789 454 841 470
rect 876 607 942 649
rect 876 573 892 607
rect 926 573 942 607
rect 876 493 942 573
rect 876 459 892 493
rect 926 459 942 493
rect 876 454 942 459
rect 977 599 1201 615
rect 977 565 993 599
rect 1027 581 1165 599
rect 1027 565 1029 581
rect 977 504 1029 565
rect 1163 565 1165 581
rect 1199 565 1201 599
rect 977 470 993 504
rect 1027 470 1029 504
rect 977 454 1029 470
rect 1063 541 1129 547
rect 1063 507 1079 541
rect 1113 507 1129 541
rect 689 420 705 436
rect 430 385 432 413
rect 294 379 432 385
rect 466 379 468 413
rect 17 351 468 379
rect 502 402 705 420
rect 739 420 755 436
rect 1063 436 1129 507
rect 1063 420 1079 436
rect 739 402 1079 420
rect 1113 402 1129 436
rect 502 386 1129 402
rect 1163 514 1201 565
rect 1163 480 1165 514
rect 1199 480 1201 514
rect 1163 438 1201 480
rect 1163 404 1165 438
rect 1199 404 1201 438
rect 1163 388 1201 404
rect 1235 607 1301 649
rect 1235 573 1251 607
rect 1285 573 1301 607
rect 1235 510 1301 573
rect 1235 476 1251 510
rect 1285 476 1301 510
rect 1235 422 1301 476
rect 1235 388 1251 422
rect 1285 388 1301 422
rect 17 245 101 351
rect 502 315 536 386
rect 155 281 171 315
rect 205 281 239 315
rect 273 281 307 315
rect 341 281 375 315
rect 409 281 443 315
rect 477 281 536 315
rect 691 319 780 352
rect 572 289 657 305
rect 17 211 343 245
rect 125 205 163 211
rect 25 173 91 177
rect 25 139 41 173
rect 75 139 91 173
rect 25 95 91 139
rect 25 61 41 95
rect 75 61 91 95
rect 25 17 91 61
rect 125 171 127 205
rect 161 171 163 205
rect 297 205 343 211
rect 125 101 163 171
rect 125 67 127 101
rect 161 67 163 101
rect 125 51 163 67
rect 197 173 263 177
rect 197 139 213 173
rect 247 139 263 173
rect 197 91 263 139
rect 197 57 213 91
rect 247 57 263 91
rect 197 17 263 57
rect 297 171 299 205
rect 333 171 343 205
rect 297 101 343 171
rect 297 67 299 101
rect 333 67 343 101
rect 297 51 343 67
rect 377 205 425 221
rect 377 171 385 205
rect 419 171 425 205
rect 377 95 425 171
rect 377 61 385 95
rect 419 61 425 95
rect 377 17 425 61
rect 459 103 493 281
rect 606 255 657 289
rect 691 285 730 319
rect 764 285 780 319
rect 1038 319 1136 352
rect 691 283 780 285
rect 822 287 888 303
rect 572 249 657 255
rect 822 253 838 287
rect 872 253 888 287
rect 822 249 888 253
rect 572 239 888 249
rect 607 215 888 239
rect 930 287 996 303
rect 930 253 946 287
rect 980 253 996 287
rect 1038 285 1054 319
rect 1088 285 1136 319
rect 1170 287 1325 354
rect 930 249 996 253
rect 1170 253 1226 287
rect 1260 253 1325 287
rect 1170 249 1325 253
rect 930 237 1325 249
rect 930 215 1211 237
rect 527 187 573 203
rect 527 153 533 187
rect 567 181 573 187
rect 1245 187 1301 203
rect 1245 181 1251 187
rect 567 175 893 181
rect 567 153 705 175
rect 527 141 705 153
rect 739 147 893 175
rect 927 147 1079 181
rect 1113 153 1251 181
rect 1285 153 1301 187
rect 1113 147 1301 153
rect 739 141 935 147
rect 527 137 935 141
rect 459 97 841 103
rect 459 63 619 97
rect 653 63 791 97
rect 825 63 841 97
rect 459 51 841 63
rect 877 101 935 137
rect 877 67 893 101
rect 927 67 935 101
rect 877 51 935 67
rect 969 105 1035 113
rect 969 71 985 105
rect 1019 71 1035 105
rect 969 17 1035 71
rect 1069 101 1115 147
rect 1069 67 1079 101
rect 1113 67 1115 101
rect 1069 51 1115 67
rect 1149 105 1215 113
rect 1149 71 1165 105
rect 1199 71 1215 105
rect 1149 17 1215 71
rect 1249 101 1301 147
rect 1249 67 1251 101
rect 1285 67 1301 101
rect 1249 51 1301 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o22a_4
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 945302
string GDS_START 934076
<< end >>
