magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 752 247
rect 0 0 768 49
<< scnmos >>
rect 80 137 110 221
rect 204 53 234 221
rect 290 53 320 221
rect 459 137 489 221
rect 531 137 561 221
rect 639 137 669 221
<< scpmoshvt >>
rect 92 367 122 451
rect 204 367 234 619
rect 290 367 320 619
rect 456 367 486 451
rect 542 367 572 451
rect 645 367 675 451
<< ndiff >>
rect 27 196 80 221
rect 27 162 35 196
rect 69 162 80 196
rect 27 137 80 162
rect 110 137 204 221
rect 132 73 204 137
rect 132 39 140 73
rect 174 53 204 73
rect 234 213 290 221
rect 234 179 245 213
rect 279 179 290 213
rect 234 53 290 179
rect 320 137 459 221
rect 489 137 531 221
rect 561 137 639 221
rect 669 196 726 221
rect 669 162 684 196
rect 718 162 726 196
rect 669 137 726 162
rect 320 73 400 137
rect 320 53 354 73
rect 174 39 182 53
rect 132 27 182 39
rect 342 39 354 53
rect 388 39 400 73
rect 342 31 400 39
<< pdiff >>
rect 145 607 204 619
rect 145 573 153 607
rect 187 573 204 607
rect 145 519 204 573
rect 145 485 153 519
rect 187 485 204 519
rect 145 451 204 485
rect 39 424 92 451
rect 39 390 47 424
rect 81 390 92 424
rect 39 367 92 390
rect 122 436 204 451
rect 122 402 133 436
rect 167 402 204 436
rect 122 367 204 402
rect 234 599 290 619
rect 234 565 245 599
rect 279 565 290 599
rect 234 503 290 565
rect 234 469 245 503
rect 279 469 290 503
rect 234 413 290 469
rect 234 379 245 413
rect 279 379 290 413
rect 234 367 290 379
rect 320 607 377 619
rect 320 573 335 607
rect 369 573 377 607
rect 320 539 377 573
rect 320 505 335 539
rect 369 505 377 539
rect 320 469 377 505
rect 320 435 335 469
rect 369 451 377 469
rect 369 435 456 451
rect 320 367 456 435
rect 486 424 542 451
rect 486 390 497 424
rect 531 390 542 424
rect 486 367 542 390
rect 572 439 645 451
rect 572 405 595 439
rect 629 405 645 439
rect 572 367 645 405
rect 675 424 728 451
rect 675 390 686 424
rect 720 390 728 424
rect 675 367 728 390
<< ndiffc >>
rect 35 162 69 196
rect 140 39 174 73
rect 245 179 279 213
rect 684 162 718 196
rect 354 39 388 73
<< pdiffc >>
rect 153 573 187 607
rect 153 485 187 519
rect 47 390 81 424
rect 133 402 167 436
rect 245 565 279 599
rect 245 469 279 503
rect 245 379 279 413
rect 335 573 369 607
rect 335 505 369 539
rect 335 435 369 469
rect 497 390 531 424
rect 595 405 629 439
rect 686 390 720 424
<< poly >>
rect 204 619 234 645
rect 290 619 320 645
rect 92 451 122 477
rect 456 451 486 477
rect 542 451 572 477
rect 645 451 675 477
rect 92 309 122 367
rect 204 325 234 367
rect 290 325 320 367
rect 204 309 381 325
rect 456 309 486 367
rect 542 309 572 367
rect 80 293 151 309
rect 80 259 101 293
rect 135 259 151 293
rect 80 243 151 259
rect 204 295 331 309
rect 80 221 110 243
rect 204 221 234 295
rect 290 275 331 295
rect 365 275 381 309
rect 290 259 381 275
rect 423 293 489 309
rect 423 259 439 293
rect 473 259 489 293
rect 290 221 320 259
rect 423 243 489 259
rect 459 221 489 243
rect 531 293 597 309
rect 531 259 547 293
rect 581 259 597 293
rect 645 273 675 367
rect 531 243 597 259
rect 639 243 675 273
rect 531 221 561 243
rect 639 221 669 243
rect 80 111 110 137
rect 459 111 489 137
rect 531 111 561 137
rect 639 115 669 137
rect 204 27 234 53
rect 290 27 320 53
rect 609 99 675 115
rect 609 65 625 99
rect 659 65 675 99
rect 609 49 675 65
<< polycont >>
rect 101 259 135 293
rect 331 275 365 309
rect 439 259 473 293
rect 547 259 581 293
rect 625 65 659 99
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 131 607 189 649
rect 131 573 153 607
rect 187 573 189 607
rect 131 519 189 573
rect 131 485 153 519
rect 187 485 189 519
rect 19 424 97 440
rect 19 390 47 424
rect 81 390 97 424
rect 19 386 97 390
rect 131 436 189 485
rect 131 402 133 436
rect 167 402 189 436
rect 131 386 189 402
rect 223 599 295 615
rect 223 565 245 599
rect 279 565 295 599
rect 223 503 295 565
rect 223 469 245 503
rect 279 469 295 503
rect 223 413 295 469
rect 329 607 385 649
rect 329 573 335 607
rect 369 573 385 607
rect 329 539 385 573
rect 329 505 335 539
rect 369 505 385 539
rect 329 469 385 505
rect 329 435 335 469
rect 369 435 385 469
rect 329 419 385 435
rect 481 424 543 440
rect 19 208 65 386
rect 223 379 245 413
rect 279 379 295 413
rect 481 390 497 424
rect 531 390 543 424
rect 579 439 645 649
rect 579 405 595 439
rect 629 405 645 439
rect 579 399 645 405
rect 682 424 734 440
rect 481 385 543 390
rect 101 293 184 352
rect 135 259 184 293
rect 101 242 184 259
rect 223 213 295 379
rect 329 365 543 385
rect 682 390 686 424
rect 720 390 734 424
rect 682 365 734 390
rect 329 343 734 365
rect 329 309 371 343
rect 509 331 734 343
rect 329 275 331 309
rect 365 275 371 309
rect 329 259 371 275
rect 405 293 473 309
rect 405 259 439 293
rect 405 226 473 259
rect 507 293 646 297
rect 507 259 547 293
rect 581 259 646 293
rect 507 226 646 259
rect 19 196 85 208
rect 19 162 35 196
rect 69 162 85 196
rect 223 179 245 213
rect 279 179 295 213
rect 223 177 295 179
rect 680 196 734 331
rect 19 143 85 162
rect 329 143 646 174
rect 680 162 684 196
rect 718 162 734 196
rect 680 146 734 162
rect 19 112 646 143
rect 19 109 675 112
rect 609 99 675 109
rect 124 73 190 75
rect 124 39 140 73
rect 174 39 190 73
rect 124 17 190 39
rect 338 73 404 75
rect 338 39 354 73
rect 388 39 404 73
rect 609 65 625 99
rect 659 65 675 99
rect 609 51 675 65
rect 338 17 404 39
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and3b_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6379858
string GDS_START 6373092
<< end >>
