magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 738 241
rect 0 0 768 49
<< scnmos >>
rect 80 47 110 215
rect 318 47 348 215
rect 408 47 438 215
rect 515 47 545 215
rect 629 47 659 215
<< scpmoshvt >>
rect 183 367 213 619
rect 318 367 348 619
rect 396 367 426 619
rect 515 367 545 619
rect 629 367 659 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 135 80 169
rect 27 101 35 135
rect 69 101 80 135
rect 27 47 80 101
rect 110 161 163 215
rect 110 127 121 161
rect 155 127 163 161
rect 110 93 163 127
rect 110 59 121 93
rect 155 59 163 93
rect 110 47 163 59
rect 265 175 318 215
rect 265 141 273 175
rect 307 141 318 175
rect 265 107 318 141
rect 265 73 273 107
rect 307 73 318 107
rect 265 47 318 73
rect 348 203 408 215
rect 348 169 363 203
rect 397 169 408 203
rect 348 47 408 169
rect 438 187 515 215
rect 438 153 449 187
rect 483 153 515 187
rect 438 119 515 153
rect 438 85 449 119
rect 483 85 515 119
rect 438 47 515 85
rect 545 161 629 215
rect 545 127 556 161
rect 590 127 629 161
rect 545 93 629 127
rect 545 59 556 93
rect 590 59 629 93
rect 545 47 629 59
rect 659 203 712 215
rect 659 169 670 203
rect 704 169 712 203
rect 659 135 712 169
rect 659 101 670 135
rect 704 101 712 135
rect 659 47 712 101
<< pdiff >>
rect 130 549 183 619
rect 130 515 138 549
rect 172 515 183 549
rect 130 481 183 515
rect 130 447 138 481
rect 172 447 183 481
rect 130 413 183 447
rect 130 379 138 413
rect 172 379 183 413
rect 130 367 183 379
rect 213 607 318 619
rect 213 573 224 607
rect 258 573 318 607
rect 213 539 318 573
rect 213 505 224 539
rect 258 505 318 539
rect 213 367 318 505
rect 348 367 396 619
rect 426 572 515 619
rect 426 538 437 572
rect 471 538 515 572
rect 426 504 515 538
rect 426 470 437 504
rect 471 470 515 504
rect 426 436 515 470
rect 426 402 437 436
rect 471 402 515 436
rect 426 367 515 402
rect 545 367 629 619
rect 659 607 723 619
rect 659 573 681 607
rect 715 573 723 607
rect 659 539 723 573
rect 659 505 681 539
rect 715 505 723 539
rect 659 471 723 505
rect 659 437 681 471
rect 715 437 723 471
rect 659 367 723 437
<< ndiffc >>
rect 35 169 69 203
rect 35 101 69 135
rect 121 127 155 161
rect 121 59 155 93
rect 273 141 307 175
rect 273 73 307 107
rect 363 169 397 203
rect 449 153 483 187
rect 449 85 483 119
rect 556 127 590 161
rect 556 59 590 93
rect 670 169 704 203
rect 670 101 704 135
<< pdiffc >>
rect 138 515 172 549
rect 138 447 172 481
rect 138 379 172 413
rect 224 573 258 607
rect 224 505 258 539
rect 437 538 471 572
rect 437 470 471 504
rect 437 402 471 436
rect 681 573 715 607
rect 681 505 715 539
rect 681 437 715 471
<< poly >>
rect 183 619 213 645
rect 318 619 348 645
rect 396 619 426 645
rect 515 619 545 645
rect 629 619 659 645
rect 183 303 213 367
rect 318 335 348 367
rect 80 287 213 303
rect 80 253 126 287
rect 160 253 213 287
rect 282 319 348 335
rect 282 285 298 319
rect 332 285 348 319
rect 282 269 348 285
rect 396 335 426 367
rect 515 335 545 367
rect 396 319 462 335
rect 396 285 412 319
rect 446 285 462 319
rect 396 269 462 285
rect 515 319 581 335
rect 515 285 531 319
rect 565 285 581 319
rect 515 269 581 285
rect 629 325 659 367
rect 629 309 743 325
rect 629 275 693 309
rect 727 275 743 309
rect 80 237 213 253
rect 80 215 110 237
rect 318 215 348 269
rect 408 215 438 269
rect 515 215 545 269
rect 629 259 743 275
rect 629 215 659 259
rect 80 21 110 47
rect 318 21 348 47
rect 408 21 438 47
rect 515 21 545 47
rect 629 21 659 47
<< polycont >>
rect 126 253 160 287
rect 298 285 332 319
rect 412 285 446 319
rect 531 285 565 319
rect 693 275 727 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 220 607 262 649
rect 220 573 224 607
rect 258 573 262 607
rect 677 607 719 649
rect 31 397 73 572
rect 134 549 176 565
rect 134 515 138 549
rect 172 515 176 549
rect 134 481 176 515
rect 220 539 262 573
rect 220 505 224 539
rect 258 505 262 539
rect 220 489 262 505
rect 433 572 475 588
rect 677 573 681 607
rect 715 573 719 607
rect 433 538 437 572
rect 471 538 475 572
rect 433 504 475 538
rect 134 447 138 481
rect 172 447 176 481
rect 134 413 176 447
rect 433 470 437 504
rect 471 470 475 504
rect 433 436 475 470
rect 433 420 437 436
rect 134 397 138 413
rect 31 379 138 397
rect 172 379 176 413
rect 31 363 176 379
rect 212 402 437 420
rect 471 402 475 436
rect 212 386 475 402
rect 31 203 73 363
rect 110 253 126 287
rect 160 253 176 287
rect 110 249 176 253
rect 212 249 246 386
rect 282 319 353 350
rect 282 285 298 319
rect 332 285 353 319
rect 396 319 462 350
rect 396 285 412 319
rect 446 285 462 319
rect 511 319 641 572
rect 677 539 719 573
rect 677 505 681 539
rect 715 505 719 539
rect 677 471 719 505
rect 677 437 681 471
rect 715 437 719 471
rect 677 421 719 437
rect 511 285 531 319
rect 565 285 641 319
rect 677 309 743 350
rect 677 275 693 309
rect 727 275 743 309
rect 110 215 401 249
rect 31 169 35 203
rect 69 169 73 203
rect 359 203 401 215
rect 31 135 73 169
rect 31 101 35 135
rect 69 101 73 135
rect 31 85 73 101
rect 117 161 159 177
rect 117 127 121 161
rect 155 127 159 161
rect 117 93 159 127
rect 117 59 121 93
rect 155 59 159 93
rect 257 175 323 179
rect 257 141 273 175
rect 307 141 323 175
rect 359 169 363 203
rect 397 169 401 203
rect 359 153 401 169
rect 445 203 708 235
rect 445 201 670 203
rect 445 187 487 201
rect 445 153 449 187
rect 483 153 487 187
rect 666 169 670 201
rect 704 169 708 203
rect 257 107 323 141
rect 257 73 273 107
rect 307 103 323 107
rect 445 119 487 153
rect 445 103 449 119
rect 307 85 449 103
rect 483 85 487 119
rect 307 73 487 85
rect 257 69 487 73
rect 540 161 606 165
rect 540 127 556 161
rect 590 127 606 161
rect 540 93 606 127
rect 117 17 159 59
rect 540 59 556 93
rect 590 59 606 93
rect 666 135 708 169
rect 666 101 670 135
rect 704 101 708 135
rect 666 85 708 101
rect 540 17 606 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o22a_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 953350
string GDS_START 945358
<< end >>
