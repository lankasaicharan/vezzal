magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2126 1852
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 778 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 277 47 307 177
rect 382 47 412 177
rect 510 47 540 177
rect 652 47 682 177
<< scpmoshvt >>
rect 81 297 117 497
rect 279 297 315 497
rect 384 297 420 497
rect 512 297 548 497
rect 654 297 690 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 161 171 177
rect 109 127 129 161
rect 163 127 171 161
rect 109 93 171 127
rect 109 59 129 93
rect 163 59 171 93
rect 109 47 171 59
rect 225 161 277 177
rect 225 127 233 161
rect 267 127 277 161
rect 225 93 277 127
rect 225 59 233 93
rect 267 59 277 93
rect 225 47 277 59
rect 307 93 382 177
rect 307 59 333 93
rect 367 59 382 93
rect 307 47 382 59
rect 412 161 510 177
rect 412 127 432 161
rect 466 127 510 161
rect 412 93 510 127
rect 412 59 432 93
rect 466 59 510 93
rect 412 47 510 59
rect 540 47 652 177
rect 682 161 752 177
rect 682 127 710 161
rect 744 127 752 161
rect 682 93 752 127
rect 682 59 710 93
rect 744 59 752 93
rect 682 47 752 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 171 497
rect 117 451 129 485
rect 163 451 171 485
rect 117 417 171 451
rect 117 383 129 417
rect 163 383 171 417
rect 117 349 171 383
rect 117 315 129 349
rect 163 315 171 349
rect 117 297 171 315
rect 225 485 279 497
rect 225 451 233 485
rect 267 451 279 485
rect 225 417 279 451
rect 225 383 233 417
rect 267 383 279 417
rect 225 297 279 383
rect 315 297 384 497
rect 420 485 512 497
rect 420 451 443 485
rect 477 451 512 485
rect 420 417 512 451
rect 420 383 443 417
rect 477 383 512 417
rect 420 349 512 383
rect 420 315 443 349
rect 477 315 512 349
rect 420 297 512 315
rect 548 485 654 497
rect 548 451 568 485
rect 602 451 654 485
rect 548 417 654 451
rect 548 383 568 417
rect 602 383 654 417
rect 548 297 654 383
rect 690 485 752 497
rect 690 451 710 485
rect 744 451 752 485
rect 690 417 752 451
rect 690 383 710 417
rect 744 383 752 417
rect 690 349 752 383
rect 690 315 710 349
rect 744 315 752 349
rect 690 297 752 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 127 163 161
rect 129 59 163 93
rect 233 127 267 161
rect 233 59 267 93
rect 333 59 367 93
rect 432 127 466 161
rect 432 59 466 93
rect 710 127 744 161
rect 710 59 744 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 233 451 267 485
rect 233 383 267 417
rect 443 451 477 485
rect 443 383 477 417
rect 443 315 477 349
rect 568 451 602 485
rect 568 383 602 417
rect 710 451 744 485
rect 710 383 744 417
rect 710 315 744 349
<< poly >>
rect 81 497 117 523
rect 279 497 315 523
rect 384 497 420 523
rect 512 497 548 523
rect 654 497 690 523
rect 81 282 117 297
rect 279 282 315 297
rect 384 282 420 297
rect 512 282 548 297
rect 654 282 690 297
rect 79 259 119 282
rect 277 265 317 282
rect 382 265 422 282
rect 510 265 550 282
rect 652 265 692 282
rect 79 249 162 259
rect 79 215 102 249
rect 136 215 162 249
rect 79 205 162 215
rect 277 249 340 265
rect 277 215 288 249
rect 322 215 340 249
rect 79 177 109 205
rect 277 199 340 215
rect 382 249 468 265
rect 382 215 424 249
rect 458 215 468 249
rect 382 199 468 215
rect 510 249 578 265
rect 510 215 524 249
rect 558 215 578 249
rect 510 199 578 215
rect 652 249 797 265
rect 652 215 747 249
rect 781 215 797 249
rect 652 199 797 215
rect 277 177 307 199
rect 382 177 412 199
rect 510 177 540 199
rect 652 177 682 199
rect 79 21 109 47
rect 277 21 307 47
rect 382 21 412 47
rect 510 21 540 47
rect 652 21 682 47
<< polycont >>
rect 102 215 136 249
rect 288 215 322 249
rect 424 215 458 249
rect 524 215 558 249
rect 747 215 781 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 485 85 493
rect 17 451 35 485
rect 69 451 85 485
rect 17 417 85 451
rect 17 383 35 417
rect 69 383 85 417
rect 17 349 85 383
rect 17 315 35 349
rect 69 315 85 349
rect 17 299 85 315
rect 129 485 163 527
rect 129 417 163 451
rect 129 349 163 383
rect 217 485 267 527
rect 217 451 233 485
rect 217 417 267 451
rect 217 383 233 417
rect 217 367 267 383
rect 417 485 493 493
rect 417 451 443 485
rect 477 451 493 485
rect 417 417 493 451
rect 417 383 443 417
rect 477 383 493 417
rect 417 349 493 383
rect 552 485 618 527
rect 552 451 568 485
rect 602 451 618 485
rect 552 417 618 451
rect 552 383 568 417
rect 602 383 618 417
rect 552 367 618 383
rect 694 485 760 493
rect 694 451 710 485
rect 744 451 760 485
rect 694 417 760 451
rect 694 383 710 417
rect 744 383 760 417
rect 417 333 443 349
rect 129 299 163 315
rect 201 315 443 333
rect 477 333 493 349
rect 694 349 760 383
rect 694 333 710 349
rect 477 315 710 333
rect 744 315 760 349
rect 201 299 760 315
rect 17 177 52 299
rect 201 249 235 299
rect 86 215 102 249
rect 136 215 235 249
rect 270 249 363 255
rect 270 215 288 249
rect 322 215 363 249
rect 397 249 474 255
rect 397 215 424 249
rect 458 215 474 249
rect 508 249 616 255
rect 508 215 524 249
rect 558 215 616 249
rect 17 161 85 177
rect 17 127 35 161
rect 69 127 85 161
rect 17 93 85 127
rect 17 59 35 93
rect 69 59 85 93
rect 17 51 85 59
rect 129 161 179 177
rect 163 127 179 161
rect 129 93 179 127
rect 163 59 179 93
rect 129 17 179 59
rect 217 161 482 181
rect 217 127 233 161
rect 267 147 432 161
rect 267 127 283 147
rect 217 93 283 127
rect 406 127 432 147
rect 466 127 482 161
rect 217 59 233 93
rect 267 59 283 93
rect 217 51 283 59
rect 327 93 372 109
rect 327 59 333 93
rect 367 59 372 93
rect 327 17 372 59
rect 406 93 482 127
rect 406 59 432 93
rect 466 59 482 93
rect 563 87 616 215
rect 650 173 694 299
rect 728 249 801 265
rect 728 215 747 249
rect 781 215 801 249
rect 650 161 760 173
rect 650 127 710 161
rect 744 127 760 161
rect 650 93 760 127
rect 406 51 482 59
rect 650 59 710 93
rect 744 59 760 93
rect 650 51 760 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 755 221 789 255 0 FreeSans 250 0 0 0 C1
port 4 nsew signal input
flabel locali s 524 221 568 255 0 FreeSans 250 0 0 0 B1
port 3 nsew signal input
flabel locali s 432 221 466 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 304 221 338 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 30 85 64 119 0 FreeSans 250 0 0 0 X
port 9 nsew signal output
flabel locali s 30 425 64 459 0 FreeSans 250 0 0 0 X
port 9 nsew signal output
flabel locali s 30 357 64 391 0 FreeSans 250 0 0 0 X
port 9 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o211a_1
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1034664
string GDS_START 1027576
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
