magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 4 49 767 248
rect 0 0 768 49
<< scpmos >>
rect 84 368 114 568
rect 192 368 222 568
rect 284 368 314 568
rect 378 368 408 568
rect 552 368 582 592
rect 642 368 672 592
<< nmoslvt >>
rect 87 74 117 222
rect 165 74 195 222
rect 267 74 297 222
rect 379 74 409 222
rect 571 74 601 222
rect 657 74 687 222
<< ndiff >>
rect 30 199 87 222
rect 30 165 42 199
rect 76 165 87 199
rect 30 120 87 165
rect 30 86 42 120
rect 76 86 87 120
rect 30 74 87 86
rect 117 74 165 222
rect 195 136 267 222
rect 195 102 221 136
rect 255 102 267 136
rect 195 74 267 102
rect 297 84 379 222
rect 297 74 321 84
rect 312 50 321 74
rect 355 74 379 84
rect 409 136 463 222
rect 409 102 420 136
rect 454 102 463 136
rect 409 74 463 102
rect 517 136 571 222
rect 517 102 526 136
rect 560 102 571 136
rect 517 74 571 102
rect 601 210 657 222
rect 601 176 612 210
rect 646 176 657 210
rect 601 120 657 176
rect 601 86 612 120
rect 646 86 657 120
rect 601 74 657 86
rect 687 210 741 222
rect 687 176 698 210
rect 732 176 741 210
rect 687 120 741 176
rect 687 86 698 120
rect 732 86 741 120
rect 687 74 741 86
rect 355 50 364 74
rect 312 38 364 50
<< pdiff >>
rect 499 568 552 592
rect 27 556 84 568
rect 27 522 37 556
rect 71 522 84 556
rect 27 485 84 522
rect 27 451 37 485
rect 71 451 84 485
rect 27 414 84 451
rect 27 380 37 414
rect 71 380 84 414
rect 27 368 84 380
rect 114 560 192 568
rect 114 526 137 560
rect 171 526 192 560
rect 114 492 192 526
rect 114 458 137 492
rect 171 458 192 492
rect 114 368 192 458
rect 222 560 284 568
rect 222 526 237 560
rect 271 526 284 560
rect 222 492 284 526
rect 222 458 237 492
rect 271 458 284 492
rect 222 424 284 458
rect 222 390 237 424
rect 271 390 284 424
rect 222 368 284 390
rect 314 368 378 568
rect 408 560 552 568
rect 408 526 421 560
rect 455 526 495 560
rect 529 526 552 560
rect 408 492 552 526
rect 408 458 421 492
rect 455 458 495 492
rect 529 458 552 492
rect 408 368 552 458
rect 582 580 642 592
rect 582 546 595 580
rect 629 546 642 580
rect 582 497 642 546
rect 582 463 595 497
rect 629 463 642 497
rect 582 414 642 463
rect 582 380 595 414
rect 629 380 642 414
rect 582 368 642 380
rect 672 580 741 592
rect 672 546 695 580
rect 729 546 741 580
rect 672 497 741 546
rect 672 463 695 497
rect 729 463 741 497
rect 672 414 741 463
rect 672 380 695 414
rect 729 380 741 414
rect 672 368 741 380
<< ndiffc >>
rect 42 165 76 199
rect 42 86 76 120
rect 221 102 255 136
rect 321 50 355 84
rect 420 102 454 136
rect 526 102 560 136
rect 612 176 646 210
rect 612 86 646 120
rect 698 176 732 210
rect 698 86 732 120
<< pdiffc >>
rect 37 522 71 556
rect 37 451 71 485
rect 37 380 71 414
rect 137 526 171 560
rect 137 458 171 492
rect 237 526 271 560
rect 237 458 271 492
rect 237 390 271 424
rect 421 526 455 560
rect 495 526 529 560
rect 421 458 455 492
rect 495 458 529 492
rect 595 546 629 580
rect 595 463 629 497
rect 595 380 629 414
rect 695 546 729 580
rect 695 463 729 497
rect 695 380 729 414
<< poly >>
rect 84 568 114 594
rect 192 568 222 594
rect 284 568 314 594
rect 378 568 408 594
rect 552 592 582 618
rect 642 592 672 618
rect 84 353 114 368
rect 192 353 222 368
rect 284 353 314 368
rect 378 353 408 368
rect 552 353 582 368
rect 642 353 672 368
rect 81 310 117 353
rect 189 336 225 353
rect 281 336 317 353
rect 375 336 411 353
rect 549 345 585 353
rect 21 294 117 310
rect 21 260 37 294
rect 71 260 117 294
rect 159 320 225 336
rect 159 286 175 320
rect 209 286 225 320
rect 159 270 225 286
rect 267 320 333 336
rect 267 286 283 320
rect 317 286 333 320
rect 267 270 333 286
rect 375 320 459 336
rect 375 286 409 320
rect 443 286 459 320
rect 375 270 459 286
rect 501 315 585 345
rect 639 315 675 353
rect 501 310 675 315
rect 501 276 517 310
rect 551 276 675 310
rect 21 244 117 260
rect 87 222 117 244
rect 165 222 195 270
rect 267 222 297 270
rect 379 222 409 270
rect 501 267 675 276
rect 501 237 687 267
rect 571 222 601 237
rect 657 222 687 237
rect 87 48 117 74
rect 165 48 195 74
rect 267 48 297 74
rect 379 48 409 74
rect 571 48 601 74
rect 657 48 687 74
<< polycont >>
rect 37 260 71 294
rect 175 286 209 320
rect 283 286 317 320
rect 409 286 443 320
rect 517 276 551 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 21 556 87 572
rect 21 522 37 556
rect 71 522 87 556
rect 21 485 87 522
rect 21 451 37 485
rect 71 451 87 485
rect 121 560 187 649
rect 121 526 137 560
rect 171 526 187 560
rect 121 492 187 526
rect 121 458 137 492
rect 171 458 187 492
rect 221 560 287 572
rect 221 526 237 560
rect 271 526 287 560
rect 221 492 287 526
rect 221 458 237 492
rect 271 458 287 492
rect 405 560 545 649
rect 405 526 421 560
rect 455 526 495 560
rect 529 526 545 560
rect 405 492 545 526
rect 405 458 421 492
rect 455 458 495 492
rect 529 458 545 492
rect 579 580 645 596
rect 579 546 595 580
rect 629 546 645 580
rect 579 497 645 546
rect 579 463 595 497
rect 629 463 645 497
rect 21 424 87 451
rect 221 424 287 458
rect 21 414 237 424
rect 21 380 37 414
rect 71 390 237 414
rect 271 390 535 424
rect 71 380 87 390
rect 21 364 87 380
rect 121 320 225 356
rect 21 294 87 310
rect 21 260 37 294
rect 71 260 87 294
rect 121 286 175 320
rect 209 286 225 320
rect 121 270 225 286
rect 267 320 359 356
rect 267 286 283 320
rect 317 286 359 320
rect 267 270 359 286
rect 393 320 459 356
rect 393 286 409 320
rect 443 286 459 320
rect 393 270 459 286
rect 501 326 535 390
rect 579 414 645 463
rect 579 380 595 414
rect 629 380 645 414
rect 579 364 645 380
rect 679 580 745 649
rect 679 546 695 580
rect 729 546 745 580
rect 679 497 745 546
rect 679 463 695 497
rect 729 463 745 497
rect 679 414 745 463
rect 679 380 695 414
rect 729 380 745 414
rect 679 364 745 380
rect 501 310 567 326
rect 501 276 517 310
rect 551 276 567 310
rect 21 236 87 260
rect 501 260 567 276
rect 601 282 645 364
rect 501 236 535 260
rect 121 202 535 236
rect 601 226 647 282
rect 596 210 647 226
rect 26 199 155 202
rect 26 165 42 199
rect 76 165 155 199
rect 596 176 612 210
rect 646 176 647 210
rect 26 120 155 165
rect 26 86 42 120
rect 76 86 155 120
rect 26 70 155 86
rect 205 136 470 168
rect 205 102 221 136
rect 255 134 420 136
rect 255 102 271 134
rect 205 70 271 102
rect 404 102 420 134
rect 454 102 470 136
rect 305 84 355 100
rect 305 50 321 84
rect 404 70 470 102
rect 510 136 560 168
rect 510 102 526 136
rect 305 17 355 50
rect 510 17 560 102
rect 596 120 647 176
rect 596 86 612 120
rect 646 86 647 120
rect 596 70 647 86
rect 682 210 748 226
rect 682 176 698 210
rect 732 176 748 210
rect 682 120 748 176
rect 682 86 698 120
rect 732 86 748 120
rect 682 17 748 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o211a_2
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 1654436
string GDS_START 1647156
<< end >>
