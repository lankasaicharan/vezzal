magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 191 159 551 168
rect 1 49 551 159
rect 0 0 576 49
<< scnmos >>
rect 80 49 110 133
rect 270 58 300 142
rect 356 58 386 142
rect 442 58 472 142
<< scpmoshvt >>
rect 113 483 143 611
rect 210 483 240 611
rect 307 483 337 611
rect 379 483 409 611
<< ndiff >>
rect 27 105 80 133
rect 27 71 35 105
rect 69 71 80 105
rect 27 49 80 71
rect 110 105 163 133
rect 110 71 121 105
rect 155 71 163 105
rect 110 49 163 71
rect 217 117 270 142
rect 217 83 225 117
rect 259 83 270 117
rect 217 58 270 83
rect 300 117 356 142
rect 300 83 311 117
rect 345 83 356 117
rect 300 58 356 83
rect 386 117 442 142
rect 386 83 397 117
rect 431 83 442 117
rect 386 58 442 83
rect 472 117 525 142
rect 472 83 483 117
rect 517 83 525 117
rect 472 58 525 83
<< pdiff >>
rect 60 599 113 611
rect 60 565 68 599
rect 102 565 113 599
rect 60 529 113 565
rect 60 495 68 529
rect 102 495 113 529
rect 60 483 113 495
rect 143 599 210 611
rect 143 565 163 599
rect 197 565 210 599
rect 143 529 210 565
rect 143 495 163 529
rect 197 495 210 529
rect 143 483 210 495
rect 240 599 307 611
rect 240 565 251 599
rect 285 565 307 599
rect 240 529 307 565
rect 240 495 251 529
rect 285 495 307 529
rect 240 483 307 495
rect 337 483 379 611
rect 409 599 462 611
rect 409 565 420 599
rect 454 565 462 599
rect 409 529 462 565
rect 409 495 420 529
rect 454 495 462 529
rect 409 483 462 495
<< ndiffc >>
rect 35 71 69 105
rect 121 71 155 105
rect 225 83 259 117
rect 311 83 345 117
rect 397 83 431 117
rect 483 83 517 117
<< pdiffc >>
rect 68 565 102 599
rect 68 495 102 529
rect 163 565 197 599
rect 163 495 197 529
rect 251 565 285 599
rect 251 495 285 529
rect 420 565 454 599
rect 420 495 454 529
<< poly >>
rect 113 611 143 637
rect 210 611 240 637
rect 307 611 337 637
rect 379 611 409 637
rect 113 289 143 483
rect 210 359 240 483
rect 307 376 337 483
rect 379 454 409 483
rect 379 429 500 454
rect 379 424 450 429
rect 434 395 450 424
rect 484 395 500 429
rect 307 360 386 376
rect 199 343 265 359
rect 199 309 215 343
rect 249 309 265 343
rect 80 273 151 289
rect 80 239 101 273
rect 135 239 151 273
rect 80 205 151 239
rect 199 275 265 309
rect 199 241 215 275
rect 249 241 265 275
rect 307 326 329 360
rect 363 326 386 360
rect 307 292 386 326
rect 434 361 500 395
rect 434 327 450 361
rect 484 327 500 361
rect 434 311 500 327
rect 307 258 329 292
rect 363 258 386 292
rect 307 242 386 258
rect 199 225 265 241
rect 80 171 101 205
rect 135 171 151 205
rect 80 155 151 171
rect 235 194 265 225
rect 235 164 300 194
rect 80 133 110 155
rect 270 142 300 164
rect 356 142 386 242
rect 442 142 472 311
rect 80 23 110 49
rect 270 32 300 58
rect 356 32 386 58
rect 442 32 472 58
<< polycont >>
rect 450 395 484 429
rect 215 309 249 343
rect 101 239 135 273
rect 215 241 249 275
rect 329 326 363 360
rect 450 327 484 361
rect 329 258 363 292
rect 101 171 135 205
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 17 599 113 615
rect 17 565 68 599
rect 102 565 113 599
rect 17 529 113 565
rect 17 495 68 529
rect 102 495 113 529
rect 17 479 113 495
rect 147 599 201 649
rect 147 565 163 599
rect 197 565 201 599
rect 147 529 201 565
rect 147 495 163 529
rect 197 495 201 529
rect 147 479 201 495
rect 235 599 285 615
rect 235 565 251 599
rect 404 599 470 649
rect 235 529 285 565
rect 235 495 251 529
rect 17 121 67 479
rect 235 443 285 495
rect 101 409 285 443
rect 101 273 151 409
rect 319 360 368 594
rect 404 565 420 599
rect 454 565 470 599
rect 404 529 470 565
rect 404 495 420 529
rect 454 495 470 529
rect 404 479 470 495
rect 135 239 151 273
rect 101 205 151 239
rect 199 343 273 359
rect 199 309 215 343
rect 249 309 273 343
rect 199 275 273 309
rect 199 241 215 275
rect 249 241 273 275
rect 199 225 273 241
rect 319 326 329 360
rect 363 326 368 360
rect 319 292 368 326
rect 319 258 329 292
rect 363 258 368 292
rect 319 235 368 258
rect 402 429 511 445
rect 402 395 450 429
rect 484 395 511 429
rect 402 361 511 395
rect 402 327 450 361
rect 484 327 511 361
rect 402 235 511 327
rect 135 191 151 205
rect 135 171 269 191
rect 101 155 269 171
rect 17 105 80 121
rect 17 71 35 105
rect 69 71 80 105
rect 17 55 80 71
rect 114 105 171 121
rect 114 71 121 105
rect 155 71 171 105
rect 114 17 171 71
rect 221 117 269 155
rect 221 83 225 117
rect 259 83 269 117
rect 221 67 269 83
rect 303 167 533 201
rect 303 117 353 167
rect 303 83 311 117
rect 345 83 353 117
rect 303 67 353 83
rect 387 117 441 133
rect 387 83 397 117
rect 431 83 441 117
rect 387 17 441 83
rect 475 117 533 167
rect 475 83 483 117
rect 517 83 533 117
rect 475 67 533 83
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21a_0
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 832866
string GDS_START 825988
<< end >>
