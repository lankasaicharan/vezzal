magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 72 49 671 241
rect 0 0 672 49
<< scnmos >>
rect 151 47 181 215
rect 240 47 270 215
rect 331 47 361 215
rect 445 47 475 215
rect 562 47 592 215
<< scpmoshvt >>
rect 151 367 181 619
rect 242 367 272 619
rect 373 367 403 619
rect 490 367 520 619
rect 562 367 592 619
<< ndiff >>
rect 98 202 151 215
rect 98 168 106 202
rect 140 168 151 202
rect 98 93 151 168
rect 98 59 106 93
rect 140 59 151 93
rect 98 47 151 59
rect 181 47 240 215
rect 270 47 331 215
rect 361 186 445 215
rect 361 152 398 186
rect 432 152 445 186
rect 361 118 445 152
rect 361 84 398 118
rect 432 84 445 118
rect 361 47 445 84
rect 475 126 562 215
rect 475 92 501 126
rect 535 92 562 126
rect 475 47 562 92
rect 592 201 645 215
rect 592 167 603 201
rect 637 167 645 201
rect 592 93 645 167
rect 592 59 603 93
rect 637 59 645 93
rect 592 47 645 59
<< pdiff >>
rect 98 607 151 619
rect 98 573 106 607
rect 140 573 151 607
rect 98 507 151 573
rect 98 473 106 507
rect 140 473 151 507
rect 98 413 151 473
rect 98 379 106 413
rect 140 379 151 413
rect 98 367 151 379
rect 181 599 242 619
rect 181 565 197 599
rect 231 565 242 599
rect 181 501 242 565
rect 181 467 197 501
rect 231 467 242 501
rect 181 413 242 467
rect 181 379 197 413
rect 231 379 242 413
rect 181 367 242 379
rect 272 607 373 619
rect 272 573 308 607
rect 342 573 373 607
rect 272 522 373 573
rect 272 488 308 522
rect 342 488 373 522
rect 272 440 373 488
rect 272 406 308 440
rect 342 406 373 440
rect 272 367 373 406
rect 403 599 490 619
rect 403 565 431 599
rect 465 565 490 599
rect 403 506 490 565
rect 403 472 431 506
rect 465 472 490 506
rect 403 413 490 472
rect 403 379 431 413
rect 465 379 490 413
rect 403 367 490 379
rect 520 367 562 619
rect 592 599 645 619
rect 592 565 603 599
rect 637 565 645 599
rect 592 506 645 565
rect 592 472 603 506
rect 637 472 645 506
rect 592 413 645 472
rect 592 379 603 413
rect 637 379 645 413
rect 592 367 645 379
<< ndiffc >>
rect 106 168 140 202
rect 106 59 140 93
rect 398 152 432 186
rect 398 84 432 118
rect 501 92 535 126
rect 603 167 637 201
rect 603 59 637 93
<< pdiffc >>
rect 106 573 140 607
rect 106 473 140 507
rect 106 379 140 413
rect 197 565 231 599
rect 197 467 231 501
rect 197 379 231 413
rect 308 573 342 607
rect 308 488 342 522
rect 308 406 342 440
rect 431 565 465 599
rect 431 472 465 506
rect 431 379 465 413
rect 603 565 637 599
rect 603 472 637 506
rect 603 379 637 413
<< poly >>
rect 151 619 181 645
rect 242 619 272 645
rect 373 619 403 645
rect 490 619 520 645
rect 562 619 592 645
rect 151 304 181 367
rect 242 304 272 367
rect 373 304 403 367
rect 115 288 181 304
rect 115 254 131 288
rect 165 254 181 288
rect 115 238 181 254
rect 223 288 289 304
rect 223 254 239 288
rect 273 254 289 288
rect 223 238 289 254
rect 331 288 403 304
rect 490 303 520 367
rect 331 254 347 288
rect 381 254 403 288
rect 331 238 403 254
rect 445 287 520 303
rect 445 253 461 287
rect 495 253 520 287
rect 151 215 181 238
rect 240 215 270 238
rect 331 215 361 238
rect 445 237 520 253
rect 562 303 592 367
rect 562 287 647 303
rect 562 253 597 287
rect 631 253 647 287
rect 562 237 647 253
rect 445 215 475 237
rect 562 215 592 237
rect 151 21 181 47
rect 240 21 270 47
rect 331 21 361 47
rect 445 21 475 47
rect 562 21 592 47
<< polycont >>
rect 131 254 165 288
rect 239 254 273 288
rect 347 254 381 288
rect 461 253 495 287
rect 597 253 631 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 90 607 156 649
rect 90 573 106 607
rect 140 573 156 607
rect 90 507 156 573
rect 90 473 106 507
rect 140 473 156 507
rect 90 413 156 473
rect 90 379 106 413
rect 140 379 156 413
rect 90 363 156 379
rect 190 599 247 615
rect 190 565 197 599
rect 231 565 247 599
rect 190 501 247 565
rect 190 467 197 501
rect 231 467 247 501
rect 190 413 247 467
rect 190 379 197 413
rect 231 379 247 413
rect 292 607 358 649
rect 292 573 308 607
rect 342 573 358 607
rect 292 522 358 573
rect 292 488 308 522
rect 342 488 358 522
rect 292 440 358 488
rect 292 406 308 440
rect 342 406 358 440
rect 415 599 481 615
rect 415 565 431 599
rect 465 565 481 599
rect 415 506 481 565
rect 415 472 431 506
rect 465 472 481 506
rect 415 413 481 472
rect 190 372 247 379
rect 415 379 431 413
rect 465 379 481 413
rect 415 372 481 379
rect 594 599 653 615
rect 594 565 603 599
rect 637 565 653 599
rect 594 506 653 565
rect 594 472 603 506
rect 637 472 653 506
rect 594 413 653 472
rect 594 379 603 413
rect 637 379 653 413
rect 594 375 653 379
rect 190 338 481 372
rect 529 341 653 375
rect 17 288 178 304
rect 17 254 131 288
rect 165 254 178 288
rect 17 238 178 254
rect 212 288 275 304
rect 212 254 239 288
rect 273 254 275 288
rect 212 237 275 254
rect 309 288 381 304
rect 309 254 347 288
rect 309 237 381 254
rect 415 287 495 303
rect 415 253 461 287
rect 415 237 495 253
rect 90 202 156 204
rect 529 203 563 341
rect 597 287 647 303
rect 631 253 647 287
rect 597 237 647 253
rect 90 168 106 202
rect 140 168 156 202
rect 90 93 156 168
rect 90 59 106 93
rect 140 59 156 93
rect 90 17 156 59
rect 207 201 653 203
rect 207 186 603 201
rect 207 152 398 186
rect 432 168 603 186
rect 432 152 449 168
rect 207 118 449 152
rect 587 167 603 168
rect 637 167 653 201
rect 207 84 398 118
rect 432 84 449 118
rect 207 51 449 84
rect 485 126 551 134
rect 485 92 501 126
rect 535 92 551 126
rect 485 17 551 92
rect 587 93 653 167
rect 587 59 603 93
rect 637 59 653 93
rect 587 51 653 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a311oi_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3244080
string GDS_START 3237384
<< end >>
