magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
rect 427 303 663 331
<< pwell >>
rect 31 49 1141 157
rect 0 0 1152 49
<< scnmos >>
rect 114 47 144 131
rect 186 47 216 131
rect 272 47 302 131
rect 344 47 374 131
rect 430 47 460 131
rect 502 47 532 131
rect 594 47 624 131
rect 666 47 696 131
rect 752 47 782 131
rect 836 47 866 131
rect 950 47 980 131
rect 1028 47 1058 131
<< scpmoshvt >>
rect 84 409 134 609
rect 302 409 352 609
rect 520 339 570 539
rect 738 409 788 609
rect 836 409 886 609
rect 950 409 1000 609
<< ndiff >>
rect 57 111 114 131
rect 57 77 69 111
rect 103 77 114 111
rect 57 47 114 77
rect 144 47 186 131
rect 216 103 272 131
rect 216 69 227 103
rect 261 69 272 103
rect 216 47 272 69
rect 302 47 344 131
rect 374 111 430 131
rect 374 77 385 111
rect 419 77 430 111
rect 374 47 430 77
rect 460 47 502 131
rect 532 102 594 131
rect 532 68 543 102
rect 577 68 594 102
rect 532 47 594 68
rect 624 47 666 131
rect 696 111 752 131
rect 696 77 707 111
rect 741 77 752 111
rect 696 47 752 77
rect 782 47 836 131
rect 866 103 950 131
rect 866 69 877 103
rect 911 69 950 103
rect 866 47 950 69
rect 980 47 1028 131
rect 1058 108 1115 131
rect 1058 74 1069 108
rect 1103 74 1115 108
rect 1058 47 1115 74
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 191 609
rect 134 563 145 597
rect 179 563 191 597
rect 134 526 191 563
rect 134 492 145 526
rect 179 492 191 526
rect 134 455 191 492
rect 134 421 145 455
rect 179 421 191 455
rect 134 409 191 421
rect 245 597 302 609
rect 245 563 257 597
rect 291 563 302 597
rect 245 526 302 563
rect 245 492 257 526
rect 291 492 302 526
rect 245 455 302 492
rect 245 421 257 455
rect 291 421 302 455
rect 245 409 302 421
rect 352 577 409 609
rect 352 543 363 577
rect 397 543 409 577
rect 681 597 738 609
rect 352 409 409 543
rect 681 563 693 597
rect 727 563 738 597
rect 463 385 520 539
rect 463 351 475 385
rect 509 351 520 385
rect 463 339 520 351
rect 570 527 627 539
rect 570 493 581 527
rect 615 493 627 527
rect 570 455 627 493
rect 570 421 581 455
rect 615 421 627 455
rect 570 339 627 421
rect 681 526 738 563
rect 681 492 693 526
rect 727 492 738 526
rect 681 455 738 492
rect 681 421 693 455
rect 727 421 738 455
rect 681 409 738 421
rect 788 409 836 609
rect 886 597 950 609
rect 886 563 897 597
rect 931 563 950 597
rect 886 526 950 563
rect 886 492 897 526
rect 931 492 950 526
rect 886 455 950 492
rect 886 421 897 455
rect 931 421 950 455
rect 886 409 950 421
rect 1000 597 1057 609
rect 1000 563 1011 597
rect 1045 563 1057 597
rect 1000 526 1057 563
rect 1000 492 1011 526
rect 1045 492 1057 526
rect 1000 455 1057 492
rect 1000 421 1011 455
rect 1045 421 1057 455
rect 1000 409 1057 421
<< ndiffc >>
rect 69 77 103 111
rect 227 69 261 103
rect 385 77 419 111
rect 543 68 577 102
rect 707 77 741 111
rect 877 69 911 103
rect 1069 74 1103 108
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 492 179 526
rect 145 421 179 455
rect 257 563 291 597
rect 257 492 291 526
rect 257 421 291 455
rect 363 543 397 577
rect 693 563 727 597
rect 475 351 509 385
rect 581 493 615 527
rect 581 421 615 455
rect 693 492 727 526
rect 693 421 727 455
rect 897 563 931 597
rect 897 492 931 526
rect 897 421 931 455
rect 1011 563 1045 597
rect 1011 492 1045 526
rect 1011 421 1045 455
<< poly >>
rect 84 609 134 635
rect 302 609 352 635
rect 738 609 788 635
rect 836 609 886 635
rect 950 609 1000 635
rect 520 539 570 565
rect 84 369 134 409
rect 84 353 159 369
rect 302 358 352 409
rect 84 319 109 353
rect 143 319 159 353
rect 84 285 159 319
rect 84 251 109 285
rect 143 251 159 285
rect 84 235 159 251
rect 211 342 374 358
rect 211 308 227 342
rect 261 308 374 342
rect 211 274 374 308
rect 520 299 570 339
rect 738 299 788 409
rect 211 240 227 274
rect 261 240 374 274
rect 502 283 570 299
rect 502 263 520 283
rect 114 176 144 235
rect 211 224 374 240
rect 114 146 216 176
rect 114 131 144 146
rect 186 131 216 146
rect 272 131 302 224
rect 344 131 374 224
rect 430 249 520 263
rect 554 249 570 283
rect 430 233 570 249
rect 666 283 788 299
rect 666 249 693 283
rect 727 249 788 283
rect 666 233 788 249
rect 836 299 886 409
rect 950 299 1000 409
rect 836 283 902 299
rect 836 249 852 283
rect 886 249 902 283
rect 430 131 460 233
rect 502 131 532 233
rect 666 176 696 233
rect 836 215 902 249
rect 836 181 852 215
rect 886 181 902 215
rect 836 176 902 181
rect 594 146 696 176
rect 594 131 624 146
rect 666 131 696 146
rect 752 165 902 176
rect 950 283 1058 299
rect 950 249 987 283
rect 1021 249 1058 283
rect 950 215 1058 249
rect 950 181 987 215
rect 1021 181 1058 215
rect 950 165 1058 181
rect 752 146 866 165
rect 752 131 782 146
rect 836 131 866 146
rect 950 131 980 165
rect 1028 131 1058 165
rect 114 21 144 47
rect 186 21 216 47
rect 272 21 302 47
rect 344 21 374 47
rect 430 21 460 47
rect 502 21 532 47
rect 594 21 624 47
rect 666 21 696 47
rect 752 21 782 47
rect 836 21 866 47
rect 950 21 980 47
rect 1028 21 1058 47
<< polycont >>
rect 109 319 143 353
rect 109 251 143 285
rect 227 308 261 342
rect 227 240 261 274
rect 520 249 554 283
rect 693 249 727 283
rect 852 249 886 283
rect 852 181 886 215
rect 987 249 1021 283
rect 987 181 1021 215
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 597 73 613
rect 23 563 39 597
rect 23 526 73 563
rect 23 492 39 526
rect 23 455 73 492
rect 23 421 39 455
rect 23 405 73 421
rect 129 597 195 649
rect 129 563 145 597
rect 179 563 195 597
rect 129 526 195 563
rect 129 492 145 526
rect 179 492 195 526
rect 129 455 195 492
rect 129 421 145 455
rect 179 421 195 455
rect 129 405 195 421
rect 241 597 307 613
rect 241 563 257 597
rect 291 563 307 597
rect 241 526 307 563
rect 241 492 257 526
rect 291 492 307 526
rect 347 597 743 613
rect 347 579 693 597
rect 347 577 413 579
rect 347 543 363 577
rect 397 543 413 577
rect 677 563 693 579
rect 727 563 743 597
rect 347 507 413 543
rect 565 527 631 543
rect 241 471 307 492
rect 565 493 581 527
rect 615 493 631 527
rect 565 471 631 493
rect 241 455 631 471
rect 241 421 257 455
rect 291 437 581 455
rect 291 421 307 437
rect 241 405 307 421
rect 565 421 581 437
rect 615 421 631 455
rect 565 405 631 421
rect 677 526 743 563
rect 677 492 693 526
rect 727 492 743 526
rect 677 455 743 492
rect 677 421 693 455
rect 727 421 743 455
rect 677 405 743 421
rect 881 597 947 649
rect 881 563 897 597
rect 931 563 947 597
rect 881 526 947 563
rect 881 492 897 526
rect 931 492 947 526
rect 881 455 947 492
rect 881 421 897 455
rect 931 421 947 455
rect 881 405 947 421
rect 995 597 1119 613
rect 995 563 1011 597
rect 1045 563 1119 597
rect 995 526 1119 563
rect 995 492 1011 526
rect 1045 492 1119 526
rect 995 455 1119 492
rect 995 421 1011 455
rect 1045 421 1119 455
rect 23 199 57 405
rect 421 385 525 401
rect 93 353 167 369
rect 93 319 109 353
rect 143 319 167 353
rect 93 285 167 319
rect 93 251 109 285
rect 143 251 167 285
rect 93 235 167 251
rect 211 342 277 358
rect 421 356 475 385
rect 211 308 227 342
rect 261 308 277 342
rect 211 274 277 308
rect 211 240 227 274
rect 261 240 277 274
rect 211 199 277 240
rect 23 165 277 199
rect 313 351 475 356
rect 509 351 525 385
rect 995 369 1119 421
rect 313 335 525 351
rect 561 335 1119 369
rect 313 197 455 335
rect 561 299 595 335
rect 504 283 595 299
rect 504 249 520 283
rect 554 249 595 283
rect 504 233 595 249
rect 677 283 743 299
rect 677 249 693 283
rect 727 249 743 283
rect 677 233 743 249
rect 793 283 935 299
rect 793 249 852 283
rect 886 249 935 283
rect 793 215 935 249
rect 23 111 119 165
rect 313 163 757 197
rect 793 181 852 215
rect 886 181 935 215
rect 793 165 935 181
rect 971 283 1037 299
rect 971 249 987 283
rect 1021 249 1037 283
rect 971 215 1037 249
rect 971 181 987 215
rect 1021 181 1037 215
rect 971 165 1037 181
rect 23 77 69 111
rect 103 77 119 111
rect 23 53 119 77
rect 211 103 277 129
rect 211 69 227 103
rect 261 69 277 103
rect 211 17 277 69
rect 313 111 435 163
rect 313 77 385 111
rect 419 77 435 111
rect 313 53 435 77
rect 527 102 593 127
rect 527 68 543 102
rect 577 68 593 102
rect 527 17 593 68
rect 691 111 757 163
rect 1085 129 1119 335
rect 691 77 707 111
rect 741 77 757 111
rect 691 53 757 77
rect 861 103 927 129
rect 861 69 877 103
rect 911 69 927 103
rect 861 17 927 69
rect 1053 108 1119 129
rect 1053 74 1069 108
rect 1103 74 1119 108
rect 1053 53 1119 74
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4bb_lp
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3385604
string GDS_START 3376322
<< end >>
