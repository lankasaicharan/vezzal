magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 37 241 839 259
rect 37 49 1631 241
rect 0 0 1632 49
<< scnmos >>
rect 116 65 146 233
rect 202 65 232 233
rect 288 65 318 233
rect 374 65 404 233
rect 472 65 502 233
rect 558 65 588 233
rect 644 65 674 233
rect 730 65 760 233
rect 920 47 950 215
rect 1006 47 1036 215
rect 1092 47 1122 215
rect 1178 47 1208 215
rect 1264 47 1294 215
rect 1350 47 1380 215
rect 1436 47 1466 215
rect 1522 47 1552 215
<< scpmoshvt >>
rect 142 367 172 619
rect 228 367 258 619
rect 314 367 344 619
rect 400 367 430 619
rect 486 367 516 619
rect 572 367 602 619
rect 674 367 704 619
rect 760 367 790 619
rect 867 367 897 619
rect 953 367 983 619
rect 1039 367 1069 619
rect 1134 367 1164 619
rect 1220 367 1250 619
rect 1306 367 1336 619
rect 1392 367 1422 619
rect 1478 367 1508 619
<< ndiff >>
rect 63 192 116 233
rect 63 158 71 192
rect 105 158 116 192
rect 63 113 116 158
rect 63 79 71 113
rect 105 79 116 113
rect 63 65 116 79
rect 146 132 202 233
rect 146 98 157 132
rect 191 98 202 132
rect 146 65 202 98
rect 232 192 288 233
rect 232 158 243 192
rect 277 158 288 192
rect 232 113 288 158
rect 232 79 243 113
rect 277 79 288 113
rect 232 65 288 79
rect 318 132 374 233
rect 318 98 329 132
rect 363 98 374 132
rect 318 65 374 98
rect 404 190 472 233
rect 404 156 415 190
rect 449 156 472 190
rect 404 111 472 156
rect 404 77 415 111
rect 449 77 472 111
rect 404 65 472 77
rect 502 225 558 233
rect 502 191 513 225
rect 547 191 558 225
rect 502 157 558 191
rect 502 123 513 157
rect 547 123 558 157
rect 502 65 558 123
rect 588 111 644 233
rect 588 77 599 111
rect 633 77 644 111
rect 588 65 644 77
rect 674 201 730 233
rect 674 167 685 201
rect 719 167 730 201
rect 674 65 730 167
rect 760 111 813 233
rect 760 77 771 111
rect 805 77 813 111
rect 760 65 813 77
rect 867 93 920 215
rect 867 59 875 93
rect 909 59 920 93
rect 867 47 920 59
rect 950 201 1006 215
rect 950 167 961 201
rect 995 167 1006 201
rect 950 47 1006 167
rect 1036 93 1092 215
rect 1036 59 1047 93
rect 1081 59 1092 93
rect 1036 47 1092 59
rect 1122 189 1178 215
rect 1122 155 1133 189
rect 1167 155 1178 189
rect 1122 47 1178 155
rect 1208 192 1264 215
rect 1208 158 1219 192
rect 1253 158 1264 192
rect 1208 105 1264 158
rect 1208 71 1219 105
rect 1253 71 1264 105
rect 1208 47 1264 71
rect 1294 113 1350 215
rect 1294 79 1305 113
rect 1339 79 1350 113
rect 1294 47 1350 79
rect 1380 203 1436 215
rect 1380 169 1391 203
rect 1425 169 1436 203
rect 1380 101 1436 169
rect 1380 67 1391 101
rect 1425 67 1436 101
rect 1380 47 1436 67
rect 1466 175 1522 215
rect 1466 141 1477 175
rect 1511 141 1522 175
rect 1466 93 1522 141
rect 1466 59 1477 93
rect 1511 59 1522 93
rect 1466 47 1522 59
rect 1552 203 1605 215
rect 1552 169 1563 203
rect 1597 169 1605 203
rect 1552 101 1605 169
rect 1552 67 1563 101
rect 1597 67 1605 101
rect 1552 47 1605 67
<< pdiff >>
rect 89 599 142 619
rect 89 565 97 599
rect 131 565 142 599
rect 89 507 142 565
rect 89 473 97 507
rect 131 473 142 507
rect 89 415 142 473
rect 89 381 97 415
rect 131 381 142 415
rect 89 367 142 381
rect 172 538 228 619
rect 172 504 183 538
rect 217 504 228 538
rect 172 413 228 504
rect 172 379 183 413
rect 217 379 228 413
rect 172 367 228 379
rect 258 599 314 619
rect 258 565 269 599
rect 303 565 314 599
rect 258 529 314 565
rect 258 495 269 529
rect 303 495 314 529
rect 258 459 314 495
rect 258 425 269 459
rect 303 425 314 459
rect 258 367 314 425
rect 344 538 400 619
rect 344 504 355 538
rect 389 504 400 538
rect 344 413 400 504
rect 344 379 355 413
rect 389 379 400 413
rect 344 367 400 379
rect 430 597 486 619
rect 430 563 441 597
rect 475 563 486 597
rect 430 529 486 563
rect 430 495 441 529
rect 475 495 486 529
rect 430 459 486 495
rect 430 425 441 459
rect 475 425 486 459
rect 430 367 486 425
rect 516 538 572 619
rect 516 504 527 538
rect 561 504 572 538
rect 516 413 572 504
rect 516 379 527 413
rect 561 379 572 413
rect 516 367 572 379
rect 602 597 674 619
rect 602 563 623 597
rect 657 563 674 597
rect 602 529 674 563
rect 602 495 623 529
rect 657 495 674 529
rect 602 459 674 495
rect 602 425 623 459
rect 657 425 674 459
rect 602 367 674 425
rect 704 538 760 619
rect 704 504 715 538
rect 749 504 760 538
rect 704 413 760 504
rect 704 379 715 413
rect 749 379 760 413
rect 704 367 760 379
rect 790 599 867 619
rect 790 565 811 599
rect 845 565 867 599
rect 790 509 867 565
rect 790 475 811 509
rect 845 475 867 509
rect 790 413 867 475
rect 790 379 811 413
rect 845 379 867 413
rect 790 367 867 379
rect 897 607 953 619
rect 897 573 908 607
rect 942 573 953 607
rect 897 528 953 573
rect 897 494 908 528
rect 942 494 953 528
rect 897 453 953 494
rect 897 419 908 453
rect 942 419 953 453
rect 897 367 953 419
rect 983 599 1039 619
rect 983 565 994 599
rect 1028 565 1039 599
rect 983 509 1039 565
rect 983 475 994 509
rect 1028 475 1039 509
rect 983 413 1039 475
rect 983 379 994 413
rect 1028 379 1039 413
rect 983 367 1039 379
rect 1069 607 1134 619
rect 1069 573 1080 607
rect 1114 573 1134 607
rect 1069 528 1134 573
rect 1069 494 1080 528
rect 1114 494 1134 528
rect 1069 453 1134 494
rect 1069 419 1080 453
rect 1114 419 1134 453
rect 1069 367 1134 419
rect 1164 599 1220 619
rect 1164 565 1175 599
rect 1209 565 1220 599
rect 1164 509 1220 565
rect 1164 475 1175 509
rect 1209 475 1220 509
rect 1164 413 1220 475
rect 1164 379 1175 413
rect 1209 379 1220 413
rect 1164 367 1220 379
rect 1250 607 1306 619
rect 1250 573 1261 607
rect 1295 573 1306 607
rect 1250 494 1306 573
rect 1250 460 1261 494
rect 1295 460 1306 494
rect 1250 367 1306 460
rect 1336 599 1392 619
rect 1336 565 1347 599
rect 1381 565 1392 599
rect 1336 516 1392 565
rect 1336 482 1347 516
rect 1381 482 1392 516
rect 1336 436 1392 482
rect 1336 402 1347 436
rect 1381 402 1392 436
rect 1336 367 1392 402
rect 1422 607 1478 619
rect 1422 573 1433 607
rect 1467 573 1478 607
rect 1422 494 1478 573
rect 1422 460 1433 494
rect 1467 460 1478 494
rect 1422 367 1478 460
rect 1508 599 1561 619
rect 1508 565 1519 599
rect 1553 565 1561 599
rect 1508 516 1561 565
rect 1508 482 1519 516
rect 1553 482 1561 516
rect 1508 436 1561 482
rect 1508 402 1519 436
rect 1553 402 1561 436
rect 1508 367 1561 402
<< ndiffc >>
rect 71 158 105 192
rect 71 79 105 113
rect 157 98 191 132
rect 243 158 277 192
rect 243 79 277 113
rect 329 98 363 132
rect 415 156 449 190
rect 415 77 449 111
rect 513 191 547 225
rect 513 123 547 157
rect 599 77 633 111
rect 685 167 719 201
rect 771 77 805 111
rect 875 59 909 93
rect 961 167 995 201
rect 1047 59 1081 93
rect 1133 155 1167 189
rect 1219 158 1253 192
rect 1219 71 1253 105
rect 1305 79 1339 113
rect 1391 169 1425 203
rect 1391 67 1425 101
rect 1477 141 1511 175
rect 1477 59 1511 93
rect 1563 169 1597 203
rect 1563 67 1597 101
<< pdiffc >>
rect 97 565 131 599
rect 97 473 131 507
rect 97 381 131 415
rect 183 504 217 538
rect 183 379 217 413
rect 269 565 303 599
rect 269 495 303 529
rect 269 425 303 459
rect 355 504 389 538
rect 355 379 389 413
rect 441 563 475 597
rect 441 495 475 529
rect 441 425 475 459
rect 527 504 561 538
rect 527 379 561 413
rect 623 563 657 597
rect 623 495 657 529
rect 623 425 657 459
rect 715 504 749 538
rect 715 379 749 413
rect 811 565 845 599
rect 811 475 845 509
rect 811 379 845 413
rect 908 573 942 607
rect 908 494 942 528
rect 908 419 942 453
rect 994 565 1028 599
rect 994 475 1028 509
rect 994 379 1028 413
rect 1080 573 1114 607
rect 1080 494 1114 528
rect 1080 419 1114 453
rect 1175 565 1209 599
rect 1175 475 1209 509
rect 1175 379 1209 413
rect 1261 573 1295 607
rect 1261 460 1295 494
rect 1347 565 1381 599
rect 1347 482 1381 516
rect 1347 402 1381 436
rect 1433 573 1467 607
rect 1433 460 1467 494
rect 1519 565 1553 599
rect 1519 482 1553 516
rect 1519 402 1553 436
<< poly >>
rect 142 619 172 645
rect 228 619 258 645
rect 314 619 344 645
rect 400 619 430 645
rect 486 619 516 645
rect 572 619 602 645
rect 674 619 704 645
rect 760 619 790 645
rect 867 619 897 645
rect 953 619 983 645
rect 1039 619 1069 645
rect 1134 619 1164 645
rect 1220 619 1250 645
rect 1306 619 1336 645
rect 1392 619 1422 645
rect 1478 619 1508 645
rect 142 321 172 367
rect 228 321 258 367
rect 314 321 344 367
rect 400 321 430 367
rect 24 305 430 321
rect 24 271 40 305
rect 74 271 108 305
rect 142 271 176 305
rect 210 271 244 305
rect 278 271 312 305
rect 346 271 380 305
rect 414 271 430 305
rect 486 321 516 367
rect 572 321 602 367
rect 674 321 704 367
rect 760 321 790 367
rect 486 305 825 321
rect 486 285 571 305
rect 24 255 430 271
rect 472 271 571 285
rect 605 271 639 305
rect 673 271 707 305
rect 741 271 775 305
rect 809 271 825 305
rect 472 255 825 271
rect 867 303 897 367
rect 953 303 983 367
rect 1039 303 1069 367
rect 1134 303 1164 367
rect 1220 345 1250 367
rect 1306 345 1336 367
rect 1392 345 1422 367
rect 1478 345 1508 367
rect 1220 319 1552 345
rect 1220 315 1366 319
rect 867 287 1178 303
rect 116 233 146 255
rect 202 233 232 255
rect 288 233 318 255
rect 374 233 404 255
rect 472 233 502 255
rect 558 233 588 255
rect 644 233 674 255
rect 730 233 760 255
rect 867 253 992 287
rect 1026 253 1060 287
rect 1094 253 1128 287
rect 1162 267 1178 287
rect 1264 285 1366 315
rect 1400 285 1434 319
rect 1468 285 1502 319
rect 1536 285 1552 319
rect 1264 269 1552 285
rect 1162 253 1208 267
rect 867 237 1208 253
rect 920 215 950 237
rect 1006 215 1036 237
rect 1092 215 1122 237
rect 1178 215 1208 237
rect 1264 215 1294 269
rect 1350 215 1380 269
rect 1436 215 1466 269
rect 1522 215 1552 269
rect 116 39 146 65
rect 202 39 232 65
rect 288 39 318 65
rect 374 39 404 65
rect 472 39 502 65
rect 558 39 588 65
rect 644 39 674 65
rect 730 39 760 65
rect 920 21 950 47
rect 1006 21 1036 47
rect 1092 21 1122 47
rect 1178 21 1208 47
rect 1264 21 1294 47
rect 1350 21 1380 47
rect 1436 21 1466 47
rect 1522 21 1552 47
<< polycont >>
rect 40 271 74 305
rect 108 271 142 305
rect 176 271 210 305
rect 244 271 278 305
rect 312 271 346 305
rect 380 271 414 305
rect 571 271 605 305
rect 639 271 673 305
rect 707 271 741 305
rect 775 271 809 305
rect 992 253 1026 287
rect 1060 253 1094 287
rect 1128 253 1162 287
rect 1366 285 1400 319
rect 1434 285 1468 319
rect 1502 285 1536 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 81 599 858 615
rect 81 565 97 599
rect 131 581 269 599
rect 131 565 133 581
rect 81 507 133 565
rect 267 565 269 581
rect 303 597 811 599
rect 303 581 441 597
rect 303 565 305 581
rect 81 473 97 507
rect 131 473 133 507
rect 81 415 133 473
rect 81 381 97 415
rect 131 381 133 415
rect 81 365 133 381
rect 167 538 233 547
rect 167 504 183 538
rect 217 504 233 538
rect 167 413 233 504
rect 167 379 183 413
rect 217 379 233 413
rect 267 529 305 565
rect 439 563 441 581
rect 475 581 623 597
rect 475 563 477 581
rect 267 495 269 529
rect 303 495 305 529
rect 267 459 305 495
rect 267 425 269 459
rect 303 425 305 459
rect 267 409 305 425
rect 339 538 405 547
rect 339 504 355 538
rect 389 504 405 538
rect 339 413 405 504
rect 167 375 233 379
rect 339 379 355 413
rect 389 379 405 413
rect 439 529 477 563
rect 611 563 623 581
rect 657 581 811 597
rect 657 563 665 581
rect 439 495 441 529
rect 475 495 477 529
rect 439 459 477 495
rect 439 425 441 459
rect 475 425 477 459
rect 439 409 477 425
rect 511 538 577 547
rect 511 504 527 538
rect 561 504 577 538
rect 511 413 577 504
rect 339 375 405 379
rect 511 379 527 413
rect 561 379 577 413
rect 611 529 665 563
rect 799 565 811 581
rect 845 565 858 599
rect 611 495 623 529
rect 657 495 665 529
rect 611 459 665 495
rect 611 425 623 459
rect 657 425 665 459
rect 611 409 665 425
rect 699 538 765 547
rect 699 504 715 538
rect 749 504 765 538
rect 699 413 765 504
rect 511 375 577 379
rect 699 379 715 413
rect 749 379 765 413
rect 699 375 765 379
rect 167 341 765 375
rect 799 509 858 565
rect 799 475 811 509
rect 845 475 858 509
rect 799 413 858 475
rect 892 607 958 649
rect 892 573 908 607
rect 942 573 958 607
rect 892 528 958 573
rect 892 494 908 528
rect 942 494 958 528
rect 892 453 958 494
rect 892 419 908 453
rect 942 419 958 453
rect 992 599 1030 615
rect 992 565 994 599
rect 1028 565 1030 599
rect 992 509 1030 565
rect 992 475 994 509
rect 1028 475 1030 509
rect 799 379 811 413
rect 845 385 858 413
rect 992 413 1030 475
rect 1064 607 1130 649
rect 1064 573 1080 607
rect 1114 573 1130 607
rect 1064 528 1130 573
rect 1064 494 1080 528
rect 1114 494 1130 528
rect 1064 453 1130 494
rect 1064 419 1080 453
rect 1114 419 1130 453
rect 1164 599 1211 615
rect 1164 565 1175 599
rect 1209 565 1211 599
rect 1164 509 1211 565
rect 1164 475 1175 509
rect 1209 475 1211 509
rect 1164 420 1211 475
rect 1245 607 1311 649
rect 1245 573 1261 607
rect 1295 573 1311 607
rect 1245 494 1311 573
rect 1245 460 1261 494
rect 1295 460 1311 494
rect 1245 454 1311 460
rect 1345 599 1383 615
rect 1345 565 1347 599
rect 1381 565 1383 599
rect 1345 516 1383 565
rect 1345 482 1347 516
rect 1381 482 1383 516
rect 1345 436 1383 482
rect 1417 607 1483 649
rect 1417 573 1433 607
rect 1467 573 1483 607
rect 1417 494 1483 573
rect 1417 460 1433 494
rect 1467 460 1483 494
rect 1417 454 1483 460
rect 1517 599 1569 615
rect 1517 565 1519 599
rect 1553 565 1569 599
rect 1517 516 1569 565
rect 1517 482 1519 516
rect 1553 482 1569 516
rect 1345 420 1347 436
rect 992 385 994 413
rect 845 379 994 385
rect 1028 385 1030 413
rect 1164 413 1347 420
rect 1164 385 1175 413
rect 1028 379 1175 385
rect 1209 402 1347 413
rect 1381 420 1383 436
rect 1517 436 1569 482
rect 1517 420 1519 436
rect 1381 402 1519 420
rect 1553 402 1569 436
rect 1209 386 1569 402
rect 799 351 1209 379
rect 24 271 40 305
rect 74 271 108 305
rect 142 271 176 305
rect 210 271 244 305
rect 278 271 312 305
rect 346 271 380 305
rect 414 271 449 305
rect 24 242 449 271
rect 485 229 519 341
rect 1350 319 1601 352
rect 555 271 571 305
rect 605 271 639 305
rect 673 271 707 305
rect 741 271 775 305
rect 809 271 929 305
rect 597 242 929 271
rect 976 253 992 287
rect 1026 253 1060 287
rect 1094 253 1128 287
rect 1162 253 1316 287
rect 1350 285 1366 319
rect 1400 285 1434 319
rect 1468 285 1502 319
rect 1536 285 1601 319
rect 976 242 1316 253
rect 485 225 563 229
rect 55 192 449 208
rect 55 158 71 192
rect 105 174 243 192
rect 105 158 107 174
rect 55 113 107 158
rect 241 158 243 174
rect 277 190 449 192
rect 277 174 415 190
rect 277 158 279 174
rect 55 79 71 113
rect 105 79 107 113
rect 55 63 107 79
rect 141 132 207 140
rect 141 98 157 132
rect 191 98 207 132
rect 141 17 207 98
rect 241 113 279 158
rect 413 156 415 174
rect 241 79 243 113
rect 277 79 279 113
rect 241 63 279 79
rect 313 132 379 140
rect 313 98 329 132
rect 363 98 379 132
rect 313 17 379 98
rect 413 111 449 156
rect 485 191 513 225
rect 547 208 563 225
rect 1371 213 1613 251
rect 1371 208 1427 213
rect 547 201 1169 208
rect 547 191 685 201
rect 485 167 685 191
rect 719 167 961 201
rect 995 189 1169 201
rect 995 167 1133 189
rect 485 163 1133 167
rect 485 157 563 163
rect 485 123 513 157
rect 547 123 563 157
rect 1129 155 1133 163
rect 1167 155 1169 189
rect 1129 139 1169 155
rect 1203 203 1427 208
rect 1203 192 1391 203
rect 1203 158 1219 192
rect 1253 169 1391 192
rect 1425 169 1427 203
rect 1561 203 1613 213
rect 1253 158 1427 169
rect 1203 155 1427 158
rect 485 119 563 123
rect 413 77 415 111
rect 599 111 809 127
rect 449 77 599 85
rect 633 77 771 111
rect 805 77 809 111
rect 1203 105 1255 155
rect 413 51 809 77
rect 859 93 1219 105
rect 859 59 875 93
rect 909 59 1047 93
rect 1081 71 1219 93
rect 1253 71 1255 105
rect 1081 59 1255 71
rect 859 55 1255 59
rect 1289 113 1355 121
rect 1289 79 1305 113
rect 1339 79 1355 113
rect 1289 17 1355 79
rect 1389 101 1427 155
rect 1389 67 1391 101
rect 1425 67 1427 101
rect 1389 51 1427 67
rect 1461 175 1527 179
rect 1461 141 1477 175
rect 1511 141 1527 175
rect 1461 93 1527 141
rect 1461 59 1477 93
rect 1511 59 1527 93
rect 1461 17 1527 59
rect 1561 169 1563 203
rect 1597 169 1613 203
rect 1561 101 1613 169
rect 1561 67 1563 101
rect 1597 67 1613 101
rect 1561 51 1613 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a22oi_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 437958
string GDS_START 423362
<< end >>
