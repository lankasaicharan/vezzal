magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 23 243 297 273
rect 23 49 940 243
rect 0 0 960 49
<< scnmos >>
rect 102 79 132 247
rect 188 79 218 247
rect 435 49 465 217
rect 530 49 560 217
rect 637 49 667 217
rect 723 49 753 217
rect 831 49 861 217
<< scpmoshvt >>
rect 102 367 132 619
rect 188 367 218 619
rect 389 367 419 619
rect 543 367 573 619
rect 615 367 645 619
rect 723 367 753 619
rect 831 367 861 619
<< ndiff >>
rect 49 235 102 247
rect 49 201 57 235
rect 91 201 102 235
rect 49 125 102 201
rect 49 91 57 125
rect 91 91 102 125
rect 49 79 102 91
rect 132 235 188 247
rect 132 201 143 235
rect 177 201 188 235
rect 132 125 188 201
rect 132 91 143 125
rect 177 91 188 125
rect 132 79 188 91
rect 218 235 271 247
rect 218 201 229 235
rect 263 201 271 235
rect 218 125 271 201
rect 218 91 229 125
rect 263 91 271 125
rect 218 79 271 91
rect 382 205 435 217
rect 382 171 390 205
rect 424 171 435 205
rect 382 95 435 171
rect 382 61 390 95
rect 424 61 435 95
rect 382 49 435 61
rect 465 205 530 217
rect 465 171 485 205
rect 519 171 530 205
rect 465 101 530 171
rect 465 67 485 101
rect 519 67 530 101
rect 465 49 530 67
rect 560 167 637 217
rect 560 133 582 167
rect 616 133 637 167
rect 560 91 637 133
rect 560 57 582 91
rect 616 57 637 91
rect 560 49 637 57
rect 667 205 723 217
rect 667 171 678 205
rect 712 171 723 205
rect 667 101 723 171
rect 667 67 678 101
rect 712 67 723 101
rect 667 49 723 67
rect 753 167 831 217
rect 753 133 776 167
rect 810 133 831 167
rect 753 91 831 133
rect 753 57 776 91
rect 810 57 831 91
rect 753 49 831 57
rect 861 205 914 217
rect 861 171 872 205
rect 906 171 914 205
rect 861 101 914 171
rect 861 67 872 101
rect 906 67 914 101
rect 861 49 914 67
<< pdiff >>
rect 49 607 102 619
rect 49 573 57 607
rect 91 573 102 607
rect 49 512 102 573
rect 49 478 57 512
rect 91 478 102 512
rect 49 413 102 478
rect 49 379 57 413
rect 91 379 102 413
rect 49 367 102 379
rect 132 599 188 619
rect 132 565 143 599
rect 177 565 188 599
rect 132 509 188 565
rect 132 475 143 509
rect 177 475 188 509
rect 132 413 188 475
rect 132 379 143 413
rect 177 379 188 413
rect 132 367 188 379
rect 218 607 389 619
rect 218 573 229 607
rect 263 573 344 607
rect 378 573 389 607
rect 218 512 389 573
rect 218 478 229 512
rect 263 478 344 512
rect 378 478 389 512
rect 218 413 389 478
rect 218 379 229 413
rect 263 379 389 413
rect 218 367 389 379
rect 419 607 543 619
rect 419 573 430 607
rect 464 573 498 607
rect 532 573 543 607
rect 419 516 543 573
rect 419 482 430 516
rect 464 482 498 516
rect 532 482 543 516
rect 419 442 543 482
rect 419 408 430 442
rect 464 408 543 442
rect 419 367 543 408
rect 573 367 615 619
rect 645 367 723 619
rect 753 367 831 619
rect 861 607 915 619
rect 861 573 873 607
rect 907 573 915 607
rect 861 519 915 573
rect 861 485 873 519
rect 907 485 915 519
rect 861 435 915 485
rect 861 401 873 435
rect 907 401 915 435
rect 861 367 915 401
<< ndiffc >>
rect 57 201 91 235
rect 57 91 91 125
rect 143 201 177 235
rect 143 91 177 125
rect 229 201 263 235
rect 229 91 263 125
rect 390 171 424 205
rect 390 61 424 95
rect 485 171 519 205
rect 485 67 519 101
rect 582 133 616 167
rect 582 57 616 91
rect 678 171 712 205
rect 678 67 712 101
rect 776 133 810 167
rect 776 57 810 91
rect 872 171 906 205
rect 872 67 906 101
<< pdiffc >>
rect 57 573 91 607
rect 57 478 91 512
rect 57 379 91 413
rect 143 565 177 599
rect 143 475 177 509
rect 143 379 177 413
rect 229 573 263 607
rect 344 573 378 607
rect 229 478 263 512
rect 344 478 378 512
rect 229 379 263 413
rect 430 573 464 607
rect 498 573 532 607
rect 430 482 464 516
rect 498 482 532 516
rect 430 408 464 442
rect 873 573 907 607
rect 873 485 907 519
rect 873 401 907 435
<< poly >>
rect 102 619 132 645
rect 188 619 218 645
rect 389 619 419 645
rect 543 619 573 645
rect 615 619 645 645
rect 723 619 753 645
rect 831 619 861 645
rect 102 335 132 367
rect 188 335 218 367
rect 102 319 332 335
rect 102 285 214 319
rect 248 285 282 319
rect 316 285 332 319
rect 102 269 332 285
rect 389 308 419 367
rect 543 335 573 367
rect 507 319 573 335
rect 389 292 465 308
rect 102 247 132 269
rect 188 247 218 269
rect 389 258 415 292
rect 449 258 465 292
rect 507 285 523 319
rect 557 285 573 319
rect 507 269 573 285
rect 615 335 645 367
rect 723 335 753 367
rect 615 319 681 335
rect 615 285 631 319
rect 665 285 681 319
rect 615 269 681 285
rect 723 319 789 335
rect 723 285 739 319
rect 773 285 789 319
rect 723 269 789 285
rect 831 325 861 367
rect 831 309 935 325
rect 831 275 885 309
rect 919 275 935 309
rect 389 242 465 258
rect 435 217 465 242
rect 530 217 560 269
rect 637 217 667 269
rect 723 217 753 269
rect 831 259 935 275
rect 831 217 861 259
rect 102 53 132 79
rect 188 53 218 79
rect 435 23 465 49
rect 530 23 560 49
rect 637 23 667 49
rect 723 23 753 49
rect 831 23 861 49
<< polycont >>
rect 214 285 248 319
rect 282 285 316 319
rect 415 258 449 292
rect 523 285 557 319
rect 631 285 665 319
rect 739 285 773 319
rect 885 275 919 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 41 607 93 649
rect 41 573 57 607
rect 91 573 93 607
rect 41 512 93 573
rect 41 478 57 512
rect 91 478 93 512
rect 41 413 93 478
rect 41 379 57 413
rect 91 379 93 413
rect 41 363 93 379
rect 127 599 179 615
rect 127 565 143 599
rect 177 565 179 599
rect 127 509 179 565
rect 127 475 143 509
rect 177 475 179 509
rect 127 413 179 475
rect 127 379 143 413
rect 177 379 179 413
rect 41 235 93 251
rect 41 201 57 235
rect 91 201 93 235
rect 41 125 93 201
rect 41 91 57 125
rect 91 91 93 125
rect 41 17 93 91
rect 127 235 179 379
rect 213 607 380 649
rect 213 573 229 607
rect 263 573 344 607
rect 378 573 380 607
rect 213 512 380 573
rect 213 478 229 512
rect 263 478 344 512
rect 378 478 380 512
rect 213 462 380 478
rect 414 607 548 615
rect 414 573 430 607
rect 464 573 498 607
rect 532 573 548 607
rect 869 607 923 649
rect 414 516 548 573
rect 414 482 430 516
rect 464 482 498 516
rect 532 482 548 516
rect 414 466 548 482
rect 213 413 290 462
rect 414 442 465 466
rect 414 428 430 442
rect 213 379 229 413
rect 263 379 290 413
rect 213 369 290 379
rect 324 408 430 428
rect 464 408 465 442
rect 324 392 465 408
rect 324 335 379 392
rect 213 319 379 335
rect 213 285 214 319
rect 248 285 282 319
rect 316 285 379 319
rect 213 269 379 285
rect 127 201 143 235
rect 177 201 179 235
rect 127 125 179 201
rect 127 91 143 125
rect 177 91 179 125
rect 127 75 179 91
rect 213 201 229 235
rect 263 201 279 235
rect 213 125 279 201
rect 213 91 229 125
rect 263 91 279 125
rect 213 17 279 91
rect 324 208 379 269
rect 413 292 451 350
rect 413 258 415 292
rect 449 258 451 292
rect 499 319 563 432
rect 499 285 523 319
rect 557 285 563 319
rect 499 269 563 285
rect 597 319 665 593
rect 597 285 631 319
rect 597 269 665 285
rect 699 319 835 593
rect 869 573 873 607
rect 907 573 923 607
rect 869 519 923 573
rect 869 485 873 519
rect 907 485 923 519
rect 869 435 923 485
rect 869 401 873 435
rect 907 401 923 435
rect 869 385 923 401
rect 699 285 739 319
rect 773 285 835 319
rect 699 269 835 285
rect 869 309 935 350
rect 869 275 885 309
rect 919 275 935 309
rect 869 269 935 275
rect 413 242 451 258
rect 324 205 440 208
rect 324 171 390 205
rect 424 171 440 205
rect 324 95 440 171
rect 324 61 390 95
rect 424 61 440 95
rect 324 51 440 61
rect 485 205 922 235
rect 519 201 678 205
rect 519 171 532 201
rect 485 101 532 171
rect 666 171 678 201
rect 712 201 872 205
rect 712 171 726 201
rect 519 67 532 101
rect 485 51 532 67
rect 566 133 582 167
rect 616 133 632 167
rect 566 91 632 133
rect 566 57 582 91
rect 616 57 632 91
rect 566 17 632 57
rect 666 101 726 171
rect 860 171 872 201
rect 906 171 922 205
rect 666 67 678 101
rect 712 67 726 101
rect 666 51 726 67
rect 760 133 776 167
rect 810 133 826 167
rect 760 91 826 133
rect 760 57 776 91
rect 810 57 826 91
rect 760 17 826 57
rect 860 101 922 171
rect 860 67 872 101
rect 906 67 922 101
rect 860 51 922 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o41a_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 538 833 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 512076
string GDS_START 501776
<< end >>
