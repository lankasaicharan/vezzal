magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4274 1975
<< nwell >>
rect -38 331 3014 704
rect 2195 306 2600 331
<< pwell >>
rect 1094 273 1304 281
rect 197 214 679 229
rect 1094 222 2099 273
rect 2308 222 2975 241
rect 1094 214 2975 222
rect 197 167 2975 214
rect 1 49 2975 167
rect 0 0 2976 49
<< scnmos >>
rect 83 57 113 141
rect 279 119 309 203
rect 464 119 494 203
rect 550 119 580 203
rect 675 104 705 188
rect 789 104 819 188
rect 988 60 1018 188
rect 1075 60 1105 188
rect 1191 127 1221 255
rect 1417 119 1447 247
rect 1519 119 1549 247
rect 1668 163 1698 247
rect 1746 163 1776 247
rect 1881 119 1911 247
rect 1970 119 2000 247
rect 2088 68 2118 196
rect 2289 47 2319 131
rect 2391 47 2421 215
rect 2477 47 2507 215
rect 2675 131 2705 215
rect 2777 47 2807 215
rect 2863 47 2893 215
<< scpmoshvt >>
rect 105 481 135 609
rect 303 449 333 577
rect 433 449 463 533
rect 519 449 549 533
rect 679 449 709 533
rect 789 449 819 533
rect 1003 379 1033 547
rect 1089 379 1119 547
rect 1191 379 1221 547
rect 1417 379 1447 547
rect 1512 428 1542 596
rect 1614 506 1644 590
rect 1783 506 1813 590
rect 1932 428 1962 596
rect 2018 428 2048 596
rect 2090 428 2120 596
rect 2287 342 2317 470
rect 2389 342 2419 594
rect 2475 342 2505 594
rect 2675 367 2705 495
rect 2777 367 2807 619
rect 2863 367 2893 619
<< ndiff >>
rect 223 174 279 203
rect 27 116 83 141
rect 27 82 38 116
rect 72 82 83 116
rect 27 57 83 82
rect 113 116 169 141
rect 223 140 234 174
rect 268 140 279 174
rect 223 119 279 140
rect 309 174 464 203
rect 309 140 336 174
rect 370 140 464 174
rect 309 119 464 140
rect 494 178 550 203
rect 494 144 505 178
rect 539 144 550 178
rect 494 119 550 144
rect 580 188 653 203
rect 1120 243 1191 255
rect 1120 209 1131 243
rect 1165 209 1191 243
rect 1120 188 1191 209
rect 580 162 675 188
rect 580 128 607 162
rect 641 128 675 162
rect 580 119 675 128
rect 113 82 124 116
rect 158 82 169 116
rect 113 57 169 82
rect 595 104 675 119
rect 705 104 789 188
rect 819 132 988 188
rect 819 104 857 132
rect 845 98 857 104
rect 891 98 988 132
rect 845 60 988 98
rect 1018 166 1075 188
rect 1018 132 1029 166
rect 1063 132 1075 166
rect 1018 60 1075 132
rect 1105 127 1191 188
rect 1221 173 1278 255
rect 1221 139 1232 173
rect 1266 139 1278 173
rect 1221 127 1278 139
rect 1360 165 1417 247
rect 1360 131 1372 165
rect 1406 131 1417 165
rect 1105 60 1176 127
rect 1360 119 1417 131
rect 1447 119 1519 247
rect 1549 235 1668 247
rect 1549 201 1607 235
rect 1641 201 1668 235
rect 1549 165 1668 201
rect 1549 131 1607 165
rect 1641 163 1668 165
rect 1698 163 1746 247
rect 1776 168 1881 247
rect 1776 163 1823 168
rect 1641 131 1653 163
rect 1549 119 1653 131
rect 1811 134 1823 163
rect 1857 134 1881 168
rect 1811 119 1881 134
rect 1911 168 1970 247
rect 1911 134 1925 168
rect 1959 134 1970 168
rect 1911 119 1970 134
rect 2000 196 2073 247
rect 2000 195 2088 196
rect 2000 161 2027 195
rect 2061 161 2088 195
rect 2000 119 2088 161
rect 2015 68 2088 119
rect 2118 114 2177 196
rect 2334 184 2391 215
rect 2334 150 2346 184
rect 2380 150 2391 184
rect 2334 131 2391 150
rect 2118 80 2131 114
rect 2165 80 2177 114
rect 2118 68 2177 80
rect 2232 111 2289 131
rect 2232 77 2244 111
rect 2278 77 2289 111
rect 2232 47 2289 77
rect 2319 93 2391 131
rect 2319 59 2346 93
rect 2380 59 2391 93
rect 2319 47 2391 59
rect 2421 185 2477 215
rect 2421 151 2432 185
rect 2466 151 2477 185
rect 2421 103 2477 151
rect 2421 69 2432 103
rect 2466 69 2477 103
rect 2421 47 2477 69
rect 2507 203 2564 215
rect 2507 169 2518 203
rect 2552 169 2564 203
rect 2507 93 2564 169
rect 2618 190 2675 215
rect 2618 156 2630 190
rect 2664 156 2675 190
rect 2618 131 2675 156
rect 2705 203 2777 215
rect 2705 169 2732 203
rect 2766 169 2777 203
rect 2705 131 2777 169
rect 2507 59 2518 93
rect 2552 59 2564 93
rect 2507 47 2564 59
rect 2720 93 2777 131
rect 2720 59 2732 93
rect 2766 59 2777 93
rect 2720 47 2777 59
rect 2807 203 2863 215
rect 2807 169 2818 203
rect 2852 169 2863 203
rect 2807 103 2863 169
rect 2807 69 2818 103
rect 2852 69 2863 103
rect 2807 47 2863 69
rect 2893 113 2949 215
rect 2893 79 2904 113
rect 2938 79 2949 113
rect 2893 47 2949 79
<< pdiff >>
rect 32 597 105 609
rect 32 563 44 597
rect 78 563 105 597
rect 32 527 105 563
rect 32 493 44 527
rect 78 493 105 527
rect 32 481 105 493
rect 135 597 192 609
rect 135 563 146 597
rect 180 563 192 597
rect 135 527 192 563
rect 135 493 146 527
rect 180 493 192 527
rect 135 481 192 493
rect 246 565 303 577
rect 246 531 258 565
rect 292 531 303 565
rect 246 495 303 531
rect 246 461 258 495
rect 292 461 303 495
rect 246 449 303 461
rect 333 565 406 577
rect 333 531 360 565
rect 394 533 406 565
rect 930 582 988 594
rect 930 548 942 582
rect 976 548 988 582
rect 930 547 988 548
rect 1462 547 1512 596
rect 930 533 1003 547
rect 394 531 433 533
rect 333 495 433 531
rect 333 461 360 495
rect 394 461 433 495
rect 333 449 433 461
rect 463 508 519 533
rect 463 474 474 508
rect 508 474 519 508
rect 463 449 519 474
rect 549 508 679 533
rect 549 474 634 508
rect 668 474 679 508
rect 549 449 679 474
rect 709 449 789 533
rect 819 449 1003 533
rect 930 379 1003 449
rect 1033 523 1089 547
rect 1033 489 1044 523
rect 1078 489 1089 523
rect 1033 379 1089 489
rect 1119 379 1191 547
rect 1221 535 1417 547
rect 1221 501 1263 535
rect 1297 501 1417 535
rect 1221 425 1417 501
rect 1221 391 1263 425
rect 1297 391 1417 425
rect 1221 379 1417 391
rect 1447 428 1512 547
rect 1542 590 1592 596
rect 1875 590 1932 596
rect 1542 506 1614 590
rect 1644 506 1783 590
rect 1813 572 1932 590
rect 1813 538 1887 572
rect 1921 538 1932 572
rect 1813 506 1932 538
rect 1542 500 1599 506
rect 1542 466 1553 500
rect 1587 466 1599 500
rect 1542 428 1599 466
rect 1447 379 1497 428
rect 1875 428 1932 506
rect 1962 584 2018 596
rect 1962 550 1973 584
rect 2007 550 2018 584
rect 1962 490 2018 550
rect 1962 456 1973 490
rect 2007 456 2018 490
rect 1962 428 2018 456
rect 2048 428 2090 596
rect 2120 572 2177 596
rect 2720 607 2777 619
rect 2120 538 2131 572
rect 2165 538 2177 572
rect 2120 428 2177 538
rect 2332 571 2389 594
rect 2332 537 2344 571
rect 2378 537 2389 571
rect 2332 470 2389 537
rect 2231 388 2287 470
rect 2231 354 2242 388
rect 2276 354 2287 388
rect 2231 342 2287 354
rect 2317 342 2389 470
rect 2419 582 2475 594
rect 2419 548 2430 582
rect 2464 548 2475 582
rect 2419 485 2475 548
rect 2419 451 2430 485
rect 2464 451 2475 485
rect 2419 389 2475 451
rect 2419 355 2430 389
rect 2464 355 2475 389
rect 2419 342 2475 355
rect 2505 582 2564 594
rect 2505 548 2518 582
rect 2552 548 2564 582
rect 2505 485 2564 548
rect 2720 573 2732 607
rect 2766 573 2777 607
rect 2720 510 2777 573
rect 2720 495 2732 510
rect 2505 451 2518 485
rect 2552 451 2564 485
rect 2505 388 2564 451
rect 2505 354 2518 388
rect 2552 354 2564 388
rect 2618 483 2675 495
rect 2618 449 2630 483
rect 2664 449 2675 483
rect 2618 413 2675 449
rect 2618 379 2630 413
rect 2664 379 2675 413
rect 2618 367 2675 379
rect 2705 476 2732 495
rect 2766 476 2777 510
rect 2705 413 2777 476
rect 2705 379 2732 413
rect 2766 379 2777 413
rect 2705 367 2777 379
rect 2807 597 2863 619
rect 2807 563 2818 597
rect 2852 563 2863 597
rect 2807 505 2863 563
rect 2807 471 2818 505
rect 2852 471 2863 505
rect 2807 413 2863 471
rect 2807 379 2818 413
rect 2852 379 2863 413
rect 2807 367 2863 379
rect 2893 607 2949 619
rect 2893 573 2904 607
rect 2938 573 2949 607
rect 2893 477 2949 573
rect 2893 443 2904 477
rect 2938 443 2949 477
rect 2893 367 2949 443
rect 2505 342 2564 354
<< ndiffc >>
rect 38 82 72 116
rect 234 140 268 174
rect 336 140 370 174
rect 505 144 539 178
rect 1131 209 1165 243
rect 607 128 641 162
rect 124 82 158 116
rect 857 98 891 132
rect 1029 132 1063 166
rect 1232 139 1266 173
rect 1372 131 1406 165
rect 1607 201 1641 235
rect 1607 131 1641 165
rect 1823 134 1857 168
rect 1925 134 1959 168
rect 2027 161 2061 195
rect 2346 150 2380 184
rect 2131 80 2165 114
rect 2244 77 2278 111
rect 2346 59 2380 93
rect 2432 151 2466 185
rect 2432 69 2466 103
rect 2518 169 2552 203
rect 2630 156 2664 190
rect 2732 169 2766 203
rect 2518 59 2552 93
rect 2732 59 2766 93
rect 2818 169 2852 203
rect 2818 69 2852 103
rect 2904 79 2938 113
<< pdiffc >>
rect 44 563 78 597
rect 44 493 78 527
rect 146 563 180 597
rect 146 493 180 527
rect 258 531 292 565
rect 258 461 292 495
rect 360 531 394 565
rect 942 548 976 582
rect 360 461 394 495
rect 474 474 508 508
rect 634 474 668 508
rect 1044 489 1078 523
rect 1263 501 1297 535
rect 1263 391 1297 425
rect 1887 538 1921 572
rect 1553 466 1587 500
rect 1973 550 2007 584
rect 1973 456 2007 490
rect 2131 538 2165 572
rect 2344 537 2378 571
rect 2242 354 2276 388
rect 2430 548 2464 582
rect 2430 451 2464 485
rect 2430 355 2464 389
rect 2518 548 2552 582
rect 2732 573 2766 607
rect 2518 451 2552 485
rect 2518 354 2552 388
rect 2630 449 2664 483
rect 2630 379 2664 413
rect 2732 476 2766 510
rect 2732 379 2766 413
rect 2818 563 2852 597
rect 2818 471 2852 505
rect 2818 379 2852 413
rect 2904 573 2938 607
rect 2904 443 2938 477
<< poly >>
rect 105 609 135 635
rect 303 601 549 631
rect 303 577 333 601
rect 105 466 135 481
rect 57 436 135 466
rect 433 533 463 559
rect 519 533 549 601
rect 679 615 1542 645
rect 679 533 709 615
rect 1512 596 1542 615
rect 789 533 819 559
rect 1003 547 1033 573
rect 1089 547 1119 573
rect 1191 547 1221 573
rect 1417 547 1447 573
rect 57 316 87 436
rect 303 394 333 449
rect 433 434 463 449
rect 21 300 87 316
rect 21 266 37 300
rect 71 266 87 300
rect 21 232 87 266
rect 135 378 333 394
rect 135 344 151 378
rect 185 364 333 378
rect 381 404 463 434
rect 519 423 549 449
rect 679 430 709 449
rect 185 344 201 364
rect 135 310 201 344
rect 135 276 151 310
rect 185 290 201 310
rect 381 302 411 404
rect 597 400 709 430
rect 789 417 819 449
rect 789 401 887 417
rect 597 362 627 400
rect 459 346 627 362
rect 789 367 837 401
rect 871 367 887 401
rect 1614 590 1644 616
rect 1783 590 1813 616
rect 1932 596 1962 622
rect 2018 596 2048 622
rect 2090 596 2120 622
rect 1614 491 1644 506
rect 1614 461 1735 491
rect 1783 474 1813 506
rect 1669 458 1735 461
rect 1512 413 1542 428
rect 1669 424 1685 458
rect 1719 424 1735 458
rect 1512 383 1627 413
rect 459 312 475 346
rect 509 332 627 346
rect 675 336 741 352
rect 509 312 580 332
rect 185 276 309 290
rect 135 260 309 276
rect 21 198 37 232
rect 71 212 87 232
rect 71 198 113 212
rect 279 203 309 260
rect 351 286 417 302
rect 459 296 580 312
rect 351 252 367 286
rect 401 252 417 286
rect 351 248 417 252
rect 351 218 494 248
rect 464 203 494 218
rect 550 203 580 296
rect 675 302 691 336
rect 725 302 741 336
rect 675 268 741 302
rect 675 234 691 268
rect 725 234 741 268
rect 675 218 741 234
rect 789 351 887 367
rect 21 182 113 198
rect 83 141 113 182
rect 675 188 705 218
rect 789 188 819 351
rect 1003 347 1033 379
rect 1089 347 1119 379
rect 967 331 1033 347
rect 967 297 983 331
rect 1017 297 1033 331
rect 967 281 1033 297
rect 1075 331 1141 347
rect 1075 297 1091 331
rect 1125 297 1141 331
rect 1075 281 1141 297
rect 988 188 1018 281
rect 1075 188 1105 281
rect 1191 255 1221 379
rect 1417 347 1447 379
rect 1365 331 1447 347
rect 1365 297 1381 331
rect 1415 297 1447 331
rect 1365 281 1447 297
rect 83 31 113 57
rect 279 51 309 119
rect 464 93 494 119
rect 550 93 580 119
rect 675 51 705 104
rect 789 78 819 104
rect 1417 247 1447 281
rect 1489 319 1555 335
rect 1489 285 1505 319
rect 1539 285 1555 319
rect 1489 269 1555 285
rect 1597 292 1627 383
rect 1669 390 1735 424
rect 1669 356 1685 390
rect 1719 356 1735 390
rect 1669 340 1735 356
rect 1777 458 1843 474
rect 1777 424 1793 458
rect 1827 424 1843 458
rect 2389 594 2419 620
rect 2475 594 2505 620
rect 2777 619 2807 645
rect 2863 619 2893 645
rect 2287 470 2317 496
rect 1777 408 1843 424
rect 1932 413 1962 428
rect 2018 413 2048 428
rect 1777 292 1807 408
rect 1885 383 1962 413
rect 2010 383 2048 413
rect 1885 360 1915 383
rect 1849 344 1915 360
rect 1849 310 1865 344
rect 1899 310 1915 344
rect 2010 335 2040 383
rect 2090 335 2120 428
rect 2675 495 2705 521
rect 1849 294 1915 310
rect 1959 319 2040 335
rect 1519 247 1549 269
rect 1597 262 1698 292
rect 1668 247 1698 262
rect 1746 262 1807 292
rect 1746 247 1776 262
rect 1881 247 1911 294
rect 1959 285 1975 319
rect 2009 285 2040 319
rect 1959 269 2040 285
rect 2088 319 2197 335
rect 2088 285 2147 319
rect 2181 285 2197 319
rect 2287 302 2317 342
rect 2389 303 2419 342
rect 2088 269 2197 285
rect 2246 286 2317 302
rect 1970 247 2000 269
rect 279 21 705 51
rect 988 34 1018 60
rect 1075 34 1105 60
rect 1191 51 1221 127
rect 1668 137 1698 163
rect 1746 137 1776 163
rect 2088 196 2118 269
rect 2246 252 2262 286
rect 2296 252 2317 286
rect 2246 236 2317 252
rect 2359 287 2425 303
rect 2359 253 2375 287
rect 2409 267 2425 287
rect 2475 267 2505 342
rect 2675 267 2705 367
rect 2777 321 2807 367
rect 2409 253 2705 267
rect 2753 305 2819 321
rect 2753 271 2769 305
rect 2803 285 2819 305
rect 2863 285 2893 367
rect 2803 271 2893 285
rect 2753 255 2893 271
rect 2359 237 2705 253
rect 1417 93 1447 119
rect 1519 93 1549 119
rect 1881 93 1911 119
rect 1970 93 2000 119
rect 2246 189 2276 236
rect 2391 215 2421 237
rect 2477 215 2507 237
rect 2675 215 2705 237
rect 2777 215 2807 255
rect 2863 215 2893 255
rect 2246 159 2319 189
rect 2289 131 2319 159
rect 2088 51 2118 68
rect 1191 21 2118 51
rect 2675 105 2705 131
rect 2289 21 2319 47
rect 2391 21 2421 47
rect 2477 21 2507 47
rect 2777 21 2807 47
rect 2863 21 2893 47
<< polycont >>
rect 37 266 71 300
rect 151 344 185 378
rect 151 276 185 310
rect 837 367 871 401
rect 1685 424 1719 458
rect 475 312 509 346
rect 37 198 71 232
rect 367 252 401 286
rect 691 302 725 336
rect 691 234 725 268
rect 983 297 1017 331
rect 1091 297 1125 331
rect 1381 297 1415 331
rect 1505 285 1539 319
rect 1685 356 1719 390
rect 1793 424 1827 458
rect 1865 310 1899 344
rect 1975 285 2009 319
rect 2147 285 2181 319
rect 2262 252 2296 286
rect 2375 253 2409 287
rect 2769 271 2803 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 28 597 94 649
rect 28 563 44 597
rect 78 563 94 597
rect 28 527 94 563
rect 28 493 44 527
rect 78 493 94 527
rect 28 477 94 493
rect 130 597 201 613
rect 130 563 146 597
rect 180 563 201 597
rect 130 527 201 563
rect 130 493 146 527
rect 180 493 201 527
rect 21 300 87 430
rect 21 266 37 300
rect 71 266 87 300
rect 21 232 87 266
rect 21 198 37 232
rect 71 198 87 232
rect 21 182 87 198
rect 130 378 201 493
rect 130 344 151 378
rect 185 344 201 378
rect 130 310 201 344
rect 130 276 151 310
rect 185 276 201 310
rect 130 260 201 276
rect 242 565 308 581
rect 242 531 258 565
rect 292 531 308 565
rect 242 495 308 531
rect 242 461 258 495
rect 292 461 308 495
rect 242 409 308 461
rect 344 565 410 649
rect 344 531 360 565
rect 394 531 410 565
rect 926 582 992 649
rect 926 548 942 582
rect 976 548 992 582
rect 344 495 410 531
rect 344 461 360 495
rect 394 461 410 495
rect 458 508 524 537
rect 458 474 474 508
rect 508 495 524 508
rect 618 508 684 537
rect 926 532 992 548
rect 508 474 582 495
rect 458 461 582 474
rect 344 445 410 461
rect 242 375 512 409
rect 130 145 174 260
rect 242 200 276 375
rect 459 346 512 375
rect 459 312 475 346
rect 509 312 512 346
rect 313 286 417 302
rect 459 296 512 312
rect 313 252 367 286
rect 401 252 417 286
rect 548 260 582 461
rect 313 236 417 252
rect 489 226 582 260
rect 618 474 634 508
rect 668 479 684 508
rect 1028 523 1094 551
rect 1028 496 1044 523
rect 834 489 1044 496
rect 1078 496 1094 523
rect 1247 535 1313 649
rect 1247 501 1263 535
rect 1297 501 1313 535
rect 1078 489 1211 496
rect 668 474 798 479
rect 618 445 798 474
rect 22 116 72 145
rect 22 82 38 116
rect 22 17 72 82
rect 108 116 174 145
rect 108 82 124 116
rect 158 82 174 116
rect 218 174 284 200
rect 218 140 234 174
rect 268 140 284 174
rect 218 115 284 140
rect 320 174 386 200
rect 320 140 336 174
rect 370 140 386 174
rect 108 53 174 82
rect 320 17 386 140
rect 489 178 555 226
rect 618 190 652 445
rect 688 336 728 352
rect 688 302 691 336
rect 725 302 728 336
rect 688 268 728 302
rect 764 315 798 445
rect 834 462 1211 489
rect 834 401 874 462
rect 834 367 837 401
rect 871 367 874 401
rect 834 351 874 367
rect 910 392 1141 426
rect 910 315 944 392
rect 764 281 944 315
rect 980 350 1033 356
rect 980 331 991 350
rect 980 297 983 331
rect 1025 316 1033 350
rect 1017 297 1033 316
rect 980 281 1033 297
rect 1075 331 1141 392
rect 1075 297 1091 331
rect 1125 297 1141 331
rect 1075 295 1141 297
rect 1177 321 1211 462
rect 1247 425 1313 501
rect 1247 391 1263 425
rect 1297 391 1313 425
rect 1247 375 1313 391
rect 1467 579 1723 613
rect 1365 331 1431 347
rect 1365 321 1381 331
rect 1177 297 1381 321
rect 1415 297 1431 331
rect 1177 287 1431 297
rect 1467 335 1501 579
rect 1537 500 1625 543
rect 1537 466 1553 500
rect 1587 466 1625 500
rect 1537 424 1625 466
rect 1467 319 1555 335
rect 688 234 691 268
rect 725 245 728 268
rect 1177 259 1211 287
rect 725 234 977 245
rect 688 211 977 234
rect 489 144 505 178
rect 539 144 555 178
rect 489 115 555 144
rect 607 162 652 190
rect 641 128 652 162
rect 607 100 652 128
rect 841 132 907 175
rect 841 98 857 132
rect 891 98 907 132
rect 841 17 907 98
rect 943 87 977 211
rect 1115 243 1211 259
rect 1467 285 1505 319
rect 1539 285 1555 319
rect 1467 251 1555 285
rect 1115 209 1131 243
rect 1165 225 1211 243
rect 1165 209 1181 225
rect 1115 193 1181 209
rect 1302 217 1555 251
rect 1591 258 1625 424
rect 1669 458 1723 579
rect 1871 572 1921 649
rect 1871 538 1887 572
rect 1871 510 1921 538
rect 1957 584 2023 600
rect 1957 550 1973 584
rect 2007 550 2023 584
rect 1957 490 2023 550
rect 2115 572 2181 649
rect 2115 538 2131 572
rect 2165 538 2181 572
rect 2115 510 2181 538
rect 2328 571 2394 649
rect 2328 537 2344 571
rect 2378 537 2394 571
rect 2328 510 2394 537
rect 2430 582 2482 598
rect 2464 548 2482 582
rect 1957 474 1973 490
rect 1669 424 1685 458
rect 1719 424 1723 458
rect 1669 390 1723 424
rect 1777 458 1973 474
rect 1777 424 1793 458
rect 1827 456 1973 458
rect 2007 474 2023 490
rect 2430 485 2482 548
rect 2007 456 2393 474
rect 1827 440 2393 456
rect 1827 424 1843 440
rect 1777 408 1843 424
rect 1669 356 1685 390
rect 1719 356 1723 390
rect 1669 340 1723 356
rect 1759 350 1915 360
rect 1793 344 1915 350
rect 1793 316 1865 344
rect 1759 310 1865 316
rect 1899 310 1915 344
rect 1759 294 1915 310
rect 1957 319 2025 335
rect 1957 285 1975 319
rect 2009 285 2025 319
rect 1957 269 2025 285
rect 1957 258 1991 269
rect 1591 235 1991 258
rect 1013 166 1079 192
rect 1013 132 1029 166
rect 1063 157 1079 166
rect 1232 173 1266 189
rect 1063 139 1232 157
rect 1063 132 1266 139
rect 1013 123 1266 132
rect 1302 87 1336 217
rect 1591 201 1607 235
rect 1641 224 1991 235
rect 2061 233 2095 440
rect 2163 388 2292 404
rect 2163 354 2242 388
rect 2276 354 2292 388
rect 2163 338 2292 354
rect 1641 201 1657 224
rect 943 53 1336 87
rect 1372 165 1422 181
rect 1406 131 1422 165
rect 1372 17 1422 131
rect 1591 165 1657 201
rect 2027 195 2095 233
rect 1591 131 1607 165
rect 1641 131 1657 165
rect 1591 115 1657 131
rect 1807 168 1873 188
rect 1807 134 1823 168
rect 1857 134 1873 168
rect 1807 17 1873 134
rect 1909 168 1975 188
rect 1909 134 1925 168
rect 1959 134 1975 168
rect 1909 87 1975 134
rect 2061 161 2095 195
rect 2131 319 2197 338
rect 2131 285 2147 319
rect 2181 285 2197 319
rect 2359 303 2393 440
rect 2464 451 2482 485
rect 2430 389 2482 451
rect 2464 355 2482 389
rect 2430 339 2482 355
rect 2131 200 2197 285
rect 2233 286 2312 302
rect 2233 252 2262 286
rect 2296 252 2312 286
rect 2233 236 2312 252
rect 2359 287 2412 303
rect 2359 253 2375 287
rect 2409 253 2412 287
rect 2359 237 2412 253
rect 2448 201 2482 339
rect 2518 582 2568 649
rect 2552 548 2568 582
rect 2518 485 2568 548
rect 2716 607 2766 649
rect 2716 573 2732 607
rect 2716 510 2766 573
rect 2552 451 2568 485
rect 2518 388 2568 451
rect 2552 354 2568 388
rect 2518 338 2568 354
rect 2614 483 2680 499
rect 2614 449 2630 483
rect 2664 449 2680 483
rect 2614 413 2680 449
rect 2614 379 2630 413
rect 2664 379 2680 413
rect 2614 321 2680 379
rect 2716 476 2732 510
rect 2716 413 2766 476
rect 2716 379 2732 413
rect 2716 363 2766 379
rect 2802 597 2868 613
rect 2802 563 2818 597
rect 2852 563 2868 597
rect 2802 505 2868 563
rect 2802 471 2818 505
rect 2852 471 2868 505
rect 2802 413 2868 471
rect 2904 607 2954 649
rect 2938 573 2954 607
rect 2904 477 2954 573
rect 2938 443 2954 477
rect 2904 427 2954 443
rect 2802 379 2818 413
rect 2852 391 2868 413
rect 2852 379 2889 391
rect 2802 357 2889 379
rect 2614 305 2819 321
rect 2614 271 2769 305
rect 2803 271 2819 305
rect 2614 255 2819 271
rect 2131 166 2294 200
rect 2027 123 2095 161
rect 2131 114 2181 130
rect 1909 80 2131 87
rect 2165 80 2181 114
rect 1909 53 2181 80
rect 2244 111 2294 166
rect 2278 77 2294 111
rect 2244 53 2294 77
rect 2330 184 2380 200
rect 2330 150 2346 184
rect 2330 93 2380 150
rect 2330 59 2346 93
rect 2330 17 2380 59
rect 2416 185 2482 201
rect 2416 151 2432 185
rect 2466 151 2482 185
rect 2416 103 2482 151
rect 2416 69 2432 103
rect 2466 69 2482 103
rect 2416 53 2482 69
rect 2518 203 2568 219
rect 2552 169 2568 203
rect 2518 93 2568 169
rect 2614 190 2680 255
rect 2855 219 2889 357
rect 2614 156 2630 190
rect 2664 156 2680 190
rect 2614 127 2680 156
rect 2716 203 2766 219
rect 2716 169 2732 203
rect 2552 59 2568 93
rect 2518 17 2568 59
rect 2716 93 2766 169
rect 2716 59 2732 93
rect 2716 17 2766 59
rect 2802 203 2889 219
rect 2802 169 2818 203
rect 2852 185 2889 203
rect 2852 169 2868 185
rect 2802 103 2868 169
rect 2802 69 2818 103
rect 2852 69 2868 103
rect 2802 53 2868 69
rect 2904 113 2954 149
rect 2938 79 2954 113
rect 2904 17 2954 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 991 331 1025 350
rect 991 316 1017 331
rect 1017 316 1025 331
rect 1759 316 1793 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
<< metal1 >>
rect 0 683 2976 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 2976 683
rect 0 617 2976 649
rect 979 350 1037 356
rect 979 316 991 350
rect 1025 347 1037 350
rect 1747 350 1805 356
rect 1747 347 1759 350
rect 1025 319 1759 347
rect 1025 316 1037 319
rect 979 310 1037 316
rect 1747 316 1759 319
rect 1793 316 1805 350
rect 1747 310 1805 316
rect 0 17 2976 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 2976 17
rect 0 -49 2976 -17
<< labels >>
flabel pwell s 0 0 2976 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2976 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfbbn_2
flabel comment s 486 39 486 39 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 617 2976 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2976 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 2239 242 2273 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 SET_B
port 4 nsew signal input
flabel locali s 2815 94 2849 128 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2815 168 2849 202 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2431 94 2465 128 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2976 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2153020
string GDS_START 2133292
<< end >>
