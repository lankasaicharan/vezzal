magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 1 49 911 263
rect 0 0 960 49
<< scnmos >>
rect 80 69 110 237
rect 166 69 196 237
rect 252 69 282 237
rect 338 69 368 237
rect 529 69 559 237
rect 630 69 660 237
rect 716 69 746 237
rect 802 69 832 237
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 252 367 282 619
rect 354 367 384 619
rect 440 367 470 619
rect 630 367 660 619
rect 716 367 746 619
rect 802 367 832 619
<< ndiff >>
rect 27 208 80 237
rect 27 174 35 208
rect 69 174 80 208
rect 27 117 80 174
rect 27 83 35 117
rect 69 83 80 117
rect 27 69 80 83
rect 110 132 166 237
rect 110 98 121 132
rect 155 98 166 132
rect 110 69 166 98
rect 196 208 252 237
rect 196 174 207 208
rect 241 174 252 208
rect 196 117 252 174
rect 196 83 207 117
rect 241 83 252 117
rect 196 69 252 83
rect 282 124 338 237
rect 282 90 293 124
rect 327 90 338 124
rect 282 69 338 90
rect 368 225 421 237
rect 368 191 379 225
rect 413 191 421 225
rect 368 157 421 191
rect 368 123 379 157
rect 413 123 421 157
rect 368 69 421 123
rect 475 225 529 237
rect 475 191 483 225
rect 517 191 529 225
rect 475 155 529 191
rect 475 121 483 155
rect 517 121 529 155
rect 475 69 529 121
rect 559 183 630 237
rect 559 149 585 183
rect 619 149 630 183
rect 559 111 630 149
rect 559 77 585 111
rect 619 77 630 111
rect 559 69 630 77
rect 660 225 716 237
rect 660 191 671 225
rect 705 191 716 225
rect 660 115 716 191
rect 660 81 671 115
rect 705 81 716 115
rect 660 69 716 81
rect 746 183 802 237
rect 746 149 757 183
rect 791 149 802 183
rect 746 111 802 149
rect 746 77 757 111
rect 791 77 802 111
rect 746 69 802 77
rect 832 225 885 237
rect 832 191 843 225
rect 877 191 885 225
rect 832 115 885 191
rect 832 81 843 115
rect 877 81 885 115
rect 832 69 885 81
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 510 80 565
rect 27 476 35 510
rect 69 476 80 510
rect 27 413 80 476
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 607 166 619
rect 110 573 121 607
rect 155 573 166 607
rect 110 527 166 573
rect 110 493 121 527
rect 155 493 166 527
rect 110 445 166 493
rect 110 411 121 445
rect 155 411 166 445
rect 110 367 166 411
rect 196 599 252 619
rect 196 565 207 599
rect 241 565 252 599
rect 196 510 252 565
rect 196 476 207 510
rect 241 476 252 510
rect 196 413 252 476
rect 196 379 207 413
rect 241 379 252 413
rect 196 367 252 379
rect 282 607 354 619
rect 282 573 302 607
rect 336 573 354 607
rect 282 527 354 573
rect 282 493 302 527
rect 336 493 354 527
rect 282 445 354 493
rect 282 411 302 445
rect 336 411 354 445
rect 282 367 354 411
rect 384 599 440 619
rect 384 565 395 599
rect 429 565 440 599
rect 384 510 440 565
rect 384 476 395 510
rect 429 476 440 510
rect 384 409 440 476
rect 384 375 395 409
rect 429 375 440 409
rect 384 367 440 375
rect 470 571 630 619
rect 470 537 481 571
rect 515 537 585 571
rect 619 537 630 571
rect 470 367 630 537
rect 660 599 716 619
rect 660 565 671 599
rect 705 565 716 599
rect 660 510 716 565
rect 660 476 671 510
rect 705 476 716 510
rect 660 367 716 476
rect 746 537 802 619
rect 746 503 757 537
rect 791 503 802 537
rect 746 428 802 503
rect 746 394 757 428
rect 791 394 802 428
rect 746 367 802 394
rect 832 599 885 619
rect 832 565 843 599
rect 877 565 885 599
rect 832 512 885 565
rect 832 478 843 512
rect 877 478 885 512
rect 832 434 885 478
rect 832 400 843 434
rect 877 400 885 434
rect 832 367 885 400
<< ndiffc >>
rect 35 174 69 208
rect 35 83 69 117
rect 121 98 155 132
rect 207 174 241 208
rect 207 83 241 117
rect 293 90 327 124
rect 379 191 413 225
rect 379 123 413 157
rect 483 191 517 225
rect 483 121 517 155
rect 585 149 619 183
rect 585 77 619 111
rect 671 191 705 225
rect 671 81 705 115
rect 757 149 791 183
rect 757 77 791 111
rect 843 191 877 225
rect 843 81 877 115
<< pdiffc >>
rect 35 565 69 599
rect 35 476 69 510
rect 35 379 69 413
rect 121 573 155 607
rect 121 493 155 527
rect 121 411 155 445
rect 207 565 241 599
rect 207 476 241 510
rect 207 379 241 413
rect 302 573 336 607
rect 302 493 336 527
rect 302 411 336 445
rect 395 565 429 599
rect 395 476 429 510
rect 395 375 429 409
rect 481 537 515 571
rect 585 537 619 571
rect 671 565 705 599
rect 671 476 705 510
rect 757 503 791 537
rect 757 394 791 428
rect 843 565 877 599
rect 843 478 877 512
rect 843 400 877 434
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 252 619 282 645
rect 354 619 384 645
rect 440 619 470 645
rect 630 619 660 645
rect 716 619 746 645
rect 802 619 832 645
rect 80 325 110 367
rect 25 309 110 325
rect 25 275 41 309
rect 75 289 110 309
rect 166 289 196 367
rect 75 275 196 289
rect 25 259 196 275
rect 80 237 110 259
rect 166 237 196 259
rect 252 325 282 367
rect 354 325 384 367
rect 252 309 384 325
rect 252 275 277 309
rect 311 275 384 309
rect 252 259 384 275
rect 440 299 470 367
rect 630 335 660 367
rect 716 335 746 367
rect 802 335 832 367
rect 601 319 667 335
rect 601 299 617 319
rect 440 285 617 299
rect 651 285 667 319
rect 440 269 667 285
rect 716 319 832 335
rect 716 285 782 319
rect 816 285 832 319
rect 716 269 832 285
rect 252 237 282 259
rect 338 237 368 259
rect 529 237 559 269
rect 630 237 660 269
rect 716 237 746 269
rect 802 237 832 269
rect 80 43 110 69
rect 166 43 196 69
rect 252 43 282 69
rect 338 43 368 69
rect 529 43 559 69
rect 630 43 660 69
rect 716 43 746 69
rect 802 43 832 69
<< polycont >>
rect 41 275 75 309
rect 277 275 311 309
rect 617 285 651 319
rect 782 285 816 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 19 599 71 615
rect 19 565 35 599
rect 69 565 71 599
rect 19 510 71 565
rect 19 476 35 510
rect 69 476 71 510
rect 19 413 71 476
rect 19 379 35 413
rect 69 379 71 413
rect 105 607 171 649
rect 105 573 121 607
rect 155 573 171 607
rect 105 527 171 573
rect 105 493 121 527
rect 155 493 171 527
rect 105 445 171 493
rect 105 411 121 445
rect 155 411 171 445
rect 205 599 252 615
rect 205 565 207 599
rect 241 565 252 599
rect 205 510 252 565
rect 205 476 207 510
rect 241 476 252 510
rect 205 413 252 476
rect 19 377 71 379
rect 205 379 207 413
rect 241 379 252 413
rect 286 607 352 649
rect 286 573 302 607
rect 336 573 352 607
rect 286 527 352 573
rect 286 493 302 527
rect 336 493 352 527
rect 286 445 352 493
rect 286 411 302 445
rect 336 411 352 445
rect 386 599 431 615
rect 386 565 395 599
rect 429 565 431 599
rect 386 510 431 565
rect 465 571 635 649
rect 465 537 481 571
rect 515 537 585 571
rect 619 537 635 571
rect 465 528 635 537
rect 669 599 893 615
rect 669 565 671 599
rect 705 581 843 599
rect 705 565 707 581
rect 386 476 395 510
rect 429 494 431 510
rect 669 510 707 565
rect 841 565 843 581
rect 877 565 893 599
rect 669 494 671 510
rect 429 476 671 494
rect 705 476 707 510
rect 386 460 707 476
rect 741 537 807 547
rect 741 503 757 537
rect 791 503 807 537
rect 205 377 252 379
rect 386 409 433 460
rect 741 428 807 503
rect 741 426 757 428
rect 386 377 395 409
rect 19 375 395 377
rect 429 375 433 409
rect 19 343 433 375
rect 467 394 757 426
rect 791 394 807 428
rect 467 390 807 394
rect 841 512 893 565
rect 841 478 843 512
rect 877 478 893 512
rect 841 434 893 478
rect 841 400 843 434
rect 877 400 893 434
rect 18 275 41 309
rect 75 275 91 309
rect 18 242 91 275
rect 125 275 277 309
rect 311 275 327 309
rect 125 242 327 275
rect 467 251 558 390
rect 841 384 893 400
rect 592 319 667 350
rect 592 285 617 319
rect 651 285 667 319
rect 701 319 943 350
rect 701 285 782 319
rect 816 285 943 319
rect 363 225 429 241
rect 363 208 379 225
rect 19 174 35 208
rect 69 174 207 208
rect 241 191 379 208
rect 413 191 429 225
rect 241 174 429 191
rect 19 117 69 174
rect 19 83 35 117
rect 19 67 69 83
rect 105 132 171 140
rect 105 98 121 132
rect 155 98 171 132
rect 105 17 171 98
rect 205 117 251 174
rect 363 157 429 174
rect 205 83 207 117
rect 241 83 251 117
rect 205 67 251 83
rect 285 124 329 140
rect 285 90 293 124
rect 327 90 329 124
rect 363 123 379 157
rect 413 123 429 157
rect 363 121 429 123
rect 467 225 893 251
rect 467 191 483 225
rect 517 217 671 225
rect 517 191 535 217
rect 467 155 535 191
rect 669 191 671 217
rect 705 217 843 225
rect 705 191 707 217
rect 467 121 483 155
rect 517 121 535 155
rect 569 149 585 183
rect 619 149 635 183
rect 285 87 329 90
rect 569 111 635 149
rect 569 87 585 111
rect 285 77 585 87
rect 619 77 635 111
rect 285 51 635 77
rect 669 115 707 191
rect 841 191 843 217
rect 877 191 893 225
rect 669 81 671 115
rect 705 81 707 115
rect 669 65 707 81
rect 741 149 757 183
rect 791 149 807 183
rect 741 111 807 149
rect 741 77 757 111
rect 791 77 807 111
rect 741 17 807 77
rect 841 115 893 191
rect 841 81 843 115
rect 877 81 893 115
rect 841 65 893 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a31oi_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3449032
string GDS_START 3440444
<< end >>
