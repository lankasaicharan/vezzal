magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 10 241 386 261
rect 10 49 849 241
rect 0 0 864 49
<< scnmos >>
rect 89 67 119 235
rect 175 67 205 235
rect 277 67 307 235
rect 467 47 497 215
rect 568 47 598 215
rect 654 47 684 215
rect 740 47 770 215
<< scpmoshvt >>
rect 97 367 127 619
rect 205 367 235 619
rect 277 367 307 619
rect 431 367 461 619
rect 503 367 533 619
rect 657 367 687 619
rect 743 367 773 619
<< ndiff >>
rect 36 206 89 235
rect 36 172 44 206
rect 78 172 89 206
rect 36 113 89 172
rect 36 79 44 113
rect 78 79 89 113
rect 36 67 89 79
rect 119 130 175 235
rect 119 96 130 130
rect 164 96 175 130
rect 119 67 175 96
rect 205 227 277 235
rect 205 193 230 227
rect 264 193 277 227
rect 205 153 277 193
rect 205 119 230 153
rect 264 119 277 153
rect 205 67 277 119
rect 307 149 360 235
rect 307 115 318 149
rect 352 115 360 149
rect 307 67 360 115
rect 414 165 467 215
rect 414 131 422 165
rect 456 131 467 165
rect 414 93 467 131
rect 414 59 422 93
rect 456 59 467 93
rect 414 47 467 59
rect 497 203 568 215
rect 497 169 519 203
rect 553 169 568 203
rect 497 101 568 169
rect 497 67 519 101
rect 553 67 568 101
rect 497 47 568 67
rect 598 203 654 215
rect 598 169 609 203
rect 643 169 654 203
rect 598 93 654 169
rect 598 59 609 93
rect 643 59 654 93
rect 598 47 654 59
rect 684 203 740 215
rect 684 169 695 203
rect 729 169 740 203
rect 684 101 740 169
rect 684 67 695 101
rect 729 67 740 101
rect 684 47 740 67
rect 770 163 823 215
rect 770 129 781 163
rect 815 129 823 163
rect 770 93 823 129
rect 770 59 781 93
rect 815 59 823 93
rect 770 47 823 59
<< pdiff >>
rect 44 599 97 619
rect 44 565 52 599
rect 86 565 97 599
rect 44 510 97 565
rect 44 476 52 510
rect 86 476 97 510
rect 44 420 97 476
rect 44 386 52 420
rect 86 386 97 420
rect 44 367 97 386
rect 127 607 205 619
rect 127 573 149 607
rect 183 573 205 607
rect 127 492 205 573
rect 127 458 149 492
rect 183 458 205 492
rect 127 367 205 458
rect 235 367 277 619
rect 307 599 431 619
rect 307 565 318 599
rect 352 565 386 599
rect 420 565 431 599
rect 307 515 431 565
rect 307 481 318 515
rect 352 481 386 515
rect 420 481 431 515
rect 307 420 431 481
rect 307 386 318 420
rect 352 386 386 420
rect 420 386 431 420
rect 307 367 431 386
rect 461 367 503 619
rect 533 607 657 619
rect 533 573 544 607
rect 578 573 612 607
rect 646 573 657 607
rect 533 492 657 573
rect 533 458 544 492
rect 578 458 612 492
rect 646 458 657 492
rect 533 367 657 458
rect 687 599 743 619
rect 687 565 698 599
rect 732 565 743 599
rect 687 505 743 565
rect 687 471 698 505
rect 732 471 743 505
rect 687 413 743 471
rect 687 379 698 413
rect 732 379 743 413
rect 687 367 743 379
rect 773 607 826 619
rect 773 573 784 607
rect 818 573 826 607
rect 773 538 826 573
rect 773 504 784 538
rect 818 504 826 538
rect 773 467 826 504
rect 773 433 784 467
rect 818 433 826 467
rect 773 367 826 433
<< ndiffc >>
rect 44 172 78 206
rect 44 79 78 113
rect 130 96 164 130
rect 230 193 264 227
rect 230 119 264 153
rect 318 115 352 149
rect 422 131 456 165
rect 422 59 456 93
rect 519 169 553 203
rect 519 67 553 101
rect 609 169 643 203
rect 609 59 643 93
rect 695 169 729 203
rect 695 67 729 101
rect 781 129 815 163
rect 781 59 815 93
<< pdiffc >>
rect 52 565 86 599
rect 52 476 86 510
rect 52 386 86 420
rect 149 573 183 607
rect 149 458 183 492
rect 318 565 352 599
rect 386 565 420 599
rect 318 481 352 515
rect 386 481 420 515
rect 318 386 352 420
rect 386 386 420 420
rect 544 573 578 607
rect 612 573 646 607
rect 544 458 578 492
rect 612 458 646 492
rect 698 565 732 599
rect 698 471 732 505
rect 698 379 732 413
rect 784 573 818 607
rect 784 504 818 538
rect 784 433 818 467
<< poly >>
rect 97 619 127 645
rect 205 619 235 645
rect 277 619 307 645
rect 431 619 461 645
rect 503 619 533 645
rect 657 619 687 645
rect 743 619 773 645
rect 97 323 127 367
rect 205 344 235 367
rect 23 307 127 323
rect 23 273 39 307
rect 73 293 127 307
rect 169 319 235 344
rect 73 273 119 293
rect 23 257 119 273
rect 169 285 185 319
rect 219 285 235 319
rect 169 269 235 285
rect 277 333 307 367
rect 277 317 343 333
rect 431 317 461 367
rect 277 283 293 317
rect 327 283 343 317
rect 89 235 119 257
rect 175 235 205 269
rect 277 266 343 283
rect 395 301 461 317
rect 503 345 533 367
rect 503 319 605 345
rect 657 335 687 367
rect 743 335 773 367
rect 503 315 555 319
rect 395 267 411 301
rect 445 267 461 301
rect 539 285 555 315
rect 589 285 605 319
rect 539 269 605 285
rect 654 319 773 335
rect 654 285 670 319
rect 704 287 773 319
rect 704 285 770 287
rect 654 269 770 285
rect 277 235 307 266
rect 395 237 497 267
rect 467 215 497 237
rect 568 215 598 269
rect 654 215 684 269
rect 740 215 770 269
rect 89 41 119 67
rect 175 41 205 67
rect 277 41 307 67
rect 467 21 497 47
rect 568 21 598 47
rect 654 21 684 47
rect 740 21 770 47
<< polycont >>
rect 39 273 73 307
rect 185 285 219 319
rect 293 283 327 317
rect 411 267 445 301
rect 555 285 589 319
rect 670 285 704 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 36 599 99 615
rect 36 565 52 599
rect 86 565 99 599
rect 36 510 99 565
rect 36 476 52 510
rect 86 476 99 510
rect 36 420 99 476
rect 133 607 199 649
rect 133 573 149 607
rect 183 573 199 607
rect 133 492 199 573
rect 133 458 149 492
rect 183 458 199 492
rect 133 454 199 458
rect 302 599 439 615
rect 302 565 318 599
rect 352 565 386 599
rect 420 565 439 599
rect 302 515 439 565
rect 302 481 318 515
rect 352 481 386 515
rect 420 481 439 515
rect 302 420 439 481
rect 528 607 662 649
rect 528 573 544 607
rect 578 573 612 607
rect 646 573 662 607
rect 528 492 662 573
rect 528 458 544 492
rect 578 458 612 492
rect 646 458 662 492
rect 528 454 662 458
rect 696 599 734 615
rect 696 565 698 599
rect 732 565 734 599
rect 696 505 734 565
rect 696 471 698 505
rect 732 471 734 505
rect 36 386 52 420
rect 86 386 318 420
rect 352 386 386 420
rect 420 386 659 420
rect 17 307 75 352
rect 17 273 39 307
rect 73 273 75 307
rect 17 242 75 273
rect 109 206 143 386
rect 177 319 259 352
rect 177 285 185 319
rect 219 285 259 319
rect 177 269 259 285
rect 293 317 361 350
rect 327 283 361 317
rect 293 267 361 283
rect 395 301 475 352
rect 395 267 411 301
rect 445 267 475 301
rect 509 319 591 352
rect 509 285 555 319
rect 589 285 591 319
rect 509 269 591 285
rect 625 329 659 386
rect 696 413 734 471
rect 768 607 834 649
rect 768 573 784 607
rect 818 573 834 607
rect 768 538 834 573
rect 768 504 784 538
rect 818 504 834 538
rect 768 467 834 504
rect 768 433 784 467
rect 818 433 834 467
rect 696 379 698 413
rect 732 397 734 413
rect 732 379 844 397
rect 696 363 844 379
rect 625 319 720 329
rect 625 285 670 319
rect 704 285 720 319
rect 625 281 720 285
rect 754 247 844 363
rect 28 172 44 206
rect 78 172 143 206
rect 214 227 568 233
rect 214 193 230 227
rect 264 203 568 227
rect 264 199 519 203
rect 264 193 280 199
rect 28 113 80 172
rect 214 153 280 193
rect 506 169 519 199
rect 553 169 568 203
rect 28 79 44 113
rect 78 79 80 113
rect 28 63 80 79
rect 114 130 180 138
rect 114 96 130 130
rect 164 96 180 130
rect 214 119 230 153
rect 264 119 280 153
rect 314 149 368 165
rect 114 85 180 96
rect 314 115 318 149
rect 352 115 368 149
rect 314 85 368 115
rect 114 51 368 85
rect 406 131 422 165
rect 456 131 472 165
rect 406 93 472 131
rect 406 59 422 93
rect 456 59 472 93
rect 406 17 472 59
rect 506 101 568 169
rect 506 67 519 101
rect 553 67 568 101
rect 506 51 568 67
rect 602 203 651 219
rect 602 169 609 203
rect 643 169 651 203
rect 602 93 651 169
rect 602 59 609 93
rect 643 59 651 93
rect 602 17 651 59
rect 685 213 844 247
rect 685 203 737 213
rect 685 169 695 203
rect 729 169 737 203
rect 685 101 737 169
rect 685 67 695 101
rect 729 67 737 101
rect 685 51 737 67
rect 771 163 831 179
rect 771 129 781 163
rect 815 129 831 163
rect 771 93 831 129
rect 771 59 781 93
rect 815 59 831 93
rect 771 17 831 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221a_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4874650
string GDS_START 4866144
<< end >>
