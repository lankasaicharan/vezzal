magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 77 49 608 160
rect 0 0 672 49
<< scnmos >>
rect 183 50 213 134
rect 255 50 285 134
rect 327 50 357 134
rect 413 50 443 134
rect 499 50 529 134
<< scpmoshvt >>
rect 155 535 185 619
rect 241 535 271 619
rect 327 535 357 619
rect 413 535 443 619
rect 485 535 515 619
<< ndiff >>
rect 103 104 183 134
rect 103 70 111 104
rect 145 70 183 104
rect 103 50 183 70
rect 213 50 255 134
rect 285 50 327 134
rect 357 122 413 134
rect 357 88 368 122
rect 402 88 413 122
rect 357 50 413 88
rect 443 96 499 134
rect 443 62 454 96
rect 488 62 499 96
rect 443 50 499 62
rect 529 122 582 134
rect 529 88 540 122
rect 574 88 582 122
rect 529 50 582 88
<< pdiff >>
rect 49 607 155 619
rect 49 573 57 607
rect 91 573 155 607
rect 49 535 155 573
rect 185 581 241 619
rect 185 547 196 581
rect 230 547 241 581
rect 185 535 241 547
rect 271 611 327 619
rect 271 577 282 611
rect 316 577 327 611
rect 271 535 327 577
rect 357 577 413 619
rect 357 543 368 577
rect 402 543 413 577
rect 357 535 413 543
rect 443 535 485 619
rect 515 607 568 619
rect 515 573 526 607
rect 560 573 568 607
rect 515 535 568 573
<< ndiffc >>
rect 111 70 145 104
rect 368 88 402 122
rect 454 62 488 96
rect 540 88 574 122
<< pdiffc >>
rect 57 573 91 607
rect 196 547 230 581
rect 282 577 316 611
rect 368 543 402 577
rect 526 573 560 607
<< poly >>
rect 155 619 185 645
rect 241 619 271 645
rect 327 619 357 645
rect 413 619 443 645
rect 485 619 515 645
rect 155 446 185 535
rect 241 512 271 535
rect 119 416 185 446
rect 227 482 271 512
rect 119 290 149 416
rect 227 368 257 482
rect 327 440 357 535
rect 305 424 371 440
rect 305 390 321 424
rect 355 390 371 424
rect 83 274 149 290
rect 83 240 99 274
rect 133 240 149 274
rect 83 206 149 240
rect 197 352 263 368
rect 197 318 213 352
rect 247 318 263 352
rect 197 284 263 318
rect 305 356 371 390
rect 305 322 321 356
rect 355 322 371 356
rect 305 306 371 322
rect 413 376 443 535
rect 485 454 515 535
rect 485 438 593 454
rect 485 424 543 438
rect 527 404 543 424
rect 577 404 593 438
rect 413 360 479 376
rect 413 326 429 360
rect 463 326 479 360
rect 197 250 213 284
rect 247 258 263 284
rect 247 250 285 258
rect 197 228 285 250
rect 83 172 99 206
rect 133 186 149 206
rect 133 172 213 186
rect 83 156 213 172
rect 183 134 213 156
rect 255 134 285 228
rect 327 134 357 306
rect 413 292 479 326
rect 413 258 429 292
rect 463 258 479 292
rect 413 242 479 258
rect 527 370 593 404
rect 527 336 543 370
rect 577 336 593 370
rect 527 320 593 336
rect 413 134 443 242
rect 527 194 557 320
rect 499 164 557 194
rect 499 134 529 164
rect 183 24 213 50
rect 255 24 285 50
rect 327 24 357 50
rect 413 24 443 50
rect 499 24 529 50
<< polycont >>
rect 321 390 355 424
rect 99 240 133 274
rect 213 318 247 352
rect 321 322 355 356
rect 543 404 577 438
rect 429 326 463 360
rect 213 250 247 284
rect 99 172 133 206
rect 429 258 463 292
rect 543 336 577 370
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 53 607 91 649
rect 53 573 57 607
rect 278 611 320 649
rect 53 557 91 573
rect 127 581 234 597
rect 127 547 196 581
rect 230 547 234 581
rect 278 577 282 611
rect 316 577 320 611
rect 510 607 576 649
rect 278 561 320 577
rect 364 577 449 593
rect 127 525 234 547
rect 364 543 368 577
rect 402 543 449 577
rect 510 573 526 607
rect 560 573 576 607
rect 510 569 576 573
rect 364 525 449 543
rect 127 498 449 525
rect 29 464 449 498
rect 29 120 63 464
rect 511 438 577 498
rect 99 274 161 424
rect 133 240 161 274
rect 99 206 161 240
rect 133 172 161 206
rect 99 156 161 172
rect 213 352 257 424
rect 247 318 257 352
rect 213 284 257 318
rect 247 250 257 284
rect 29 104 149 120
rect 29 70 111 104
rect 145 70 149 104
rect 213 94 257 250
rect 305 390 321 424
rect 355 390 371 424
rect 305 356 371 390
rect 305 322 321 356
rect 355 322 371 356
rect 305 242 371 322
rect 415 360 463 424
rect 415 326 429 360
rect 415 292 463 326
rect 415 258 429 292
rect 415 242 463 258
rect 511 404 543 438
rect 511 370 577 404
rect 511 336 543 370
rect 511 242 577 336
rect 364 148 578 182
rect 364 122 406 148
rect 364 88 368 122
rect 402 88 406 122
rect 536 122 578 148
rect 364 72 406 88
rect 450 96 492 112
rect 29 54 149 70
rect 450 62 454 96
rect 488 62 492 96
rect 536 88 540 122
rect 574 88 578 122
rect 536 72 578 88
rect 450 17 492 62
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2111ai_m
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4735716
string GDS_START 4727666
<< end >>
