magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1336 -1345 414140 2582
<< locali >>
rect 407485 1035 407543 1071
rect 407485 561 407543 597
rect 366545 491 366603 527
rect 407485 491 407543 527
rect 366545 17 366603 53
rect 407485 17 407543 53
<< metal1 >>
rect -76 1074 0 1102
rect 412804 1074 412880 1102
rect -76 14 -48 1074
rect 33244 592 33272 623
rect 33336 592 33364 691
rect 29 527 63 561
rect -76 -14 0 14
rect 29 -17 63 17
rect 412852 14 412880 1074
rect 412804 -14 412880 14
use sky130_fd_sc_hdll__a211o_1  sky130_fd_sc_hdll__a211o_1_0
timestamp 1627202621
transform 1 0 0 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__a211o_2  sky130_fd_sc_hdll__a211o_2_0
timestamp 1627202621
transform 1 0 828 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__a211o_4  sky130_fd_sc_hdll__a211o_4_0
timestamp 1627202621
transform 1 0 1748 0 1 0
box -38 -48 1510 592
use sky130_fd_sc_hdll__a211oi_1  sky130_fd_sc_hdll__a211oi_1_0
timestamp 1627202621
transform 1 0 3312 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__a211oi_2  sky130_fd_sc_hdll__a211oi_2_0
timestamp 1627202621
transform 1 0 3956 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__a211oi_4  sky130_fd_sc_hdll__a211oi_4_0
timestamp 1627202621
transform 1 0 5060 0 1 0
box -38 -48 1694 592
use sky130_fd_sc_hdll__a21bo_1  sky130_fd_sc_hdll__a21bo_1_0
timestamp 1627202621
transform 1 0 6808 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__a21bo_2  sky130_fd_sc_hdll__a21bo_2_0
timestamp 1627202621
transform 1 0 7728 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__a21bo_4  sky130_fd_sc_hdll__a21bo_4_0
timestamp 1627202621
transform 1 0 8648 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__a21boi_1  sky130_fd_sc_hdll__a21boi_1_0
timestamp 1627202621
transform 1 0 10028 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__a21boi_2  sky130_fd_sc_hdll__a21boi_2_0
timestamp 1627202621
transform 1 0 10764 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__a21boi_4  sky130_fd_sc_hdll__a21boi_4_0
timestamp 1627202621
transform 1 0 11776 0 1 0
box -38 -48 1510 592
use sky130_fd_sc_hdll__a21o_1  sky130_fd_sc_hdll__a21o_1_0
timestamp 1627202621
transform 1 0 13340 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__a21o_2  sky130_fd_sc_hdll__a21o_2_0
timestamp 1627202621
transform 1 0 14076 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__a21o_4  sky130_fd_sc_hdll__a21o_4_0
timestamp 1627202621
transform 1 0 14904 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__a21oi_1  sky130_fd_sc_hdll__a21oi_1_0
timestamp 1627202621
transform 1 0 16192 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__a21oi_2  sky130_fd_sc_hdll__a21oi_2_0
timestamp 1627202621
transform 1 0 16744 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__a21oi_4  sky130_fd_sc_hdll__a21oi_4_0
timestamp 1627202621
transform 1 0 17572 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__a221oi_1  sky130_fd_sc_hdll__a221oi_1_0
timestamp 1627202621
transform 1 0 18952 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__a221oi_2  sky130_fd_sc_hdll__a221oi_2_0
timestamp 1627202621
transform 1 0 19780 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__a221oi_4  sky130_fd_sc_hdll__a221oi_4_0
timestamp 1627202621
transform 1 0 21068 0 1 0
box -38 -48 2154 592
use sky130_fd_sc_hdll__a222oi_1  sky130_fd_sc_hdll__a222oi_1_0
timestamp 1627202621
transform 1 0 23276 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__a22o_1  sky130_fd_sc_hdll__a22o_1_0
timestamp 1627202621
transform 1 0 24196 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__a22o_2  sky130_fd_sc_hdll__a22o_2_0
timestamp 1627202621
transform 1 0 25024 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__a22o_4  sky130_fd_sc_hdll__a22o_4_0
timestamp 1627202621
transform 1 0 25944 0 1 0
box -38 -48 1418 592
use sky130_fd_sc_hdll__a22oi_1  sky130_fd_sc_hdll__a22oi_1_0
timestamp 1627202621
transform 1 0 27416 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__a22oi_2  sky130_fd_sc_hdll__a22oi_2_0
timestamp 1627202621
transform 1 0 28152 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__a22oi_4  sky130_fd_sc_hdll__a22oi_4_0
timestamp 1627202621
transform 1 0 29256 0 1 0
box -38 -48 1786 592
use sky130_fd_sc_hdll__a2bb2o_1  sky130_fd_sc_hdll__a2bb2o_1_0
timestamp 1627202621
transform 1 0 31096 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__a2bb2o_2  sky130_fd_sc_hdll__a2bb2o_2_0
timestamp 1627202621
transform 1 0 32016 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__a2bb2o_4  sky130_fd_sc_hdll__a2bb2o_4_0
timestamp 1627202621
transform 1 0 33028 0 1 0
box -38 -48 1602 592
use sky130_fd_sc_hdll__a2bb2oi_1  sky130_fd_sc_hdll__a2bb2oi_1_0
timestamp 1627202621
transform 1 0 34684 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__a2bb2oi_2  sky130_fd_sc_hdll__a2bb2oi_2_0
timestamp 1627202621
transform 1 0 35512 0 1 0
box -65 -48 1234 592
use sky130_fd_sc_hdll__a2bb2oi_4  sky130_fd_sc_hdll__a2bb2oi_4_0
timestamp 1627202621
transform 1 0 36800 0 1 0
box -38 -48 2154 592
use sky130_fd_sc_hdll__a31o_1  sky130_fd_sc_hdll__a31o_1_0
timestamp 1627202621
transform 1 0 39008 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__a31o_2  sky130_fd_sc_hdll__a31o_2_0
timestamp 1627202621
transform 1 0 39744 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__a31o_4  sky130_fd_sc_hdll__a31o_4_0
timestamp 1627202621
transform 1 0 40572 0 1 0
box -38 -48 1418 592
use sky130_fd_sc_hdll__a31oi_1  sky130_fd_sc_hdll__a31oi_1_0
timestamp 1627202621
transform 1 0 42044 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__a31oi_2  sky130_fd_sc_hdll__a31oi_2_0
timestamp 1627202621
transform 1 0 42688 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__a31oi_4  sky130_fd_sc_hdll__a31oi_4_0
timestamp 1627202621
transform 1 0 43792 0 1 0
box -38 -48 1786 592
use sky130_fd_sc_hdll__a32o_1  sky130_fd_sc_hdll__a32o_1_0
timestamp 1627202621
transform 1 0 45632 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__a32o_2  sky130_fd_sc_hdll__a32o_2_0
timestamp 1627202621
transform 1 0 46552 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__a32o_4  sky130_fd_sc_hdll__a32o_4_0
timestamp 1627202621
transform 1 0 47564 0 1 0
box -38 -48 1694 592
use sky130_fd_sc_hdll__a32oi_1  sky130_fd_sc_hdll__a32oi_1_0
timestamp 1627202621
transform 1 0 49312 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__a32oi_2  sky130_fd_sc_hdll__a32oi_2_0
timestamp 1627202621
transform 1 0 50048 0 1 0
box -39 -48 1326 592
use sky130_fd_sc_hdll__a32oi_4  sky130_fd_sc_hdll__a32oi_4_0
timestamp 1627202621
transform 1 0 51428 0 1 0
box -38 -48 2338 592
use sky130_fd_sc_hdll__and2_1  sky130_fd_sc_hdll__and2_1_0
timestamp 1627202621
transform 1 0 53820 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__and2_2  sky130_fd_sc_hdll__and2_2_0
timestamp 1627202621
transform 1 0 54372 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__and2_4  sky130_fd_sc_hdll__and2_4_0
timestamp 1627202621
transform 1 0 55016 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__and2b_1  sky130_fd_sc_hdll__and2b_1_0
timestamp 1627202621
transform 1 0 55844 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__and2b_2  sky130_fd_sc_hdll__and2b_2_0
timestamp 1627202621
transform 1 0 56580 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__and2b_4  sky130_fd_sc_hdll__and2b_4_0
timestamp 1627202621
transform 1 0 57408 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__and3_1  sky130_fd_sc_hdll__and3_1_0
timestamp 1627202621
transform 1 0 58328 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__and3_2  sky130_fd_sc_hdll__and3_2_0
timestamp 1627202621
transform 1 0 58972 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__and3_4  sky130_fd_sc_hdll__and3_4_0
timestamp 1627202621
transform 1 0 59708 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__and3b_1  sky130_fd_sc_hdll__and3b_1_0
timestamp 1627202621
transform 1 0 60720 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__and3b_2  sky130_fd_sc_hdll__and3b_2_0
timestamp 1627202621
transform 1 0 61548 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__and3b_4  sky130_fd_sc_hdll__and3b_4_0
timestamp 1627202621
transform 1 0 62468 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__and4_1  sky130_fd_sc_hdll__and4_1_0
timestamp 1627202621
transform 1 0 63572 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__and4_2  sky130_fd_sc_hdll__and4_2_0
timestamp 1627202621
transform 1 0 64308 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__and4_4  sky130_fd_sc_hdll__and4_4_0
timestamp 1627202621
transform 1 0 65136 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__and4b_1  sky130_fd_sc_hdll__and4b_1_0
timestamp 1627202621
transform 1 0 66148 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__and4b_2  sky130_fd_sc_hdll__and4b_2_0
timestamp 1627202621
transform 1 0 67068 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__and4b_4  sky130_fd_sc_hdll__and4b_4_0
timestamp 1627202621
transform 1 0 68080 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__and4bb_1  sky130_fd_sc_hdll__and4bb_1_0
timestamp 1627202621
transform 1 0 69184 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__and4bb_2  sky130_fd_sc_hdll__and4bb_2_0
timestamp 1627202621
transform 1 0 70196 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__and4bb_4  sky130_fd_sc_hdll__and4bb_4_0
timestamp 1627202621
transform 1 0 71300 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__buf_1  sky130_fd_sc_hdll__buf_1_0
timestamp 1627202621
transform 1 0 72680 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hdll__buf_12  sky130_fd_sc_hdll__buf_12_0
timestamp 1627202621
transform 1 0 73140 0 1 0
box -38 -48 1694 592
use sky130_fd_sc_hdll__buf_16  sky130_fd_sc_hdll__buf_16_0
timestamp 1627202621
transform 1 0 74888 0 1 0
box -38 -48 2338 592
use sky130_fd_sc_hdll__buf_2  sky130_fd_sc_hdll__buf_2_0
timestamp 1627202621
transform 1 0 77280 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__buf_4  sky130_fd_sc_hdll__buf_4_0
timestamp 1627202621
transform 1 0 77832 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__buf_6  sky130_fd_sc_hdll__buf_6_0
timestamp 1627202621
transform 1 0 78568 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__buf_8  sky130_fd_sc_hdll__buf_8_0
timestamp 1627202621
transform 1 0 79580 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__bufbuf_16  sky130_fd_sc_hdll__bufbuf_16_0
timestamp 1627202621
transform 1 0 80868 0 1 0
box -38 -48 2706 592
use sky130_fd_sc_hdll__bufbuf_8  sky130_fd_sc_hdll__bufbuf_8_0
timestamp 1627202621
transform 1 0 83628 0 1 0
box -38 -48 1510 592
use sky130_fd_sc_hdll__bufinv_16  sky130_fd_sc_hdll__bufinv_16_0
timestamp 1627202621
transform 1 0 85192 0 1 0
box -38 -48 2522 592
use sky130_fd_sc_hdll__bufinv_8  sky130_fd_sc_hdll__bufinv_8_0
timestamp 1627202621
transform 1 0 87768 0 1 0
box -38 -48 1418 592
use sky130_fd_sc_hdll__clkbuf_1  sky130_fd_sc_hdll__clkbuf_1_0
timestamp 1627202621
transform 1 0 89240 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hdll__clkbuf_16  sky130_fd_sc_hdll__clkbuf_16_0
timestamp 1627202621
transform 1 0 89700 0 1 0
box -38 -48 2062 592
use sky130_fd_sc_hdll__clkbuf_2  sky130_fd_sc_hdll__clkbuf_2_0
timestamp 1627202621
transform 1 0 91816 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__clkbuf_4  sky130_fd_sc_hdll__clkbuf_4_0
timestamp 1627202621
transform 1 0 92368 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__clkbuf_8  sky130_fd_sc_hdll__clkbuf_8_0
timestamp 1627202621
transform 1 0 93104 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hdll__clkinv_1  sky130_fd_sc_hdll__clkinv_1_0
timestamp 1627202621
transform 1 0 94300 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hdll__clkinv_16  sky130_fd_sc_hdll__clkinv_16_0
timestamp 1627202621
transform 1 0 94760 0 1 0
box -38 -48 2522 592
use sky130_fd_sc_hdll__clkinv_2  sky130_fd_sc_hdll__clkinv_2_0
timestamp 1627202621
transform 1 0 97336 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__clkinv_4  sky130_fd_sc_hdll__clkinv_4_0
timestamp 1627202621
transform 1 0 97888 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__clkinv_8  sky130_fd_sc_hdll__clkinv_8_0
timestamp 1627202621
transform 1 0 98716 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__clkinvlp_2  sky130_fd_sc_hdll__clkinvlp_2_0
timestamp 1627202621
transform 1 0 100096 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hdll__clkinvlp_4  sky130_fd_sc_hdll__clkinvlp_4_0
timestamp 1627202621
transform 1 0 100556 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__conb_1  sky130_fd_sc_hdll__conb_1_0
timestamp 1627202621
transform 1 0 101200 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hdll__dfrtp_1  sky130_fd_sc_hdll__dfrtp_1_0
timestamp 1627202621
transform 1 0 101568 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hdll__dfrtp_2  sky130_fd_sc_hdll__dfrtp_2_0
timestamp 1627202621
transform 1 0 103592 0 1 0
box -38 -48 2062 592
use sky130_fd_sc_hdll__dfrtp_4  sky130_fd_sc_hdll__dfrtp_4_0
timestamp 1627202621
transform 1 0 105708 0 1 0
box -38 -48 2338 592
use sky130_fd_sc_hdll__dfstp_1  sky130_fd_sc_hdll__dfstp_1_0
timestamp 1627202621
transform 1 0 108100 0 1 0
box -38 -48 2062 592
use sky130_fd_sc_hdll__dfstp_2  sky130_fd_sc_hdll__dfstp_2_0
timestamp 1627202621
transform 1 0 110216 0 1 0
box -38 -48 2154 592
use sky130_fd_sc_hdll__dfstp_4  sky130_fd_sc_hdll__dfstp_4_0
timestamp 1627202621
transform 1 0 112424 0 1 0
box -38 -48 2430 592
use sky130_fd_sc_hdll__dlxtn_1  sky130_fd_sc_hdll__dlxtn_1_0
timestamp 1627202621
transform 1 0 114908 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__dlxtn_2  sky130_fd_sc_hdll__dlxtn_2_0
timestamp 1627202621
transform 1 0 116196 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__dlxtn_4  sky130_fd_sc_hdll__dlxtn_4_0
timestamp 1627202621
transform 1 0 117576 0 1 0
box -38 -48 1510 592
use sky130_fd_sc_hdll__dlygate4sd1_1  sky130_fd_sc_hdll__dlygate4sd1_1_0
timestamp 1627202621
transform 1 0 119140 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__ebufn_1  sky130_fd_sc_hdll__ebufn_1_0
timestamp 1627202621
transform 1 0 121440 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__ebufn_2  sky130_fd_sc_hdll__ebufn_2_0
timestamp 1627202621
transform 1 0 122268 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__ebufn_4  sky130_fd_sc_hdll__ebufn_4_0
timestamp 1627202621
transform 1 0 123280 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__ebufn_8  sky130_fd_sc_hdll__ebufn_8_0
timestamp 1627202621
transform 1 0 124660 0 1 0
box -38 -48 2246 592
use sky130_fd_sc_hdll__einvn_1  sky130_fd_sc_hdll__einvn_1_0
timestamp 1627202621
transform 1 0 126960 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__einvn_2  sky130_fd_sc_hdll__einvn_2_0
timestamp 1627202621
transform 1 0 127604 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__einvn_4  sky130_fd_sc_hdll__einvn_4_0
timestamp 1627202621
transform 1 0 128432 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hdll__einvn_8  sky130_fd_sc_hdll__einvn_8_0
timestamp 1627202621
transform 1 0 129628 0 1 0
box -38 -48 1878 592
use sky130_fd_sc_hdll__einvp_1  sky130_fd_sc_hdll__einvp_1_0
timestamp 1627202621
transform 1 0 131560 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__einvp_2  sky130_fd_sc_hdll__einvp_2_0
timestamp 1627202621
transform 1 0 132204 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__einvp_4  sky130_fd_sc_hdll__einvp_4_0
timestamp 1627202621
transform 1 0 133032 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hdll__einvp_8  sky130_fd_sc_hdll__einvp_8_0
timestamp 1627202621
transform 1 0 134228 0 1 0
box -38 -48 1878 592
use sky130_fd_sc_hdll__inv_1  sky130_fd_sc_hdll__inv_1_0
timestamp 1627202621
transform 1 0 136160 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hdll__inv_12  sky130_fd_sc_hdll__inv_12_0
timestamp 1627202621
transform 1 0 136528 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__inv_16  sky130_fd_sc_hdll__inv_16_0
timestamp 1627202621
transform 1 0 137908 0 1 0
box -38 -48 1694 592
use sky130_fd_sc_hdll__inv_2  sky130_fd_sc_hdll__inv_2_0
timestamp 1627202621
transform 1 0 139656 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hdll__inv_4  sky130_fd_sc_hdll__inv_4_0
timestamp 1627202621
transform 1 0 140116 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__inv_6  sky130_fd_sc_hdll__inv_6_0
timestamp 1627202621
transform 1 0 140760 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__inv_8  sky130_fd_sc_hdll__inv_8_0
timestamp 1627202621
transform 1 0 141588 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__mux2_1  sky130_fd_sc_hdll__mux2_1_0
timestamp 1627202621
transform 1 0 142600 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__mux2_2  sky130_fd_sc_hdll__mux2_2_0
timestamp 1627202621
transform 1 0 143612 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__mux2_4  sky130_fd_sc_hdll__mux2_4_0
timestamp 1627202621
transform 1 0 144624 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__mux2_8  sky130_fd_sc_hdll__mux2_8_0
timestamp 1627202621
transform 1 0 145912 0 1 0
box -38 -48 2154 592
use sky130_fd_sc_hdll__mux2i_1  sky130_fd_sc_hdll__mux2i_1_0
timestamp 1627202621
transform 1 0 148120 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__mux2i_2  sky130_fd_sc_hdll__mux2i_2_0
timestamp 1627202621
transform 1 0 149040 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hdll__mux2i_4  sky130_fd_sc_hdll__mux2i_4_0
timestamp 1627202621
transform 1 0 150236 0 1 0
box -38 -48 1878 592
use sky130_fd_sc_hdll__nand2_1  sky130_fd_sc_hdll__nand2_1_0
timestamp 1627202621
transform 1 0 152168 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hdll__nand2_2  sky130_fd_sc_hdll__nand2_2_0
timestamp 1627202621
transform 1 0 152628 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__nand2_4  sky130_fd_sc_hdll__nand2_4_0
timestamp 1627202621
transform 1 0 153272 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__nand2_8  sky130_fd_sc_hdll__nand2_8_0
timestamp 1627202621
transform 1 0 154284 0 1 0
box -38 -48 1694 592
use sky130_fd_sc_hdll__nand2b_1  sky130_fd_sc_hdll__nand2b_1_0
timestamp 1627202621
transform 1 0 156032 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__nand2b_2  sky130_fd_sc_hdll__nand2b_2_0
timestamp 1627202621
transform 1 0 156584 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__nand2b_4  sky130_fd_sc_hdll__nand2b_4_0
timestamp 1627202621
transform 1 0 157320 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hdll__nand3_1  sky130_fd_sc_hdll__nand3_1_0
timestamp 1627202621
transform 1 0 158516 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__nand3_2  sky130_fd_sc_hdll__nand3_2_0
timestamp 1627202621
transform 1 0 159068 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__nand3_4  sky130_fd_sc_hdll__nand3_4_0
timestamp 1627202621
transform 1 0 159988 0 1 0
box -38 -48 1418 592
use sky130_fd_sc_hdll__nand3b_1  sky130_fd_sc_hdll__nand3b_1_0
timestamp 1627202621
transform 1 0 161460 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__nand3b_2  sky130_fd_sc_hdll__nand3b_2_0
timestamp 1627202621
transform 1 0 162104 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__nand3b_4  sky130_fd_sc_hdll__nand3b_4_0
timestamp 1627202621
transform 1 0 163116 0 1 0
box -38 -48 1602 592
use sky130_fd_sc_hdll__nand4_1  sky130_fd_sc_hdll__nand4_1_0
timestamp 1627202621
transform 1 0 164772 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__nand4_2  sky130_fd_sc_hdll__nand4_2_0
timestamp 1627202621
transform 1 0 165416 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__nand4_4  sky130_fd_sc_hdll__nand4_4_0
timestamp 1627202621
transform 1 0 166520 0 1 0
box -38 -48 1785 592
use sky130_fd_sc_hdll__nand4b_1  sky130_fd_sc_hdll__nand4b_1_0
timestamp 1627202621
transform 1 0 168360 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__nand4b_2  sky130_fd_sc_hdll__nand4b_2_0
timestamp 1627202621
transform 1 0 169096 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__nand4b_4  sky130_fd_sc_hdll__nand4b_4_0
timestamp 1627202621
transform 1 0 170384 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hdll__nand4bb_1  sky130_fd_sc_hdll__nand4bb_1_0
timestamp 1627202621
transform 1 0 172408 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__nand4bb_2  sky130_fd_sc_hdll__nand4bb_2_0
timestamp 1627202621
transform 1 0 173328 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__nand4bb_4  sky130_fd_sc_hdll__nand4bb_4_0
timestamp 1627202621
transform 1 0 174708 0 1 0
box -38 -48 2154 592
use sky130_fd_sc_hdll__nor2_1  sky130_fd_sc_hdll__nor2_1_0
timestamp 1627202621
transform 1 0 176916 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hdll__nor2_2  sky130_fd_sc_hdll__nor2_2_0
timestamp 1627202621
transform 1 0 177376 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__nor2_4  sky130_fd_sc_hdll__nor2_4_0
timestamp 1627202621
transform 1 0 178020 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__nor2_8  sky130_fd_sc_hdll__nor2_8_0
timestamp 1627202621
transform 1 0 179032 0 1 0
box -38 -48 1694 592
use sky130_fd_sc_hdll__nor2b_1  sky130_fd_sc_hdll__nor2b_1_0
timestamp 1627202621
transform 1 0 180780 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__nor2b_2  sky130_fd_sc_hdll__nor2b_2_0
timestamp 1627202621
transform 1 0 181332 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__nor2b_4  sky130_fd_sc_hdll__nor2b_4_0
timestamp 1627202621
transform 1 0 182160 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hdll__nor3_1  sky130_fd_sc_hdll__nor3_1_0
timestamp 1627202621
transform 1 0 183356 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__nor3_2  sky130_fd_sc_hdll__nor3_2_0
timestamp 1627202621
transform 1 0 183908 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__nor3_4  sky130_fd_sc_hdll__nor3_4_0
timestamp 1627202621
transform 1 0 184828 0 1 0
box -38 -85 1326 592
use sky130_fd_sc_hdll__nor3b_1  sky130_fd_sc_hdll__nor3b_1_0
timestamp 1627202621
transform 1 0 186208 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__nor3b_2  sky130_fd_sc_hdll__nor3b_2_0
timestamp 1627202621
transform 1 0 186852 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__nor3b_4  sky130_fd_sc_hdll__nor3b_4_0
timestamp 1627202621
transform 1 0 187956 0 1 0
box -38 -48 1510 592
use sky130_fd_sc_hdll__nor4_1  sky130_fd_sc_hdll__nor4_1_0
timestamp 1627202621
transform 1 0 189520 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__nor4_2  sky130_fd_sc_hdll__nor4_2_0
timestamp 1627202621
transform 1 0 190164 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__nor4_4  sky130_fd_sc_hdll__nor4_4_0
timestamp 1627202621
transform 1 0 191268 0 1 0
box -38 -48 1786 592
use sky130_fd_sc_hdll__nor4b_1  sky130_fd_sc_hdll__nor4b_1_0
timestamp 1627202621
transform 1 0 193108 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__nor4b_2  sky130_fd_sc_hdll__nor4b_2_0
timestamp 1627202621
transform 1 0 193936 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__nor4b_4  sky130_fd_sc_hdll__nor4b_4_0
timestamp 1627202621
transform 1 0 195224 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hdll__nor4bb_1  sky130_fd_sc_hdll__nor4bb_1_0
timestamp 1627202621
transform 1 0 197248 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__nor4bb_2  sky130_fd_sc_hdll__nor4bb_2_0
timestamp 1627202621
transform 1 0 198168 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__nor4bb_4  sky130_fd_sc_hdll__nor4bb_4_0
timestamp 1627202621
transform 1 0 199548 0 1 0
box -38 -48 2062 592
use sky130_fd_sc_hdll__o211a_1  sky130_fd_sc_hdll__o211a_1_0
timestamp 1627202621
transform 1 0 201664 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__o211a_2  sky130_fd_sc_hdll__o211a_2_0
timestamp 1627202621
transform 1 0 202584 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__o211a_4  sky130_fd_sc_hdll__o211a_4_0
timestamp 1627202621
transform 1 0 203504 0 1 0
box -38 -48 1418 592
use sky130_fd_sc_hdll__o211ai_1  sky130_fd_sc_hdll__o211ai_1_0
timestamp 1627202621
transform 1 0 204976 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__o211ai_2  sky130_fd_sc_hdll__o211ai_2_0
timestamp 1627202621
transform 1 0 205620 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__o211ai_4  sky130_fd_sc_hdll__o211ai_4_0
timestamp 1627202621
transform 1 0 206724 0 1 0
box -38 -48 1786 592
use sky130_fd_sc_hdll__o21a_1  sky130_fd_sc_hdll__o21a_1_0
timestamp 1627202621
transform 1 0 208564 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__o21a_2  sky130_fd_sc_hdll__o21a_2_0
timestamp 1627202621
transform 1 0 209300 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__o21a_4  sky130_fd_sc_hdll__o21a_4_0
timestamp 1627202621
transform 1 0 210128 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__o21ai_1  sky130_fd_sc_hdll__o21ai_1_0
timestamp 1627202621
transform 1 0 211416 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__o21ai_2  sky130_fd_sc_hdll__o21ai_2_0
timestamp 1627202621
transform 1 0 211968 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__o21ai_4  sky130_fd_sc_hdll__o21ai_4_0
timestamp 1627202621
transform 1 0 212796 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__o21ba_1  sky130_fd_sc_hdll__o21ba_1_0
timestamp 1627202621
transform 1 0 214176 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__o21ba_2  sky130_fd_sc_hdll__o21ba_2_0
timestamp 1627202621
transform 1 0 215004 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__o21ba_4  sky130_fd_sc_hdll__o21ba_4_0
timestamp 1627202621
transform 1 0 215924 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__o21bai_1  sky130_fd_sc_hdll__o21bai_1_0
timestamp 1627202621
transform 1 0 217304 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__o21bai_2  sky130_fd_sc_hdll__o21bai_2_0
timestamp 1627202621
transform 1 0 218040 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__o21bai_4  sky130_fd_sc_hdll__o21bai_4_0
timestamp 1627202621
transform 1 0 219052 0 1 0
box -38 -48 1510 592
use sky130_fd_sc_hdll__o221a_1  sky130_fd_sc_hdll__o221a_1_0
timestamp 1627202621
transform 1 0 220616 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__o221a_2  sky130_fd_sc_hdll__o221a_2_0
timestamp 1627202621
transform 1 0 221536 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__o221a_4  sky130_fd_sc_hdll__o221a_4_0
timestamp 1627202621
transform 1 0 222548 0 1 0
box -38 -48 1602 592
use sky130_fd_sc_hdll__o221ai_1  sky130_fd_sc_hdll__o221ai_1_0
timestamp 1627202621
transform 1 0 224204 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__o221ai_2  sky130_fd_sc_hdll__o221ai_2_0
timestamp 1627202621
transform 1 0 225032 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__o221ai_4  sky130_fd_sc_hdll__o221ai_4_0
timestamp 1627202621
transform 1 0 226320 0 1 0
box -38 -48 2154 592
use sky130_fd_sc_hdll__o22a_1  sky130_fd_sc_hdll__o22a_1_0
timestamp 1627202621
transform 1 0 228528 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__o22a_2  sky130_fd_sc_hdll__o22a_2_0
timestamp 1627202621
transform 1 0 229356 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__o22a_4  sky130_fd_sc_hdll__o22a_4_0
timestamp 1627202621
transform 1 0 230276 0 1 0
box -38 -48 1418 592
use sky130_fd_sc_hdll__o22ai_1  sky130_fd_sc_hdll__o22ai_1_0
timestamp 1627202621
transform 1 0 231748 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__o22ai_2  sky130_fd_sc_hdll__o22ai_2_0
timestamp 1627202621
transform 1 0 232392 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__o22ai_4  sky130_fd_sc_hdll__o22ai_4_0
timestamp 1627202621
transform 1 0 233496 0 1 0
box -38 -48 1694 592
use sky130_fd_sc_hdll__o2bb2a_1  sky130_fd_sc_hdll__o2bb2a_1_0
timestamp 1627202621
transform 1 0 235244 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__o2bb2a_2  sky130_fd_sc_hdll__o2bb2a_2_0
timestamp 1627202621
transform 1 0 236164 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__o2bb2a_4  sky130_fd_sc_hdll__o2bb2a_4_0
timestamp 1627202621
transform 1 0 237176 0 1 0
box -38 -48 1602 592
use sky130_fd_sc_hdll__o2bb2ai_1  sky130_fd_sc_hdll__o2bb2ai_1_0
timestamp 1627202621
transform 1 0 238832 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__o2bb2ai_2  sky130_fd_sc_hdll__o2bb2ai_2_0
timestamp 1627202621
transform 1 0 239660 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__o2bb2ai_4  sky130_fd_sc_hdll__o2bb2ai_4_0
timestamp 1627202621
transform 1 0 240948 0 1 0
box -38 -48 2246 592
use sky130_fd_sc_hdll__o31ai_1  sky130_fd_sc_hdll__o31ai_1_0
timestamp 1627202621
transform 1 0 243248 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__o31ai_2  sky130_fd_sc_hdll__o31ai_2_0
timestamp 1627202621
transform 1 0 243892 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__o31ai_4  sky130_fd_sc_hdll__o31ai_4_0
timestamp 1627202621
transform 1 0 244996 0 1 0
box -38 -48 1786 592
use sky130_fd_sc_hdll__o32ai_1  sky130_fd_sc_hdll__o32ai_1_0
timestamp 1627202621
transform 1 0 246836 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__o32ai_2  sky130_fd_sc_hdll__o32ai_2_0
timestamp 1627202621
transform 1 0 247572 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__o32ai_4  sky130_fd_sc_hdll__o32ai_4_0
timestamp 1627202621
transform 1 0 248952 0 1 0
box -38 -48 2246 592
use sky130_fd_sc_hdll__or2_1  sky130_fd_sc_hdll__or2_1_0
timestamp 1627202621
transform 1 0 251252 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__or2_2  sky130_fd_sc_hdll__or2_2_0
timestamp 1627202621
transform 1 0 251804 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__or2_4  sky130_fd_sc_hdll__or2_4_0
timestamp 1627202621
transform 1 0 252448 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__or2b_1  sky130_fd_sc_hdll__or2b_1_0
timestamp 1627202621
transform 1 0 253276 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__or2b_2  sky130_fd_sc_hdll__or2b_2_0
timestamp 1627202621
transform 1 0 254012 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__or2b_4  sky130_fd_sc_hdll__or2b_4_0
timestamp 1627202621
transform 1 0 254840 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__or3_1  sky130_fd_sc_hdll__or3_1_0
timestamp 1627202621
transform 1 0 255852 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__or3_2  sky130_fd_sc_hdll__or3_2_0
timestamp 1627202621
transform 1 0 256496 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__or3_4  sky130_fd_sc_hdll__or3_4_0
timestamp 1627202621
transform 1 0 257232 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__or3b_1  sky130_fd_sc_hdll__or3b_1_0
timestamp 1627202621
transform 1 0 258244 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__or3b_2  sky130_fd_sc_hdll__or3b_2_0
timestamp 1627202621
transform 1 0 259072 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__or3b_4  sky130_fd_sc_hdll__or3b_4_0
timestamp 1627202621
transform 1 0 259900 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__or4_1  sky130_fd_sc_hdll__or4_1_0
timestamp 1627202621
transform 1 0 260912 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__or4_2  sky130_fd_sc_hdll__or4_2_0
timestamp 1627202621
transform 1 0 261648 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__or4_4  sky130_fd_sc_hdll__or4_4_0
timestamp 1627202621
transform 1 0 262476 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__or4b_1  sky130_fd_sc_hdll__or4b_1_0
timestamp 1627202621
transform 1 0 263488 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__or4b_2  sky130_fd_sc_hdll__or4b_2_0
timestamp 1627202621
transform 1 0 264408 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hdll__or4b_4  sky130_fd_sc_hdll__or4b_4_0
timestamp 1627202621
transform 1 0 265328 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hdll__or4bb_1  sky130_fd_sc_hdll__or4bb_1_0
timestamp 1627202621
transform 1 0 266524 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__or4bb_2  sky130_fd_sc_hdll__or4bb_2_0
timestamp 1627202621
transform 1 0 267536 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__or4bb_4  sky130_fd_sc_hdll__or4bb_4_0
timestamp 1627202621
transform 1 0 268640 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__sdfbbp_1  sky130_fd_sc_hdll__sdfbbp_1_0
timestamp 1627202621
transform 1 0 269928 0 1 0
box -38 -48 3166 592
use sky130_fd_sc_hdll__sdfrbp_1  sky130_fd_sc_hdll__sdfrbp_1_0
timestamp 1627202621
transform 1 0 273148 0 1 0
box -38 -48 2890 592
use sky130_fd_sc_hdll__sdfrbp_2  sky130_fd_sc_hdll__sdfrbp_2_0
timestamp 1627202621
transform 1 0 276092 0 1 0
box -38 -48 2982 592
use sky130_fd_sc_hdll__sdfrtn_1  sky130_fd_sc_hdll__sdfrtn_1_0
timestamp 1627202621
transform 1 0 279128 0 1 0
box -38 -48 2614 592
use sky130_fd_sc_hdll__sdfrtp_1  sky130_fd_sc_hdll__sdfrtp_1_0
timestamp 1627202621
transform 1 0 281796 0 1 0
box -38 -48 2614 592
use sky130_fd_sc_hdll__sdfrtp_2  sky130_fd_sc_hdll__sdfrtp_2_0
timestamp 1627202621
transform 1 0 284464 0 1 0
box -38 -48 2706 592
use sky130_fd_sc_hdll__sdfsbp_1  sky130_fd_sc_hdll__sdfsbp_1_0
timestamp 1627202621
transform 1 0 287224 0 1 0
box -38 -48 2982 592
use sky130_fd_sc_hdll__sdfsbp_2  sky130_fd_sc_hdll__sdfsbp_2_0
timestamp 1627202621
transform 1 0 290260 0 1 0
box -38 -48 3166 592
use sky130_fd_sc_hdll__sdfstp_1  sky130_fd_sc_hdll__sdfstp_1_0
timestamp 1627202621
transform 1 0 293480 0 1 0
box -38 -48 2706 592
use sky130_fd_sc_hdll__sdfstp_2  sky130_fd_sc_hdll__sdfstp_2_0
timestamp 1627202621
transform 1 0 296240 0 1 0
box -38 -48 2890 592
use sky130_fd_sc_hdll__sdfstp_4  sky130_fd_sc_hdll__sdfstp_4_0
timestamp 1627202621
transform 1 0 299184 0 1 0
box -38 -48 3074 592
use sky130_fd_sc_hdll__sdfxbp_1  sky130_fd_sc_hdll__sdfxbp_1_0
timestamp 1627202621
transform 1 0 302312 0 1 0
box -38 -48 2430 592
use sky130_fd_sc_hdll__sdfxbp_2  sky130_fd_sc_hdll__sdfxbp_2_0
timestamp 1627202621
transform 1 0 304796 0 1 0
box -38 -48 2706 592
use sky130_fd_sc_hdll__sdfxtp_1  sky130_fd_sc_hdll__sdfxtp_1_0
timestamp 1627202621
transform 1 0 307556 0 1 0
box -38 -48 2154 592
use sky130_fd_sc_hdll__sdfxtp_2  sky130_fd_sc_hdll__sdfxtp_2_0
timestamp 1627202621
transform 1 0 309764 0 1 0
box -38 -48 2246 592
use sky130_fd_sc_hdll__sdfxtp_4  sky130_fd_sc_hdll__sdfxtp_4_0
timestamp 1627202621
transform 1 0 312064 0 1 0
box -38 -48 2430 592
use sky130_fd_sc_hdll__sdlclkp_1  sky130_fd_sc_hdll__sdlclkp_1_0
timestamp 1627202621
transform 1 0 314548 0 1 0
box -38 -48 1510 592
use sky130_fd_sc_hdll__sdlclkp_2  sky130_fd_sc_hdll__sdlclkp_2_0
timestamp 1627202621
transform 1 0 316112 0 1 0
box -38 -48 1602 592
use sky130_fd_sc_hdll__sdlclkp_4  sky130_fd_sc_hdll__sdlclkp_4_0
timestamp 1627202621
transform 1 0 317768 0 1 0
box -38 -48 1878 592
use sky130_fd_sc_hdll__sedfxbp_1  sky130_fd_sc_hdll__sedfxbp_1_0
timestamp 1627202621
transform 1 0 319700 0 1 0
box -38 -48 3074 592
use sky130_fd_sc_hdll__sedfxbp_2  sky130_fd_sc_hdll__sedfxbp_2_0
timestamp 1627202621
transform 1 0 322828 0 1 0
box -38 -48 3350 592
use sky130_fd_sc_hdll__xnor2_1  sky130_fd_sc_hdll__xnor2_1_0
timestamp 1627202621
transform 1 0 326232 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__xnor2_2  sky130_fd_sc_hdll__xnor2_2_0
timestamp 1627202621
transform 1 0 327060 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__xnor2_4  sky130_fd_sc_hdll__xnor2_4_0
timestamp 1627202621
transform 1 0 328440 0 1 0
box -38 -48 2246 592
use sky130_fd_sc_hdll__xnor3_1  sky130_fd_sc_hdll__xnor3_1_0
timestamp 1627202621
transform 1 0 330740 0 1 0
box -38 -48 1878 592
use sky130_fd_sc_hdll__xnor3_2  sky130_fd_sc_hdll__xnor3_2_0
timestamp 1627202621
transform 1 0 332672 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hdll__xnor3_4  sky130_fd_sc_hdll__xnor3_4_0
timestamp 1627202621
transform 1 0 334696 0 1 0
box -38 -48 2154 592
use sky130_fd_sc_hdll__xor2_1  sky130_fd_sc_hdll__xor2_1_0
timestamp 1627202621
transform 1 0 336904 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__xor2_2  sky130_fd_sc_hdll__xor2_2_0
timestamp 1627202621
transform 1 0 337732 0 1 0
box -38 -48 1326 592
use sky130_fd_sc_hdll__xor2_4  sky130_fd_sc_hdll__xor2_4_0
timestamp 1627202621
transform 1 0 339112 0 1 0
box -38 -48 2246 592
use sky130_fd_sc_hdll__xor3_1  sky130_fd_sc_hdll__xor3_1_0
timestamp 1627202621
transform 1 0 341412 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hdll__xor3_2  sky130_fd_sc_hdll__xor3_2_0
timestamp 1627202621
transform 1 0 343436 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hdll__xor3_4  sky130_fd_sc_hdll__xor3_4_0
timestamp 1627202621
transform 1 0 345460 0 1 0
box -38 -48 2154 592
use sky130_fd_sc_hdll__sdfrtp_4  sky130_fd_sc_hdll__sdfrtp_4_0
timestamp 1627202621
transform 1 0 347668 0 1 0
box -38 -48 2890 592
use sky130_fd_sc_hdll__inputiso0n_1  sky130_fd_sc_hdll__inputiso0n_1_0
timestamp 1627202621
transform 1 0 350612 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__inputiso0p_1  sky130_fd_sc_hdll__inputiso0p_1_0
timestamp 1627202621
transform 1 0 351164 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__inputiso1n_1  sky130_fd_sc_hdll__inputiso1n_1_0
timestamp 1627202621
transform 1 0 351900 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__inputiso1p_1  sky130_fd_sc_hdll__inputiso1p_1_0
timestamp 1627202621
transform 1 0 352636 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__isobufsrc_1  sky130_fd_sc_hdll__isobufsrc_1_0
timestamp 1627202621
transform 1 0 353188 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hdll__isobufsrc_2  sky130_fd_sc_hdll__isobufsrc_2_0
timestamp 1627202621
transform 1 0 353740 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__isobufsrc_4  sky130_fd_sc_hdll__isobufsrc_4_0
timestamp 1627202621
transform 1 0 354568 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hdll__isobufsrc_8  sky130_fd_sc_hdll__isobufsrc_8_0
timestamp 1627202621
transform 1 0 355764 0 1 0
box -38 -48 1970 592
use sky130_fd_sc_hdll__isobufsrc_16  sky130_fd_sc_hdll__isobufsrc_16_0
timestamp 1627202621
transform 1 0 357788 0 1 0
box -38 -48 3718 592
use sky130_fd_sc_hdll__fill_8  sky130_fd_sc_hdll__fill_8_0
timestamp 1627202621
transform 1 0 365700 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__fill_4  sky130_fd_sc_hdll__fill_4_0
timestamp 1627202621
transform 1 0 365332 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hdll__fill_2  sky130_fd_sc_hdll__fill_2_0
timestamp 1627202621
transform 1 0 365148 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hdll__fill_1  sky130_fd_sc_hdll__fill_1_0
timestamp 1627202621
transform 1 0 365056 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__decap_12  sky130_fd_sc_hdll__decap_12_0
timestamp 1627202621
transform 1 0 363860 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hdll__decap_8  sky130_fd_sc_hdll__decap_8_0
timestamp 1627202621
transform 1 0 363032 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__decap_6  sky130_fd_sc_hdll__decap_6_0
timestamp 1627202621
transform 1 0 362388 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hdll__decap_4  sky130_fd_sc_hdll__decap_4_0
timestamp 1627202621
transform 1 0 361928 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hdll__decap_3  sky130_fd_sc_hdll__decap_3_0
timestamp 1627202621
transform 1 0 361560 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_0
timestamp 1627202621
transform 1 0 46828 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_1
timestamp 1627202621
transform 1 0 44896 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_2
timestamp 1627202621
transform 1 0 43240 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_3
timestamp 1627202621
transform 1 0 41584 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_4
timestamp 1627202621
transform 1 0 40112 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_5
timestamp 1627202621
transform 1 0 38640 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_6
timestamp 1627202621
transform 1 0 37260 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_7
timestamp 1627202621
transform 1 0 35880 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_8
timestamp 1627202621
transform 1 0 34592 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_9
timestamp 1627202621
transform 1 0 31740 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_10
timestamp 1627202621
transform 1 0 30452 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_11
timestamp 1627202621
transform 1 0 27140 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_12
timestamp 1627202621
transform 1 0 24564 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_13
timestamp 1627202621
transform 1 0 21344 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_14
timestamp 1627202621
transform 1 0 18860 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_15
timestamp 1627202621
transform 1 0 17480 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_16
timestamp 1627202621
transform 1 0 13708 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_17
timestamp 1627202621
transform 1 0 10304 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_18
timestamp 1627202621
transform 1 0 8372 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_19
timestamp 1627202621
transform 1 0 6624 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_20
timestamp 1627202621
transform 1 0 5612 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_21
timestamp 1627202621
transform 1 0 4232 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_22
timestamp 1627202621
transform 1 0 3036 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_23
timestamp 1627202621
transform 1 0 1380 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_24
timestamp 1627202621
transform 1 0 120520 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_25
timestamp 1627202621
transform 1 0 119784 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_26
timestamp 1627202621
transform 1 0 412712 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_27
timestamp 1627202621
transform 1 0 412712 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_28
timestamp 1627202621
transform 1 0 402224 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_29
timestamp 1627202621
transform 1 0 396980 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_30
timestamp 1627202621
transform 1 0 388424 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_31
timestamp 1627202621
transform 1 0 393484 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_32
timestamp 1627202621
transform 1 0 387136 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_33
timestamp 1627202621
transform 1 0 386032 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_34
timestamp 1627202621
transform 1 0 385020 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_35
timestamp 1627202621
transform 1 0 402224 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_36
timestamp 1627202621
transform 1 0 396980 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_37
timestamp 1627202621
transform 1 0 393484 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_38
timestamp 1627202621
transform 1 0 388424 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_39
timestamp 1627202621
transform 1 0 379776 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_40
timestamp 1627202621
transform 1 0 376280 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_41
timestamp 1627202621
transform 1 0 368368 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_42
timestamp 1627202621
transform 1 0 371036 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_43
timestamp 1627202621
transform 1 0 361836 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_44
timestamp 1627202621
transform 1 0 362296 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_45
timestamp 1627202621
transform 1 0 362940 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_46
timestamp 1627202621
transform 1 0 363768 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_47
timestamp 1627202621
transform 1 0 366436 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_48
timestamp 1627202621
transform 1 0 364964 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_49
timestamp 1627202621
transform 1 0 361468 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_50
timestamp 1627202621
transform 1 0 357696 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_51
timestamp 1627202621
transform 1 0 355672 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_52
timestamp 1627202621
transform 1 0 354476 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_53
timestamp 1627202621
transform 1 0 353648 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_54
timestamp 1627202621
transform 1 0 353096 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_55
timestamp 1627202621
transform 1 0 352544 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_56
timestamp 1627202621
transform 1 0 351808 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_57
timestamp 1627202621
transform 1 0 351072 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_58
timestamp 1627202621
transform 1 0 350520 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_59
timestamp 1627202621
transform 1 0 347576 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_60
timestamp 1627202621
transform 1 0 345368 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_61
timestamp 1627202621
transform 1 0 343344 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_62
timestamp 1627202621
transform 1 0 341320 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_63
timestamp 1627202621
transform 1 0 339020 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_64
timestamp 1627202621
transform 1 0 337640 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_65
timestamp 1627202621
transform 1 0 336812 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_66
timestamp 1627202621
transform 1 0 334604 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_67
timestamp 1627202621
transform 1 0 332580 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_68
timestamp 1627202621
transform 1 0 330648 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_69
timestamp 1627202621
transform 1 0 328348 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_70
timestamp 1627202621
transform 1 0 326968 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_71
timestamp 1627202621
transform 1 0 326140 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_72
timestamp 1627202621
transform 1 0 322736 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_73
timestamp 1627202621
transform 1 0 319608 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_74
timestamp 1627202621
transform 1 0 317676 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_75
timestamp 1627202621
transform 1 0 316020 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_76
timestamp 1627202621
transform 1 0 314456 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_77
timestamp 1627202621
transform 1 0 311972 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_78
timestamp 1627202621
transform 1 0 309672 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_79
timestamp 1627202621
transform 1 0 307464 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_80
timestamp 1627202621
transform 1 0 304704 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_81
timestamp 1627202621
transform 1 0 302220 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_82
timestamp 1627202621
transform 1 0 299092 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_83
timestamp 1627202621
transform 1 0 296148 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_84
timestamp 1627202621
transform 1 0 293388 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_85
timestamp 1627202621
transform 1 0 290168 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_86
timestamp 1627202621
transform 1 0 287132 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_87
timestamp 1627202621
transform 1 0 284372 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_88
timestamp 1627202621
transform 1 0 281704 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_89
timestamp 1627202621
transform 1 0 279036 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_90
timestamp 1627202621
transform 1 0 276000 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_91
timestamp 1627202621
transform 1 0 273056 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_92
timestamp 1627202621
transform 1 0 269836 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_93
timestamp 1627202621
transform 1 0 268548 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_94
timestamp 1627202621
transform 1 0 267444 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_95
timestamp 1627202621
transform 1 0 266432 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_96
timestamp 1627202621
transform 1 0 265236 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_97
timestamp 1627202621
transform 1 0 264316 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_98
timestamp 1627202621
transform 1 0 263396 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_99
timestamp 1627202621
transform 1 0 262384 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_100
timestamp 1627202621
transform 1 0 261556 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_101
timestamp 1627202621
transform 1 0 260820 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_102
timestamp 1627202621
transform 1 0 259808 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_103
timestamp 1627202621
transform 1 0 258980 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_104
timestamp 1627202621
transform 1 0 258152 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_105
timestamp 1627202621
transform 1 0 257140 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_106
timestamp 1627202621
transform 1 0 256404 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_107
timestamp 1627202621
transform 1 0 255760 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_108
timestamp 1627202621
transform 1 0 254748 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_109
timestamp 1627202621
transform 1 0 253920 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_110
timestamp 1627202621
transform 1 0 253184 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_111
timestamp 1627202621
transform 1 0 252356 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_112
timestamp 1627202621
transform 1 0 251712 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_113
timestamp 1627202621
transform 1 0 251160 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_114
timestamp 1627202621
transform 1 0 248860 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_115
timestamp 1627202621
transform 1 0 247480 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_116
timestamp 1627202621
transform 1 0 246744 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_117
timestamp 1627202621
transform 1 0 244904 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_118
timestamp 1627202621
transform 1 0 243800 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_119
timestamp 1627202621
transform 1 0 243156 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_120
timestamp 1627202621
transform 1 0 240856 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_121
timestamp 1627202621
transform 1 0 239568 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_122
timestamp 1627202621
transform 1 0 238740 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_123
timestamp 1627202621
transform 1 0 237084 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_124
timestamp 1627202621
transform 1 0 236072 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_125
timestamp 1627202621
transform 1 0 235152 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_126
timestamp 1627202621
transform 1 0 233404 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_127
timestamp 1627202621
transform 1 0 232300 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_128
timestamp 1627202621
transform 1 0 231656 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_129
timestamp 1627202621
transform 1 0 230184 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_130
timestamp 1627202621
transform 1 0 229264 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_131
timestamp 1627202621
transform 1 0 228436 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_132
timestamp 1627202621
transform 1 0 226228 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_133
timestamp 1627202621
transform 1 0 224940 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_134
timestamp 1627202621
transform 1 0 224112 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_135
timestamp 1627202621
transform 1 0 222456 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_136
timestamp 1627202621
transform 1 0 221444 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_137
timestamp 1627202621
transform 1 0 220524 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_138
timestamp 1627202621
transform 1 0 218960 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_139
timestamp 1627202621
transform 1 0 217948 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_140
timestamp 1627202621
transform 1 0 217212 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_141
timestamp 1627202621
transform 1 0 215832 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_142
timestamp 1627202621
transform 1 0 214912 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_143
timestamp 1627202621
transform 1 0 214084 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_144
timestamp 1627202621
transform 1 0 212704 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_145
timestamp 1627202621
transform 1 0 211876 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_146
timestamp 1627202621
transform 1 0 211324 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_147
timestamp 1627202621
transform 1 0 210036 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_148
timestamp 1627202621
transform 1 0 209208 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_149
timestamp 1627202621
transform 1 0 208472 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_150
timestamp 1627202621
transform 1 0 206632 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_151
timestamp 1627202621
transform 1 0 205528 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_152
timestamp 1627202621
transform 1 0 204884 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_153
timestamp 1627202621
transform 1 0 203412 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_154
timestamp 1627202621
transform 1 0 202492 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_155
timestamp 1627202621
transform 1 0 201572 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_156
timestamp 1627202621
transform 1 0 199456 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_157
timestamp 1627202621
transform 1 0 198076 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_158
timestamp 1627202621
transform 1 0 197156 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_159
timestamp 1627202621
transform 1 0 195132 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_160
timestamp 1627202621
transform 1 0 193844 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_161
timestamp 1627202621
transform 1 0 193016 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_162
timestamp 1627202621
transform 1 0 191176 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_163
timestamp 1627202621
transform 1 0 190072 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_164
timestamp 1627202621
transform 1 0 189428 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_165
timestamp 1627202621
transform 1 0 187864 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_166
timestamp 1627202621
transform 1 0 186760 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_167
timestamp 1627202621
transform 1 0 186116 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_168
timestamp 1627202621
transform 1 0 184736 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_169
timestamp 1627202621
transform 1 0 183816 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_170
timestamp 1627202621
transform 1 0 183264 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_171
timestamp 1627202621
transform 1 0 182068 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_172
timestamp 1627202621
transform 1 0 181240 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_173
timestamp 1627202621
transform 1 0 180688 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_174
timestamp 1627202621
transform 1 0 178940 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_175
timestamp 1627202621
transform 1 0 177928 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_176
timestamp 1627202621
transform 1 0 177284 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_177
timestamp 1627202621
transform 1 0 176824 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_178
timestamp 1627202621
transform 1 0 174616 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_179
timestamp 1627202621
transform 1 0 173236 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_180
timestamp 1627202621
transform 1 0 172316 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_181
timestamp 1627202621
transform 1 0 170292 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_182
timestamp 1627202621
transform 1 0 169004 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_183
timestamp 1627202621
transform 1 0 168268 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_184
timestamp 1627202621
transform 1 0 166428 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_185
timestamp 1627202621
transform 1 0 165324 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_186
timestamp 1627202621
transform 1 0 164680 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_187
timestamp 1627202621
transform 1 0 163024 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_188
timestamp 1627202621
transform 1 0 162012 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_189
timestamp 1627202621
transform 1 0 161368 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_190
timestamp 1627202621
transform 1 0 159896 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_191
timestamp 1627202621
transform 1 0 158976 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_192
timestamp 1627202621
transform 1 0 158424 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_193
timestamp 1627202621
transform 1 0 157228 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_194
timestamp 1627202621
transform 1 0 156492 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_195
timestamp 1627202621
transform 1 0 155940 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_196
timestamp 1627202621
transform 1 0 154192 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_197
timestamp 1627202621
transform 1 0 153180 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_198
timestamp 1627202621
transform 1 0 152536 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_199
timestamp 1627202621
transform 1 0 152076 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_200
timestamp 1627202621
transform 1 0 150144 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_201
timestamp 1627202621
transform 1 0 148948 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_202
timestamp 1627202621
transform 1 0 148028 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_203
timestamp 1627202621
transform 1 0 145820 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_204
timestamp 1627202621
transform 1 0 144532 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_205
timestamp 1627202621
transform 1 0 143520 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_206
timestamp 1627202621
transform 1 0 142508 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_207
timestamp 1627202621
transform 1 0 141496 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_208
timestamp 1627202621
transform 1 0 140668 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_209
timestamp 1627202621
transform 1 0 140024 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_210
timestamp 1627202621
transform 1 0 139564 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_211
timestamp 1627202621
transform 1 0 137816 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_212
timestamp 1627202621
transform 1 0 136436 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_213
timestamp 1627202621
transform 1 0 136068 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_214
timestamp 1627202621
transform 1 0 134136 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_215
timestamp 1627202621
transform 1 0 132940 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_216
timestamp 1627202621
transform 1 0 132112 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_217
timestamp 1627202621
transform 1 0 131468 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_218
timestamp 1627202621
transform 1 0 129536 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_219
timestamp 1627202621
transform 1 0 128340 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_220
timestamp 1627202621
transform 1 0 127512 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_221
timestamp 1627202621
transform 1 0 126868 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_222
timestamp 1627202621
transform 1 0 124568 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_223
timestamp 1627202621
transform 1 0 123188 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_224
timestamp 1627202621
transform 1 0 122176 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_225
timestamp 1627202621
transform 1 0 121348 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_226
timestamp 1627202621
transform 1 0 119048 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_227
timestamp 1627202621
transform 1 0 117484 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_228
timestamp 1627202621
transform 1 0 116104 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_229
timestamp 1627202621
transform 1 0 114816 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_230
timestamp 1627202621
transform 1 0 110124 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_231
timestamp 1627202621
transform 1 0 108008 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_232
timestamp 1627202621
transform 1 0 105616 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_233
timestamp 1627202621
transform 1 0 103500 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_234
timestamp 1627202621
transform 1 0 101476 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_235
timestamp 1627202621
transform 1 0 101108 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_236
timestamp 1627202621
transform 1 0 100464 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_237
timestamp 1627202621
transform 1 0 100004 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_238
timestamp 1627202621
transform 1 0 98624 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_239
timestamp 1627202621
transform 1 0 97796 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_240
timestamp 1627202621
transform 1 0 97244 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_241
timestamp 1627202621
transform 1 0 94668 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_242
timestamp 1627202621
transform 1 0 94208 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_243
timestamp 1627202621
transform 1 0 93012 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_244
timestamp 1627202621
transform 1 0 92276 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_245
timestamp 1627202621
transform 1 0 91724 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_246
timestamp 1627202621
transform 1 0 89608 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_247
timestamp 1627202621
transform 1 0 89148 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_248
timestamp 1627202621
transform 1 0 87676 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_249
timestamp 1627202621
transform 1 0 85100 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_250
timestamp 1627202621
transform 1 0 83536 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_251
timestamp 1627202621
transform 1 0 80776 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_252
timestamp 1627202621
transform 1 0 79488 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_253
timestamp 1627202621
transform 1 0 78476 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_254
timestamp 1627202621
transform 1 0 77740 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_255
timestamp 1627202621
transform 1 0 77188 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_256
timestamp 1627202621
transform 1 0 74796 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_257
timestamp 1627202621
transform 1 0 73048 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_258
timestamp 1627202621
transform 1 0 72588 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_259
timestamp 1627202621
transform 1 0 71208 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_260
timestamp 1627202621
transform 1 0 70104 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_261
timestamp 1627202621
transform 1 0 69092 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_262
timestamp 1627202621
transform 1 0 67988 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_263
timestamp 1627202621
transform 1 0 66976 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_264
timestamp 1627202621
transform 1 0 66056 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_265
timestamp 1627202621
transform 1 0 65044 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_266
timestamp 1627202621
transform 1 0 112332 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_267
timestamp 1627202621
transform 1 0 64216 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_268
timestamp 1627202621
transform 1 0 63480 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_269
timestamp 1627202621
transform 1 0 62376 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_270
timestamp 1627202621
transform 1 0 61456 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_271
timestamp 1627202621
transform 1 0 60628 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_272
timestamp 1627202621
transform 1 0 59616 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_273
timestamp 1627202621
transform 1 0 58880 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_274
timestamp 1627202621
transform 1 0 58236 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_275
timestamp 1627202621
transform 1 0 57316 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_276
timestamp 1627202621
transform 1 0 56488 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_277
timestamp 1627202621
transform 1 0 55752 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_278
timestamp 1627202621
transform 1 0 54924 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_279
timestamp 1627202621
transform 1 0 54280 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_280
timestamp 1627202621
transform 1 0 53728 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_281
timestamp 1627202621
transform 1 0 51336 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_282
timestamp 1627202621
transform 1 0 49956 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_283
timestamp 1627202621
transform 1 0 49220 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_284
timestamp 1627202621
transform 1 0 47472 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_285
timestamp 1627202621
transform 1 0 45540 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_286
timestamp 1627202621
transform 1 0 43700 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_287
timestamp 1627202621
transform 1 0 42596 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_288
timestamp 1627202621
transform 1 0 41952 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_289
timestamp 1627202621
transform 1 0 40480 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_290
timestamp 1627202621
transform 1 0 39652 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_291
timestamp 1627202621
transform 1 0 38916 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_292
timestamp 1627202621
transform 1 0 36708 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_293
timestamp 1627202621
transform 1 0 35420 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_294
timestamp 1627202621
transform 1 0 34592 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_295
timestamp 1627202621
transform 1 0 32936 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_296
timestamp 1627202621
transform 1 0 31924 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_297
timestamp 1627202621
transform 1 0 31004 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_298
timestamp 1627202621
transform 1 0 29164 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_299
timestamp 1627202621
transform 1 0 28060 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_300
timestamp 1627202621
transform 1 0 27324 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_301
timestamp 1627202621
transform 1 0 25852 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_302
timestamp 1627202621
transform 1 0 24932 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_303
timestamp 1627202621
transform 1 0 24104 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_304
timestamp 1627202621
transform 1 0 23184 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_305
timestamp 1627202621
transform 1 0 20976 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_306
timestamp 1627202621
transform 1 0 19688 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_307
timestamp 1627202621
transform 1 0 18860 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_308
timestamp 1627202621
transform 1 0 17480 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_309
timestamp 1627202621
transform 1 0 16652 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_310
timestamp 1627202621
transform 1 0 16100 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_311
timestamp 1627202621
transform 1 0 14812 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_312
timestamp 1627202621
transform 1 0 13984 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_313
timestamp 1627202621
transform 1 0 13248 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_314
timestamp 1627202621
transform 1 0 11684 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_315
timestamp 1627202621
transform 1 0 10672 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_316
timestamp 1627202621
transform 1 0 9936 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_317
timestamp 1627202621
transform 1 0 8556 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_318
timestamp 1627202621
transform 1 0 7636 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_319
timestamp 1627202621
transform 1 0 6716 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_320
timestamp 1627202621
transform 1 0 4968 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_321
timestamp 1627202621
transform 1 0 46460 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_322
timestamp 1627202621
transform 1 0 3864 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_323
timestamp 1627202621
transform 1 0 3220 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_324
timestamp 1627202621
transform 1 0 1656 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvpwrvgnd_1  sky130_fd_sc_hdll__tapvpwrvgnd_1_325
timestamp 1627202621
transform 1 0 736 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__tap_1  sky130_fd_sc_hdll__tap_1_0
timestamp 1627202621
transform 1 0 366528 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hdll__muxb4to1_1  sky130_fd_sc_hdll__muxb4to1_1_0
timestamp 1627202621
transform 1 0 366620 0 1 0
box -38 -48 1786 592
use sky130_fd_sc_hdll__muxb4to1_2  sky130_fd_sc_hdll__muxb4to1_2_0
timestamp 1627202621
transform 1 0 368460 0 1 0
box -38 -48 2614 592
use sky130_fd_sc_hdll__muxb4to1_4  sky130_fd_sc_hdll__muxb4to1_4_0
timestamp 1627202621
transform 1 0 371128 0 1 0
box -38 -48 5190 592
use sky130_fd_sc_hdll__muxb8to1_1  sky130_fd_sc_hdll__muxb8to1_1_0
timestamp 1627202621
transform 1 0 376372 0 1 0
box -38 -48 3442 592
use sky130_fd_sc_hdll__muxb8to1_2  sky130_fd_sc_hdll__muxb8to1_2_0
timestamp 1627202621
transform 1 0 379868 0 1 0
box -38 -48 5190 592
use sky130_fd_sc_hdll__muxb8to1_4  sky130_fd_sc_hdll__muxb8to1_4_0
timestamp 1627202621
transform 1 0 388516 0 1 0
box -38 -48 5006 1136
use sky130_fd_sc_hdll__muxb16to1_1  sky130_fd_sc_hdll__muxb16to1_1_0
timestamp 1627202621
transform 1 0 393576 0 1 0
box -38 -48 3442 1136
use sky130_fd_sc_hdll__muxb16to1_2  sky130_fd_sc_hdll__muxb16to1_2_0
timestamp 1627202621
transform 1 0 397072 0 1 0
box -38 -48 5190 1136
use sky130_fd_sc_hdll__muxb16to1_4  sky130_fd_sc_hdll__muxb16to1_4_0
timestamp 1627202621
transform 1 0 402316 0 1 0
box -38 -48 10434 1136
use sky130_fd_sc_hdll__clkmux2_1  sky130_fd_sc_hdll__clkmux2_1_0
timestamp 1627202621
transform 1 0 385112 0 1 0
box -38 -48 958 592
use sky130_fd_sc_hdll__clkmux2_2  sky130_fd_sc_hdll__clkmux2_2_0
timestamp 1627202621
transform 1 0 386124 0 1 0
box -38 -48 1050 592
use sky130_fd_sc_hdll__clkmux2_4  sky130_fd_sc_hdll__clkmux2_4_0
timestamp 1627202621
transform 1 0 387228 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hdll__dlygate4sd2_1  sky130_fd_sc_hdll__dlygate4sd2_1_0
timestamp 1627202621
transform 1 0 119876 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hdll__dlygate4sd3_1  sky130_fd_sc_hdll__dlygate4sd3_1_0
timestamp 1627202621
transform 1 0 120612 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hdll__a21o_6  sky130_fd_sc_hdll__a21o_6_0
timestamp 1627202621
transform 1 0 0 0 -1 1088
box -38 -48 1418 592
use sky130_fd_sc_hdll__a21o_8  sky130_fd_sc_hdll__a21o_8_0
timestamp 1627202621
transform 1 0 1472 0 -1 1088
box -38 -48 1602 592
use sky130_fd_sc_hdll__and2_6  sky130_fd_sc_hdll__and2_6_0
timestamp 1627202621
transform 1 0 3128 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hdll__and2_8  sky130_fd_sc_hdll__and2_8_0
timestamp 1627202621
transform 1 0 4324 0 -1 1088
box -38 -48 1326 592
use sky130_fd_sc_hdll__clkbuf_6  sky130_fd_sc_hdll__clkbuf_6_0
timestamp 1627202621
transform 1 0 5704 0 -1 1088
box -38 -48 958 592
use sky130_fd_sc_hdll__clkbuf_12  sky130_fd_sc_hdll__clkbuf_12_0
timestamp 1627202621
transform 1 0 6716 0 -1 1088
box -38 -48 1694 592
use sky130_fd_sc_hdll__clkinv_12  sky130_fd_sc_hdll__clkinv_12_0
timestamp 1627202621
transform 1 0 8464 0 -1 1088
box -38 -48 1878 592
use sky130_fd_sc_hdll__mux2_12  sky130_fd_sc_hdll__mux2_12_0
timestamp 1627202621
transform 1 0 10396 0 -1 1088
box -38 -48 3350 592
use sky130_fd_sc_hdll__mux2_16  sky130_fd_sc_hdll__mux2_16_0
timestamp 1627202621
transform 1 0 13800 0 -1 1088
box -38 -48 3718 592
use sky130_fd_sc_hdll__nand2_6  sky130_fd_sc_hdll__nand2_6_0
timestamp 1627202621
transform 1 0 17572 0 -1 1088
box -38 -48 1326 592
use sky130_fd_sc_hdll__nand2_12  sky130_fd_sc_hdll__nand2_12_0
timestamp 1627202621
transform 1 0 18952 0 -1 1088
box -38 -48 2430 592
use sky130_fd_sc_hdll__nand2_16  sky130_fd_sc_hdll__nand2_16_0
timestamp 1627202621
transform 1 0 21436 0 -1 1088
box -38 -48 3166 592
use sky130_fd_sc_hdll__nor4_6  sky130_fd_sc_hdll__nor4_6_0
timestamp 1627202621
transform 1 0 24656 0 -1 1088
box -38 -48 2522 592
use sky130_fd_sc_hdll__nor4_8  sky130_fd_sc_hdll__nor4_8_0
timestamp 1627202621
transform 1 0 27232 0 -1 1088
box -38 -48 3258 592
use sky130_fd_sc_hdll__or2_6  sky130_fd_sc_hdll__or2_6_0
timestamp 1627202621
transform 1 0 33396 0 -1 1088
box -38 -48 1234 592
use sky130_fd_sc_hdll__or2_8  sky130_fd_sc_hdll__or2_8_0
timestamp 1627202621
transform 1 0 31832 0 -1 1088
box -38 -48 1418 592
use sky130_fd_sc_hdll__tapvgnd_1  sky130_fd_sc_hdll__tapvgnd_1_0
timestamp 1627202621
transform 1 0 33212 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__tapvgnd2_1  sky130_fd_sc_hdll__tapvgnd2_1_0
timestamp 1627202621
transform 1 0 33304 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hdll__probe_p_8  sky130_fd_sc_hdll__probe_p_8_0
timestamp 1627202621
transform 1 0 30544 0 -1 1088
box -38 -48 1234 592
use sky130_fd_sc_hdll__probec_p_8  sky130_fd_sc_hdll__probec_p_8_0
timestamp 1627202621
transform 1 0 34684 0 -1 1088
box -252 -234 1335 778
use sky130_fd_sc_hdll__dlrtn_1  sky130_fd_sc_hdll__dlrtn_1_0
timestamp 1627202621
transform 1 0 35972 0 -1 1088
box -38 -48 1326 592
use sky130_fd_sc_hdll__dlrtp_1  sky130_fd_sc_hdll__dlrtp_1_0
timestamp 1627202621
transform 1 0 37352 0 -1 1088
box -38 -48 1326 592
use sky130_fd_sc_hdll__dlrtn_2  sky130_fd_sc_hdll__dlrtn_2_0
timestamp 1627202621
transform 1 0 38732 0 -1 1088
box -38 -48 1418 592
use sky130_fd_sc_hdll__dlrtp_2  sky130_fd_sc_hdll__dlrtp_2_0
timestamp 1627202621
transform 1 0 40204 0 -1 1088
box -38 -48 1418 592
use sky130_fd_sc_hdll__dlrtn_4  sky130_fd_sc_hdll__dlrtn_4_0
timestamp 1627202621
transform 1 0 41676 0 -1 1088
box -38 -48 1602 592
use sky130_fd_sc_hdll__dlrtp_4  sky130_fd_sc_hdll__dlrtp_4_0
timestamp 1627202621
transform 1 0 43332 0 -1 1088
box -38 -48 1602 592
use sky130_fd_sc_hdll__diode_2  sky130_fd_sc_hdll__diode_2_0
timestamp 1627202621
transform 1 0 44988 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hdll__diode_4  sky130_fd_sc_hdll__diode_4_0
timestamp 1627202621
transform 1 0 45172 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hdll__diode_6  sky130_fd_sc_hdll__diode_6_0
timestamp 1627202621
transform 1 0 45540 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hdll__diode_8  sky130_fd_sc_hdll__diode_8_0
timestamp 1627202621
transform 1 0 46092 0 -1 1088
box -38 -48 774 592
<< labels >>
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 1 nsew power default
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground default
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -2976 -3165 415786 3725
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3646290
string GDS_START 3609774
<< end >>
