magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 331 1478 704
<< pwell >>
rect 9 241 197 268
rect 9 49 1437 241
rect 0 0 1440 49
<< scnmos >>
rect 88 74 118 242
rect 278 47 308 215
rect 364 47 394 215
rect 450 47 480 215
rect 536 47 566 215
rect 622 47 652 215
rect 708 47 738 215
rect 794 47 824 215
rect 880 47 910 215
rect 1070 47 1100 215
rect 1156 47 1186 215
rect 1242 47 1272 215
rect 1328 47 1358 215
<< scpmoshvt >>
rect 143 367 173 619
rect 242 367 272 619
rect 328 367 358 619
rect 414 367 444 619
rect 500 367 530 619
rect 592 367 622 619
rect 678 367 708 619
rect 780 367 810 619
rect 866 367 896 619
rect 989 367 1019 619
rect 1075 367 1105 619
rect 1161 367 1191 619
rect 1247 367 1277 619
<< ndiff >>
rect 35 230 88 242
rect 35 196 43 230
rect 77 196 88 230
rect 35 122 88 196
rect 35 88 43 122
rect 77 88 88 122
rect 35 74 88 88
rect 118 134 171 242
rect 118 100 129 134
rect 163 100 171 134
rect 118 74 171 100
rect 225 124 278 215
rect 225 90 233 124
rect 267 90 278 124
rect 225 47 278 90
rect 308 169 364 215
rect 308 135 319 169
rect 353 135 364 169
rect 308 47 364 135
rect 394 161 450 215
rect 394 127 405 161
rect 439 127 450 161
rect 394 89 450 127
rect 394 55 405 89
rect 439 55 450 89
rect 394 47 450 55
rect 480 169 536 215
rect 480 135 491 169
rect 525 135 536 169
rect 480 47 536 135
rect 566 161 622 215
rect 566 127 577 161
rect 611 127 622 161
rect 566 89 622 127
rect 566 55 577 89
rect 611 55 622 89
rect 566 47 622 55
rect 652 173 708 215
rect 652 139 663 173
rect 697 139 708 173
rect 652 47 708 139
rect 738 157 794 215
rect 738 123 749 157
rect 783 123 794 157
rect 738 89 794 123
rect 738 55 749 89
rect 783 55 794 89
rect 738 47 794 55
rect 824 173 880 215
rect 824 139 835 173
rect 869 139 880 173
rect 824 47 880 139
rect 910 176 963 215
rect 910 142 921 176
rect 955 142 963 176
rect 910 93 963 142
rect 910 59 921 93
rect 955 59 963 93
rect 910 47 963 59
rect 1017 177 1070 215
rect 1017 143 1025 177
rect 1059 143 1070 177
rect 1017 93 1070 143
rect 1017 59 1025 93
rect 1059 59 1070 93
rect 1017 47 1070 59
rect 1100 207 1156 215
rect 1100 173 1111 207
rect 1145 173 1156 207
rect 1100 101 1156 173
rect 1100 67 1111 101
rect 1145 67 1156 101
rect 1100 47 1156 67
rect 1186 179 1242 215
rect 1186 145 1197 179
rect 1231 145 1242 179
rect 1186 89 1242 145
rect 1186 55 1197 89
rect 1231 55 1242 89
rect 1186 47 1242 55
rect 1272 207 1328 215
rect 1272 173 1283 207
rect 1317 173 1328 207
rect 1272 101 1328 173
rect 1272 67 1283 101
rect 1317 67 1328 101
rect 1272 47 1328 67
rect 1358 203 1411 215
rect 1358 169 1369 203
rect 1403 169 1411 203
rect 1358 93 1411 169
rect 1358 59 1369 93
rect 1403 59 1411 93
rect 1358 47 1411 59
<< pdiff >>
rect 90 599 143 619
rect 90 565 98 599
rect 132 565 143 599
rect 90 507 143 565
rect 90 473 98 507
rect 132 473 143 507
rect 90 418 143 473
rect 90 384 98 418
rect 132 384 143 418
rect 90 367 143 384
rect 173 611 242 619
rect 173 577 195 611
rect 229 577 242 611
rect 173 517 242 577
rect 173 483 195 517
rect 229 483 242 517
rect 173 427 242 483
rect 173 393 195 427
rect 229 393 242 427
rect 173 367 242 393
rect 272 599 328 619
rect 272 565 283 599
rect 317 565 328 599
rect 272 512 328 565
rect 272 478 283 512
rect 317 478 328 512
rect 272 409 328 478
rect 272 375 283 409
rect 317 375 328 409
rect 272 367 328 375
rect 358 611 414 619
rect 358 577 369 611
rect 403 577 414 611
rect 358 531 414 577
rect 358 497 369 531
rect 403 497 414 531
rect 358 457 414 497
rect 358 423 369 457
rect 403 423 414 457
rect 358 367 414 423
rect 444 599 500 619
rect 444 565 455 599
rect 489 565 500 599
rect 444 512 500 565
rect 444 478 455 512
rect 489 478 500 512
rect 444 409 500 478
rect 444 375 455 409
rect 489 375 500 409
rect 444 367 500 375
rect 530 573 592 619
rect 530 539 541 573
rect 575 539 592 573
rect 530 367 592 539
rect 622 599 678 619
rect 622 565 633 599
rect 667 565 678 599
rect 622 523 678 565
rect 622 489 633 523
rect 667 489 678 523
rect 622 436 678 489
rect 622 402 633 436
rect 667 402 678 436
rect 622 367 678 402
rect 708 611 780 619
rect 708 577 726 611
rect 760 577 780 611
rect 708 493 780 577
rect 708 459 726 493
rect 760 459 780 493
rect 708 367 780 459
rect 810 599 866 619
rect 810 565 821 599
rect 855 565 866 599
rect 810 523 866 565
rect 810 489 821 523
rect 855 489 866 523
rect 810 436 866 489
rect 810 402 821 436
rect 855 402 866 436
rect 810 367 866 402
rect 896 611 989 619
rect 896 577 923 611
rect 957 577 989 611
rect 896 492 989 577
rect 896 458 923 492
rect 957 458 989 492
rect 896 367 989 458
rect 1019 599 1075 619
rect 1019 565 1030 599
rect 1064 565 1075 599
rect 1019 523 1075 565
rect 1019 489 1030 523
rect 1064 489 1075 523
rect 1019 436 1075 489
rect 1019 402 1030 436
rect 1064 402 1075 436
rect 1019 367 1075 402
rect 1105 611 1161 619
rect 1105 577 1116 611
rect 1150 577 1161 611
rect 1105 494 1161 577
rect 1105 460 1116 494
rect 1150 460 1161 494
rect 1105 367 1161 460
rect 1191 599 1247 619
rect 1191 565 1202 599
rect 1236 565 1247 599
rect 1191 523 1247 565
rect 1191 489 1202 523
rect 1236 489 1247 523
rect 1191 436 1247 489
rect 1191 402 1202 436
rect 1236 402 1247 436
rect 1191 367 1247 402
rect 1277 607 1330 619
rect 1277 573 1288 607
rect 1322 573 1330 607
rect 1277 509 1330 573
rect 1277 475 1288 509
rect 1322 475 1330 509
rect 1277 420 1330 475
rect 1277 386 1288 420
rect 1322 386 1330 420
rect 1277 367 1330 386
<< ndiffc >>
rect 43 196 77 230
rect 43 88 77 122
rect 129 100 163 134
rect 233 90 267 124
rect 319 135 353 169
rect 405 127 439 161
rect 405 55 439 89
rect 491 135 525 169
rect 577 127 611 161
rect 577 55 611 89
rect 663 139 697 173
rect 749 123 783 157
rect 749 55 783 89
rect 835 139 869 173
rect 921 142 955 176
rect 921 59 955 93
rect 1025 143 1059 177
rect 1025 59 1059 93
rect 1111 173 1145 207
rect 1111 67 1145 101
rect 1197 145 1231 179
rect 1197 55 1231 89
rect 1283 173 1317 207
rect 1283 67 1317 101
rect 1369 169 1403 203
rect 1369 59 1403 93
<< pdiffc >>
rect 98 565 132 599
rect 98 473 132 507
rect 98 384 132 418
rect 195 577 229 611
rect 195 483 229 517
rect 195 393 229 427
rect 283 565 317 599
rect 283 478 317 512
rect 283 375 317 409
rect 369 577 403 611
rect 369 497 403 531
rect 369 423 403 457
rect 455 565 489 599
rect 455 478 489 512
rect 455 375 489 409
rect 541 539 575 573
rect 633 565 667 599
rect 633 489 667 523
rect 633 402 667 436
rect 726 577 760 611
rect 726 459 760 493
rect 821 565 855 599
rect 821 489 855 523
rect 821 402 855 436
rect 923 577 957 611
rect 923 458 957 492
rect 1030 565 1064 599
rect 1030 489 1064 523
rect 1030 402 1064 436
rect 1116 577 1150 611
rect 1116 460 1150 494
rect 1202 565 1236 599
rect 1202 489 1236 523
rect 1202 402 1236 436
rect 1288 573 1322 607
rect 1288 475 1322 509
rect 1288 386 1322 420
<< poly >>
rect 143 619 173 645
rect 242 619 272 645
rect 328 619 358 645
rect 414 619 444 645
rect 500 619 530 645
rect 592 619 622 645
rect 678 619 708 645
rect 780 619 810 645
rect 866 619 896 645
rect 989 619 1019 645
rect 1075 619 1105 645
rect 1161 619 1191 645
rect 1247 619 1277 645
rect 143 344 173 367
rect 88 330 173 344
rect 88 314 170 330
rect 88 280 120 314
rect 154 280 170 314
rect 242 313 272 367
rect 328 313 358 367
rect 414 313 444 367
rect 500 313 530 367
rect 592 345 622 367
rect 678 345 708 367
rect 780 345 810 367
rect 866 345 896 367
rect 592 319 947 345
rect 592 315 693 319
rect 88 264 170 280
rect 212 297 550 313
rect 88 242 118 264
rect 212 263 228 297
rect 262 263 296 297
rect 330 263 364 297
rect 398 263 432 297
rect 466 263 500 297
rect 534 267 550 297
rect 622 285 693 315
rect 727 285 761 319
rect 795 285 829 319
rect 863 285 897 319
rect 931 285 947 319
rect 622 269 947 285
rect 989 335 1019 367
rect 1075 335 1105 367
rect 1161 335 1191 367
rect 1247 335 1277 367
rect 989 319 1396 335
rect 989 285 1006 319
rect 1040 285 1074 319
rect 1108 285 1142 319
rect 1176 285 1210 319
rect 1244 285 1278 319
rect 1312 285 1346 319
rect 1380 285 1396 319
rect 989 269 1396 285
rect 534 263 566 267
rect 212 237 566 263
rect 278 215 308 237
rect 364 215 394 237
rect 450 215 480 237
rect 536 215 566 237
rect 622 215 652 269
rect 708 215 738 269
rect 794 215 824 269
rect 880 215 910 269
rect 1070 215 1100 269
rect 1156 215 1186 269
rect 1242 215 1272 269
rect 1328 215 1358 269
rect 88 48 118 74
rect 278 21 308 47
rect 364 21 394 47
rect 450 21 480 47
rect 536 21 566 47
rect 622 21 652 47
rect 708 21 738 47
rect 794 21 824 47
rect 880 21 910 47
rect 1070 21 1100 47
rect 1156 21 1186 47
rect 1242 21 1272 47
rect 1328 21 1358 47
<< polycont >>
rect 120 280 154 314
rect 228 263 262 297
rect 296 263 330 297
rect 364 263 398 297
rect 432 263 466 297
rect 500 263 534 297
rect 693 285 727 319
rect 761 285 795 319
rect 829 285 863 319
rect 897 285 931 319
rect 1006 285 1040 319
rect 1074 285 1108 319
rect 1142 285 1176 319
rect 1210 285 1244 319
rect 1278 285 1312 319
rect 1346 285 1380 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 27 599 148 615
rect 27 565 98 599
rect 132 565 148 599
rect 27 507 148 565
rect 27 473 98 507
rect 132 473 148 507
rect 27 418 148 473
rect 27 384 98 418
rect 132 384 148 418
rect 182 611 237 649
rect 182 577 195 611
rect 229 577 237 611
rect 182 517 237 577
rect 182 483 195 517
rect 229 483 237 517
rect 182 427 237 483
rect 182 393 195 427
rect 229 393 237 427
rect 27 230 81 384
rect 182 377 237 393
rect 271 599 319 615
rect 271 565 283 599
rect 317 565 319 599
rect 271 512 319 565
rect 271 478 283 512
rect 317 478 319 512
rect 271 409 319 478
rect 353 611 419 649
rect 353 577 369 611
rect 403 577 419 611
rect 353 531 419 577
rect 353 497 369 531
rect 403 497 419 531
rect 353 457 419 497
rect 353 423 369 457
rect 403 423 419 457
rect 453 599 491 615
rect 453 565 455 599
rect 489 565 491 599
rect 453 512 491 565
rect 525 573 591 649
rect 525 539 541 573
rect 575 539 591 573
rect 525 532 591 539
rect 629 599 676 615
rect 629 565 633 599
rect 667 565 676 599
rect 453 478 455 512
rect 489 498 491 512
rect 629 523 676 565
rect 629 498 633 523
rect 489 489 633 498
rect 667 489 676 523
rect 489 478 676 489
rect 453 436 676 478
rect 710 611 776 649
rect 710 577 726 611
rect 760 577 776 611
rect 710 493 776 577
rect 710 459 726 493
rect 760 459 776 493
rect 710 454 776 459
rect 810 599 873 615
rect 810 565 821 599
rect 855 565 873 599
rect 810 523 873 565
rect 810 489 821 523
rect 855 489 873 523
rect 271 375 283 409
rect 317 389 319 409
rect 453 409 633 436
rect 453 389 455 409
rect 317 375 455 389
rect 489 402 633 409
rect 667 420 676 436
rect 810 436 873 489
rect 907 611 973 649
rect 907 577 923 611
rect 957 577 973 611
rect 907 492 973 577
rect 907 458 923 492
rect 957 458 973 492
rect 907 454 973 458
rect 1007 599 1066 615
rect 1007 565 1030 599
rect 1064 565 1066 599
rect 1007 523 1066 565
rect 1007 489 1030 523
rect 1064 489 1066 523
rect 810 420 821 436
rect 667 402 821 420
rect 855 420 873 436
rect 1007 436 1066 489
rect 1100 611 1166 649
rect 1100 577 1116 611
rect 1150 577 1166 611
rect 1100 494 1166 577
rect 1100 460 1116 494
rect 1150 460 1166 494
rect 1100 454 1166 460
rect 1200 599 1238 615
rect 1200 565 1202 599
rect 1236 565 1238 599
rect 1200 523 1238 565
rect 1200 489 1202 523
rect 1236 489 1238 523
rect 1007 420 1030 436
rect 855 402 1030 420
rect 1064 420 1066 436
rect 1200 436 1238 489
rect 1200 420 1202 436
rect 1064 402 1202 420
rect 1236 402 1238 436
rect 489 386 1238 402
rect 1272 607 1338 649
rect 1272 573 1288 607
rect 1322 573 1338 607
rect 1272 509 1338 573
rect 1272 475 1288 509
rect 1322 475 1338 509
rect 1272 420 1338 475
rect 1272 386 1288 420
rect 1322 386 1338 420
rect 489 375 641 386
rect 120 314 161 350
rect 271 338 641 375
rect 154 280 161 314
rect 120 242 161 280
rect 195 297 550 304
rect 195 263 228 297
rect 262 263 296 297
rect 330 263 364 297
rect 398 263 432 297
rect 466 263 500 297
rect 534 263 550 297
rect 27 196 43 230
rect 77 208 81 230
rect 195 208 264 263
rect 584 242 641 338
rect 677 319 947 352
rect 677 285 693 319
rect 727 285 761 319
rect 795 285 829 319
rect 863 285 897 319
rect 931 285 947 319
rect 677 281 947 285
rect 990 319 1409 352
rect 990 285 1006 319
rect 1040 285 1074 319
rect 1108 285 1142 319
rect 1176 285 1210 319
rect 1244 285 1278 319
rect 1312 285 1346 319
rect 1380 285 1409 319
rect 990 281 1409 285
rect 584 229 618 242
rect 77 196 264 208
rect 27 174 264 196
rect 303 195 618 229
rect 675 217 1326 247
rect 666 213 1326 217
rect 27 122 79 174
rect 303 169 355 195
rect 27 88 43 122
rect 77 88 79 122
rect 27 72 79 88
rect 113 134 179 140
rect 113 100 129 134
rect 163 100 179 134
rect 113 17 179 100
rect 217 124 269 140
rect 217 90 233 124
rect 267 90 269 124
rect 303 135 319 169
rect 353 135 355 169
rect 489 169 527 195
rect 303 119 355 135
rect 389 127 405 161
rect 439 127 455 161
rect 217 85 269 90
rect 389 89 455 127
rect 489 135 491 169
rect 525 135 527 169
rect 661 191 871 213
rect 661 173 699 191
rect 489 119 527 135
rect 561 127 577 161
rect 611 127 627 161
rect 389 85 405 89
rect 217 55 405 85
rect 439 85 455 89
rect 561 89 627 127
rect 661 139 663 173
rect 697 139 699 173
rect 833 173 871 191
rect 1109 207 1147 213
rect 661 123 699 139
rect 733 123 749 157
rect 783 123 799 157
rect 833 139 835 173
rect 869 139 871 173
rect 833 123 871 139
rect 905 176 971 179
rect 905 142 921 176
rect 955 142 971 176
rect 733 89 799 123
rect 905 93 971 142
rect 905 89 921 93
rect 561 85 577 89
rect 439 55 577 85
rect 611 55 749 89
rect 783 59 921 89
rect 955 59 971 93
rect 783 55 971 59
rect 217 51 971 55
rect 1009 143 1025 177
rect 1059 143 1075 177
rect 1009 93 1075 143
rect 1009 59 1025 93
rect 1059 59 1075 93
rect 1009 17 1075 59
rect 1109 173 1111 207
rect 1145 173 1147 207
rect 1281 207 1326 213
rect 1109 101 1147 173
rect 1109 67 1111 101
rect 1145 67 1147 101
rect 1109 51 1147 67
rect 1181 145 1197 179
rect 1231 145 1247 179
rect 1181 89 1247 145
rect 1181 55 1197 89
rect 1231 55 1247 89
rect 1181 17 1247 55
rect 1281 173 1283 207
rect 1317 173 1326 207
rect 1281 101 1326 173
rect 1281 67 1283 101
rect 1317 67 1326 101
rect 1281 51 1326 67
rect 1360 203 1419 219
rect 1360 169 1369 203
rect 1403 169 1419 203
rect 1360 93 1419 169
rect 1360 59 1369 93
rect 1403 59 1419 93
rect 1360 17 1419 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand3b_4
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3722990
string GDS_START 3710136
<< end >>
