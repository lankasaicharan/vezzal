magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 4082 1975
<< nwell >>
rect -38 449 2822 704
rect -38 335 426 449
rect -38 332 207 335
rect 1040 332 2822 449
rect 2047 316 2477 332
<< pwell >>
rect 676 314 998 342
rect 217 191 417 293
rect 647 272 998 314
rect 647 259 1414 272
rect 647 191 1775 259
rect 217 184 1775 191
rect 2131 184 2783 248
rect 44 49 2783 184
rect 0 0 2784 49
<< scpmos >>
rect 106 392 142 476
rect 196 392 232 476
rect 298 392 334 592
rect 497 485 533 569
rect 650 485 686 569
rect 728 485 764 569
rect 818 485 854 569
rect 1151 368 1187 592
rect 1311 368 1347 592
rect 1586 389 1622 589
rect 1722 389 1758 473
rect 1806 389 1842 473
rect 1936 389 1972 473
rect 2026 389 2062 473
rect 2133 352 2169 576
rect 2223 352 2259 576
rect 2330 352 2366 552
rect 2565 368 2601 592
rect 2655 368 2691 592
<< nmoslvt >>
rect 126 74 156 158
rect 198 74 228 158
rect 304 119 334 267
rect 752 232 782 316
rect 838 232 868 316
rect 506 81 536 165
rect 584 81 614 165
rect 1080 98 1110 246
rect 1301 98 1331 246
rect 1556 149 1586 233
rect 1651 85 1681 233
rect 1858 74 1888 158
rect 1944 74 1974 158
rect 2016 74 2046 158
rect 2214 74 2244 222
rect 2300 74 2330 222
rect 2395 74 2425 202
rect 2587 74 2617 222
rect 2673 74 2703 222
<< ndiff >>
rect 243 158 304 267
rect 70 128 126 158
rect 70 94 81 128
rect 115 94 126 128
rect 70 74 126 94
rect 156 74 198 158
rect 228 146 304 158
rect 228 112 245 146
rect 279 119 304 146
rect 334 255 391 267
rect 334 221 345 255
rect 379 221 391 255
rect 334 165 391 221
rect 702 288 752 316
rect 673 277 752 288
rect 673 243 689 277
rect 723 243 752 277
rect 673 232 752 243
rect 782 305 838 316
rect 782 271 793 305
rect 827 271 838 305
rect 782 232 838 271
rect 868 291 972 316
rect 868 257 929 291
rect 963 257 972 291
rect 868 232 972 257
rect 1026 234 1080 246
rect 334 131 345 165
rect 379 131 391 165
rect 334 119 391 131
rect 445 140 506 165
rect 279 112 289 119
rect 228 74 289 112
rect 445 106 457 140
rect 491 106 506 140
rect 445 81 506 106
rect 536 81 584 165
rect 614 153 675 165
rect 614 119 625 153
rect 659 119 675 153
rect 614 81 675 119
rect 1026 200 1035 234
rect 1069 200 1080 234
rect 1026 98 1080 200
rect 1110 98 1301 246
rect 1331 177 1388 246
rect 1331 143 1342 177
rect 1376 143 1388 177
rect 1499 208 1556 233
rect 1499 174 1511 208
rect 1545 174 1556 208
rect 1499 149 1556 174
rect 1586 221 1651 233
rect 1586 187 1601 221
rect 1635 187 1651 221
rect 1586 149 1651 187
rect 1331 98 1388 143
rect 1125 82 1183 98
rect 1125 48 1137 82
rect 1171 48 1183 82
rect 1601 85 1651 149
rect 1681 85 1749 233
rect 2157 204 2214 222
rect 2157 170 2169 204
rect 2203 170 2214 204
rect 1125 36 1183 48
rect 1696 51 1706 85
rect 1740 51 1749 85
rect 1803 128 1858 158
rect 1803 94 1813 128
rect 1847 94 1858 128
rect 1803 74 1858 94
rect 1888 128 1944 158
rect 1888 94 1899 128
rect 1933 94 1944 128
rect 1888 74 1944 94
rect 1974 74 2016 158
rect 2046 128 2103 158
rect 2046 94 2057 128
rect 2091 94 2103 128
rect 2046 74 2103 94
rect 2157 120 2214 170
rect 2157 86 2169 120
rect 2203 86 2214 120
rect 2157 74 2214 86
rect 2244 204 2300 222
rect 2244 170 2255 204
rect 2289 170 2300 204
rect 2244 120 2300 170
rect 2244 86 2255 120
rect 2289 86 2300 120
rect 2244 74 2300 86
rect 2330 202 2380 222
rect 2533 210 2587 222
rect 2330 120 2395 202
rect 2330 86 2342 120
rect 2376 86 2395 120
rect 2330 74 2395 86
rect 2425 190 2479 202
rect 2425 156 2436 190
rect 2470 156 2479 190
rect 2425 120 2479 156
rect 2425 86 2436 120
rect 2470 86 2479 120
rect 2425 74 2479 86
rect 2533 176 2542 210
rect 2576 176 2587 210
rect 2533 120 2587 176
rect 2533 86 2542 120
rect 2576 86 2587 120
rect 2533 74 2587 86
rect 2617 207 2673 222
rect 2617 173 2628 207
rect 2662 173 2673 207
rect 2617 116 2673 173
rect 2617 82 2628 116
rect 2662 82 2673 116
rect 2617 74 2673 82
rect 2703 210 2757 222
rect 2703 176 2714 210
rect 2748 176 2757 210
rect 2703 120 2757 176
rect 2703 86 2714 120
rect 2748 86 2757 120
rect 2703 74 2757 86
rect 1696 39 1749 51
<< pdiff >>
rect 27 627 283 639
rect 27 593 39 627
rect 73 593 138 627
rect 172 593 237 627
rect 271 593 283 627
rect 27 592 283 593
rect 27 562 298 592
rect 248 476 298 562
rect 40 451 106 476
rect 40 417 52 451
rect 86 417 106 451
rect 40 392 106 417
rect 142 452 196 476
rect 142 418 152 452
rect 186 418 196 452
rect 142 392 196 418
rect 232 392 298 476
rect 334 491 390 592
rect 577 575 635 586
rect 577 569 589 575
rect 334 457 344 491
rect 378 457 390 491
rect 444 531 497 569
rect 444 497 453 531
rect 487 497 497 531
rect 444 485 497 497
rect 533 541 589 569
rect 623 569 635 575
rect 1202 592 1296 599
rect 1095 580 1151 592
rect 623 541 650 569
rect 533 485 650 541
rect 686 485 728 569
rect 764 531 818 569
rect 764 497 774 531
rect 808 497 818 531
rect 764 485 818 497
rect 854 547 984 569
rect 854 513 874 547
rect 908 513 942 547
rect 976 513 984 547
rect 854 485 984 513
rect 1095 546 1107 580
rect 1141 546 1151 580
rect 1095 499 1151 546
rect 334 392 390 457
rect 1095 465 1107 499
rect 1141 465 1151 499
rect 1095 418 1151 465
rect 1095 384 1107 418
rect 1141 384 1151 418
rect 1095 368 1151 384
rect 1187 587 1311 592
rect 1187 553 1232 587
rect 1266 553 1311 587
rect 1187 368 1311 553
rect 1347 426 1403 592
rect 1533 531 1586 589
rect 1533 497 1542 531
rect 1576 497 1586 531
rect 1533 435 1586 497
rect 1347 392 1357 426
rect 1391 392 1403 426
rect 1347 368 1403 392
rect 1533 401 1542 435
rect 1576 401 1586 435
rect 1533 389 1586 401
rect 1622 473 1672 589
rect 2499 580 2565 592
rect 2077 560 2133 576
rect 2077 526 2089 560
rect 2123 526 2133 560
rect 1857 508 1921 520
rect 1857 474 1872 508
rect 1906 474 1921 508
rect 1857 473 1921 474
rect 2077 492 2133 526
rect 2077 473 2089 492
rect 1622 448 1722 473
rect 1622 414 1678 448
rect 1712 414 1722 448
rect 1622 389 1722 414
rect 1758 389 1806 473
rect 1842 389 1936 473
rect 1972 450 2026 473
rect 1972 416 1982 450
rect 2016 416 2026 450
rect 1972 389 2026 416
rect 2062 458 2089 473
rect 2123 458 2133 492
rect 2062 389 2133 458
rect 2083 352 2133 389
rect 2169 564 2223 576
rect 2169 530 2179 564
rect 2213 530 2223 564
rect 2169 484 2223 530
rect 2169 450 2179 484
rect 2213 450 2223 484
rect 2169 404 2223 450
rect 2169 370 2179 404
rect 2213 370 2223 404
rect 2169 352 2223 370
rect 2259 564 2315 576
rect 2259 530 2269 564
rect 2303 552 2315 564
rect 2303 530 2330 552
rect 2259 472 2330 530
rect 2259 438 2269 472
rect 2303 438 2330 472
rect 2259 398 2330 438
rect 2259 364 2269 398
rect 2303 364 2330 398
rect 2259 352 2330 364
rect 2366 540 2441 552
rect 2366 506 2395 540
rect 2429 506 2441 540
rect 2366 469 2441 506
rect 2366 435 2395 469
rect 2429 435 2441 469
rect 2366 398 2441 435
rect 2366 364 2395 398
rect 2429 364 2441 398
rect 2499 546 2511 580
rect 2545 546 2565 580
rect 2499 497 2565 546
rect 2499 463 2511 497
rect 2545 463 2565 497
rect 2499 414 2565 463
rect 2499 380 2511 414
rect 2545 380 2565 414
rect 2499 368 2565 380
rect 2601 580 2655 592
rect 2601 546 2611 580
rect 2645 546 2655 580
rect 2601 497 2655 546
rect 2601 463 2611 497
rect 2645 463 2655 497
rect 2601 414 2655 463
rect 2601 380 2611 414
rect 2645 380 2655 414
rect 2601 368 2655 380
rect 2691 580 2757 592
rect 2691 546 2711 580
rect 2745 546 2757 580
rect 2691 497 2757 546
rect 2691 463 2711 497
rect 2745 463 2757 497
rect 2691 414 2757 463
rect 2691 380 2711 414
rect 2745 380 2757 414
rect 2691 368 2757 380
rect 2366 352 2441 364
<< ndiffc >>
rect 81 94 115 128
rect 245 112 279 146
rect 345 221 379 255
rect 689 243 723 277
rect 793 271 827 305
rect 929 257 963 291
rect 345 131 379 165
rect 457 106 491 140
rect 625 119 659 153
rect 1035 200 1069 234
rect 1342 143 1376 177
rect 1511 174 1545 208
rect 1601 187 1635 221
rect 1137 48 1171 82
rect 2169 170 2203 204
rect 1706 51 1740 85
rect 1813 94 1847 128
rect 1899 94 1933 128
rect 2057 94 2091 128
rect 2169 86 2203 120
rect 2255 170 2289 204
rect 2255 86 2289 120
rect 2342 86 2376 120
rect 2436 156 2470 190
rect 2436 86 2470 120
rect 2542 176 2576 210
rect 2542 86 2576 120
rect 2628 173 2662 207
rect 2628 82 2662 116
rect 2714 176 2748 210
rect 2714 86 2748 120
<< pdiffc >>
rect 39 593 73 627
rect 138 593 172 627
rect 237 593 271 627
rect 52 417 86 451
rect 152 418 186 452
rect 344 457 378 491
rect 453 497 487 531
rect 589 541 623 575
rect 774 497 808 531
rect 874 513 908 547
rect 942 513 976 547
rect 1107 546 1141 580
rect 1107 465 1141 499
rect 1107 384 1141 418
rect 1232 553 1266 587
rect 1542 497 1576 531
rect 1357 392 1391 426
rect 1542 401 1576 435
rect 2089 526 2123 560
rect 1872 474 1906 508
rect 1678 414 1712 448
rect 1982 416 2016 450
rect 2089 458 2123 492
rect 2179 530 2213 564
rect 2179 450 2213 484
rect 2179 370 2213 404
rect 2269 530 2303 564
rect 2269 438 2303 472
rect 2269 364 2303 398
rect 2395 506 2429 540
rect 2395 435 2429 469
rect 2395 364 2429 398
rect 2511 546 2545 580
rect 2511 463 2545 497
rect 2511 380 2545 414
rect 2611 546 2645 580
rect 2611 463 2645 497
rect 2611 380 2645 414
rect 2711 546 2745 580
rect 2711 463 2745 497
rect 2711 380 2745 414
<< poly >>
rect 298 592 334 618
rect 106 476 142 502
rect 196 476 232 502
rect 497 569 533 595
rect 650 569 686 595
rect 728 569 764 595
rect 818 569 854 595
rect 1151 592 1187 618
rect 1311 592 1347 618
rect 106 314 142 392
rect 196 356 232 392
rect 298 360 334 392
rect 44 298 142 314
rect 44 264 60 298
rect 94 264 142 298
rect 190 340 256 356
rect 190 306 206 340
rect 240 306 256 340
rect 190 290 256 306
rect 298 344 431 360
rect 497 355 533 485
rect 650 369 686 485
rect 298 310 381 344
rect 415 310 431 344
rect 298 294 431 310
rect 477 339 543 355
rect 477 305 493 339
rect 527 305 543 339
rect 44 230 142 264
rect 44 196 60 230
rect 94 210 142 230
rect 94 196 156 210
rect 44 180 156 196
rect 126 158 156 180
rect 198 158 228 290
rect 304 267 334 294
rect 477 289 543 305
rect 585 353 686 369
rect 585 319 601 353
rect 635 319 686 353
rect 728 361 764 485
rect 818 448 854 485
rect 818 432 1063 448
rect 818 418 945 432
rect 728 331 782 361
rect 585 303 686 319
rect 752 316 782 331
rect 838 316 868 418
rect 929 398 945 418
rect 979 398 1013 432
rect 1047 398 1063 432
rect 929 382 1063 398
rect 1586 589 1622 615
rect 1435 418 1501 434
rect 1435 384 1451 418
rect 1485 384 1501 418
rect 2133 576 2169 602
rect 2223 576 2259 602
rect 2565 592 2601 618
rect 2655 592 2691 618
rect 1722 473 1758 499
rect 1806 473 1842 499
rect 1936 473 1972 499
rect 2026 473 2062 499
rect 1435 374 1501 384
rect 1586 374 1622 389
rect 1151 334 1187 368
rect 1311 334 1347 368
rect 1435 344 1622 374
rect 1080 318 1253 334
rect 506 165 536 289
rect 591 210 621 303
rect 1080 284 1135 318
rect 1169 284 1203 318
rect 1237 284 1253 318
rect 1311 318 1393 334
rect 1311 298 1343 318
rect 1080 268 1253 284
rect 1301 284 1343 298
rect 1377 284 1393 318
rect 1301 268 1393 284
rect 1080 246 1110 268
rect 1301 246 1331 268
rect 584 180 621 210
rect 584 165 614 180
rect 304 93 334 119
rect 752 83 782 232
rect 838 206 868 232
rect 1556 233 1586 344
rect 1722 321 1758 389
rect 1806 357 1842 389
rect 1658 305 1758 321
rect 1658 285 1674 305
rect 1651 271 1674 285
rect 1708 271 1758 305
rect 1800 341 1866 357
rect 1936 356 1972 389
rect 1800 307 1816 341
rect 1850 307 1866 341
rect 1800 291 1866 307
rect 1908 340 1974 356
rect 1908 306 1924 340
rect 1958 306 1974 340
rect 1651 255 1758 271
rect 1651 233 1681 255
rect 1556 123 1586 149
rect 1080 83 1110 98
rect 126 48 156 74
rect 198 51 228 74
rect 506 51 536 81
rect 584 55 614 81
rect 752 53 1110 83
rect 198 21 536 51
rect 1301 72 1331 98
rect 1830 203 1860 291
rect 1908 290 1974 306
rect 1830 173 1888 203
rect 1858 158 1888 173
rect 1944 158 1974 290
rect 2026 320 2062 389
rect 2330 552 2366 578
rect 2133 320 2169 352
rect 2223 320 2259 352
rect 2330 320 2366 352
rect 2565 326 2601 368
rect 2655 326 2691 368
rect 2026 267 2425 320
rect 2016 237 2425 267
rect 2527 310 2691 326
rect 2527 276 2543 310
rect 2577 290 2691 310
rect 2577 276 2703 290
rect 2527 260 2703 276
rect 2016 203 2032 237
rect 2066 203 2082 237
rect 2214 222 2244 237
rect 2300 222 2330 237
rect 2016 187 2082 203
rect 2016 158 2046 187
rect 1651 59 1681 85
rect 2395 202 2425 237
rect 2587 222 2617 260
rect 2673 222 2703 260
rect 1858 48 1888 74
rect 1944 48 1974 74
rect 2016 48 2046 74
rect 2214 48 2244 74
rect 2300 48 2330 74
rect 2395 48 2425 74
rect 2587 48 2617 74
rect 2673 48 2703 74
<< polycont >>
rect 60 264 94 298
rect 206 306 240 340
rect 381 310 415 344
rect 493 305 527 339
rect 60 196 94 230
rect 601 319 635 353
rect 945 398 979 432
rect 1013 398 1047 432
rect 1451 384 1485 418
rect 1135 284 1169 318
rect 1203 284 1237 318
rect 1343 284 1377 318
rect 1674 271 1708 305
rect 1816 307 1850 341
rect 1924 306 1958 340
rect 2543 276 2577 310
rect 2032 203 2066 237
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 23 627 287 649
rect 23 593 39 627
rect 73 593 138 627
rect 172 593 237 627
rect 271 593 287 627
rect 23 451 102 593
rect 321 581 555 615
rect 321 559 355 581
rect 23 417 52 451
rect 86 417 102 451
rect 23 388 102 417
rect 136 525 355 559
rect 437 531 487 547
rect 136 452 202 525
rect 437 497 453 531
rect 136 418 152 452
rect 186 418 202 452
rect 136 390 202 418
rect 297 457 344 491
rect 378 457 394 491
rect 25 298 103 314
rect 25 264 60 298
rect 94 264 103 298
rect 25 230 103 264
rect 25 196 60 230
rect 94 196 103 230
rect 25 162 103 196
rect 137 128 171 390
rect 205 350 263 356
rect 205 340 223 350
rect 205 306 206 340
rect 257 316 263 350
rect 240 306 263 316
rect 205 290 263 306
rect 297 260 331 457
rect 437 423 487 497
rect 521 491 555 581
rect 589 575 639 649
rect 623 541 639 575
rect 589 525 639 541
rect 673 581 892 615
rect 673 491 707 581
rect 858 563 892 581
rect 1085 580 1157 596
rect 858 547 992 563
rect 521 457 707 491
rect 758 531 824 547
rect 758 497 774 531
rect 808 497 824 531
rect 758 423 824 497
rect 858 513 874 547
rect 908 513 942 547
rect 976 513 992 547
rect 858 497 992 513
rect 1085 546 1107 580
rect 1141 546 1157 580
rect 1198 587 1300 649
rect 1198 553 1232 587
rect 1266 553 1300 587
rect 1463 581 1644 615
rect 1085 519 1157 546
rect 1463 519 1501 581
rect 1085 499 1501 519
rect 858 482 895 497
rect 365 389 824 423
rect 365 344 431 389
rect 365 310 381 344
rect 415 310 431 344
rect 365 294 431 310
rect 477 350 551 355
rect 477 339 511 350
rect 477 305 493 339
rect 545 316 551 350
rect 527 305 551 316
rect 477 289 551 305
rect 585 353 651 355
rect 585 319 601 353
rect 635 319 651 353
rect 585 311 651 319
rect 777 322 824 389
rect 297 255 431 260
rect 297 221 345 255
rect 379 237 431 255
rect 585 237 619 311
rect 777 305 827 322
rect 379 221 619 237
rect 297 215 619 221
rect 329 203 619 215
rect 669 243 689 277
rect 723 243 743 277
rect 777 271 793 305
rect 777 255 827 271
rect 669 221 743 243
rect 861 221 895 482
rect 1085 465 1107 499
rect 1141 485 1501 499
rect 1542 531 1576 547
rect 1141 465 1157 485
rect 1085 448 1157 465
rect 929 432 1157 448
rect 1341 434 1407 451
rect 1542 435 1576 497
rect 929 398 945 432
rect 979 398 1013 432
rect 1047 418 1157 432
rect 1047 398 1107 418
rect 929 384 1107 398
rect 1141 384 1157 418
rect 929 382 1157 384
rect 1019 368 1157 382
rect 1219 426 1501 434
rect 1219 392 1357 426
rect 1391 418 1501 426
rect 1391 392 1451 418
rect 1219 384 1451 392
rect 1485 384 1501 418
rect 1219 368 1501 384
rect 65 94 81 128
rect 115 94 171 128
rect 65 78 171 94
rect 229 146 295 181
rect 229 112 245 146
rect 279 112 295 146
rect 229 17 295 112
rect 329 165 395 203
rect 329 131 345 165
rect 379 131 395 165
rect 329 70 395 131
rect 441 140 507 156
rect 441 106 457 140
rect 491 106 507 140
rect 441 17 507 106
rect 541 85 575 203
rect 669 187 895 221
rect 929 291 979 320
rect 963 257 979 291
rect 929 153 979 257
rect 1019 234 1085 368
rect 1219 334 1253 368
rect 1119 318 1307 334
rect 1119 284 1135 318
rect 1169 284 1203 318
rect 1237 284 1307 318
rect 1119 268 1307 284
rect 1019 200 1035 234
rect 1069 200 1085 234
rect 1273 193 1307 268
rect 1341 318 1409 334
rect 1341 284 1343 318
rect 1377 284 1409 318
rect 1542 305 1576 401
rect 1341 236 1409 284
rect 1443 271 1576 305
rect 1610 321 1644 581
rect 1853 508 1925 649
rect 1678 448 1728 477
rect 1853 474 1872 508
rect 1906 474 1925 508
rect 2073 560 2139 649
rect 2073 526 2089 560
rect 2123 526 2139 560
rect 2073 492 2139 526
rect 1853 458 1925 474
rect 1712 419 1728 448
rect 1966 450 2032 477
rect 2073 458 2089 492
rect 2123 458 2139 492
rect 2179 564 2213 580
rect 2179 484 2213 530
rect 1966 424 1982 450
rect 1712 414 1779 419
rect 1678 385 1779 414
rect 1610 305 1711 321
rect 1610 271 1674 305
rect 1708 271 1711 305
rect 1273 177 1392 193
rect 609 119 625 153
rect 659 119 979 153
rect 1013 132 1239 166
rect 1013 85 1047 132
rect 541 51 1047 85
rect 1121 82 1171 98
rect 1121 48 1137 82
rect 1205 85 1239 132
rect 1273 143 1342 177
rect 1376 143 1392 177
rect 1273 127 1392 143
rect 1443 85 1477 271
rect 1610 255 1711 271
rect 1745 253 1779 385
rect 1813 416 1982 424
rect 2016 424 2032 450
rect 2016 416 2135 424
rect 1813 390 2135 416
rect 1813 341 1866 390
rect 1813 307 1816 341
rect 1850 307 1866 341
rect 1813 291 1866 307
rect 1908 350 1991 356
rect 1908 340 1951 350
rect 1908 306 1924 340
rect 1985 316 1991 350
rect 1958 306 1991 316
rect 1908 290 1991 306
rect 1745 237 2067 253
rect 1511 208 1545 237
rect 1745 221 2032 237
rect 1581 187 1601 221
rect 1635 203 2032 221
rect 2066 203 2067 237
rect 1635 187 2067 203
rect 1511 153 1545 174
rect 2101 153 2135 390
rect 2179 404 2213 450
rect 2179 308 2213 370
rect 2253 564 2319 649
rect 2253 530 2269 564
rect 2303 530 2319 564
rect 2495 580 2561 649
rect 2253 472 2319 530
rect 2253 438 2269 472
rect 2303 438 2319 472
rect 2253 398 2319 438
rect 2253 364 2269 398
rect 2303 364 2319 398
rect 2253 348 2319 364
rect 2379 540 2461 556
rect 2379 506 2395 540
rect 2429 506 2461 540
rect 2379 469 2461 506
rect 2379 435 2395 469
rect 2429 435 2461 469
rect 2379 398 2461 435
rect 2379 364 2395 398
rect 2429 364 2461 398
rect 2495 546 2511 580
rect 2545 546 2561 580
rect 2495 497 2561 546
rect 2495 463 2511 497
rect 2545 463 2561 497
rect 2495 414 2561 463
rect 2495 380 2511 414
rect 2545 380 2561 414
rect 2495 364 2561 380
rect 2595 580 2661 596
rect 2595 546 2611 580
rect 2645 546 2661 580
rect 2595 497 2661 546
rect 2595 463 2611 497
rect 2645 463 2661 497
rect 2595 414 2661 463
rect 2595 380 2611 414
rect 2645 380 2661 414
rect 2595 364 2661 380
rect 2695 580 2761 649
rect 2695 546 2711 580
rect 2745 546 2761 580
rect 2695 497 2761 546
rect 2695 463 2711 497
rect 2745 463 2761 497
rect 2695 414 2761 463
rect 2695 380 2711 414
rect 2745 380 2761 414
rect 2695 364 2761 380
rect 2379 348 2461 364
rect 2427 326 2461 348
rect 2427 310 2593 326
rect 2179 282 2345 308
rect 2179 264 2375 282
rect 1511 128 1847 153
rect 1511 119 1813 128
rect 1797 94 1813 119
rect 1205 51 1706 85
rect 1740 51 1756 85
rect 1797 70 1847 94
rect 1883 128 1949 144
rect 1883 94 1899 128
rect 1933 94 1949 128
rect 1121 17 1171 48
rect 1883 17 1949 94
rect 2041 128 2135 153
rect 2041 94 2057 128
rect 2091 94 2135 128
rect 2041 70 2135 94
rect 2169 204 2203 220
rect 2169 120 2203 170
rect 2169 17 2203 86
rect 2239 204 2375 264
rect 2239 170 2255 204
rect 2289 170 2375 204
rect 2239 154 2375 170
rect 2427 276 2543 310
rect 2577 276 2593 310
rect 2427 260 2593 276
rect 2427 190 2486 260
rect 2627 226 2661 364
rect 2427 156 2436 190
rect 2470 156 2486 190
rect 2239 120 2291 154
rect 2427 120 2486 156
rect 2239 86 2255 120
rect 2289 86 2291 120
rect 2239 70 2291 86
rect 2325 86 2342 120
rect 2376 86 2393 120
rect 2325 17 2393 86
rect 2427 86 2436 120
rect 2470 86 2486 120
rect 2427 70 2486 86
rect 2526 210 2576 226
rect 2526 176 2542 210
rect 2526 120 2576 176
rect 2526 86 2542 120
rect 2526 17 2576 86
rect 2612 207 2678 226
rect 2612 173 2628 207
rect 2662 173 2678 207
rect 2612 116 2678 173
rect 2612 82 2628 116
rect 2662 82 2678 116
rect 2612 66 2678 82
rect 2712 210 2764 226
rect 2712 176 2714 210
rect 2748 176 2764 210
rect 2712 120 2764 176
rect 2712 86 2714 120
rect 2748 86 2764 120
rect 2712 17 2764 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 223 340 257 350
rect 223 316 240 340
rect 240 316 257 340
rect 511 339 545 350
rect 511 316 527 339
rect 527 316 545 339
rect 1951 340 1985 350
rect 1951 316 1958 340
rect 1958 316 1985 340
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 211 350 269 356
rect 211 316 223 350
rect 257 347 269 350
rect 499 350 557 356
rect 499 347 511 350
rect 257 319 511 347
rect 257 316 269 319
rect 211 310 269 316
rect 499 316 511 319
rect 545 347 557 350
rect 1939 350 1997 356
rect 1939 347 1951 350
rect 545 319 1951 347
rect 545 316 557 319
rect 499 310 557 316
rect 1939 316 1951 319
rect 1985 316 1997 350
rect 1939 310 1997 316
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel comment s 936 68 936 68 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 361 36 361 36 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfrbp_2
flabel metal1 s 511 316 545 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 2623 168 2657 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2335 168 2369 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2335 242 2369 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y R90
string GDS_END 2581840
string GDS_START 2562092
<< end >>
