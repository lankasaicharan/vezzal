magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3698 1975
<< nwell >>
rect -38 343 2438 704
rect -38 331 249 343
rect 1049 340 2438 343
rect 1440 331 2438 340
rect 1440 292 2003 331
<< pwell >>
rect 291 282 1041 301
rect 291 238 1398 282
rect 2119 244 2393 263
rect 1735 238 2393 244
rect 291 189 2393 238
rect 1 49 2393 189
rect 0 0 2400 49
<< scnmos >>
rect 397 191 427 275
rect 469 191 499 275
rect 607 191 637 275
rect 754 191 784 275
rect 831 191 861 275
rect 916 191 946 275
rect 80 79 110 163
rect 166 79 196 163
rect 1133 128 1163 256
rect 1242 128 1272 256
rect 1394 128 1424 212
rect 1466 128 1496 212
rect 1552 128 1582 212
rect 1624 128 1654 212
rect 1814 50 1844 218
rect 1900 50 1930 218
rect 2093 69 2123 153
rect 2198 69 2228 237
rect 2284 69 2314 237
<< scpmoshvt >>
rect 85 472 115 600
rect 171 472 201 600
rect 361 463 391 547
rect 475 463 505 547
rect 677 463 707 547
rect 763 463 793 547
rect 835 463 865 547
rect 945 463 975 547
rect 1135 379 1165 547
rect 1267 412 1297 580
rect 1372 496 1402 580
rect 1444 496 1474 580
rect 1607 496 1637 580
rect 1693 496 1723 580
rect 1798 328 1828 580
rect 1884 328 1914 580
rect 2081 367 2111 495
rect 2198 367 2228 619
rect 2284 367 2314 619
<< ndiff >>
rect 317 191 397 275
rect 427 191 469 275
rect 499 248 607 275
rect 499 214 562 248
rect 596 214 607 248
rect 499 191 607 214
rect 637 244 754 275
rect 637 210 709 244
rect 743 210 754 244
rect 637 191 754 210
rect 784 191 831 275
rect 861 191 916 275
rect 946 256 1015 275
rect 946 191 1133 256
rect 27 135 80 163
rect 27 101 35 135
rect 69 101 80 135
rect 27 79 80 101
rect 110 135 166 163
rect 110 101 121 135
rect 155 101 166 135
rect 110 79 166 101
rect 196 135 249 163
rect 196 101 207 135
rect 241 101 249 135
rect 196 79 249 101
rect 317 135 375 191
rect 317 101 331 135
rect 365 101 375 135
rect 317 86 375 101
rect 961 172 1133 191
rect 1053 128 1133 172
rect 1163 248 1242 256
rect 1163 214 1174 248
rect 1208 214 1242 248
rect 1163 128 1242 214
rect 1272 212 1372 256
rect 1272 198 1394 212
rect 1272 164 1330 198
rect 1364 164 1394 198
rect 1272 128 1394 164
rect 1424 128 1466 212
rect 1496 187 1552 212
rect 1496 153 1507 187
rect 1541 153 1552 187
rect 1496 128 1552 153
rect 1582 128 1624 212
rect 1654 198 1707 212
rect 1654 164 1665 198
rect 1699 164 1707 198
rect 1654 128 1707 164
rect 1053 108 1111 128
rect 1053 74 1065 108
rect 1099 74 1111 108
rect 1053 66 1111 74
rect 1761 121 1814 218
rect 1761 87 1769 121
rect 1803 87 1814 121
rect 1761 50 1814 87
rect 1844 210 1900 218
rect 1844 176 1855 210
rect 1889 176 1900 210
rect 1844 101 1900 176
rect 1844 67 1855 101
rect 1889 67 1900 101
rect 1844 50 1900 67
rect 1930 206 1983 218
rect 1930 172 1941 206
rect 1975 172 1983 206
rect 2145 221 2198 237
rect 1930 96 1983 172
rect 2145 187 2153 221
rect 2187 187 2198 221
rect 2145 153 2198 187
rect 1930 62 1941 96
rect 1975 62 1983 96
rect 2040 127 2093 153
rect 2040 93 2048 127
rect 2082 93 2093 127
rect 2040 69 2093 93
rect 2123 115 2198 153
rect 2123 81 2134 115
rect 2168 81 2198 115
rect 2123 69 2198 81
rect 2228 225 2284 237
rect 2228 191 2239 225
rect 2273 191 2284 225
rect 2228 117 2284 191
rect 2228 83 2239 117
rect 2273 83 2284 117
rect 2228 69 2284 83
rect 2314 225 2367 237
rect 2314 191 2325 225
rect 2359 191 2367 225
rect 2314 115 2367 191
rect 2314 81 2325 115
rect 2359 81 2367 115
rect 2314 69 2367 81
rect 1930 50 1983 62
<< pdiff >>
rect 32 588 85 600
rect 32 554 40 588
rect 74 554 85 588
rect 32 520 85 554
rect 32 486 40 520
rect 74 486 85 520
rect 32 472 85 486
rect 115 588 171 600
rect 115 554 126 588
rect 160 554 171 588
rect 115 520 171 554
rect 115 486 126 520
rect 160 486 171 520
rect 115 472 171 486
rect 201 588 254 600
rect 201 554 212 588
rect 246 554 254 588
rect 201 520 254 554
rect 406 567 460 583
rect 406 547 416 567
rect 201 486 212 520
rect 246 486 254 520
rect 201 472 254 486
rect 308 515 361 547
rect 308 481 316 515
rect 350 481 361 515
rect 308 463 361 481
rect 391 533 416 547
rect 450 547 460 567
rect 450 533 475 547
rect 391 463 475 533
rect 505 521 562 547
rect 505 487 516 521
rect 550 487 562 521
rect 505 463 562 487
rect 880 567 930 583
rect 2145 607 2198 619
rect 880 547 888 567
rect 622 521 677 547
rect 622 487 632 521
rect 666 487 677 521
rect 622 463 677 487
rect 707 524 763 547
rect 707 490 718 524
rect 752 490 763 524
rect 707 463 763 490
rect 793 463 835 547
rect 865 533 888 547
rect 922 547 930 567
rect 1180 566 1267 580
rect 1180 547 1195 566
rect 922 533 945 547
rect 865 463 945 533
rect 975 523 1028 547
rect 975 489 986 523
rect 1020 489 1028 523
rect 975 463 1028 489
rect 1082 493 1135 547
rect 1082 459 1090 493
rect 1124 459 1135 493
rect 1082 379 1135 459
rect 1165 532 1195 547
rect 1229 532 1267 566
rect 1165 498 1267 532
rect 1165 464 1195 498
rect 1229 464 1267 498
rect 1165 430 1267 464
rect 1165 396 1195 430
rect 1229 412 1267 430
rect 1297 566 1372 580
rect 1297 532 1308 566
rect 1342 532 1372 566
rect 1297 496 1372 532
rect 1402 496 1444 580
rect 1474 555 1607 580
rect 1474 521 1485 555
rect 1519 521 1562 555
rect 1596 521 1607 555
rect 1474 496 1607 521
rect 1637 555 1693 580
rect 1637 521 1648 555
rect 1682 521 1693 555
rect 1637 496 1693 521
rect 1723 568 1798 580
rect 1723 534 1753 568
rect 1787 534 1798 568
rect 1723 500 1798 534
rect 1723 496 1753 500
rect 1297 458 1350 496
rect 1297 424 1308 458
rect 1342 424 1350 458
rect 1297 412 1350 424
rect 1229 396 1245 412
rect 1165 379 1245 396
rect 1745 466 1753 496
rect 1787 466 1798 500
rect 1745 422 1798 466
rect 1745 388 1753 422
rect 1787 388 1798 422
rect 1745 328 1798 388
rect 1828 568 1884 580
rect 1828 534 1839 568
rect 1873 534 1884 568
rect 1828 467 1884 534
rect 1828 433 1839 467
rect 1873 433 1884 467
rect 1828 374 1884 433
rect 1828 340 1839 374
rect 1873 340 1884 374
rect 1828 328 1884 340
rect 1914 568 1967 580
rect 1914 534 1925 568
rect 1959 534 1967 568
rect 1914 467 1967 534
rect 2145 573 2153 607
rect 2187 573 2198 607
rect 2145 511 2198 573
rect 2145 495 2153 511
rect 1914 433 1925 467
rect 1959 433 1967 467
rect 1914 374 1967 433
rect 1914 340 1925 374
rect 1959 340 1967 374
rect 2028 481 2081 495
rect 2028 447 2036 481
rect 2070 447 2081 481
rect 2028 413 2081 447
rect 2028 379 2036 413
rect 2070 379 2081 413
rect 2028 367 2081 379
rect 2111 477 2153 495
rect 2187 477 2198 511
rect 2111 413 2198 477
rect 2111 379 2122 413
rect 2156 379 2198 413
rect 2111 367 2198 379
rect 2228 599 2284 619
rect 2228 565 2239 599
rect 2273 565 2284 599
rect 2228 508 2284 565
rect 2228 474 2239 508
rect 2273 474 2284 508
rect 2228 413 2284 474
rect 2228 379 2239 413
rect 2273 379 2284 413
rect 2228 367 2284 379
rect 2314 607 2367 619
rect 2314 573 2325 607
rect 2359 573 2367 607
rect 2314 511 2367 573
rect 2314 477 2325 511
rect 2359 477 2367 511
rect 2314 413 2367 477
rect 2314 379 2325 413
rect 2359 379 2367 413
rect 2314 367 2367 379
rect 1914 328 1967 340
<< ndiffc >>
rect 562 214 596 248
rect 709 210 743 244
rect 35 101 69 135
rect 121 101 155 135
rect 207 101 241 135
rect 331 101 365 135
rect 1174 214 1208 248
rect 1330 164 1364 198
rect 1507 153 1541 187
rect 1665 164 1699 198
rect 1065 74 1099 108
rect 1769 87 1803 121
rect 1855 176 1889 210
rect 1855 67 1889 101
rect 1941 172 1975 206
rect 2153 187 2187 221
rect 1941 62 1975 96
rect 2048 93 2082 127
rect 2134 81 2168 115
rect 2239 191 2273 225
rect 2239 83 2273 117
rect 2325 191 2359 225
rect 2325 81 2359 115
<< pdiffc >>
rect 40 554 74 588
rect 40 486 74 520
rect 126 554 160 588
rect 126 486 160 520
rect 212 554 246 588
rect 212 486 246 520
rect 316 481 350 515
rect 416 533 450 567
rect 516 487 550 521
rect 632 487 666 521
rect 718 490 752 524
rect 888 533 922 567
rect 986 489 1020 523
rect 1090 459 1124 493
rect 1195 532 1229 566
rect 1195 464 1229 498
rect 1195 396 1229 430
rect 1308 532 1342 566
rect 1485 521 1519 555
rect 1562 521 1596 555
rect 1648 521 1682 555
rect 1753 534 1787 568
rect 1308 424 1342 458
rect 1753 466 1787 500
rect 1753 388 1787 422
rect 1839 534 1873 568
rect 1839 433 1873 467
rect 1839 340 1873 374
rect 1925 534 1959 568
rect 2153 573 2187 607
rect 1925 433 1959 467
rect 1925 340 1959 374
rect 2036 447 2070 481
rect 2036 379 2070 413
rect 2153 477 2187 511
rect 2122 379 2156 413
rect 2239 565 2273 599
rect 2239 474 2273 508
rect 2239 379 2273 413
rect 2325 573 2359 607
rect 2325 477 2359 511
rect 2325 379 2359 413
<< poly >>
rect 85 600 115 626
rect 171 615 1297 645
rect 2198 619 2228 645
rect 2284 619 2314 645
rect 171 600 201 615
rect 361 547 391 573
rect 85 394 115 472
rect 171 457 201 472
rect 475 547 505 573
rect 171 436 232 457
rect 178 432 232 436
rect 182 430 232 432
rect 361 431 391 463
rect 475 431 505 463
rect 186 427 232 430
rect 190 424 232 427
rect 85 378 160 394
rect 85 344 110 378
rect 144 344 160 378
rect 85 328 160 344
rect 85 307 115 328
rect 80 270 115 307
rect 80 163 110 270
rect 202 251 232 424
rect 326 415 392 431
rect 326 381 342 415
rect 376 381 392 415
rect 326 347 392 381
rect 326 313 342 347
rect 376 327 392 347
rect 469 415 535 431
rect 469 381 485 415
rect 519 381 535 415
rect 469 347 535 381
rect 577 387 607 615
rect 677 547 707 573
rect 763 547 793 615
rect 835 547 865 573
rect 1267 580 1297 615
rect 1372 580 1402 606
rect 1444 580 1474 606
rect 1607 580 1637 606
rect 1693 580 1723 606
rect 1798 580 1828 606
rect 1884 580 1914 606
rect 945 547 975 573
rect 1135 547 1165 573
rect 677 389 707 463
rect 763 437 793 463
rect 835 397 865 463
rect 945 424 975 463
rect 925 408 998 424
rect 577 357 633 387
rect 376 313 427 327
rect 326 297 427 313
rect 397 275 427 297
rect 469 313 485 347
rect 519 313 535 347
rect 469 297 535 313
rect 603 310 633 357
rect 675 373 745 389
rect 675 339 691 373
rect 725 339 745 373
rect 811 381 877 397
rect 811 347 827 381
rect 861 347 877 381
rect 811 341 877 347
rect 675 323 745 339
rect 812 337 877 341
rect 814 335 877 337
rect 816 331 877 335
rect 925 374 948 408
rect 982 374 998 408
rect 1267 386 1297 412
rect 925 358 998 374
rect 715 319 772 323
rect 715 315 774 319
rect 715 311 776 315
rect 603 308 634 310
rect 715 309 778 311
rect 603 306 635 308
rect 715 306 780 309
rect 603 304 636 306
rect 469 275 499 297
rect 603 290 637 304
rect 715 303 782 306
rect 715 290 784 303
rect 607 275 637 290
rect 754 275 784 290
rect 831 275 861 331
rect 925 312 955 358
rect 1135 344 1165 379
rect 1372 344 1402 496
rect 916 290 955 312
rect 1072 328 1165 344
rect 1072 294 1088 328
rect 1122 294 1165 328
rect 916 275 946 290
rect 1072 278 1165 294
rect 1242 328 1402 344
rect 1242 294 1260 328
rect 1294 314 1402 328
rect 1444 454 1474 496
rect 1607 456 1637 496
rect 1444 438 1510 454
rect 1444 404 1460 438
rect 1494 404 1510 438
rect 1444 370 1510 404
rect 1444 336 1460 370
rect 1494 336 1510 370
rect 1444 320 1510 336
rect 1552 440 1637 456
rect 1552 406 1568 440
rect 1602 406 1637 440
rect 1552 390 1637 406
rect 1294 294 1310 314
rect 1242 278 1310 294
rect 157 235 232 251
rect 157 201 173 235
rect 207 201 232 235
rect 157 185 232 201
rect 1133 256 1163 278
rect 1242 256 1272 278
rect 166 163 196 185
rect 397 123 427 191
rect 469 165 499 191
rect 607 165 637 191
rect 754 165 784 191
rect 831 165 861 191
rect 916 123 946 191
rect 397 93 946 123
rect 1394 212 1424 238
rect 1466 212 1496 320
rect 1552 212 1582 390
rect 1693 300 1723 496
rect 2081 495 2111 521
rect 1798 300 1828 328
rect 1884 300 1914 328
rect 2081 300 2111 367
rect 2198 325 2228 367
rect 2284 325 2314 367
rect 1647 284 2111 300
rect 1647 264 1663 284
rect 1624 250 1663 264
rect 1697 270 2111 284
rect 2153 309 2314 325
rect 2153 275 2169 309
rect 2203 295 2314 309
rect 2203 275 2228 295
rect 1697 250 1723 270
rect 1624 234 1723 250
rect 1624 212 1654 234
rect 1814 218 1844 270
rect 1900 218 1930 270
rect 80 53 110 79
rect 166 51 196 79
rect 1133 102 1163 128
rect 1242 102 1272 128
rect 1394 51 1424 128
rect 1466 102 1496 128
rect 1552 102 1582 128
rect 1624 102 1654 128
rect 166 21 1424 51
rect 2075 211 2105 270
rect 2153 259 2228 275
rect 2198 237 2228 259
rect 2284 237 2314 295
rect 2075 181 2123 211
rect 2093 153 2123 181
rect 1814 24 1844 50
rect 1900 24 1930 50
rect 2093 43 2123 69
rect 2198 43 2228 69
rect 2284 43 2314 69
<< polycont >>
rect 110 344 144 378
rect 342 381 376 415
rect 342 313 376 347
rect 485 381 519 415
rect 485 313 519 347
rect 691 339 725 373
rect 827 347 861 381
rect 948 374 982 408
rect 1088 294 1122 328
rect 1260 294 1294 328
rect 1460 404 1494 438
rect 1460 336 1494 370
rect 1568 406 1602 440
rect 173 201 207 235
rect 1663 250 1697 284
rect 2169 275 2203 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 24 588 76 604
rect 24 554 40 588
rect 74 554 76 588
rect 24 520 76 554
rect 24 486 40 520
rect 74 486 76 520
rect 24 467 76 486
rect 110 588 176 649
rect 110 554 126 588
rect 160 554 176 588
rect 110 520 176 554
rect 110 486 126 520
rect 160 486 176 520
rect 110 467 176 486
rect 210 588 276 604
rect 210 554 212 588
rect 246 554 276 588
rect 210 520 276 554
rect 398 567 468 649
rect 210 486 212 520
rect 246 486 276 520
rect 210 467 276 486
rect 24 251 71 467
rect 222 461 276 467
rect 310 515 350 547
rect 398 533 416 567
rect 450 533 468 567
rect 872 567 938 649
rect 310 481 316 515
rect 512 521 673 547
rect 512 499 516 521
rect 350 487 516 499
rect 550 487 632 521
rect 666 487 673 521
rect 350 481 673 487
rect 310 465 673 481
rect 707 524 797 547
rect 872 533 888 567
rect 922 533 938 567
rect 872 530 938 533
rect 707 490 718 524
rect 752 494 797 524
rect 974 523 1023 547
rect 974 494 986 523
rect 752 490 986 494
rect 707 489 986 490
rect 1020 489 1023 523
rect 707 474 1023 489
rect 105 378 181 433
rect 242 431 276 461
rect 562 460 673 465
rect 759 460 1023 474
rect 1074 493 1140 649
rect 242 387 283 431
rect 105 344 110 378
rect 144 344 181 378
rect 105 299 181 344
rect 24 235 211 251
rect 24 201 173 235
rect 207 201 211 235
rect 24 185 211 201
rect 247 208 283 387
rect 317 424 378 431
rect 317 390 319 424
rect 353 415 378 424
rect 317 381 342 390
rect 376 381 378 415
rect 317 347 378 381
rect 317 313 342 347
rect 376 313 378 347
rect 317 290 378 313
rect 412 415 528 431
rect 412 381 485 415
rect 519 381 528 415
rect 412 347 528 381
rect 412 313 485 347
rect 519 313 528 347
rect 412 242 528 313
rect 562 423 634 460
rect 562 248 607 423
rect 596 214 607 248
rect 24 135 80 185
rect 247 174 463 208
rect 562 196 607 214
rect 641 373 725 389
rect 641 339 691 373
rect 641 323 725 339
rect 247 151 281 174
rect 24 101 35 135
rect 69 101 80 135
rect 24 85 80 101
rect 114 135 166 151
rect 114 101 121 135
rect 155 101 166 135
rect 114 17 166 101
rect 200 135 281 151
rect 415 160 463 174
rect 641 160 675 323
rect 759 260 793 460
rect 1074 459 1090 493
rect 1124 459 1140 493
rect 1074 448 1140 459
rect 1190 566 1233 582
rect 1190 532 1195 566
rect 1229 532 1233 566
rect 1190 498 1233 532
rect 1190 464 1195 498
rect 1229 464 1233 498
rect 1190 430 1233 464
rect 827 381 861 406
rect 929 408 984 424
rect 1190 414 1195 430
rect 929 390 948 408
rect 899 374 948 390
rect 982 374 984 408
rect 899 358 984 374
rect 1018 396 1195 414
rect 1229 396 1233 430
rect 1304 566 1368 583
rect 1304 532 1308 566
rect 1342 532 1368 566
rect 1304 458 1368 532
rect 1469 555 1605 649
rect 1469 521 1485 555
rect 1519 521 1562 555
rect 1596 521 1605 555
rect 1469 505 1605 521
rect 1644 555 1698 571
rect 1644 521 1648 555
rect 1682 521 1698 555
rect 1304 424 1308 458
rect 1342 424 1368 458
rect 1304 408 1368 424
rect 1018 380 1233 396
rect 827 322 861 347
rect 1018 322 1052 380
rect 827 288 1052 322
rect 1086 328 1124 344
rect 1086 294 1088 328
rect 1122 294 1124 328
rect 709 252 793 260
rect 1086 252 1124 294
rect 1190 264 1224 380
rect 709 244 1124 252
rect 743 212 1124 244
rect 1158 248 1224 264
rect 1158 214 1174 248
rect 1208 214 1224 248
rect 1158 212 1224 214
rect 1258 328 1294 344
rect 1258 294 1260 328
rect 743 210 847 212
rect 709 194 847 210
rect 1258 178 1294 294
rect 912 160 1294 178
rect 415 144 1294 160
rect 1328 286 1368 408
rect 1444 438 1510 454
rect 1444 404 1460 438
rect 1494 404 1510 438
rect 1444 370 1510 404
rect 1552 440 1610 456
rect 1552 424 1568 440
rect 1552 390 1567 424
rect 1602 406 1610 440
rect 1601 390 1610 406
rect 1444 336 1460 370
rect 1494 356 1510 370
rect 1644 356 1698 521
rect 1737 568 1803 649
rect 1737 534 1753 568
rect 1787 534 1803 568
rect 1737 500 1803 534
rect 1737 466 1753 500
rect 1787 466 1803 500
rect 1737 422 1803 466
rect 1737 388 1753 422
rect 1787 388 1803 422
rect 1839 568 1891 584
rect 1873 534 1891 568
rect 1839 467 1891 534
rect 1873 433 1891 467
rect 1494 354 1698 356
rect 1839 374 1891 433
rect 1494 336 1805 354
rect 1444 320 1805 336
rect 1328 284 1713 286
rect 1328 250 1663 284
rect 1697 250 1713 284
rect 1328 248 1713 250
rect 1328 198 1368 248
rect 1749 214 1805 320
rect 1328 164 1330 198
rect 1364 164 1368 198
rect 200 101 207 135
rect 241 101 281 135
rect 200 79 281 101
rect 315 135 381 140
rect 315 101 331 135
rect 365 101 381 135
rect 415 126 955 144
rect 1328 126 1368 164
rect 1491 187 1557 203
rect 1491 153 1507 187
rect 1541 153 1557 187
rect 1649 198 1805 214
rect 1649 164 1665 198
rect 1699 164 1805 198
rect 1873 340 1891 374
rect 1839 210 1891 340
rect 1925 568 1975 649
rect 1959 534 1975 568
rect 1925 467 1975 534
rect 2120 607 2191 649
rect 2120 573 2153 607
rect 2187 573 2191 607
rect 2120 511 2191 573
rect 1959 433 1975 467
rect 1925 374 1975 433
rect 1959 340 1975 374
rect 1925 324 1975 340
rect 2025 481 2086 497
rect 2025 447 2036 481
rect 2070 447 2086 481
rect 2025 413 2086 447
rect 2025 379 2036 413
rect 2070 379 2086 413
rect 2025 325 2086 379
rect 2120 477 2153 511
rect 2187 477 2191 511
rect 2120 413 2191 477
rect 2120 379 2122 413
rect 2156 379 2191 413
rect 2120 363 2191 379
rect 2237 599 2282 615
rect 2237 565 2239 599
rect 2273 565 2282 599
rect 2237 508 2282 565
rect 2237 474 2239 508
rect 2273 474 2282 508
rect 2237 413 2282 474
rect 2237 379 2239 413
rect 2273 379 2282 413
rect 2025 309 2203 325
rect 2025 275 2169 309
rect 2025 259 2203 275
rect 1839 176 1855 210
rect 1889 176 1891 210
rect 1839 164 1891 176
rect 315 17 381 101
rect 1049 108 1115 110
rect 1049 74 1065 108
rect 1099 74 1115 108
rect 1049 17 1115 74
rect 1491 17 1557 153
rect 1753 121 1819 130
rect 1753 87 1769 121
rect 1803 87 1819 121
rect 1753 17 1819 87
rect 1853 101 1891 164
rect 1853 67 1855 101
rect 1889 67 1891 101
rect 1853 51 1891 67
rect 1925 206 1991 222
rect 1925 172 1941 206
rect 1975 172 1991 206
rect 1925 96 1991 172
rect 1925 62 1941 96
rect 1975 62 1991 96
rect 2025 127 2098 259
rect 2237 225 2282 379
rect 2316 607 2375 649
rect 2316 573 2325 607
rect 2359 573 2375 607
rect 2316 511 2375 573
rect 2316 477 2325 511
rect 2359 477 2375 511
rect 2316 413 2375 477
rect 2316 379 2325 413
rect 2359 379 2375 413
rect 2316 363 2375 379
rect 2025 93 2048 127
rect 2082 93 2098 127
rect 2025 77 2098 93
rect 2132 221 2203 225
rect 2132 187 2153 221
rect 2187 187 2203 221
rect 2132 115 2203 187
rect 2132 81 2134 115
rect 2168 81 2203 115
rect 1925 17 1991 62
rect 2132 17 2203 81
rect 2237 191 2239 225
rect 2273 191 2282 225
rect 2237 117 2282 191
rect 2237 83 2239 117
rect 2273 83 2282 117
rect 2237 67 2282 83
rect 2316 225 2375 241
rect 2316 191 2325 225
rect 2359 191 2375 225
rect 2316 115 2375 191
rect 2316 81 2325 115
rect 2359 81 2375 115
rect 2316 17 2375 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 319 415 353 424
rect 319 390 342 415
rect 342 390 353 415
rect 895 390 929 424
rect 1567 406 1568 424
rect 1568 406 1601 424
rect 1567 390 1601 406
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 307 424 365 430
rect 307 390 319 424
rect 353 421 365 424
rect 883 424 941 430
rect 883 421 895 424
rect 353 393 895 421
rect 353 390 365 393
rect 307 384 365 390
rect 883 390 895 393
rect 929 421 941 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 929 393 1567 421
rect 929 390 941 393
rect 883 384 941 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< labels >>
flabel pwell s 0 0 2400 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2400 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel comment s 680 36 680 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 680 108 680 108 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 680 630 680 630 0 FreeSans 300 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfrbp_2
flabel metal1 s 1567 390 1601 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 2400 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2400 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2239 94 2273 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 168 2273 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 242 2273 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 316 2273 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 390 2273 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 464 2273 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 538 2273 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1855 94 1889 128 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1855 168 1889 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1855 390 1889 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1855 464 1889 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1855 538 1889 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2400 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry R90
string GDS_END 4525022
string GDS_START 4505562
<< end >>
