magic
tech sky130A
magscale 1 2
timestamp 1627202622
<< checkpaint >>
rect -1326 -1303 4878 2157
<< nwell >>
rect -66 477 3618 897
rect -66 377 1198 477
rect 2300 377 3618 477
<< pwell >>
rect 1908 329 2018 369
rect 1463 263 1721 283
rect 1908 263 2240 329
rect 4 219 418 222
rect 4 217 1138 219
rect 1463 217 2240 263
rect 2656 217 3548 283
rect 4 43 3548 217
rect -26 -43 3578 43
<< mvnmos >>
rect 83 112 183 196
rect 239 112 339 196
rect 505 109 605 193
rect 661 109 761 193
rect 817 109 917 193
rect 959 109 1059 193
rect 1225 107 1325 191
rect 1367 107 1467 191
rect 1542 107 1642 257
rect 1812 153 1912 237
rect 2014 153 2114 303
rect 2327 107 2427 191
rect 2469 107 2569 191
rect 2739 173 2839 257
rect 2914 107 3014 257
rect 3190 173 3290 257
rect 3365 107 3465 257
<< mvpmos >>
rect 87 532 187 682
rect 243 532 343 682
rect 564 543 664 627
rect 720 543 820 627
rect 876 543 976 627
rect 1018 543 1118 627
rect 1244 543 1344 627
rect 1400 543 1500 627
rect 1632 543 1732 743
rect 1774 543 1874 743
rect 1953 543 2053 627
rect 2156 543 2256 627
rect 2312 543 2412 627
rect 2733 443 2833 527
rect 2912 443 3012 743
rect 3186 479 3286 629
rect 3365 479 3465 679
<< mvndiff >>
rect 30 171 83 196
rect 30 137 38 171
rect 72 137 83 171
rect 30 112 83 137
rect 183 171 239 196
rect 183 137 194 171
rect 228 137 239 171
rect 183 112 239 137
rect 339 171 392 196
rect 339 137 350 171
rect 384 137 392 171
rect 339 112 392 137
rect 452 168 505 193
rect 452 134 460 168
rect 494 134 505 168
rect 452 109 505 134
rect 605 171 661 193
rect 605 137 616 171
rect 650 137 661 171
rect 605 109 661 137
rect 761 171 817 193
rect 761 137 772 171
rect 806 137 817 171
rect 761 109 817 137
rect 917 109 959 193
rect 1059 168 1112 193
rect 1489 191 1542 257
rect 1059 134 1070 168
rect 1104 134 1112 168
rect 1059 109 1112 134
rect 1172 166 1225 191
rect 1172 132 1180 166
rect 1214 132 1225 166
rect 1172 107 1225 132
rect 1325 107 1367 191
rect 1467 174 1542 191
rect 1467 140 1497 174
rect 1531 140 1542 174
rect 1467 107 1542 140
rect 1642 174 1695 257
rect 1934 335 1992 343
rect 1934 301 1946 335
rect 1980 303 1992 335
rect 1980 301 2014 303
rect 1934 237 2014 301
rect 1642 140 1653 174
rect 1687 140 1695 174
rect 1755 195 1812 237
rect 1755 161 1767 195
rect 1801 161 1812 195
rect 1755 153 1812 161
rect 1912 153 2014 237
rect 2114 199 2214 303
rect 2114 165 2172 199
rect 2206 165 2214 199
rect 2682 232 2739 257
rect 2682 198 2694 232
rect 2728 198 2739 232
rect 2114 153 2214 165
rect 2274 166 2327 191
rect 1642 107 1695 140
rect 2274 132 2282 166
rect 2316 132 2327 166
rect 2274 107 2327 132
rect 2427 107 2469 191
rect 2569 166 2622 191
rect 2682 173 2739 198
rect 2839 179 2914 257
rect 2839 173 2869 179
rect 2569 132 2580 166
rect 2614 132 2622 166
rect 2569 107 2622 132
rect 2861 145 2869 173
rect 2903 145 2914 179
rect 2861 107 2914 145
rect 3014 249 3071 257
rect 3014 215 3025 249
rect 3059 215 3071 249
rect 3014 149 3071 215
rect 3133 232 3190 257
rect 3133 198 3145 232
rect 3179 198 3190 232
rect 3133 173 3190 198
rect 3290 245 3365 257
rect 3290 211 3320 245
rect 3354 211 3365 245
rect 3290 173 3365 211
rect 3014 115 3025 149
rect 3059 115 3071 149
rect 3312 153 3365 173
rect 3014 107 3071 115
rect 3312 119 3320 153
rect 3354 119 3365 153
rect 3312 107 3365 119
rect 3465 249 3522 257
rect 3465 215 3476 249
rect 3510 215 3522 249
rect 3465 149 3522 215
rect 3465 115 3476 149
rect 3510 115 3522 149
rect 3465 107 3522 115
<< mvpdiff >>
rect 30 674 87 682
rect 30 640 42 674
rect 76 640 87 674
rect 30 574 87 640
rect 30 540 42 574
rect 76 540 87 574
rect 30 532 87 540
rect 187 674 243 682
rect 187 640 198 674
rect 232 640 243 674
rect 187 574 243 640
rect 187 540 198 574
rect 232 540 243 574
rect 187 532 243 540
rect 343 674 400 682
rect 343 640 354 674
rect 388 640 400 674
rect 343 574 400 640
rect 1582 627 1632 743
rect 343 540 354 574
rect 388 540 400 574
rect 489 602 564 627
rect 489 568 501 602
rect 535 568 564 602
rect 489 543 564 568
rect 664 602 720 627
rect 664 568 675 602
rect 709 568 720 602
rect 664 543 720 568
rect 820 602 876 627
rect 820 568 831 602
rect 865 568 876 602
rect 820 543 876 568
rect 976 543 1018 627
rect 1118 617 1244 627
rect 1118 583 1152 617
rect 1186 583 1244 617
rect 1118 543 1244 583
rect 1344 602 1400 627
rect 1344 568 1355 602
rect 1389 568 1400 602
rect 1344 543 1400 568
rect 1500 616 1632 627
rect 1500 582 1587 616
rect 1621 582 1632 616
rect 1500 543 1632 582
rect 1732 543 1774 743
rect 1874 735 1931 743
rect 1874 701 1885 735
rect 1919 701 1931 735
rect 1874 660 1931 701
rect 1874 626 1885 660
rect 1919 627 1931 660
rect 2855 735 2912 743
rect 2855 701 2867 735
rect 2901 701 2912 735
rect 2855 652 2912 701
rect 1919 626 1953 627
rect 1874 585 1953 626
rect 1874 551 1885 585
rect 1919 551 1953 585
rect 1874 543 1953 551
rect 2053 543 2156 627
rect 2256 602 2312 627
rect 2256 568 2267 602
rect 2301 568 2312 602
rect 2256 543 2312 568
rect 2412 602 2469 627
rect 2412 568 2423 602
rect 2457 568 2469 602
rect 2412 543 2469 568
rect 2855 618 2867 652
rect 2901 618 2912 652
rect 2855 568 2912 618
rect 343 532 400 540
rect 2855 534 2867 568
rect 2901 534 2912 568
rect 2855 527 2912 534
rect 2676 502 2733 527
rect 2676 468 2688 502
rect 2722 468 2733 502
rect 2676 443 2733 468
rect 2833 485 2912 527
rect 2833 451 2867 485
rect 2901 451 2912 485
rect 2833 443 2912 451
rect 3012 735 3069 743
rect 3012 701 3023 735
rect 3057 701 3069 735
rect 3012 652 3069 701
rect 3308 671 3365 679
rect 3012 618 3023 652
rect 3057 618 3069 652
rect 3308 637 3320 671
rect 3354 637 3365 671
rect 3308 629 3365 637
rect 3012 568 3069 618
rect 3012 534 3023 568
rect 3057 534 3069 568
rect 3012 485 3069 534
rect 3012 451 3023 485
rect 3057 451 3069 485
rect 3129 621 3186 629
rect 3129 587 3141 621
rect 3175 587 3186 621
rect 3129 521 3186 587
rect 3129 487 3141 521
rect 3175 487 3186 521
rect 3129 479 3186 487
rect 3286 596 3365 629
rect 3286 562 3320 596
rect 3354 562 3365 596
rect 3286 521 3365 562
rect 3286 487 3320 521
rect 3354 487 3365 521
rect 3286 479 3365 487
rect 3465 671 3522 679
rect 3465 637 3476 671
rect 3510 637 3522 671
rect 3465 596 3522 637
rect 3465 562 3476 596
rect 3510 562 3522 596
rect 3465 521 3522 562
rect 3465 487 3476 521
rect 3510 487 3522 521
rect 3465 479 3522 487
rect 3012 443 3069 451
<< mvndiffc >>
rect 38 137 72 171
rect 194 137 228 171
rect 350 137 384 171
rect 460 134 494 168
rect 616 137 650 171
rect 772 137 806 171
rect 1070 134 1104 168
rect 1180 132 1214 166
rect 1497 140 1531 174
rect 1946 301 1980 335
rect 1653 140 1687 174
rect 1767 161 1801 195
rect 2172 165 2206 199
rect 2694 198 2728 232
rect 2282 132 2316 166
rect 2580 132 2614 166
rect 2869 145 2903 179
rect 3025 215 3059 249
rect 3145 198 3179 232
rect 3320 211 3354 245
rect 3025 115 3059 149
rect 3320 119 3354 153
rect 3476 215 3510 249
rect 3476 115 3510 149
<< mvpdiffc >>
rect 42 640 76 674
rect 42 540 76 574
rect 198 640 232 674
rect 198 540 232 574
rect 354 640 388 674
rect 354 540 388 574
rect 501 568 535 602
rect 675 568 709 602
rect 831 568 865 602
rect 1152 583 1186 617
rect 1355 568 1389 602
rect 1587 582 1621 616
rect 1885 701 1919 735
rect 1885 626 1919 660
rect 2867 701 2901 735
rect 1885 551 1919 585
rect 2267 568 2301 602
rect 2423 568 2457 602
rect 2867 618 2901 652
rect 2867 534 2901 568
rect 2688 468 2722 502
rect 2867 451 2901 485
rect 3023 701 3057 735
rect 3023 618 3057 652
rect 3320 637 3354 671
rect 3023 534 3057 568
rect 3023 451 3057 485
rect 3141 587 3175 621
rect 3141 487 3175 521
rect 3320 562 3354 596
rect 3320 487 3354 521
rect 3476 637 3510 671
rect 3476 562 3510 596
rect 3476 487 3510 521
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3552 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
<< poly >>
rect 1632 743 1732 769
rect 1774 743 1874 769
rect 2912 743 3012 769
rect 87 682 187 708
rect 243 682 343 708
rect 564 627 664 653
rect 720 627 820 653
rect 876 627 976 653
rect 1018 627 1118 653
rect 1244 627 1344 653
rect 1400 627 1500 653
rect 1953 627 2053 653
rect 2156 627 2256 653
rect 2312 627 2412 653
rect 87 464 187 532
rect 83 444 187 464
rect 83 410 128 444
rect 162 410 187 444
rect 83 376 187 410
rect 243 378 343 532
rect 564 517 664 543
rect 83 342 128 376
rect 162 342 187 376
rect 83 322 187 342
rect 239 358 343 378
rect 239 324 268 358
rect 302 324 343 358
rect 83 196 183 322
rect 239 290 343 324
rect 239 256 268 290
rect 302 256 343 290
rect 239 222 343 256
rect 505 417 664 517
rect 720 439 820 543
rect 876 495 976 543
rect 876 481 922 495
rect 902 461 922 481
rect 956 461 976 495
rect 902 441 976 461
rect 1018 517 1118 543
rect 1018 475 1136 517
rect 1018 441 1082 475
rect 1116 441 1136 475
rect 1244 451 1344 543
rect 1400 521 1500 543
rect 505 383 525 417
rect 559 383 605 417
rect 720 399 860 439
rect 1018 417 1136 441
rect 505 349 605 383
rect 505 315 525 349
rect 559 315 605 349
rect 239 196 339 222
rect 505 193 605 315
rect 661 339 765 357
rect 661 305 711 339
rect 745 305 765 339
rect 661 271 765 305
rect 807 333 917 399
rect 807 299 867 333
rect 901 299 917 333
rect 1018 315 1118 417
rect 807 293 917 299
rect 661 237 711 271
rect 745 237 765 271
rect 661 217 765 237
rect 817 265 917 293
rect 817 231 867 265
rect 901 231 917 265
rect 661 193 761 217
rect 817 193 917 231
rect 959 265 1118 315
rect 959 231 1005 265
rect 1039 231 1118 265
rect 959 215 1118 231
rect 1225 405 1344 451
rect 1225 371 1245 405
rect 1279 371 1344 405
rect 1225 351 1344 371
rect 959 193 1059 215
rect 83 86 183 112
rect 239 86 339 112
rect 1225 191 1325 351
rect 1386 309 1500 521
rect 1632 517 1732 543
rect 1542 473 1732 517
rect 1542 439 1562 473
rect 1596 439 1732 473
rect 1542 405 1732 439
rect 1542 371 1562 405
rect 1596 371 1732 405
rect 1542 351 1732 371
rect 1774 495 1874 543
rect 1774 461 1790 495
rect 1824 461 1874 495
rect 1774 427 1874 461
rect 1774 393 1790 427
rect 1824 393 1874 427
rect 1953 517 2053 543
rect 2156 517 2256 543
rect 2312 517 2412 543
rect 2733 527 2833 553
rect 1953 495 2114 517
rect 1953 461 1987 495
rect 2021 461 2114 495
rect 1953 417 2114 461
rect 2156 417 2270 517
rect 2312 421 2569 517
rect 3365 679 3465 705
rect 3186 629 3286 655
rect 3186 453 3286 479
rect 2312 417 2489 421
rect 1774 363 1874 393
rect 1367 265 1474 309
rect 1367 231 1413 265
rect 1447 231 1474 265
rect 1542 257 1642 351
rect 1774 263 1912 363
rect 1367 213 1474 231
rect 1367 191 1467 213
rect 505 83 605 109
rect 661 83 761 109
rect 817 83 917 109
rect 959 83 1059 109
rect 1812 237 1912 263
rect 2014 303 2114 417
rect 2229 366 2270 417
rect 2469 387 2489 417
rect 2523 387 2569 421
rect 2229 346 2427 366
rect 2229 312 2344 346
rect 2378 312 2427 346
rect 2229 278 2427 312
rect 2229 244 2344 278
rect 2378 244 2427 278
rect 2229 217 2427 244
rect 2327 191 2427 217
rect 2469 353 2569 387
rect 2469 319 2489 353
rect 2523 319 2569 353
rect 2469 191 2569 319
rect 2733 383 2833 443
rect 2912 383 3012 443
rect 3186 383 3290 453
rect 2733 345 3290 383
rect 2733 311 2759 345
rect 2793 311 3290 345
rect 2733 283 3290 311
rect 2739 257 2839 283
rect 2914 257 3014 283
rect 3190 257 3290 283
rect 3365 419 3465 479
rect 3365 385 3385 419
rect 3419 385 3465 419
rect 3365 351 3465 385
rect 3365 317 3385 351
rect 3419 317 3465 351
rect 3365 257 3465 317
rect 1812 127 1912 153
rect 2014 127 2114 153
rect 2739 147 2839 173
rect 3190 147 3290 173
rect 1225 81 1325 107
rect 1367 81 1467 107
rect 1542 81 1642 107
rect 2327 81 2427 107
rect 2469 81 2569 107
rect 2914 81 3014 107
rect 3365 81 3465 107
<< polycont >>
rect 128 410 162 444
rect 128 342 162 376
rect 268 324 302 358
rect 268 256 302 290
rect 922 461 956 495
rect 1082 441 1116 475
rect 525 383 559 417
rect 525 315 559 349
rect 711 305 745 339
rect 867 299 901 333
rect 711 237 745 271
rect 867 231 901 265
rect 1005 231 1039 265
rect 1245 371 1279 405
rect 1562 439 1596 473
rect 1562 371 1596 405
rect 1790 461 1824 495
rect 1790 393 1824 427
rect 1987 461 2021 495
rect 1413 231 1447 265
rect 2489 387 2523 421
rect 2344 312 2378 346
rect 2344 244 2378 278
rect 2489 319 2523 353
rect 2759 311 2793 345
rect 3385 385 3419 419
rect 3385 317 3419 351
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3552 831
rect 130 735 248 741
rect 130 701 136 735
rect 170 701 208 735
rect 242 701 248 735
rect 22 674 76 690
rect 22 640 42 674
rect 22 574 76 640
rect 22 540 42 574
rect 130 674 248 701
rect 130 640 198 674
rect 232 640 248 674
rect 130 574 248 640
rect 130 540 198 574
rect 232 540 248 574
rect 284 726 458 760
rect 22 274 76 540
rect 112 444 178 504
rect 112 410 128 444
rect 162 410 178 444
rect 112 376 178 410
rect 112 342 128 376
rect 162 342 178 376
rect 284 374 318 726
rect 112 310 178 342
rect 252 358 318 374
rect 252 324 268 358
rect 302 324 318 358
rect 252 290 318 324
rect 252 274 268 290
rect 22 256 268 274
rect 302 256 318 290
rect 22 240 318 256
rect 354 674 388 690
rect 354 574 388 640
rect 354 267 388 540
rect 424 499 458 726
rect 494 735 535 741
rect 494 701 498 735
rect 532 701 535 735
rect 1136 735 1249 741
rect 494 602 535 701
rect 494 568 501 602
rect 494 535 535 568
rect 571 671 1100 705
rect 571 499 605 671
rect 424 465 605 499
rect 641 602 709 635
rect 641 568 675 602
rect 641 535 709 568
rect 505 417 575 429
rect 505 383 525 417
rect 559 383 575 417
rect 505 349 575 383
rect 505 315 525 349
rect 559 315 575 349
rect 505 303 575 315
rect 22 171 72 240
rect 354 233 564 267
rect 22 137 38 171
rect 22 108 72 137
rect 108 171 298 204
rect 354 200 400 233
rect 108 137 194 171
rect 228 137 298 171
rect 108 113 298 137
rect 108 79 114 113
rect 148 79 186 113
rect 220 79 258 113
rect 292 79 298 113
rect 334 171 400 200
rect 334 137 350 171
rect 384 137 400 171
rect 334 108 400 137
rect 444 168 494 197
rect 444 134 460 168
rect 444 113 494 134
rect 108 73 298 79
rect 444 79 450 113
rect 484 79 494 113
rect 444 73 494 79
rect 530 87 564 233
rect 641 201 675 535
rect 745 479 779 671
rect 815 602 1030 635
rect 815 568 831 602
rect 865 601 1030 602
rect 865 568 881 601
rect 815 535 881 568
rect 917 495 960 511
rect 917 479 922 495
rect 711 461 922 479
rect 956 461 960 495
rect 711 445 960 461
rect 711 339 745 445
rect 996 405 1030 601
rect 1066 545 1100 671
rect 1136 701 1139 735
rect 1173 701 1211 735
rect 1245 701 1249 735
rect 1571 735 1761 741
rect 1136 617 1249 701
rect 1136 583 1152 617
rect 1186 583 1249 617
rect 1136 581 1249 583
rect 1285 671 1535 705
rect 1285 545 1319 671
rect 1066 511 1319 545
rect 1355 602 1405 635
rect 1389 568 1405 602
rect 1355 475 1405 568
rect 1501 543 1535 671
rect 1571 701 1577 735
rect 1611 701 1649 735
rect 1683 701 1721 735
rect 1755 701 1761 735
rect 1571 616 1761 701
rect 1571 582 1587 616
rect 1621 582 1761 616
rect 1571 579 1761 582
rect 1869 735 2107 751
rect 1869 701 1885 735
rect 1919 717 2107 735
rect 1919 701 1935 717
rect 1869 660 1935 701
rect 1869 626 1885 660
rect 1919 626 1935 660
rect 1869 585 1935 626
rect 1869 551 1885 585
rect 1919 551 1935 585
rect 1501 509 1824 543
rect 1869 535 1935 551
rect 1066 441 1082 475
rect 1116 441 1405 475
rect 1774 495 1824 509
rect 1971 495 2037 511
rect 1546 439 1562 473
rect 1596 439 1612 473
rect 1546 405 1612 439
rect 711 271 745 305
rect 711 221 745 237
rect 781 371 1245 405
rect 1279 371 1562 405
rect 1596 371 1612 405
rect 1774 461 1790 495
rect 1774 427 1824 461
rect 1774 393 1790 427
rect 1774 377 1824 393
rect 1860 461 1987 495
rect 2021 461 2037 495
rect 2073 499 2107 717
rect 2143 735 2333 741
rect 2143 701 2149 735
rect 2183 701 2221 735
rect 2255 701 2293 735
rect 2327 701 2333 735
rect 2143 602 2333 701
rect 2774 735 2964 751
rect 2774 701 2780 735
rect 2814 701 2852 735
rect 2901 701 2924 735
rect 2958 701 2964 735
rect 2774 652 2964 701
rect 2143 568 2267 602
rect 2301 568 2333 602
rect 2143 535 2333 568
rect 2407 602 2636 635
rect 2407 568 2423 602
rect 2457 568 2636 602
rect 2407 499 2636 568
rect 2774 618 2867 652
rect 2901 618 2964 652
rect 2774 568 2964 618
rect 2073 465 2636 499
rect 600 171 675 201
rect 781 185 815 371
rect 1860 335 1894 461
rect 2073 425 2107 465
rect 851 333 1894 335
rect 851 299 867 333
rect 901 301 1894 333
rect 1930 391 2107 425
rect 2143 421 2566 429
rect 2143 395 2489 421
rect 1930 335 1996 391
rect 2143 355 2177 395
rect 2430 387 2489 395
rect 2523 387 2566 421
rect 1930 301 1946 335
rect 1980 301 1996 335
rect 2032 321 2177 355
rect 2328 346 2394 359
rect 901 299 917 301
rect 851 265 917 299
rect 2032 265 2066 321
rect 2328 312 2344 346
rect 2378 312 2394 346
rect 851 231 867 265
rect 901 231 917 265
rect 851 221 917 231
rect 989 231 1005 265
rect 1039 231 1230 265
rect 1397 231 1413 265
rect 1447 231 2066 265
rect 2102 251 2292 285
rect 600 137 616 171
rect 650 137 675 171
rect 600 123 675 137
rect 756 171 822 185
rect 756 137 772 171
rect 806 137 822 171
rect 756 123 822 137
rect 858 87 892 221
rect 989 217 1230 231
rect 530 53 892 87
rect 930 168 1120 181
rect 930 134 1070 168
rect 1104 134 1120 168
rect 930 113 1120 134
rect 930 79 936 113
rect 970 79 1008 113
rect 1042 79 1080 113
rect 1114 79 1120 113
rect 1164 166 1230 217
rect 2102 195 2136 251
rect 1164 132 1180 166
rect 1214 132 1230 166
rect 1164 103 1230 132
rect 1357 174 1547 195
rect 1357 140 1497 174
rect 1531 140 1547 174
rect 1357 113 1547 140
rect 930 73 1120 79
rect 1357 79 1363 113
rect 1397 79 1435 113
rect 1469 79 1507 113
rect 1541 79 1547 113
rect 1357 73 1547 79
rect 1637 174 1703 195
rect 1637 140 1653 174
rect 1687 140 1703 174
rect 1751 161 1767 195
rect 1801 161 2136 195
rect 1751 145 2136 161
rect 2172 199 2222 215
rect 2206 165 2222 199
rect 1637 109 1703 140
rect 2172 109 2222 165
rect 1637 75 2222 109
rect 2258 195 2292 251
rect 2328 278 2394 312
rect 2430 353 2566 387
rect 2430 319 2489 353
rect 2523 319 2566 353
rect 2430 311 2566 319
rect 2602 345 2636 465
rect 2672 502 2738 535
rect 2672 468 2688 502
rect 2722 468 2738 502
rect 2672 415 2738 468
rect 2774 534 2867 568
rect 2901 534 2964 568
rect 2774 485 2964 534
rect 2774 451 2867 485
rect 2901 451 2964 485
rect 3003 735 3075 751
rect 3003 701 3023 735
rect 3057 701 3075 735
rect 3003 652 3075 701
rect 3003 618 3023 652
rect 3057 618 3075 652
rect 3227 735 3417 741
rect 3227 701 3233 735
rect 3267 701 3305 735
rect 3339 701 3377 735
rect 3411 701 3417 735
rect 3227 671 3417 701
rect 3227 637 3320 671
rect 3354 637 3417 671
rect 3003 568 3075 618
rect 3003 534 3023 568
rect 3057 534 3075 568
rect 3003 485 3075 534
rect 3003 451 3023 485
rect 3057 451 3075 485
rect 2672 381 2879 415
rect 2602 311 2759 345
rect 2793 311 2809 345
rect 2328 244 2344 278
rect 2378 275 2394 278
rect 2845 275 2879 381
rect 2378 244 2879 275
rect 2328 241 2879 244
rect 3003 249 3075 451
rect 2328 231 2394 241
rect 2678 232 2744 241
rect 2678 198 2694 232
rect 2728 198 2744 232
rect 3003 215 3025 249
rect 3059 215 3075 249
rect 2258 166 2332 195
rect 2258 132 2282 166
rect 2316 132 2332 166
rect 2258 103 2332 132
rect 2440 166 2630 195
rect 2440 132 2580 166
rect 2614 132 2630 166
rect 2678 165 2744 198
rect 2780 179 2967 205
rect 2440 113 2630 132
rect 2440 79 2446 113
rect 2480 79 2518 113
rect 2552 79 2590 113
rect 2624 79 2630 113
rect 2440 73 2630 79
rect 2780 145 2869 179
rect 2903 145 2967 179
rect 2780 113 2967 145
rect 2780 79 2784 113
rect 2818 79 2856 113
rect 2890 79 2928 113
rect 2962 79 2967 113
rect 3003 149 3075 215
rect 3125 621 3191 637
rect 3125 587 3141 621
rect 3175 587 3191 621
rect 3125 521 3191 587
rect 3125 487 3141 521
rect 3175 487 3191 521
rect 3125 335 3191 487
rect 3227 596 3417 637
rect 3227 562 3320 596
rect 3354 562 3417 596
rect 3227 521 3417 562
rect 3227 487 3320 521
rect 3354 487 3417 521
rect 3227 471 3417 487
rect 3460 671 3527 687
rect 3460 637 3476 671
rect 3510 637 3527 671
rect 3460 596 3527 637
rect 3460 562 3476 596
rect 3510 562 3527 596
rect 3460 521 3527 562
rect 3460 487 3476 521
rect 3510 487 3527 521
rect 3460 471 3527 487
rect 3369 419 3435 435
rect 3369 385 3385 419
rect 3419 385 3435 419
rect 3369 351 3435 385
rect 3369 335 3385 351
rect 3125 317 3385 335
rect 3419 317 3435 351
rect 3125 301 3435 317
rect 3125 232 3195 301
rect 3481 265 3527 471
rect 3125 198 3145 232
rect 3179 198 3195 232
rect 3125 165 3195 198
rect 3231 245 3421 261
rect 3231 211 3320 245
rect 3354 211 3421 245
rect 3003 115 3025 149
rect 3059 115 3075 149
rect 3003 99 3075 115
rect 3231 153 3421 211
rect 3231 119 3320 153
rect 3354 119 3421 153
rect 3231 113 3421 119
rect 2780 73 2967 79
rect 3231 79 3237 113
rect 3271 79 3309 113
rect 3343 79 3381 113
rect 3415 79 3421 113
rect 3460 249 3527 265
rect 3460 215 3476 249
rect 3510 215 3527 249
rect 3460 149 3527 215
rect 3460 115 3476 149
rect 3510 115 3527 149
rect 3460 99 3527 115
rect 3231 73 3421 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 136 701 170 735
rect 208 701 242 735
rect 498 701 532 735
rect 114 79 148 113
rect 186 79 220 113
rect 258 79 292 113
rect 450 79 484 113
rect 1139 701 1173 735
rect 1211 701 1245 735
rect 1577 701 1611 735
rect 1649 701 1683 735
rect 1721 701 1755 735
rect 2149 701 2183 735
rect 2221 701 2255 735
rect 2293 701 2327 735
rect 2780 701 2814 735
rect 2852 701 2867 735
rect 2867 701 2886 735
rect 2924 701 2958 735
rect 936 79 970 113
rect 1008 79 1042 113
rect 1080 79 1114 113
rect 1363 79 1397 113
rect 1435 79 1469 113
rect 1507 79 1541 113
rect 3233 701 3267 735
rect 3305 701 3339 735
rect 3377 701 3411 735
rect 2446 79 2480 113
rect 2518 79 2552 113
rect 2590 79 2624 113
rect 2784 79 2818 113
rect 2856 79 2890 113
rect 2928 79 2962 113
rect 3237 79 3271 113
rect 3309 79 3343 113
rect 3381 79 3415 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
<< metal1 >>
rect 0 831 3552 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3552 831
rect 0 791 3552 797
rect 0 735 3552 763
rect 0 701 136 735
rect 170 701 208 735
rect 242 701 498 735
rect 532 701 1139 735
rect 1173 701 1211 735
rect 1245 701 1577 735
rect 1611 701 1649 735
rect 1683 701 1721 735
rect 1755 701 2149 735
rect 2183 701 2221 735
rect 2255 701 2293 735
rect 2327 701 2780 735
rect 2814 701 2852 735
rect 2886 701 2924 735
rect 2958 701 3233 735
rect 3267 701 3305 735
rect 3339 701 3377 735
rect 3411 701 3552 735
rect 0 689 3552 701
rect 0 113 3552 125
rect 0 79 114 113
rect 148 79 186 113
rect 220 79 258 113
rect 292 79 450 113
rect 484 79 936 113
rect 970 79 1008 113
rect 1042 79 1080 113
rect 1114 79 1363 113
rect 1397 79 1435 113
rect 1469 79 1507 113
rect 1541 79 2446 113
rect 2480 79 2518 113
rect 2552 79 2590 113
rect 2624 79 2784 113
rect 2818 79 2856 113
rect 2890 79 2928 113
rect 2962 79 3237 113
rect 3271 79 3309 113
rect 3343 79 3381 113
rect 3415 79 3552 113
rect 0 51 3552 79
rect 0 17 3552 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
rect 0 -23 3552 -17
<< labels >>
flabel comment s 1065 353 1065 353 0 FreeSans 200 90 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 dfsbp_1
flabel metal1 s 0 51 3552 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 0 3552 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 689 3552 763 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 791 3552 814 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2431 316 2465 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 2527 316 2561 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 3487 168 3521 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3487 242 3521 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3487 316 3521 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3487 390 3521 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3487 464 3521 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3487 538 3521 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3487 612 3521 646 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 3007 168 3041 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3007 242 3041 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3007 316 3041 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3007 390 3041 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3007 464 3041 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3007 538 3041 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 3007 612 3041 646 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 3552 814
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string LEFsymmetry X Y
string GDS_END 629860
string GDS_START 596428
<< end >>
