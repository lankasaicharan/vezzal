magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2954 1852
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 1 21 1607 157
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 131
rect 173 47 203 131
rect 277 47 307 131
rect 361 47 391 131
rect 465 47 495 131
rect 549 47 579 131
rect 653 47 683 131
rect 737 47 767 131
rect 841 47 871 131
rect 925 47 955 131
rect 1029 47 1059 131
rect 1113 47 1143 131
rect 1217 47 1247 131
rect 1301 47 1331 131
rect 1405 47 1435 131
rect 1489 47 1519 131
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
rect 1209 297 1245 497
rect 1303 297 1339 497
rect 1397 297 1433 497
rect 1491 297 1527 497
<< ndiff >>
rect 27 106 89 131
rect 27 72 35 106
rect 69 72 89 106
rect 27 47 89 72
rect 119 106 173 131
rect 119 72 129 106
rect 163 72 173 106
rect 119 47 173 72
rect 203 106 277 131
rect 203 72 223 106
rect 257 72 277 106
rect 203 47 277 72
rect 307 106 361 131
rect 307 72 317 106
rect 351 72 361 106
rect 307 47 361 72
rect 391 106 465 131
rect 391 72 411 106
rect 445 72 465 106
rect 391 47 465 72
rect 495 106 549 131
rect 495 72 505 106
rect 539 72 549 106
rect 495 47 549 72
rect 579 106 653 131
rect 579 72 599 106
rect 633 72 653 106
rect 579 47 653 72
rect 683 106 737 131
rect 683 72 693 106
rect 727 72 737 106
rect 683 47 737 72
rect 767 106 841 131
rect 767 72 787 106
rect 821 72 841 106
rect 767 47 841 72
rect 871 106 925 131
rect 871 72 881 106
rect 915 72 925 106
rect 871 47 925 72
rect 955 106 1029 131
rect 955 72 975 106
rect 1009 72 1029 106
rect 955 47 1029 72
rect 1059 106 1113 131
rect 1059 72 1069 106
rect 1103 72 1113 106
rect 1059 47 1113 72
rect 1143 106 1217 131
rect 1143 72 1163 106
rect 1197 72 1217 106
rect 1143 47 1217 72
rect 1247 106 1301 131
rect 1247 72 1257 106
rect 1291 72 1301 106
rect 1247 47 1301 72
rect 1331 106 1405 131
rect 1331 72 1351 106
rect 1385 72 1405 106
rect 1331 47 1405 72
rect 1435 106 1489 131
rect 1435 72 1445 106
rect 1479 72 1489 106
rect 1435 47 1489 72
rect 1519 106 1581 131
rect 1519 72 1539 106
rect 1573 72 1581 106
rect 1519 47 1581 72
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 477 175 497
rect 117 443 129 477
rect 163 443 175 477
rect 117 409 175 443
rect 117 375 129 409
rect 163 375 175 409
rect 117 341 175 375
rect 117 307 129 341
rect 163 307 175 341
rect 117 297 175 307
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 477 363 497
rect 305 443 317 477
rect 351 443 363 477
rect 305 409 363 443
rect 305 375 317 409
rect 351 375 363 409
rect 305 341 363 375
rect 305 307 317 341
rect 351 307 363 341
rect 305 297 363 307
rect 399 481 457 497
rect 399 447 411 481
rect 445 447 457 481
rect 399 413 457 447
rect 399 379 411 413
rect 445 379 457 413
rect 399 345 457 379
rect 399 311 411 345
rect 445 311 457 345
rect 399 297 457 311
rect 493 477 551 497
rect 493 443 505 477
rect 539 443 551 477
rect 493 409 551 443
rect 493 375 505 409
rect 539 375 551 409
rect 493 341 551 375
rect 493 307 505 341
rect 539 307 551 341
rect 493 297 551 307
rect 587 477 645 497
rect 587 443 599 477
rect 633 443 645 477
rect 587 409 645 443
rect 587 375 599 409
rect 633 375 645 409
rect 587 297 645 375
rect 681 477 739 497
rect 681 443 693 477
rect 727 443 739 477
rect 681 409 739 443
rect 681 375 693 409
rect 727 375 739 409
rect 681 341 739 375
rect 681 307 693 341
rect 727 307 739 341
rect 681 297 739 307
rect 775 477 833 497
rect 775 443 787 477
rect 821 443 833 477
rect 775 409 833 443
rect 775 375 787 409
rect 821 375 833 409
rect 775 297 833 375
rect 869 477 927 497
rect 869 443 881 477
rect 915 443 927 477
rect 869 409 927 443
rect 869 375 881 409
rect 915 375 927 409
rect 869 341 927 375
rect 869 307 881 341
rect 915 307 927 341
rect 869 297 927 307
rect 963 477 1021 497
rect 963 443 975 477
rect 1009 443 1021 477
rect 963 409 1021 443
rect 963 375 975 409
rect 1009 375 1021 409
rect 963 297 1021 375
rect 1057 477 1115 497
rect 1057 443 1069 477
rect 1103 443 1115 477
rect 1057 409 1115 443
rect 1057 375 1069 409
rect 1103 375 1115 409
rect 1057 341 1115 375
rect 1057 307 1069 341
rect 1103 307 1115 341
rect 1057 297 1115 307
rect 1151 477 1209 497
rect 1151 443 1163 477
rect 1197 443 1209 477
rect 1151 409 1209 443
rect 1151 375 1163 409
rect 1197 375 1209 409
rect 1151 297 1209 375
rect 1245 477 1303 497
rect 1245 443 1257 477
rect 1291 443 1303 477
rect 1245 409 1303 443
rect 1245 375 1257 409
rect 1291 375 1303 409
rect 1245 341 1303 375
rect 1245 307 1257 341
rect 1291 307 1303 341
rect 1245 297 1303 307
rect 1339 477 1397 497
rect 1339 443 1351 477
rect 1385 443 1397 477
rect 1339 409 1397 443
rect 1339 375 1351 409
rect 1385 375 1397 409
rect 1339 297 1397 375
rect 1433 477 1491 497
rect 1433 443 1445 477
rect 1479 443 1491 477
rect 1433 409 1491 443
rect 1433 375 1445 409
rect 1479 375 1491 409
rect 1433 341 1491 375
rect 1433 307 1445 341
rect 1479 307 1491 341
rect 1433 297 1491 307
rect 1527 479 1581 497
rect 1527 445 1539 479
rect 1573 445 1581 479
rect 1527 411 1581 445
rect 1527 377 1539 411
rect 1573 377 1581 411
rect 1527 343 1581 377
rect 1527 309 1539 343
rect 1573 309 1581 343
rect 1527 297 1581 309
<< ndiffc >>
rect 35 72 69 106
rect 129 72 163 106
rect 223 72 257 106
rect 317 72 351 106
rect 411 72 445 106
rect 505 72 539 106
rect 599 72 633 106
rect 693 72 727 106
rect 787 72 821 106
rect 881 72 915 106
rect 975 72 1009 106
rect 1069 72 1103 106
rect 1163 72 1197 106
rect 1257 72 1291 106
rect 1351 72 1385 106
rect 1445 72 1479 106
rect 1539 72 1573 106
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 443 163 477
rect 129 375 163 409
rect 129 307 163 341
rect 223 451 257 485
rect 223 383 257 417
rect 317 443 351 477
rect 317 375 351 409
rect 317 307 351 341
rect 411 447 445 481
rect 411 379 445 413
rect 411 311 445 345
rect 505 443 539 477
rect 505 375 539 409
rect 505 307 539 341
rect 599 443 633 477
rect 599 375 633 409
rect 693 443 727 477
rect 693 375 727 409
rect 693 307 727 341
rect 787 443 821 477
rect 787 375 821 409
rect 881 443 915 477
rect 881 375 915 409
rect 881 307 915 341
rect 975 443 1009 477
rect 975 375 1009 409
rect 1069 443 1103 477
rect 1069 375 1103 409
rect 1069 307 1103 341
rect 1163 443 1197 477
rect 1163 375 1197 409
rect 1257 443 1291 477
rect 1257 375 1291 409
rect 1257 307 1291 341
rect 1351 443 1385 477
rect 1351 375 1385 409
rect 1445 443 1479 477
rect 1445 375 1479 409
rect 1445 307 1479 341
rect 1539 445 1573 479
rect 1539 377 1573 411
rect 1539 309 1573 343
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 1209 497 1245 523
rect 1303 497 1339 523
rect 1397 497 1433 523
rect 1491 497 1527 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 1209 282 1245 297
rect 1303 282 1339 297
rect 1397 282 1433 297
rect 1491 282 1527 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 79 249 401 265
rect 79 215 146 249
rect 180 215 214 249
rect 248 215 401 249
rect 79 180 401 215
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 831 265 871 282
rect 925 265 965 282
rect 1019 265 1059 282
rect 1113 265 1153 282
rect 1207 265 1247 282
rect 1301 265 1341 282
rect 1395 265 1435 282
rect 1489 265 1529 282
rect 455 249 1529 265
rect 455 215 471 249
rect 505 215 539 249
rect 573 215 607 249
rect 641 215 675 249
rect 709 215 743 249
rect 777 215 811 249
rect 845 215 879 249
rect 913 215 947 249
rect 981 215 1015 249
rect 1049 215 1083 249
rect 1117 215 1151 249
rect 1185 215 1219 249
rect 1253 215 1287 249
rect 1321 215 1529 249
rect 455 190 1529 215
rect 89 131 119 180
rect 173 131 203 180
rect 277 131 307 180
rect 361 131 391 180
rect 465 131 495 190
rect 549 131 579 190
rect 653 131 683 190
rect 737 131 767 190
rect 841 131 871 190
rect 925 131 955 190
rect 1029 131 1059 190
rect 1113 131 1143 190
rect 1217 131 1247 190
rect 1301 131 1331 190
rect 1405 131 1435 190
rect 1489 131 1519 190
rect 89 21 119 47
rect 173 21 203 47
rect 277 21 307 47
rect 361 21 391 47
rect 465 21 495 47
rect 549 21 579 47
rect 653 21 683 47
rect 737 21 767 47
rect 841 21 871 47
rect 925 21 955 47
rect 1029 21 1059 47
rect 1113 21 1143 47
rect 1217 21 1247 47
rect 1301 21 1331 47
rect 1405 21 1435 47
rect 1489 21 1519 47
<< polycont >>
rect 146 215 180 249
rect 214 215 248 249
rect 471 215 505 249
rect 539 215 573 249
rect 607 215 641 249
rect 675 215 709 249
rect 743 215 777 249
rect 811 215 845 249
rect 879 215 913 249
rect 947 215 981 249
rect 1015 215 1049 249
rect 1083 215 1117 249
rect 1151 215 1185 249
rect 1219 215 1253 249
rect 1287 215 1321 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 19 485 79 527
rect 19 451 35 485
rect 69 451 79 485
rect 19 417 79 451
rect 19 383 35 417
rect 69 383 79 417
rect 19 349 79 383
rect 19 315 35 349
rect 69 315 79 349
rect 19 299 79 315
rect 113 477 179 493
rect 113 443 129 477
rect 163 443 179 477
rect 113 409 179 443
rect 113 375 129 409
rect 163 375 179 409
rect 113 341 179 375
rect 213 485 267 527
rect 213 451 223 485
rect 257 451 267 485
rect 213 417 267 451
rect 213 383 223 417
rect 257 383 267 417
rect 213 367 267 383
rect 307 477 361 493
rect 307 443 317 477
rect 351 443 361 477
rect 307 409 361 443
rect 307 375 317 409
rect 351 375 361 409
rect 113 307 129 341
rect 163 333 179 341
rect 307 341 361 375
rect 307 333 317 341
rect 163 307 317 333
rect 351 307 361 341
rect 113 299 361 307
rect 114 295 361 299
rect 395 481 455 527
rect 395 447 411 481
rect 445 447 455 481
rect 395 413 455 447
rect 395 379 411 413
rect 445 379 455 413
rect 395 345 455 379
rect 395 311 411 345
rect 445 311 455 345
rect 395 295 455 311
rect 489 477 549 493
rect 489 443 505 477
rect 539 443 549 477
rect 489 409 549 443
rect 489 375 505 409
rect 539 375 549 409
rect 489 341 549 375
rect 583 477 649 527
rect 583 443 599 477
rect 633 443 649 477
rect 583 409 649 443
rect 583 375 599 409
rect 633 375 649 409
rect 583 367 649 375
rect 683 477 737 493
rect 683 443 693 477
rect 727 443 737 477
rect 683 409 737 443
rect 683 375 693 409
rect 727 375 737 409
rect 489 307 505 341
rect 539 333 549 341
rect 683 341 737 375
rect 771 477 837 527
rect 771 443 787 477
rect 821 443 837 477
rect 771 409 837 443
rect 771 375 787 409
rect 821 375 837 409
rect 771 367 837 375
rect 871 477 925 493
rect 871 443 881 477
rect 915 443 925 477
rect 871 409 925 443
rect 871 375 881 409
rect 915 375 925 409
rect 683 333 693 341
rect 539 307 693 333
rect 727 333 737 341
rect 871 341 925 375
rect 959 477 1025 527
rect 959 443 975 477
rect 1009 443 1025 477
rect 959 409 1025 443
rect 959 375 975 409
rect 1009 375 1025 409
rect 959 367 1025 375
rect 1059 477 1113 493
rect 1059 443 1069 477
rect 1103 443 1113 477
rect 1059 409 1113 443
rect 1059 375 1069 409
rect 1103 375 1113 409
rect 871 333 881 341
rect 727 307 881 333
rect 915 333 925 341
rect 1059 341 1113 375
rect 1147 477 1213 527
rect 1147 443 1163 477
rect 1197 443 1213 477
rect 1147 409 1213 443
rect 1147 375 1163 409
rect 1197 375 1213 409
rect 1147 367 1213 375
rect 1247 477 1301 493
rect 1247 443 1257 477
rect 1291 443 1301 477
rect 1247 409 1301 443
rect 1247 375 1257 409
rect 1291 375 1301 409
rect 1059 333 1069 341
rect 915 307 1069 333
rect 1103 333 1113 341
rect 1247 341 1301 375
rect 1335 477 1401 527
rect 1335 443 1351 477
rect 1385 443 1401 477
rect 1335 409 1401 443
rect 1335 375 1351 409
rect 1385 375 1401 409
rect 1335 367 1401 375
rect 1435 477 1489 493
rect 1435 443 1445 477
rect 1479 443 1489 477
rect 1435 409 1489 443
rect 1435 375 1445 409
rect 1479 375 1489 409
rect 1247 333 1257 341
rect 1103 307 1257 333
rect 1291 333 1301 341
rect 1435 341 1489 375
rect 1435 333 1445 341
rect 1291 307 1445 333
rect 1479 307 1489 341
rect 489 295 1489 307
rect 307 261 361 295
rect 105 249 264 261
rect 105 215 146 249
rect 180 215 214 249
rect 248 215 264 249
rect 307 249 1337 261
rect 307 215 471 249
rect 505 215 539 249
rect 573 215 607 249
rect 641 215 675 249
rect 709 215 743 249
rect 777 215 811 249
rect 845 215 879 249
rect 913 215 947 249
rect 981 215 1015 249
rect 1049 215 1083 249
rect 1117 215 1151 249
rect 1185 215 1219 249
rect 1253 215 1287 249
rect 1321 215 1337 249
rect 307 181 361 215
rect 1392 181 1489 295
rect 1523 479 1589 527
rect 1523 445 1539 479
rect 1573 445 1589 479
rect 1523 411 1589 445
rect 1523 377 1539 411
rect 1573 377 1589 411
rect 1523 343 1589 377
rect 1523 309 1539 343
rect 1573 309 1589 343
rect 1523 293 1589 309
rect 119 143 361 181
rect 19 106 85 122
rect 19 72 35 106
rect 69 72 85 106
rect 19 17 85 72
rect 119 106 173 143
rect 119 72 129 106
rect 163 72 173 106
rect 119 56 173 72
rect 207 106 273 109
rect 207 72 223 106
rect 257 72 273 106
rect 207 17 273 72
rect 307 106 361 143
rect 495 143 1489 181
rect 307 72 317 106
rect 351 72 361 106
rect 307 56 361 72
rect 395 106 461 109
rect 395 72 411 106
rect 445 72 461 106
rect 395 17 461 72
rect 495 106 549 143
rect 495 72 505 106
rect 539 72 549 106
rect 495 56 549 72
rect 583 106 649 109
rect 583 72 599 106
rect 633 72 649 106
rect 583 17 649 72
rect 683 106 737 143
rect 683 72 693 106
rect 727 72 737 106
rect 683 56 737 72
rect 771 106 837 109
rect 771 72 787 106
rect 821 72 837 106
rect 771 17 837 72
rect 871 106 925 143
rect 871 72 881 106
rect 915 72 925 106
rect 871 56 925 72
rect 959 106 1025 109
rect 959 72 975 106
rect 1009 72 1025 106
rect 959 17 1025 72
rect 1059 106 1113 143
rect 1059 72 1069 106
rect 1103 72 1113 106
rect 1059 56 1113 72
rect 1147 106 1213 109
rect 1147 72 1163 106
rect 1197 72 1213 106
rect 1147 17 1213 72
rect 1247 106 1301 143
rect 1247 72 1257 106
rect 1291 72 1301 106
rect 1247 56 1301 72
rect 1335 106 1401 109
rect 1335 72 1351 106
rect 1385 72 1401 106
rect 1335 17 1401 72
rect 1435 106 1489 143
rect 1435 72 1445 106
rect 1479 72 1489 106
rect 1435 56 1489 72
rect 1523 106 1589 122
rect 1523 72 1539 106
rect 1573 72 1589 106
rect 1523 17 1589 72
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1409 221 1443 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkbuf_12
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1656 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 902024
string GDS_START 890252
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
