magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
rect 209 295 445 331
<< pwell >>
rect 25 49 767 167
rect 0 0 768 49
<< scnmos >>
rect 108 57 138 141
rect 180 57 210 141
rect 266 57 296 141
rect 338 57 368 141
rect 424 57 454 141
rect 496 57 526 141
rect 582 57 612 141
rect 654 57 684 141
<< scpmoshvt >>
rect 84 409 134 609
rect 302 331 352 531
rect 520 409 570 609
rect 618 409 668 609
<< ndiff >>
rect 51 116 108 141
rect 51 82 63 116
rect 97 82 108 116
rect 51 57 108 82
rect 138 57 180 141
rect 210 116 266 141
rect 210 82 221 116
rect 255 82 266 116
rect 210 57 266 82
rect 296 57 338 141
rect 368 103 424 141
rect 368 69 379 103
rect 413 69 424 103
rect 368 57 424 69
rect 454 57 496 141
rect 526 116 582 141
rect 526 82 537 116
rect 571 82 582 116
rect 526 57 582 82
rect 612 57 654 141
rect 684 116 741 141
rect 684 82 695 116
rect 729 82 741 116
rect 684 57 741 82
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 573 191 609
rect 134 539 145 573
rect 179 539 191 573
rect 463 597 520 609
rect 463 563 475 597
rect 509 563 520 597
rect 134 409 191 539
rect 245 377 302 531
rect 245 343 257 377
rect 291 343 302 377
rect 245 331 302 343
rect 352 519 409 531
rect 352 485 363 519
rect 397 485 409 519
rect 352 448 409 485
rect 352 414 363 448
rect 397 414 409 448
rect 352 377 409 414
rect 463 526 520 563
rect 463 492 475 526
rect 509 492 520 526
rect 463 455 520 492
rect 463 421 475 455
rect 509 421 520 455
rect 463 409 520 421
rect 570 409 618 609
rect 668 597 725 609
rect 668 563 679 597
rect 713 563 725 597
rect 668 526 725 563
rect 668 492 679 526
rect 713 492 725 526
rect 668 455 725 492
rect 668 421 679 455
rect 713 421 725 455
rect 668 409 725 421
rect 352 343 363 377
rect 397 343 409 377
rect 352 331 409 343
<< ndiffc >>
rect 63 82 97 116
rect 221 82 255 116
rect 379 69 413 103
rect 537 82 571 116
rect 695 82 729 116
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 539 179 573
rect 475 563 509 597
rect 257 343 291 377
rect 363 485 397 519
rect 363 414 397 448
rect 475 492 509 526
rect 475 421 509 455
rect 679 563 713 597
rect 679 492 713 526
rect 679 421 713 455
rect 363 343 397 377
<< poly >>
rect 84 609 134 635
rect 520 609 570 635
rect 618 609 668 635
rect 302 531 352 557
rect 84 356 134 409
rect 72 340 138 356
rect 72 306 88 340
rect 122 306 138 340
rect 520 369 570 409
rect 496 353 570 369
rect 72 272 138 306
rect 72 238 88 272
rect 122 252 138 272
rect 302 291 352 331
rect 496 319 512 353
rect 546 319 570 353
rect 302 275 368 291
rect 302 255 318 275
rect 122 238 210 252
rect 72 222 210 238
rect 108 141 138 222
rect 180 141 210 222
rect 266 241 318 255
rect 352 241 368 275
rect 266 225 368 241
rect 266 141 296 225
rect 338 141 368 225
rect 496 285 570 319
rect 618 315 668 409
rect 496 251 512 285
rect 546 251 570 285
rect 496 235 570 251
rect 638 299 704 315
rect 638 265 654 299
rect 688 265 704 299
rect 496 186 526 235
rect 638 231 704 265
rect 638 197 654 231
rect 688 197 704 231
rect 638 187 704 197
rect 424 156 526 186
rect 424 141 454 156
rect 496 141 526 156
rect 582 157 704 187
rect 582 141 612 157
rect 654 141 684 157
rect 108 31 138 57
rect 180 31 210 57
rect 266 31 296 57
rect 338 31 368 57
rect 424 31 454 57
rect 496 31 526 57
rect 582 31 612 57
rect 654 31 684 57
<< polycont >>
rect 88 306 122 340
rect 88 238 122 272
rect 512 319 546 353
rect 318 241 352 275
rect 512 251 546 285
rect 654 265 688 299
rect 654 197 688 231
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 526 89 563
rect 23 492 39 526
rect 73 492 89 526
rect 129 597 525 613
rect 129 579 475 597
rect 129 573 195 579
rect 129 539 145 573
rect 179 539 195 573
rect 129 499 195 539
rect 459 563 475 579
rect 509 563 525 597
rect 347 519 413 535
rect 23 463 89 492
rect 347 485 363 519
rect 397 485 413 519
rect 347 463 413 485
rect 23 455 413 463
rect 23 421 39 455
rect 73 448 413 455
rect 73 429 363 448
rect 73 421 89 429
rect 23 405 89 421
rect 347 414 363 429
rect 397 414 413 448
rect 205 377 307 393
rect 25 340 167 356
rect 25 306 88 340
rect 122 306 167 340
rect 25 272 167 306
rect 25 238 88 272
rect 122 238 167 272
rect 25 222 167 238
rect 205 343 257 377
rect 291 343 307 377
rect 205 327 307 343
rect 347 377 413 414
rect 459 526 525 563
rect 459 492 475 526
rect 509 492 525 526
rect 459 455 525 492
rect 459 421 475 455
rect 509 421 525 455
rect 459 405 525 421
rect 663 597 729 649
rect 663 563 679 597
rect 713 563 729 597
rect 663 526 729 563
rect 663 492 679 526
rect 713 492 729 526
rect 663 455 729 492
rect 663 421 679 455
rect 713 421 729 455
rect 663 405 729 421
rect 347 343 363 377
rect 397 343 413 377
rect 347 327 413 343
rect 496 353 562 369
rect 205 189 263 327
rect 496 319 512 353
rect 546 319 562 353
rect 302 275 455 291
rect 302 241 318 275
rect 352 241 455 275
rect 302 225 455 241
rect 496 285 562 319
rect 496 251 512 285
rect 546 251 562 285
rect 496 235 562 251
rect 638 299 743 356
rect 638 265 654 299
rect 688 265 743 299
rect 638 231 743 265
rect 638 197 654 231
rect 688 197 743 231
rect 205 155 587 189
rect 638 181 743 197
rect 47 116 113 145
rect 47 82 63 116
rect 97 82 113 116
rect 47 17 113 82
rect 205 116 271 155
rect 205 82 221 116
rect 255 82 271 116
rect 205 53 271 82
rect 363 103 429 119
rect 363 69 379 103
rect 413 69 429 103
rect 363 17 429 69
rect 521 116 587 155
rect 521 82 537 116
rect 571 82 587 116
rect 521 53 587 82
rect 679 116 745 145
rect 679 82 695 116
rect 729 82 745 116
rect 679 17 745 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4_lp
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4353522
string GDS_START 4345902
<< end >>
