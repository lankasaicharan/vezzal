magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 1 157 268 289
rect 631 157 1055 235
rect 1 49 1055 157
rect 0 0 1056 49
<< scnmos >>
rect 83 179 113 263
rect 155 179 185 263
rect 339 47 369 131
rect 425 47 455 131
rect 511 47 541 131
rect 713 125 743 209
rect 785 125 815 209
rect 871 125 901 209
rect 943 125 973 209
<< scpmoshvt >>
rect 190 419 240 619
rect 296 419 346 619
rect 443 419 493 619
rect 557 419 607 619
rect 673 419 723 619
rect 779 419 829 619
rect 904 419 954 619
<< ndiff >>
rect 27 238 83 263
rect 27 204 38 238
rect 72 204 83 238
rect 27 179 83 204
rect 113 179 155 263
rect 185 241 242 263
rect 185 207 196 241
rect 230 207 242 241
rect 185 185 242 207
rect 185 179 235 185
rect 657 184 713 209
rect 289 125 339 131
rect 282 108 339 125
rect 282 74 294 108
rect 328 74 339 108
rect 282 47 339 74
rect 369 111 425 131
rect 369 77 380 111
rect 414 77 425 111
rect 369 47 425 77
rect 455 95 511 131
rect 455 61 466 95
rect 500 61 511 95
rect 455 47 511 61
rect 541 111 597 131
rect 541 77 552 111
rect 586 77 597 111
rect 541 47 597 77
rect 657 150 668 184
rect 702 150 713 184
rect 657 125 713 150
rect 743 125 785 209
rect 815 182 871 209
rect 815 148 826 182
rect 860 148 871 182
rect 815 125 871 148
rect 901 125 943 209
rect 973 182 1029 209
rect 973 148 984 182
rect 1018 148 1029 182
rect 973 125 1029 148
<< pdiff >>
rect 133 607 190 619
rect 133 573 145 607
rect 179 573 190 607
rect 133 536 190 573
rect 133 502 145 536
rect 179 502 190 536
rect 133 465 190 502
rect 133 431 145 465
rect 179 431 190 465
rect 133 419 190 431
rect 240 607 296 619
rect 240 573 251 607
rect 285 573 296 607
rect 240 536 296 573
rect 240 502 251 536
rect 285 502 296 536
rect 240 465 296 502
rect 240 431 251 465
rect 285 431 296 465
rect 240 419 296 431
rect 346 597 443 619
rect 346 563 357 597
rect 391 563 443 597
rect 346 465 443 563
rect 346 431 357 465
rect 391 431 443 465
rect 346 419 443 431
rect 493 419 557 619
rect 607 607 673 619
rect 607 573 618 607
rect 652 573 673 607
rect 607 512 673 573
rect 607 478 618 512
rect 652 478 673 512
rect 607 419 673 478
rect 723 597 779 619
rect 723 563 734 597
rect 768 563 779 597
rect 723 512 779 563
rect 723 478 734 512
rect 768 478 779 512
rect 723 419 779 478
rect 829 607 904 619
rect 829 573 859 607
rect 893 573 904 607
rect 829 536 904 573
rect 829 502 859 536
rect 893 502 904 536
rect 829 465 904 502
rect 829 431 859 465
rect 893 431 904 465
rect 829 419 904 431
rect 954 597 1011 619
rect 954 563 965 597
rect 999 563 1011 597
rect 954 465 1011 563
rect 954 431 965 465
rect 999 431 1011 465
rect 954 419 1011 431
<< ndiffc >>
rect 38 204 72 238
rect 196 207 230 241
rect 294 74 328 108
rect 380 77 414 111
rect 466 61 500 95
rect 552 77 586 111
rect 668 150 702 184
rect 826 148 860 182
rect 984 148 1018 182
<< pdiffc >>
rect 145 573 179 607
rect 145 502 179 536
rect 145 431 179 465
rect 251 573 285 607
rect 251 502 285 536
rect 251 431 285 465
rect 357 563 391 597
rect 357 431 391 465
rect 618 573 652 607
rect 618 478 652 512
rect 734 563 768 597
rect 734 478 768 512
rect 859 573 893 607
rect 859 502 893 536
rect 859 431 893 465
rect 965 563 999 597
rect 965 431 999 465
<< poly >>
rect 190 619 240 645
rect 296 619 346 645
rect 443 619 493 645
rect 557 619 607 645
rect 673 619 723 645
rect 779 619 829 645
rect 904 619 954 645
rect 190 386 240 419
rect 83 363 240 386
rect 83 356 190 363
rect 83 263 113 356
rect 155 329 190 356
rect 224 329 240 363
rect 155 313 240 329
rect 155 263 185 313
rect 296 286 346 419
rect 443 387 493 419
rect 439 371 509 387
rect 439 337 459 371
rect 493 337 509 371
rect 439 321 509 337
rect 557 356 607 419
rect 673 387 723 419
rect 671 371 737 387
rect 557 340 623 356
rect 316 270 397 286
rect 316 236 347 270
rect 381 236 397 270
rect 316 220 397 236
rect 83 153 113 179
rect 155 153 185 179
rect 339 131 369 220
rect 439 176 469 321
rect 557 306 573 340
rect 607 306 623 340
rect 671 337 687 371
rect 721 337 737 371
rect 671 321 737 337
rect 557 290 623 306
rect 557 176 587 290
rect 701 254 731 321
rect 779 302 829 419
rect 904 379 954 419
rect 799 254 829 302
rect 701 224 743 254
rect 713 209 743 224
rect 785 224 829 254
rect 871 363 973 379
rect 871 329 887 363
rect 921 329 973 363
rect 871 295 973 329
rect 871 261 887 295
rect 921 261 973 295
rect 871 245 973 261
rect 785 209 815 224
rect 871 209 901 245
rect 943 209 973 245
rect 425 146 469 176
rect 511 146 642 176
rect 425 131 455 146
rect 511 131 541 146
rect 612 51 642 146
rect 713 99 743 125
rect 785 51 815 125
rect 871 99 901 125
rect 943 99 973 125
rect 339 21 369 47
rect 425 21 455 47
rect 511 21 541 47
rect 612 21 815 51
<< polycont >>
rect 190 329 224 363
rect 459 337 493 371
rect 347 236 381 270
rect 573 306 607 340
rect 687 337 721 371
rect 887 329 921 363
rect 887 261 921 295
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 235 607 301 649
rect 22 573 145 607
rect 179 573 195 607
rect 22 238 88 573
rect 129 536 195 573
rect 129 502 145 536
rect 179 502 195 536
rect 129 465 195 502
rect 129 431 145 465
rect 179 431 195 465
rect 235 573 251 607
rect 285 573 301 607
rect 235 536 301 573
rect 235 502 251 536
rect 285 502 301 536
rect 235 465 301 502
rect 235 431 251 465
rect 285 431 301 465
rect 235 415 301 431
rect 341 597 407 613
rect 341 563 357 597
rect 391 563 407 597
rect 602 607 668 649
rect 341 465 407 563
rect 341 431 357 465
rect 391 431 407 465
rect 341 379 407 431
rect 174 363 407 379
rect 174 329 190 363
rect 224 345 407 363
rect 443 426 551 578
rect 602 573 618 607
rect 652 573 668 607
rect 602 512 668 573
rect 602 478 618 512
rect 652 478 668 512
rect 602 462 668 478
rect 718 597 807 613
rect 718 563 734 597
rect 768 563 807 597
rect 718 512 807 563
rect 718 478 734 512
rect 768 478 807 512
rect 718 462 807 478
rect 443 392 737 426
rect 443 371 509 392
rect 224 329 300 345
rect 174 313 300 329
rect 443 337 459 371
rect 493 337 509 371
rect 677 371 737 392
rect 443 321 509 337
rect 557 340 641 356
rect 22 204 38 238
rect 72 204 88 238
rect 22 88 88 204
rect 180 241 230 267
rect 180 207 196 241
rect 180 17 230 207
rect 266 129 300 313
rect 557 306 573 340
rect 607 306 641 340
rect 677 337 687 371
rect 721 337 737 371
rect 677 321 737 337
rect 557 290 641 306
rect 336 270 397 286
rect 773 279 807 462
rect 843 607 909 649
rect 843 573 859 607
rect 893 573 909 607
rect 843 536 909 573
rect 843 502 859 536
rect 893 502 909 536
rect 843 465 909 502
rect 843 431 859 465
rect 893 431 909 465
rect 843 415 909 431
rect 949 597 1034 613
rect 949 563 965 597
rect 999 563 1034 597
rect 949 465 1034 563
rect 949 431 965 465
rect 999 431 1034 465
rect 949 415 1034 431
rect 871 363 937 379
rect 871 329 887 363
rect 921 329 937 363
rect 871 295 937 329
rect 871 279 887 295
rect 336 236 347 270
rect 381 254 397 270
rect 684 261 887 279
rect 921 261 937 295
rect 684 254 937 261
rect 381 245 937 254
rect 381 236 718 245
rect 336 220 718 236
rect 652 184 718 220
rect 985 209 1034 415
rect 364 150 602 184
rect 266 108 328 129
rect 266 74 294 108
rect 266 53 328 74
rect 364 111 414 150
rect 364 77 380 111
rect 364 53 414 77
rect 450 95 516 114
rect 450 61 466 95
rect 500 61 516 95
rect 450 17 516 61
rect 552 111 602 150
rect 652 150 668 184
rect 702 150 718 184
rect 652 121 718 150
rect 810 182 876 209
rect 810 148 826 182
rect 860 148 876 182
rect 586 77 602 111
rect 552 53 602 77
rect 810 17 876 148
rect 968 182 1034 209
rect 968 148 984 182
rect 1018 148 1034 182
rect 968 88 1034 148
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ha_lp
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 991 94 1025 128 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 991 168 1025 202 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 991 464 1025 498 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 991 538 1025 572 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6704376
string GDS_START 6694866
<< end >>
