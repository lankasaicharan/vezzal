magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4178 1975
<< nwell >>
rect -38 331 2918 704
<< pwell >>
rect 741 231 1007 275
rect 2118 235 2314 279
rect 15 49 541 229
rect 741 49 1270 231
rect 1845 229 2314 235
rect 1452 199 2314 229
rect 2568 199 2859 273
rect 1452 49 2859 199
rect 0 0 2880 49
<< scnmos >>
rect 94 119 124 203
rect 166 119 196 203
rect 274 119 304 203
rect 346 119 376 203
rect 432 119 462 203
rect 824 121 854 249
rect 1003 121 1033 205
rect 1075 121 1105 205
rect 1161 121 1191 205
rect 1531 119 1561 203
rect 1617 119 1647 203
rect 1924 125 1954 209
rect 2010 125 2040 209
rect 2082 125 2112 209
rect 2201 125 2231 253
rect 2457 89 2487 173
rect 2647 79 2677 247
rect 2736 79 2766 247
<< scpmoshvt >>
rect 80 483 110 611
rect 166 483 196 611
rect 238 483 268 611
rect 324 483 354 611
rect 621 481 651 609
rect 839 425 869 593
rect 944 425 974 509
rect 1186 501 1216 585
rect 1272 501 1302 585
rect 1522 391 1552 519
rect 1639 391 1669 519
rect 1843 497 1873 581
rect 1967 379 1997 547
rect 2157 441 2187 525
rect 2262 379 2292 547
rect 2462 367 2492 495
rect 2567 367 2597 619
rect 2770 367 2800 619
<< ndiff >>
rect 41 178 94 203
rect 41 144 49 178
rect 83 144 94 178
rect 41 119 94 144
rect 124 119 166 203
rect 196 178 274 203
rect 196 144 218 178
rect 252 144 274 178
rect 196 119 274 144
rect 304 119 346 203
rect 376 163 432 203
rect 376 129 387 163
rect 421 129 432 163
rect 376 119 432 129
rect 462 178 515 203
rect 462 144 473 178
rect 507 144 515 178
rect 462 119 515 144
rect 767 241 824 249
rect 767 207 779 241
rect 813 207 824 241
rect 767 173 824 207
rect 767 139 779 173
rect 813 139 824 173
rect 767 121 824 139
rect 854 231 981 249
rect 854 197 931 231
rect 965 205 981 231
rect 965 197 1003 205
rect 854 163 1003 197
rect 854 129 931 163
rect 965 129 1003 163
rect 854 121 1003 129
rect 1033 121 1075 205
rect 1105 180 1161 205
rect 1105 146 1116 180
rect 1150 146 1161 180
rect 1105 121 1161 146
rect 1191 180 1244 205
rect 1191 146 1202 180
rect 1236 146 1244 180
rect 1478 173 1531 203
rect 1191 121 1244 146
rect 1478 139 1486 173
rect 1520 139 1531 173
rect 1478 119 1531 139
rect 1561 174 1617 203
rect 1561 140 1572 174
rect 1606 140 1617 174
rect 1561 119 1617 140
rect 1647 173 1700 203
rect 2144 239 2201 253
rect 2144 209 2152 239
rect 1871 184 1924 209
rect 1647 139 1658 173
rect 1692 139 1700 173
rect 1647 119 1700 139
rect 1871 150 1879 184
rect 1913 150 1924 184
rect 1871 125 1924 150
rect 1954 197 2010 209
rect 1954 163 1965 197
rect 1999 163 2010 197
rect 1954 125 2010 163
rect 2040 125 2082 209
rect 2112 205 2152 209
rect 2186 205 2201 239
rect 2112 171 2201 205
rect 2112 137 2152 171
rect 2186 137 2201 171
rect 2112 125 2201 137
rect 2231 237 2288 253
rect 2231 203 2242 237
rect 2276 203 2288 237
rect 2231 169 2288 203
rect 2231 135 2242 169
rect 2276 135 2288 169
rect 2231 125 2288 135
rect 2594 235 2647 247
rect 2594 201 2602 235
rect 2636 201 2647 235
rect 2404 145 2457 173
rect 2404 111 2412 145
rect 2446 111 2457 145
rect 2404 89 2457 111
rect 2487 145 2540 173
rect 2487 111 2498 145
rect 2532 111 2540 145
rect 2487 89 2540 111
rect 2594 125 2647 201
rect 2594 91 2602 125
rect 2636 91 2647 125
rect 2594 79 2647 91
rect 2677 219 2736 247
rect 2677 185 2691 219
rect 2725 185 2736 219
rect 2677 125 2736 185
rect 2677 91 2691 125
rect 2725 91 2736 125
rect 2677 79 2736 91
rect 2766 212 2833 247
rect 2766 178 2777 212
rect 2811 178 2833 212
rect 2766 125 2833 178
rect 2766 91 2777 125
rect 2811 91 2833 125
rect 2766 79 2833 91
<< pdiff >>
rect 27 597 80 611
rect 27 563 35 597
rect 69 563 80 597
rect 27 529 80 563
rect 27 495 35 529
rect 69 495 80 529
rect 27 483 80 495
rect 110 568 166 611
rect 110 534 121 568
rect 155 534 166 568
rect 110 483 166 534
rect 196 483 238 611
rect 268 603 324 611
rect 268 569 279 603
rect 313 569 324 603
rect 268 483 324 569
rect 354 529 407 611
rect 354 495 365 529
rect 399 495 407 529
rect 354 483 407 495
rect 517 529 621 609
rect 517 495 525 529
rect 559 495 621 529
rect 517 481 621 495
rect 651 595 707 609
rect 651 561 665 595
rect 699 561 707 595
rect 651 481 707 561
rect 767 441 839 593
rect 767 407 775 441
rect 809 425 839 441
rect 869 581 922 593
rect 869 547 880 581
rect 914 547 922 581
rect 869 509 922 547
rect 996 581 1046 593
rect 996 547 1004 581
rect 1038 547 1046 581
rect 996 509 1046 547
rect 869 425 944 509
rect 974 425 1046 509
rect 1113 543 1186 585
rect 1113 509 1125 543
rect 1159 509 1186 543
rect 1113 501 1186 509
rect 1216 543 1272 585
rect 1216 509 1227 543
rect 1261 509 1272 543
rect 1216 501 1272 509
rect 1302 573 1371 585
rect 1302 539 1329 573
rect 1363 539 1371 573
rect 1574 573 1624 585
rect 1302 501 1371 539
rect 1574 539 1582 573
rect 1616 539 1624 573
rect 1574 519 1624 539
rect 809 407 817 425
rect 767 395 817 407
rect 1465 433 1522 519
rect 1465 399 1477 433
rect 1511 399 1522 433
rect 1465 391 1522 399
rect 1552 391 1639 519
rect 1669 433 1726 519
rect 1669 399 1680 433
rect 1714 399 1726 433
rect 1669 391 1726 399
rect 1786 573 1843 581
rect 1786 539 1798 573
rect 1832 539 1843 573
rect 1786 497 1843 539
rect 1873 547 1945 581
rect 1873 497 1967 547
rect 1914 427 1967 497
rect 1914 393 1922 427
rect 1956 393 1967 427
rect 1914 379 1967 393
rect 1997 495 2050 547
rect 2209 535 2262 547
rect 2209 525 2217 535
rect 1997 461 2008 495
rect 2042 461 2050 495
rect 1997 425 2050 461
rect 2104 499 2157 525
rect 2104 465 2112 499
rect 2146 465 2157 499
rect 2104 441 2157 465
rect 2187 501 2217 525
rect 2251 501 2262 535
rect 2187 463 2262 501
rect 2187 441 2217 463
rect 1997 391 2008 425
rect 2042 391 2050 425
rect 1997 379 2050 391
rect 2209 429 2217 441
rect 2251 429 2262 463
rect 2209 379 2262 429
rect 2292 535 2349 547
rect 2292 501 2307 535
rect 2341 501 2349 535
rect 2292 425 2349 501
rect 2292 391 2307 425
rect 2341 391 2349 425
rect 2292 379 2349 391
rect 2514 571 2567 619
rect 2514 537 2522 571
rect 2556 537 2567 571
rect 2514 495 2567 537
rect 2409 483 2462 495
rect 2409 449 2417 483
rect 2451 449 2462 483
rect 2409 413 2462 449
rect 2409 379 2417 413
rect 2451 379 2462 413
rect 2409 367 2462 379
rect 2492 367 2567 495
rect 2597 413 2650 619
rect 2597 379 2608 413
rect 2642 379 2650 413
rect 2597 367 2650 379
rect 2717 571 2770 619
rect 2717 537 2725 571
rect 2759 537 2770 571
rect 2717 367 2770 537
rect 2800 599 2853 619
rect 2800 565 2811 599
rect 2845 565 2853 599
rect 2800 506 2853 565
rect 2800 472 2811 506
rect 2845 472 2853 506
rect 2800 413 2853 472
rect 2800 379 2811 413
rect 2845 379 2853 413
rect 2800 367 2853 379
<< ndiffc >>
rect 49 144 83 178
rect 218 144 252 178
rect 387 129 421 163
rect 473 144 507 178
rect 779 207 813 241
rect 779 139 813 173
rect 931 197 965 231
rect 931 129 965 163
rect 1116 146 1150 180
rect 1202 146 1236 180
rect 1486 139 1520 173
rect 1572 140 1606 174
rect 1658 139 1692 173
rect 1879 150 1913 184
rect 1965 163 1999 197
rect 2152 205 2186 239
rect 2152 137 2186 171
rect 2242 203 2276 237
rect 2242 135 2276 169
rect 2602 201 2636 235
rect 2412 111 2446 145
rect 2498 111 2532 145
rect 2602 91 2636 125
rect 2691 185 2725 219
rect 2691 91 2725 125
rect 2777 178 2811 212
rect 2777 91 2811 125
<< pdiffc >>
rect 35 563 69 597
rect 35 495 69 529
rect 121 534 155 568
rect 279 569 313 603
rect 365 495 399 529
rect 525 495 559 529
rect 665 561 699 595
rect 775 407 809 441
rect 880 547 914 581
rect 1004 547 1038 581
rect 1125 509 1159 543
rect 1227 509 1261 543
rect 1329 539 1363 573
rect 1582 539 1616 573
rect 1477 399 1511 433
rect 1680 399 1714 433
rect 1798 539 1832 573
rect 1922 393 1956 427
rect 2008 461 2042 495
rect 2112 465 2146 499
rect 2217 501 2251 535
rect 2008 391 2042 425
rect 2217 429 2251 463
rect 2307 501 2341 535
rect 2307 391 2341 425
rect 2522 537 2556 571
rect 2417 449 2451 483
rect 2417 379 2451 413
rect 2608 379 2642 413
rect 2725 537 2759 571
rect 2811 565 2845 599
rect 2811 472 2845 506
rect 2811 379 2845 413
<< poly >>
rect 80 611 110 637
rect 166 611 196 637
rect 238 611 268 637
rect 324 611 354 637
rect 621 609 651 635
rect 722 615 1098 645
rect 80 376 110 483
rect 44 360 110 376
rect 44 326 60 360
rect 94 326 110 360
rect 44 292 110 326
rect 44 258 60 292
rect 94 272 110 292
rect 94 258 124 272
rect 44 242 124 258
rect 94 203 124 242
rect 166 203 196 483
rect 238 389 268 483
rect 324 461 354 483
rect 324 433 571 461
rect 324 431 521 433
rect 346 389 384 431
rect 505 399 521 431
rect 555 399 571 433
rect 238 373 304 389
rect 238 339 254 373
rect 288 339 304 373
rect 238 305 304 339
rect 238 271 254 305
rect 288 271 304 305
rect 238 255 304 271
rect 274 203 304 255
rect 346 203 376 389
rect 505 365 571 399
rect 505 331 521 365
rect 555 331 571 365
rect 505 315 571 331
rect 432 203 462 229
rect 621 187 651 481
rect 585 171 651 187
rect 585 137 601 171
rect 635 137 651 171
rect 94 93 124 119
rect 166 51 196 119
rect 274 93 304 119
rect 346 93 376 119
rect 432 51 462 119
rect 585 103 651 137
rect 585 69 601 103
rect 635 69 651 103
rect 585 51 651 69
rect 166 21 651 51
rect 722 301 752 615
rect 839 593 869 615
rect 944 509 974 535
rect 1068 457 1098 615
rect 1186 585 1216 611
rect 1272 607 1771 637
rect 1272 585 1302 607
rect 1522 519 1552 545
rect 1639 519 1669 545
rect 1068 441 1144 457
rect 839 399 869 425
rect 944 387 974 425
rect 1068 407 1094 441
rect 1128 407 1144 441
rect 1068 391 1144 407
rect 1186 433 1216 501
rect 1272 475 1302 501
rect 1186 417 1433 433
rect 944 371 1010 387
rect 944 337 960 371
rect 994 343 1010 371
rect 1186 383 1383 417
rect 1417 383 1433 417
rect 1186 349 1433 383
rect 1522 359 1552 391
rect 994 337 1033 343
rect 944 313 1033 337
rect 1186 335 1383 349
rect 722 271 854 301
rect 722 53 752 271
rect 824 249 854 271
rect 1003 205 1033 313
rect 1075 315 1383 335
rect 1417 315 1433 349
rect 1075 305 1433 315
rect 1075 205 1105 305
rect 1216 299 1433 305
rect 1481 343 1552 359
rect 1481 309 1497 343
rect 1531 309 1552 343
rect 1481 291 1552 309
rect 1639 292 1669 391
rect 1741 313 1771 607
rect 1843 615 2394 645
rect 2567 619 2597 645
rect 2770 619 2800 645
rect 1843 581 1873 615
rect 1967 547 1997 573
rect 1843 471 1873 497
rect 2157 525 2187 551
rect 2262 547 2292 573
rect 2157 419 2187 441
rect 2082 393 2187 419
rect 1967 313 1997 379
rect 2082 359 2098 393
rect 2132 389 2187 393
rect 2132 359 2148 389
rect 2082 343 2148 359
rect 1731 297 2032 313
rect 1481 275 1561 291
rect 1481 257 1497 275
rect 1161 241 1497 257
rect 1531 241 1561 275
rect 1161 227 1561 241
rect 1161 205 1191 227
rect 1481 225 1561 227
rect 1531 203 1561 225
rect 1617 276 1683 292
rect 1617 242 1633 276
rect 1667 242 1683 276
rect 1617 226 1683 242
rect 1731 263 1747 297
rect 1781 295 2032 297
rect 1781 283 2040 295
rect 1781 263 1797 283
rect 2002 265 2040 283
rect 1731 229 1797 263
rect 1617 203 1647 226
rect 1276 155 1342 171
rect 1276 121 1292 155
rect 1326 121 1342 155
rect 824 95 854 121
rect 1003 95 1033 121
rect 1075 95 1105 121
rect 1161 95 1191 121
rect 1276 87 1342 121
rect 1276 53 1292 87
rect 1326 53 1342 87
rect 722 23 1342 53
rect 1390 157 1456 173
rect 1390 123 1406 157
rect 1440 123 1456 157
rect 1390 87 1456 123
rect 1731 195 1747 229
rect 1781 195 1797 229
rect 1924 209 1954 235
rect 2010 209 2040 265
rect 2082 209 2112 343
rect 2262 341 2292 379
rect 2201 325 2292 341
rect 2201 291 2217 325
rect 2251 291 2292 325
rect 2201 275 2292 291
rect 2201 253 2231 275
rect 1731 179 1797 195
rect 2364 218 2394 615
rect 2462 495 2492 521
rect 2462 329 2492 367
rect 2567 329 2597 367
rect 2770 335 2800 367
rect 2340 188 2394 218
rect 2442 313 2677 329
rect 2442 279 2458 313
rect 2492 299 2677 313
rect 2492 279 2508 299
rect 2442 245 2508 279
rect 2647 247 2677 299
rect 2725 319 2800 335
rect 2725 285 2741 319
rect 2775 285 2800 319
rect 2725 269 2800 285
rect 2736 247 2766 269
rect 2442 211 2458 245
rect 2492 211 2508 245
rect 2442 195 2508 211
rect 1531 93 1561 119
rect 1617 93 1647 119
rect 1390 53 1406 87
rect 1440 53 1456 87
rect 1390 51 1456 53
rect 1924 51 1954 125
rect 2010 99 2040 125
rect 2082 99 2112 125
rect 2201 99 2231 125
rect 2340 51 2370 188
rect 2457 173 2487 195
rect 2457 63 2487 89
rect 2647 53 2677 79
rect 2736 53 2766 79
rect 1390 21 2370 51
<< polycont >>
rect 60 326 94 360
rect 60 258 94 292
rect 521 399 555 433
rect 254 339 288 373
rect 254 271 288 305
rect 521 331 555 365
rect 601 137 635 171
rect 601 69 635 103
rect 1094 407 1128 441
rect 960 337 994 371
rect 1383 383 1417 417
rect 1383 315 1417 349
rect 1497 309 1531 343
rect 2098 359 2132 393
rect 1497 241 1531 275
rect 1633 242 1667 276
rect 1747 263 1781 297
rect 1292 121 1326 155
rect 1292 53 1326 87
rect 1406 123 1440 157
rect 1747 195 1781 229
rect 2217 291 2251 325
rect 2458 279 2492 313
rect 2741 285 2775 319
rect 2458 211 2492 245
rect 1406 53 1440 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 19 597 71 613
rect 19 563 35 597
rect 69 563 71 597
rect 19 529 71 563
rect 19 495 35 529
rect 69 495 71 529
rect 105 568 171 649
rect 105 534 121 568
rect 155 534 171 568
rect 263 603 629 613
rect 263 569 279 603
rect 313 579 629 603
rect 313 569 485 579
rect 263 567 485 569
rect 105 526 171 534
rect 349 529 415 533
rect 19 492 71 495
rect 349 495 365 529
rect 399 495 415 529
rect 349 492 415 495
rect 19 458 415 492
rect 17 360 110 424
rect 17 326 60 360
rect 94 326 110 360
rect 17 292 110 326
rect 17 258 60 292
rect 94 258 110 292
rect 204 373 304 424
rect 204 339 254 373
rect 288 339 304 373
rect 204 305 304 339
rect 204 271 254 305
rect 288 271 304 305
rect 451 283 485 567
rect 204 269 304 271
rect 17 228 110 258
rect 340 241 485 283
rect 519 529 561 545
rect 519 495 525 529
rect 559 495 561 529
rect 519 433 561 495
rect 519 399 521 433
rect 555 399 561 433
rect 519 365 561 399
rect 519 331 521 365
rect 555 331 561 365
rect 340 235 374 241
rect 202 201 374 235
rect 33 178 99 194
rect 33 144 49 178
rect 83 144 99 178
rect 33 17 99 144
rect 202 178 268 201
rect 519 194 561 331
rect 595 511 629 579
rect 663 595 715 649
rect 663 561 665 595
rect 699 561 715 595
rect 663 545 715 561
rect 864 581 930 649
rect 864 547 880 581
rect 914 547 930 581
rect 864 545 930 547
rect 988 581 1379 613
rect 988 547 1004 581
rect 1038 579 1379 581
rect 1038 547 1054 579
rect 988 545 1054 547
rect 1313 573 1379 579
rect 1109 543 1175 545
rect 1109 511 1125 543
rect 595 509 1125 511
rect 1159 509 1175 543
rect 595 477 1175 509
rect 1211 543 1277 545
rect 1211 509 1227 543
rect 1261 509 1277 543
rect 1313 539 1329 573
rect 1363 539 1379 573
rect 1313 537 1379 539
rect 1566 573 1632 649
rect 1566 539 1582 573
rect 1616 539 1632 573
rect 1566 537 1632 539
rect 1782 573 2162 589
rect 1782 539 1798 573
rect 1832 545 2162 573
rect 1832 539 1848 545
rect 1782 537 1848 539
rect 595 346 629 477
rect 1211 443 1277 509
rect 2004 503 2048 511
rect 759 441 1010 443
rect 759 407 775 441
rect 809 407 1010 441
rect 759 371 1010 407
rect 1078 441 1277 443
rect 1078 407 1094 441
rect 1128 407 1277 441
rect 1078 405 1277 407
rect 1313 495 2048 503
rect 1313 469 2008 495
rect 1313 371 1347 469
rect 1664 433 1783 435
rect 595 312 711 346
rect 202 144 218 178
rect 252 144 268 178
rect 471 178 561 194
rect 202 128 268 144
rect 371 163 437 167
rect 371 129 387 163
rect 421 129 437 163
rect 371 17 437 129
rect 471 144 473 178
rect 507 144 561 178
rect 471 128 561 144
rect 595 171 643 278
rect 595 137 601 171
rect 635 137 643 171
rect 595 103 643 137
rect 595 69 601 103
rect 635 69 643 103
rect 595 53 643 69
rect 677 87 711 312
rect 759 337 960 371
rect 994 337 1347 371
rect 1381 417 1477 433
rect 1381 383 1383 417
rect 1417 399 1477 417
rect 1511 399 1527 433
rect 1417 395 1527 399
rect 1664 399 1680 433
rect 1714 399 1783 433
rect 1417 383 1433 395
rect 1381 349 1433 383
rect 1664 359 1783 399
rect 759 241 813 337
rect 1381 315 1383 349
rect 1417 315 1433 349
rect 759 207 779 241
rect 759 173 813 207
rect 759 139 779 173
rect 759 123 813 139
rect 847 267 1240 301
rect 847 87 881 267
rect 677 53 881 87
rect 915 231 981 233
rect 915 197 931 231
rect 965 197 981 231
rect 915 163 981 197
rect 915 129 931 163
rect 965 129 981 163
rect 915 17 981 129
rect 1100 180 1159 196
rect 1100 146 1116 180
rect 1150 146 1159 180
rect 1100 87 1159 146
rect 1193 180 1240 267
rect 1193 146 1202 180
rect 1236 146 1240 180
rect 1381 189 1433 315
rect 1481 343 1783 359
rect 1481 309 1497 343
rect 1531 325 1783 343
rect 1481 275 1531 309
rect 1738 297 1783 325
rect 1481 241 1497 275
rect 1481 225 1531 241
rect 1565 276 1704 291
rect 1565 242 1633 276
rect 1667 242 1704 276
rect 1565 224 1704 242
rect 1738 263 1747 297
rect 1781 263 1783 297
rect 1738 229 1783 263
rect 1738 195 1747 229
rect 1781 195 1783 229
rect 1381 173 1527 189
rect 1193 130 1240 146
rect 1276 155 1342 171
rect 1276 121 1292 155
rect 1326 121 1342 155
rect 1381 157 1486 173
rect 1381 123 1406 157
rect 1440 139 1486 157
rect 1520 139 1527 173
rect 1440 123 1527 139
rect 1561 174 1616 190
rect 1738 189 1783 195
rect 1561 140 1572 174
rect 1606 140 1616 174
rect 1276 87 1342 121
rect 1100 53 1292 87
rect 1326 53 1342 87
rect 1100 51 1342 53
rect 1390 87 1456 123
rect 1390 53 1406 87
rect 1440 53 1456 87
rect 1390 51 1456 53
rect 1561 17 1616 140
rect 1650 173 1783 189
rect 1650 139 1658 173
rect 1692 139 1783 173
rect 1650 123 1783 139
rect 1817 200 1851 469
rect 2006 461 2008 469
rect 2042 461 2048 495
rect 1906 427 1972 435
rect 1906 393 1922 427
rect 1956 393 1972 427
rect 1906 323 1972 393
rect 2006 425 2048 461
rect 2096 499 2162 545
rect 2096 465 2112 499
rect 2146 465 2162 499
rect 2096 449 2162 465
rect 2196 535 2267 649
rect 2506 571 2572 649
rect 2196 501 2217 535
rect 2251 501 2267 535
rect 2196 463 2267 501
rect 2196 429 2217 463
rect 2251 429 2267 463
rect 2301 535 2357 551
rect 2301 501 2307 535
rect 2341 501 2357 535
rect 2506 537 2522 571
rect 2556 537 2572 571
rect 2506 533 2572 537
rect 2709 571 2775 649
rect 2709 537 2725 571
rect 2759 537 2775 571
rect 2709 533 2775 537
rect 2809 599 2863 615
rect 2809 565 2811 599
rect 2845 565 2863 599
rect 2006 391 2008 425
rect 2042 391 2048 425
rect 2301 425 2357 501
rect 2809 506 2863 565
rect 2301 395 2307 425
rect 2006 375 2048 391
rect 2082 393 2307 395
rect 2082 359 2098 393
rect 2132 391 2307 393
rect 2341 391 2357 425
rect 2132 361 2357 391
rect 2401 483 2775 499
rect 2401 449 2417 483
rect 2451 465 2775 483
rect 2451 449 2562 465
rect 2401 413 2562 449
rect 2401 379 2417 413
rect 2451 379 2562 413
rect 2401 363 2562 379
rect 2132 359 2148 361
rect 2082 357 2148 359
rect 2301 329 2357 361
rect 2201 325 2267 327
rect 2201 323 2217 325
rect 1906 291 2217 323
rect 2251 291 2267 325
rect 1906 289 2267 291
rect 2301 313 2492 329
rect 1817 184 1915 200
rect 1817 150 1879 184
rect 1913 150 1915 184
rect 1949 197 2015 289
rect 2301 279 2458 313
rect 2301 253 2492 279
rect 2236 245 2492 253
rect 1949 163 1965 197
rect 1999 163 2015 197
rect 1949 159 2015 163
rect 2136 239 2202 243
rect 2136 205 2152 239
rect 2186 205 2202 239
rect 2136 171 2202 205
rect 1817 134 1915 150
rect 2136 137 2152 171
rect 2186 137 2202 171
rect 2136 17 2202 137
rect 2236 237 2458 245
rect 2236 203 2242 237
rect 2276 211 2458 237
rect 2276 203 2492 211
rect 2236 195 2492 203
rect 2236 169 2337 195
rect 2236 135 2242 169
rect 2276 135 2337 169
rect 2528 161 2562 363
rect 2236 119 2337 135
rect 2396 145 2454 161
rect 2396 111 2412 145
rect 2446 111 2454 145
rect 2396 17 2454 111
rect 2488 145 2562 161
rect 2488 111 2498 145
rect 2532 111 2562 145
rect 2488 95 2562 111
rect 2598 413 2681 429
rect 2598 379 2608 413
rect 2642 379 2681 413
rect 2598 269 2681 379
rect 2725 319 2775 465
rect 2725 285 2741 319
rect 2725 269 2775 285
rect 2809 472 2811 506
rect 2845 472 2863 506
rect 2809 413 2863 472
rect 2809 379 2811 413
rect 2845 379 2863 413
rect 2598 235 2657 269
rect 2809 235 2863 379
rect 2598 201 2602 235
rect 2636 201 2657 235
rect 2598 125 2657 201
rect 2598 91 2602 125
rect 2636 91 2657 125
rect 2598 75 2657 91
rect 2691 219 2735 235
rect 2725 185 2735 219
rect 2691 125 2735 185
rect 2725 91 2735 125
rect 2691 17 2735 91
rect 2769 212 2863 235
rect 2769 178 2777 212
rect 2811 178 2863 212
rect 2769 125 2863 178
rect 2769 91 2777 125
rect 2811 91 2863 125
rect 2769 75 2863 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfxbp_1
flabel comment s 734 338 734 338 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2815 94 2849 128 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2815 168 2849 202 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2815 242 2849 276 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2815 316 2849 350 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2815 390 2849 424 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2815 464 2849 498 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2815 538 2849 572 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2623 94 2657 128 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2623 168 2657 202 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2623 242 2657 276 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2623 316 2657 350 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2623 390 2657 424 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2880 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6083620
string GDS_START 6063196
<< end >>
