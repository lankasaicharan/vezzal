magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2310 1852
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 67 989 203
rect 1 21 787 67
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 187 47 217 177
rect 271 47 301 177
rect 375 47 405 177
rect 571 47 601 177
rect 665 47 695 177
rect 871 93 901 177
<< scpmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 573 297 609 497
rect 667 297 703 497
rect 873 297 909 381
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 187 177
rect 113 129 133 163
rect 167 129 187 163
rect 113 95 187 129
rect 113 61 133 95
rect 167 61 187 95
rect 113 47 187 61
rect 217 95 271 177
rect 217 61 227 95
rect 261 61 271 95
rect 217 47 271 61
rect 301 163 375 177
rect 301 129 321 163
rect 355 129 375 163
rect 301 95 375 129
rect 301 61 321 95
rect 355 61 375 95
rect 301 47 375 61
rect 405 95 457 177
rect 405 61 415 95
rect 449 61 457 95
rect 405 47 457 61
rect 511 95 571 177
rect 511 61 519 95
rect 553 61 571 95
rect 511 47 571 61
rect 601 163 665 177
rect 601 129 621 163
rect 655 129 665 163
rect 601 95 665 129
rect 601 61 621 95
rect 655 61 665 95
rect 601 47 665 61
rect 695 163 761 177
rect 695 129 715 163
rect 749 129 761 163
rect 695 95 761 129
rect 695 61 715 95
rect 749 61 761 95
rect 819 149 871 177
rect 819 115 827 149
rect 861 115 871 149
rect 819 93 871 115
rect 901 149 963 177
rect 901 115 921 149
rect 955 115 963 149
rect 901 93 963 115
rect 695 47 761 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 409 179 443
rect 121 375 133 409
rect 167 375 179 409
rect 121 297 179 375
rect 215 477 273 497
rect 215 443 227 477
rect 261 443 273 477
rect 215 409 273 443
rect 215 375 227 409
rect 261 375 273 409
rect 215 341 273 375
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 309 477 367 497
rect 309 443 321 477
rect 355 443 367 477
rect 309 409 367 443
rect 309 375 321 409
rect 355 375 367 409
rect 309 297 367 375
rect 403 407 461 497
rect 403 373 415 407
rect 449 373 461 407
rect 403 339 461 373
rect 403 305 415 339
rect 449 305 461 339
rect 403 297 461 305
rect 515 489 573 497
rect 515 455 527 489
rect 561 455 573 489
rect 515 297 573 455
rect 609 409 667 497
rect 609 375 621 409
rect 655 375 667 409
rect 609 341 667 375
rect 609 307 621 341
rect 655 307 667 341
rect 609 297 667 307
rect 703 477 761 497
rect 703 443 715 477
rect 749 443 761 477
rect 703 409 761 443
rect 703 375 715 409
rect 749 375 761 409
rect 703 341 761 375
rect 703 307 715 341
rect 749 307 761 341
rect 703 297 761 307
rect 819 358 873 381
rect 819 324 827 358
rect 861 324 873 358
rect 819 297 873 324
rect 909 358 963 381
rect 909 324 921 358
rect 955 324 963 358
rect 909 297 963 324
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 129 167 163
rect 133 61 167 95
rect 227 61 261 95
rect 321 129 355 163
rect 321 61 355 95
rect 415 61 449 95
rect 519 61 553 95
rect 621 129 655 163
rect 621 61 655 95
rect 715 129 749 163
rect 715 61 749 95
rect 827 115 861 149
rect 921 115 955 149
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 443 167 477
rect 133 375 167 409
rect 227 443 261 477
rect 227 375 261 409
rect 227 307 261 341
rect 321 443 355 477
rect 321 375 355 409
rect 415 373 449 407
rect 415 305 449 339
rect 527 455 561 489
rect 621 375 655 409
rect 621 307 655 341
rect 715 443 749 477
rect 715 375 749 409
rect 715 307 749 341
rect 827 324 861 358
rect 921 324 955 358
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 573 497 609 523
rect 667 497 703 523
rect 873 381 909 407
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 573 282 609 297
rect 667 282 703 297
rect 873 282 909 297
rect 83 265 123 282
rect 177 265 217 282
rect 83 249 217 265
rect 83 215 112 249
rect 146 215 217 249
rect 83 199 217 215
rect 83 177 113 199
rect 187 177 217 199
rect 271 265 311 282
rect 365 265 405 282
rect 271 249 405 265
rect 271 215 318 249
rect 352 215 405 249
rect 271 199 405 215
rect 271 177 301 199
rect 375 177 405 199
rect 571 265 611 282
rect 665 265 705 282
rect 871 265 911 282
rect 571 249 767 265
rect 571 215 723 249
rect 757 215 767 249
rect 571 199 767 215
rect 871 249 936 265
rect 871 215 882 249
rect 916 215 936 249
rect 871 199 936 215
rect 571 177 601 199
rect 665 177 695 199
rect 871 177 901 199
rect 871 67 901 93
rect 83 21 113 47
rect 187 21 217 47
rect 271 21 301 47
rect 375 21 405 47
rect 571 21 601 47
rect 665 21 695 47
<< polycont >>
rect 112 215 146 249
rect 318 215 352 249
rect 723 215 757 249
rect 882 215 916 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 18 477 81 493
rect 18 443 39 477
rect 73 443 81 477
rect 18 409 81 443
rect 18 375 39 409
rect 73 375 81 409
rect 18 341 81 375
rect 125 477 175 527
rect 125 443 133 477
rect 167 443 175 477
rect 125 409 175 443
rect 125 375 133 409
rect 167 375 175 409
rect 125 359 175 375
rect 219 477 269 493
rect 219 443 227 477
rect 261 443 269 477
rect 219 409 269 443
rect 219 375 227 409
rect 261 375 269 409
rect 18 307 39 341
rect 73 325 81 341
rect 219 341 269 375
rect 313 489 756 493
rect 313 477 527 489
rect 313 443 321 477
rect 355 455 527 477
rect 561 477 756 489
rect 561 455 715 477
rect 355 443 363 455
rect 313 409 363 443
rect 707 443 715 455
rect 749 443 756 477
rect 707 409 756 443
rect 313 375 321 409
rect 355 375 363 409
rect 313 359 363 375
rect 399 373 415 407
rect 449 373 465 407
rect 219 325 227 341
rect 73 307 227 325
rect 261 325 269 341
rect 399 339 465 373
rect 399 325 415 339
rect 261 307 415 325
rect 18 305 415 307
rect 449 305 465 339
rect 18 291 465 305
rect 574 375 621 409
rect 655 375 671 409
rect 574 341 671 375
rect 574 307 621 341
rect 655 307 671 341
rect 22 249 203 257
rect 22 215 112 249
rect 146 215 203 249
rect 247 249 440 257
rect 247 215 318 249
rect 352 215 440 249
rect 574 181 671 307
rect 707 375 715 409
rect 749 375 756 409
rect 707 341 756 375
rect 707 307 715 341
rect 749 307 756 341
rect 707 291 756 307
rect 798 358 869 374
rect 798 324 827 358
rect 861 324 869 358
rect 798 291 869 324
rect 913 358 963 527
rect 913 324 921 358
rect 955 324 963 358
rect 913 308 963 324
rect 798 257 832 291
rect 707 249 832 257
rect 707 215 723 249
rect 757 215 832 249
rect 866 249 983 257
rect 866 215 882 249
rect 916 215 983 249
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 671 181
rect 798 181 832 215
rect 107 129 133 163
rect 167 145 321 163
rect 167 129 183 145
rect 107 95 183 129
rect 295 129 321 145
rect 355 145 621 163
rect 355 129 371 145
rect 107 61 133 95
rect 167 61 183 95
rect 107 51 183 61
rect 227 95 261 111
rect 227 17 261 61
rect 295 95 371 129
rect 587 129 621 145
rect 655 129 671 163
rect 295 61 321 95
rect 355 61 371 95
rect 295 51 371 61
rect 415 95 553 111
rect 449 61 519 95
rect 415 17 553 61
rect 587 95 671 129
rect 587 61 621 95
rect 655 61 671 95
rect 587 51 671 61
rect 715 163 756 179
rect 749 129 756 163
rect 715 95 756 129
rect 749 61 756 95
rect 798 149 869 181
rect 798 115 827 149
rect 861 115 869 149
rect 798 76 869 115
rect 913 149 971 165
rect 913 115 921 149
rect 955 115 971 149
rect 715 17 756 61
rect 913 17 971 115
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel locali s 927 221 961 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel locali s 587 51 671 145 0 FreeSans 400 0 0 0 Y
port 8 nsew signal output
flabel locali s 132 221 166 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 247 215 440 257 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor3b_2
rlabel locali s 574 181 671 409 1 Y
port 8 nsew signal output
rlabel locali s 295 51 371 145 1 Y
port 8 nsew signal output
rlabel locali s 107 145 671 181 1 Y
port 8 nsew signal output
rlabel locali s 107 51 183 145 1 Y
port 8 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 84682
string GDS_START 76882
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
