magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3122 1975
<< nwell >>
rect -38 331 1862 704
rect 1174 309 1382 331
<< pwell >>
rect 751 249 936 273
rect 751 229 942 249
rect 1139 229 1820 241
rect 214 180 1820 229
rect 1 49 1820 180
rect 0 0 1824 49
<< scnmos >>
rect 80 70 110 154
rect 293 119 323 203
rect 401 119 431 203
rect 507 119 537 203
rect 612 119 642 203
rect 684 119 714 203
rect 830 119 860 247
rect 939 119 969 203
rect 1040 119 1070 203
rect 1112 119 1142 203
rect 1230 47 1260 215
rect 1453 47 1483 215
rect 1539 47 1569 215
rect 1625 47 1655 215
rect 1711 47 1741 215
<< scpmoshvt >>
rect 80 468 110 596
rect 270 413 300 541
rect 410 413 440 497
rect 496 413 526 497
rect 636 413 666 497
rect 708 413 738 497
rect 825 379 855 547
rect 911 379 941 547
rect 1086 441 1116 525
rect 1158 441 1188 525
rect 1263 345 1293 597
rect 1453 367 1483 619
rect 1539 367 1569 619
rect 1625 367 1655 619
rect 1711 367 1741 619
<< ndiff >>
rect 777 203 830 247
rect 240 178 293 203
rect 27 118 80 154
rect 27 84 35 118
rect 69 84 80 118
rect 27 70 80 84
rect 110 129 163 154
rect 110 95 121 129
rect 155 95 163 129
rect 240 144 248 178
rect 282 144 293 178
rect 240 119 293 144
rect 323 178 401 203
rect 323 144 346 178
rect 380 144 401 178
rect 323 119 401 144
rect 431 175 507 203
rect 431 141 460 175
rect 494 141 507 175
rect 431 119 507 141
rect 537 178 612 203
rect 537 144 560 178
rect 594 144 612 178
rect 537 119 612 144
rect 642 119 684 203
rect 714 176 830 203
rect 714 142 757 176
rect 791 142 830 176
rect 714 119 830 142
rect 860 223 910 247
rect 860 203 916 223
rect 1165 203 1230 215
rect 860 171 939 203
rect 860 137 874 171
rect 908 137 939 171
rect 860 119 939 137
rect 969 178 1040 203
rect 969 144 995 178
rect 1029 144 1040 178
rect 969 119 1040 144
rect 1070 119 1112 203
rect 1142 169 1230 203
rect 1142 135 1173 169
rect 1207 135 1230 169
rect 1142 119 1230 135
rect 110 70 163 95
rect 1165 93 1230 119
rect 1165 59 1173 93
rect 1207 59 1230 93
rect 1165 47 1230 59
rect 1260 169 1317 215
rect 1260 135 1275 169
rect 1309 135 1317 169
rect 1260 95 1317 135
rect 1260 61 1275 95
rect 1309 61 1317 95
rect 1260 47 1317 61
rect 1400 203 1453 215
rect 1400 169 1408 203
rect 1442 169 1453 203
rect 1400 93 1453 169
rect 1400 59 1408 93
rect 1442 59 1453 93
rect 1400 47 1453 59
rect 1483 207 1539 215
rect 1483 173 1494 207
rect 1528 173 1539 207
rect 1483 101 1539 173
rect 1483 67 1494 101
rect 1528 67 1539 101
rect 1483 47 1539 67
rect 1569 177 1625 215
rect 1569 143 1580 177
rect 1614 143 1625 177
rect 1569 89 1625 143
rect 1569 55 1580 89
rect 1614 55 1625 89
rect 1569 47 1625 55
rect 1655 207 1711 215
rect 1655 173 1666 207
rect 1700 173 1711 207
rect 1655 101 1711 173
rect 1655 67 1666 101
rect 1700 67 1711 101
rect 1655 47 1711 67
rect 1741 125 1794 215
rect 1741 91 1752 125
rect 1786 91 1794 125
rect 1741 47 1794 91
<< pdiff >>
rect 27 583 80 596
rect 27 549 35 583
rect 69 549 80 583
rect 27 468 80 549
rect 110 582 163 596
rect 110 548 121 582
rect 155 548 163 582
rect 110 514 163 548
rect 110 480 121 514
rect 155 480 163 514
rect 110 468 163 480
rect 217 527 270 541
rect 217 493 225 527
rect 259 493 270 527
rect 217 459 270 493
rect 217 425 225 459
rect 259 425 270 459
rect 217 413 270 425
rect 300 529 353 541
rect 300 495 311 529
rect 345 497 353 529
rect 760 561 810 573
rect 760 527 768 561
rect 802 547 810 561
rect 1400 607 1453 619
rect 1210 585 1263 597
rect 1210 551 1218 585
rect 1252 551 1263 585
rect 802 527 825 547
rect 760 497 825 527
rect 345 495 410 497
rect 300 413 410 495
rect 440 455 496 497
rect 440 421 451 455
rect 485 421 496 455
rect 440 413 496 421
rect 526 455 636 497
rect 526 421 589 455
rect 623 421 636 455
rect 526 413 636 421
rect 666 413 708 497
rect 738 413 825 497
rect 760 379 825 413
rect 855 421 911 547
rect 855 387 866 421
rect 900 387 911 421
rect 855 379 911 387
rect 941 525 1064 547
rect 1210 525 1263 551
rect 941 524 1086 525
rect 941 490 1022 524
rect 1056 490 1086 524
rect 941 456 1086 490
rect 941 422 1022 456
rect 1056 441 1086 456
rect 1116 441 1158 525
rect 1188 517 1263 525
rect 1188 483 1218 517
rect 1252 483 1263 517
rect 1188 449 1263 483
rect 1188 441 1218 449
rect 1056 422 1064 441
rect 941 410 1064 422
rect 941 379 991 410
rect 1210 415 1218 441
rect 1252 415 1263 449
rect 1210 345 1263 415
rect 1293 585 1346 597
rect 1293 551 1304 585
rect 1338 551 1346 585
rect 1293 494 1346 551
rect 1293 460 1304 494
rect 1338 460 1346 494
rect 1293 391 1346 460
rect 1293 357 1304 391
rect 1338 357 1346 391
rect 1400 573 1408 607
rect 1442 573 1453 607
rect 1400 508 1453 573
rect 1400 474 1408 508
rect 1442 474 1453 508
rect 1400 413 1453 474
rect 1400 379 1408 413
rect 1442 379 1453 413
rect 1400 367 1453 379
rect 1483 599 1539 619
rect 1483 565 1494 599
rect 1528 565 1539 599
rect 1483 508 1539 565
rect 1483 474 1494 508
rect 1528 474 1539 508
rect 1483 409 1539 474
rect 1483 375 1494 409
rect 1528 375 1539 409
rect 1483 367 1539 375
rect 1569 611 1625 619
rect 1569 577 1580 611
rect 1614 577 1625 611
rect 1569 533 1625 577
rect 1569 499 1580 533
rect 1614 499 1625 533
rect 1569 449 1625 499
rect 1569 415 1580 449
rect 1614 415 1625 449
rect 1569 367 1625 415
rect 1655 599 1711 619
rect 1655 565 1666 599
rect 1700 565 1711 599
rect 1655 508 1711 565
rect 1655 474 1666 508
rect 1700 474 1711 508
rect 1655 409 1711 474
rect 1655 375 1666 409
rect 1700 375 1711 409
rect 1655 367 1711 375
rect 1741 576 1794 619
rect 1741 542 1752 576
rect 1786 542 1794 576
rect 1741 367 1794 542
rect 1293 345 1346 357
<< ndiffc >>
rect 35 84 69 118
rect 121 95 155 129
rect 248 144 282 178
rect 346 144 380 178
rect 460 141 494 175
rect 560 144 594 178
rect 757 142 791 176
rect 874 137 908 171
rect 995 144 1029 178
rect 1173 135 1207 169
rect 1173 59 1207 93
rect 1275 135 1309 169
rect 1275 61 1309 95
rect 1408 169 1442 203
rect 1408 59 1442 93
rect 1494 173 1528 207
rect 1494 67 1528 101
rect 1580 143 1614 177
rect 1580 55 1614 89
rect 1666 173 1700 207
rect 1666 67 1700 101
rect 1752 91 1786 125
<< pdiffc >>
rect 35 549 69 583
rect 121 548 155 582
rect 121 480 155 514
rect 225 493 259 527
rect 225 425 259 459
rect 311 495 345 529
rect 768 527 802 561
rect 1218 551 1252 585
rect 451 421 485 455
rect 589 421 623 455
rect 866 387 900 421
rect 1022 490 1056 524
rect 1022 422 1056 456
rect 1218 483 1252 517
rect 1218 415 1252 449
rect 1304 551 1338 585
rect 1304 460 1338 494
rect 1304 357 1338 391
rect 1408 573 1442 607
rect 1408 474 1442 508
rect 1408 379 1442 413
rect 1494 565 1528 599
rect 1494 474 1528 508
rect 1494 375 1528 409
rect 1580 577 1614 611
rect 1580 499 1614 533
rect 1580 415 1614 449
rect 1666 565 1700 599
rect 1666 474 1700 508
rect 1666 375 1700 409
rect 1752 542 1786 576
<< poly >>
rect 80 596 110 622
rect 270 615 941 645
rect 270 541 300 615
rect 80 310 110 468
rect 410 497 440 523
rect 496 497 526 523
rect 636 497 666 615
rect 825 547 855 573
rect 911 547 941 615
rect 1263 597 1293 623
rect 1453 619 1483 645
rect 1539 619 1569 645
rect 1625 619 1655 645
rect 1711 619 1741 645
rect 708 497 738 523
rect 31 294 110 310
rect 31 260 47 294
rect 81 260 110 294
rect 31 226 110 260
rect 156 357 222 373
rect 156 323 172 357
rect 206 323 222 357
rect 156 289 222 323
rect 156 255 172 289
rect 206 269 222 289
rect 270 269 300 413
rect 410 359 440 413
rect 365 343 440 359
rect 365 309 381 343
rect 415 309 440 343
rect 496 375 526 413
rect 636 387 666 413
rect 496 359 571 375
rect 496 325 521 359
rect 555 339 571 359
rect 708 339 738 413
rect 1086 525 1116 551
rect 1158 525 1188 551
rect 1086 395 1116 441
rect 555 325 642 339
rect 496 309 642 325
rect 365 307 440 309
rect 365 275 431 307
rect 206 255 323 269
rect 156 239 323 255
rect 31 192 47 226
rect 81 192 110 226
rect 293 203 323 239
rect 365 241 381 275
rect 415 241 431 275
rect 365 225 431 241
rect 401 203 431 225
rect 507 203 537 229
rect 612 203 642 309
rect 684 323 750 339
rect 825 335 855 379
rect 911 353 941 379
rect 1006 365 1116 395
rect 684 289 700 323
rect 734 289 750 323
rect 684 273 750 289
rect 792 319 860 335
rect 792 285 808 319
rect 842 285 860 319
rect 1006 311 1036 365
rect 1158 323 1188 441
rect 684 203 714 273
rect 792 269 860 285
rect 830 247 860 269
rect 932 295 1036 311
rect 932 261 948 295
rect 982 281 1036 295
rect 1112 307 1188 323
rect 982 261 998 281
rect 31 176 110 192
rect 80 154 110 176
rect 932 245 998 261
rect 1112 273 1128 307
rect 1162 273 1188 307
rect 1263 303 1293 345
rect 1453 329 1483 367
rect 1539 329 1569 367
rect 1625 329 1655 367
rect 1711 329 1741 367
rect 1385 313 1741 329
rect 1112 257 1188 273
rect 1230 287 1296 303
rect 939 203 969 245
rect 1040 203 1070 229
rect 1112 203 1142 257
rect 1230 253 1246 287
rect 1280 253 1296 287
rect 1385 279 1401 313
rect 1435 279 1469 313
rect 1503 279 1537 313
rect 1571 279 1605 313
rect 1639 279 1673 313
rect 1707 279 1741 313
rect 1385 263 1741 279
rect 1230 237 1296 253
rect 1230 215 1260 237
rect 1453 215 1483 263
rect 1539 215 1569 263
rect 1625 215 1655 263
rect 1711 215 1741 263
rect 80 44 110 70
rect 293 51 323 119
rect 401 93 431 119
rect 507 51 537 119
rect 612 93 642 119
rect 684 93 714 119
rect 830 93 860 119
rect 939 93 969 119
rect 1040 51 1070 119
rect 1112 93 1142 119
rect 293 21 1070 51
rect 1230 21 1260 47
rect 1453 21 1483 47
rect 1539 21 1569 47
rect 1625 21 1655 47
rect 1711 21 1741 47
<< polycont >>
rect 47 260 81 294
rect 172 323 206 357
rect 172 255 206 289
rect 381 309 415 343
rect 521 325 555 359
rect 47 192 81 226
rect 381 241 415 275
rect 700 289 734 323
rect 808 285 842 319
rect 948 261 982 295
rect 1128 273 1162 307
rect 1246 253 1280 287
rect 1401 279 1435 313
rect 1469 279 1503 313
rect 1537 279 1571 313
rect 1605 279 1639 313
rect 1673 279 1707 313
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 19 583 85 649
rect 19 549 35 583
rect 69 549 85 583
rect 19 533 85 549
rect 119 582 171 598
rect 119 548 121 582
rect 155 548 171 582
rect 119 514 171 548
rect 17 294 85 498
rect 17 260 47 294
rect 81 260 85 294
rect 17 226 85 260
rect 17 192 47 226
rect 81 192 85 226
rect 17 168 85 192
rect 119 480 121 514
rect 155 480 171 514
rect 119 373 171 480
rect 209 527 263 543
rect 209 493 225 527
rect 259 493 263 527
rect 209 459 263 493
rect 307 529 345 649
rect 752 561 818 649
rect 307 495 311 529
rect 307 479 345 495
rect 381 507 699 541
rect 752 527 768 561
rect 802 527 818 561
rect 1202 585 1268 649
rect 1392 607 1451 649
rect 1202 551 1218 585
rect 1252 551 1268 585
rect 752 525 818 527
rect 209 425 225 459
rect 259 443 263 459
rect 381 443 415 507
rect 259 425 415 443
rect 209 409 415 425
rect 449 455 485 471
rect 449 421 451 455
rect 119 357 206 373
rect 119 323 172 357
rect 119 289 206 323
rect 119 255 172 289
rect 119 239 206 255
rect 19 118 85 134
rect 19 84 35 118
rect 69 84 85 118
rect 19 17 85 84
rect 119 129 171 239
rect 119 95 121 129
rect 155 95 171 129
rect 240 192 282 409
rect 449 386 485 421
rect 316 343 415 359
rect 316 309 381 343
rect 316 275 415 309
rect 316 241 381 275
rect 316 225 415 241
rect 240 178 296 192
rect 449 191 483 386
rect 519 359 555 507
rect 665 491 699 507
rect 1022 524 1072 540
rect 519 325 521 359
rect 519 309 555 325
rect 589 455 629 471
rect 665 457 986 491
rect 623 421 629 455
rect 589 270 629 421
rect 684 421 916 423
rect 684 387 866 421
rect 900 387 916 421
rect 684 383 916 387
rect 684 371 912 383
rect 684 323 750 371
rect 684 289 700 323
rect 734 289 750 323
rect 792 319 844 335
rect 544 255 629 270
rect 792 285 808 319
rect 842 285 844 319
rect 792 255 844 285
rect 544 221 844 255
rect 240 144 248 178
rect 282 144 296 178
rect 240 128 296 144
rect 330 178 396 191
rect 330 144 346 178
rect 380 144 396 178
rect 119 79 171 95
rect 330 17 396 144
rect 444 175 510 191
rect 444 141 460 175
rect 494 141 510 175
rect 444 125 510 141
rect 544 178 610 221
rect 878 187 912 371
rect 952 311 986 457
rect 946 295 986 311
rect 946 261 948 295
rect 982 261 986 295
rect 946 245 986 261
rect 1056 490 1072 524
rect 1022 456 1072 490
rect 1056 422 1072 456
rect 1022 237 1072 422
rect 1202 517 1268 551
rect 1202 483 1218 517
rect 1252 483 1268 517
rect 1202 449 1268 483
rect 1202 415 1218 449
rect 1252 415 1268 449
rect 1202 407 1268 415
rect 1302 585 1350 601
rect 1302 551 1304 585
rect 1338 551 1350 585
rect 1302 494 1350 551
rect 1302 460 1304 494
rect 1338 460 1350 494
rect 1302 391 1350 460
rect 1302 373 1304 391
rect 1112 357 1304 373
rect 1338 357 1350 391
rect 1392 573 1408 607
rect 1442 573 1451 607
rect 1392 508 1451 573
rect 1392 474 1408 508
rect 1442 474 1451 508
rect 1392 413 1451 474
rect 1392 379 1408 413
rect 1442 379 1451 413
rect 1392 363 1451 379
rect 1485 599 1530 615
rect 1485 565 1494 599
rect 1528 565 1530 599
rect 1485 508 1530 565
rect 1485 474 1494 508
rect 1528 474 1530 508
rect 1485 409 1530 474
rect 1564 611 1630 649
rect 1564 577 1580 611
rect 1614 577 1630 611
rect 1564 533 1630 577
rect 1564 499 1580 533
rect 1614 499 1630 533
rect 1564 449 1630 499
rect 1564 415 1580 449
rect 1614 415 1630 449
rect 1664 599 1702 615
rect 1664 565 1666 599
rect 1700 565 1702 599
rect 1664 508 1702 565
rect 1736 576 1802 649
rect 1736 542 1752 576
rect 1786 542 1802 576
rect 1736 532 1802 542
rect 1664 474 1666 508
rect 1700 474 1702 508
rect 1485 375 1494 409
rect 1528 381 1530 409
rect 1664 409 1702 474
rect 1664 381 1666 409
rect 1528 375 1666 381
rect 1700 389 1702 409
rect 1759 389 1807 498
rect 1700 375 1807 389
rect 1112 339 1350 357
rect 1485 347 1807 375
rect 1112 307 1178 339
rect 1112 273 1128 307
rect 1162 273 1178 307
rect 1316 313 1350 339
rect 1112 271 1178 273
rect 1230 287 1282 303
rect 1230 253 1246 287
rect 1280 253 1282 287
rect 1230 237 1282 253
rect 1022 203 1282 237
rect 1316 279 1401 313
rect 1435 279 1469 313
rect 1503 279 1537 313
rect 1571 279 1605 313
rect 1639 279 1673 313
rect 1707 279 1723 313
rect 1022 199 1056 203
rect 544 144 560 178
rect 594 144 610 178
rect 544 128 610 144
rect 741 176 807 187
rect 741 142 757 176
rect 791 142 807 176
rect 741 17 807 142
rect 858 171 912 187
rect 858 137 874 171
rect 908 137 912 171
rect 858 117 912 137
rect 979 178 1056 199
rect 979 144 995 178
rect 1029 144 1056 178
rect 1316 169 1350 279
rect 1759 245 1807 347
rect 979 128 1056 144
rect 1157 135 1173 169
rect 1207 135 1223 169
rect 1157 93 1223 135
rect 1157 59 1173 93
rect 1207 59 1223 93
rect 1157 17 1223 59
rect 1259 135 1275 169
rect 1309 135 1350 169
rect 1259 95 1350 135
rect 1259 61 1275 95
rect 1309 61 1350 95
rect 1259 57 1350 61
rect 1392 203 1450 219
rect 1392 169 1408 203
rect 1442 169 1450 203
rect 1392 93 1450 169
rect 1392 59 1408 93
rect 1442 59 1450 93
rect 1392 17 1450 59
rect 1484 211 1807 245
rect 1484 207 1530 211
rect 1484 173 1494 207
rect 1528 173 1530 207
rect 1664 207 1807 211
rect 1484 101 1530 173
rect 1484 67 1494 101
rect 1528 67 1530 101
rect 1484 51 1530 67
rect 1564 143 1580 177
rect 1614 143 1630 177
rect 1564 89 1630 143
rect 1564 55 1580 89
rect 1614 55 1630 89
rect 1564 17 1630 55
rect 1664 173 1666 207
rect 1700 173 1807 207
rect 1664 168 1807 173
rect 1664 101 1702 168
rect 1664 67 1666 101
rect 1700 67 1702 101
rect 1664 51 1702 67
rect 1736 125 1802 134
rect 1736 91 1752 125
rect 1786 91 1802 125
rect 1736 17 1802 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfxtp_4
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1759 168 1793 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1759 316 1793 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1759 390 1793 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1759 464 1793 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 989790
string GDS_START 975630
<< end >>
