magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4082 1975
<< nwell >>
rect -38 331 2822 704
<< pwell >>
rect 2107 251 2476 288
rect 673 223 1049 249
rect 1598 223 1882 235
rect 673 157 1882 223
rect 11 49 1882 157
rect 2107 49 2783 251
rect 0 0 2784 49
<< scnmos >>
rect 756 139 786 223
rect 842 139 872 223
rect 920 139 950 223
rect 94 47 124 131
rect 180 47 210 131
rect 258 47 288 131
rect 366 47 396 131
rect 444 47 474 131
rect 540 47 570 131
rect 1081 69 1111 197
rect 1217 69 1247 197
rect 1289 69 1319 197
rect 1421 113 1451 197
rect 1493 113 1523 197
rect 1565 113 1595 197
rect 1674 125 1704 209
rect 1746 125 1776 209
rect 2213 178 2243 262
rect 2291 178 2321 262
rect 2363 178 2393 262
rect 2561 57 2591 141
rect 2670 57 2700 225
<< scpmoshvt >>
rect 88 477 118 605
rect 174 477 204 605
rect 252 477 282 605
rect 338 477 368 605
rect 432 477 462 605
rect 600 477 630 605
rect 894 530 924 614
rect 980 530 1010 614
rect 1058 530 1088 614
rect 1240 425 1270 593
rect 1342 379 1372 547
rect 1414 379 1444 547
rect 1808 419 1858 619
rect 1906 419 1956 619
rect 2035 419 2065 547
rect 2175 419 2205 547
rect 2284 419 2334 619
rect 2561 367 2591 495
rect 2670 367 2700 619
<< ndiff >>
rect 699 206 756 223
rect 699 172 711 206
rect 745 172 756 206
rect 699 139 756 172
rect 786 198 842 223
rect 786 164 797 198
rect 831 164 842 198
rect 786 139 842 164
rect 872 139 920 223
rect 950 197 1023 223
rect 1624 197 1674 209
rect 950 139 1081 197
rect 37 110 94 131
rect 37 76 49 110
rect 83 76 94 110
rect 37 47 94 76
rect 124 105 180 131
rect 124 71 135 105
rect 169 71 180 105
rect 124 47 180 71
rect 210 47 258 131
rect 288 109 366 131
rect 288 75 321 109
rect 355 75 366 109
rect 288 47 366 75
rect 396 47 444 131
rect 474 105 540 131
rect 474 71 495 105
rect 529 71 540 105
rect 474 47 540 71
rect 570 110 626 131
rect 570 76 581 110
rect 615 76 626 110
rect 570 47 626 76
rect 965 73 1081 139
rect 965 39 977 73
rect 1011 69 1081 73
rect 1111 177 1217 197
rect 1111 143 1122 177
rect 1156 143 1217 177
rect 1111 69 1217 143
rect 1247 69 1289 197
rect 1319 169 1421 197
rect 1319 135 1376 169
rect 1410 135 1421 169
rect 1319 113 1421 135
rect 1451 113 1493 197
rect 1523 113 1565 197
rect 1595 163 1674 197
rect 1595 129 1606 163
rect 1640 129 1674 163
rect 1595 125 1674 129
rect 1704 125 1746 209
rect 1776 167 1856 209
rect 1776 133 1810 167
rect 1844 133 1856 167
rect 1776 125 1856 133
rect 1595 113 1652 125
rect 1319 69 1406 113
rect 1011 39 1023 69
rect 1798 121 1856 125
rect 2133 243 2213 262
rect 2133 209 2145 243
rect 2179 209 2213 243
rect 2133 178 2213 209
rect 2243 178 2291 262
rect 2321 178 2363 262
rect 2393 237 2450 262
rect 2393 203 2404 237
rect 2438 203 2450 237
rect 2393 178 2450 203
rect 965 27 1023 39
rect 2613 213 2670 225
rect 2613 179 2625 213
rect 2659 179 2670 213
rect 2613 141 2670 179
rect 2504 116 2561 141
rect 2504 82 2516 116
rect 2550 82 2561 116
rect 2504 57 2561 82
rect 2591 103 2670 141
rect 2591 69 2625 103
rect 2659 69 2670 103
rect 2591 57 2670 69
rect 2700 213 2757 225
rect 2700 179 2711 213
rect 2745 179 2757 213
rect 2700 103 2757 179
rect 2700 69 2711 103
rect 2745 69 2757 103
rect 2700 57 2757 69
<< pdiff >>
rect 1103 627 1190 639
rect 1103 614 1115 627
rect 31 593 88 605
rect 31 559 43 593
rect 77 559 88 593
rect 31 523 88 559
rect 31 489 43 523
rect 77 489 88 523
rect 31 477 88 489
rect 118 593 174 605
rect 118 559 129 593
rect 163 559 174 593
rect 118 523 174 559
rect 118 489 129 523
rect 163 489 174 523
rect 118 477 174 489
rect 204 477 252 605
rect 282 593 338 605
rect 282 559 293 593
rect 327 559 338 593
rect 282 523 338 559
rect 282 489 293 523
rect 327 489 338 523
rect 282 477 338 489
rect 368 477 432 605
rect 462 587 600 605
rect 462 553 496 587
rect 530 553 600 587
rect 462 477 600 553
rect 630 531 687 605
rect 823 587 894 614
rect 823 553 835 587
rect 869 553 894 587
rect 630 497 641 531
rect 675 497 687 531
rect 630 477 687 497
rect 823 530 894 553
rect 924 587 980 614
rect 924 553 935 587
rect 969 553 980 587
rect 924 530 980 553
rect 1010 530 1058 614
rect 1088 593 1115 614
rect 1149 593 1190 627
rect 1088 530 1240 593
rect 1190 425 1240 530
rect 1270 547 1320 593
rect 1751 599 1808 619
rect 1751 565 1763 599
rect 1797 565 1808 599
rect 1270 501 1342 547
rect 1270 467 1283 501
rect 1317 467 1342 501
rect 1270 425 1342 467
rect 1292 379 1342 425
rect 1372 379 1414 547
rect 1444 531 1501 547
rect 1444 497 1455 531
rect 1489 497 1501 531
rect 1444 425 1501 497
rect 1444 391 1455 425
rect 1489 391 1501 425
rect 1751 503 1808 565
rect 1751 469 1763 503
rect 1797 469 1808 503
rect 1751 419 1808 469
rect 1858 419 1906 619
rect 1956 592 2013 619
rect 1956 558 1967 592
rect 2001 558 2013 592
rect 2227 592 2284 619
rect 1956 547 2013 558
rect 2227 558 2239 592
rect 2273 558 2284 592
rect 2227 547 2284 558
rect 1956 419 2035 547
rect 2065 498 2175 547
rect 2065 464 2103 498
rect 2137 464 2175 498
rect 2065 419 2175 464
rect 2205 419 2284 547
rect 2334 482 2421 619
rect 2334 448 2375 482
rect 2409 448 2421 482
rect 2334 419 2421 448
rect 2613 607 2670 619
rect 2613 573 2625 607
rect 2659 573 2670 607
rect 1444 379 1501 391
rect 2613 510 2670 573
rect 2613 495 2625 510
rect 2504 483 2561 495
rect 2504 449 2516 483
rect 2550 449 2561 483
rect 2504 413 2561 449
rect 2504 379 2516 413
rect 2550 379 2561 413
rect 2504 367 2561 379
rect 2591 476 2625 495
rect 2659 476 2670 510
rect 2591 413 2670 476
rect 2591 379 2625 413
rect 2659 379 2670 413
rect 2591 367 2670 379
rect 2700 599 2757 619
rect 2700 565 2711 599
rect 2745 565 2757 599
rect 2700 506 2757 565
rect 2700 472 2711 506
rect 2745 472 2757 506
rect 2700 413 2757 472
rect 2700 379 2711 413
rect 2745 379 2757 413
rect 2700 367 2757 379
<< ndiffc >>
rect 711 172 745 206
rect 797 164 831 198
rect 49 76 83 110
rect 135 71 169 105
rect 321 75 355 109
rect 495 71 529 105
rect 581 76 615 110
rect 977 39 1011 73
rect 1122 143 1156 177
rect 1376 135 1410 169
rect 1606 129 1640 163
rect 1810 133 1844 167
rect 2145 209 2179 243
rect 2404 203 2438 237
rect 2625 179 2659 213
rect 2516 82 2550 116
rect 2625 69 2659 103
rect 2711 179 2745 213
rect 2711 69 2745 103
<< pdiffc >>
rect 43 559 77 593
rect 43 489 77 523
rect 129 559 163 593
rect 129 489 163 523
rect 293 559 327 593
rect 293 489 327 523
rect 496 553 530 587
rect 835 553 869 587
rect 641 497 675 531
rect 935 553 969 587
rect 1115 593 1149 627
rect 1763 565 1797 599
rect 1283 467 1317 501
rect 1455 497 1489 531
rect 1455 391 1489 425
rect 1763 469 1797 503
rect 1967 558 2001 592
rect 2239 558 2273 592
rect 2103 464 2137 498
rect 2375 448 2409 482
rect 2625 573 2659 607
rect 2516 449 2550 483
rect 2516 379 2550 413
rect 2625 476 2659 510
rect 2625 379 2659 413
rect 2711 565 2745 599
rect 2711 472 2745 506
rect 2711 379 2745 413
<< poly >>
rect 88 605 118 631
rect 174 605 204 631
rect 252 605 282 631
rect 338 605 368 631
rect 432 605 462 631
rect 600 605 630 631
rect 894 614 924 640
rect 980 614 1010 640
rect 1058 614 1088 640
rect 719 531 785 547
rect 719 497 735 531
rect 769 508 785 531
rect 1240 615 1668 645
rect 1808 619 1858 645
rect 1906 619 1956 645
rect 2284 619 2334 645
rect 2670 619 2700 645
rect 1240 593 1270 615
rect 1602 599 1668 615
rect 894 508 924 530
rect 769 497 924 508
rect 719 478 924 497
rect 88 455 118 477
rect 174 455 204 477
rect 39 425 204 455
rect 39 263 69 425
rect 117 361 210 377
rect 117 327 133 361
rect 167 327 210 361
rect 117 311 210 327
rect 39 247 138 263
rect 39 213 88 247
rect 122 213 138 247
rect 39 197 138 213
rect 94 131 124 197
rect 180 131 210 311
rect 252 302 282 477
rect 338 416 368 477
rect 432 416 462 477
rect 324 400 390 416
rect 324 366 340 400
rect 374 366 390 400
rect 324 350 390 366
rect 432 400 498 416
rect 432 366 448 400
rect 482 366 498 400
rect 600 383 630 477
rect 980 390 1010 530
rect 1058 498 1088 530
rect 1058 482 1124 498
rect 1058 448 1074 482
rect 1108 448 1124 482
rect 1058 432 1124 448
rect 1342 547 1372 573
rect 1414 547 1444 573
rect 1602 565 1618 599
rect 1652 565 1668 599
rect 1602 549 1668 565
rect 1240 399 1270 425
rect 756 383 1189 390
rect 432 350 498 366
rect 252 286 318 302
rect 252 252 268 286
rect 302 252 318 286
rect 252 236 318 252
rect 360 286 426 302
rect 360 252 376 286
rect 410 252 426 286
rect 360 236 426 252
rect 258 131 288 236
rect 366 131 396 236
rect 468 194 498 350
rect 580 360 1189 383
rect 2035 547 2065 573
rect 2175 547 2205 573
rect 2453 599 2519 615
rect 2453 565 2469 599
rect 2503 565 2519 599
rect 2453 549 2519 565
rect 1602 403 1668 419
rect 580 353 786 360
rect 580 195 610 353
rect 756 223 786 353
rect 1159 357 1189 360
rect 1342 357 1372 379
rect 1414 357 1444 379
rect 1602 369 1618 403
rect 1652 369 1668 403
rect 1808 393 1858 419
rect 1906 393 1956 419
rect 1602 357 1668 369
rect 1159 327 1668 357
rect 1710 335 1776 351
rect 914 295 980 311
rect 914 261 930 295
rect 964 261 980 295
rect 842 223 872 249
rect 914 245 980 261
rect 1022 302 1111 318
rect 1022 268 1038 302
rect 1072 268 1111 302
rect 1022 252 1111 268
rect 920 223 950 245
rect 444 164 498 194
rect 540 165 610 195
rect 444 131 474 164
rect 540 131 570 165
rect 1081 197 1111 252
rect 1190 269 1328 285
rect 1190 235 1206 269
rect 1240 235 1274 269
rect 1308 235 1328 269
rect 1190 219 1328 235
rect 1217 197 1247 219
rect 1289 197 1319 219
rect 1421 197 1451 327
rect 1710 301 1726 335
rect 1760 301 1776 335
rect 1710 279 1776 301
rect 1818 345 1848 393
rect 1818 329 1884 345
rect 1818 295 1834 329
rect 1868 295 1884 329
rect 1818 279 1884 295
rect 1674 249 1776 279
rect 1493 197 1523 223
rect 1565 197 1595 223
rect 1674 209 1704 249
rect 1746 209 1776 249
rect 1926 224 1956 393
rect 648 101 714 117
rect 756 113 786 139
rect 648 67 664 101
rect 698 67 714 101
rect 648 65 714 67
rect 842 65 872 139
rect 920 113 950 139
rect 94 21 124 47
rect 180 21 210 47
rect 258 21 288 47
rect 366 21 396 47
rect 444 21 474 47
rect 540 21 570 47
rect 648 35 872 65
rect 1918 208 1984 224
rect 1918 188 1934 208
rect 1421 87 1451 113
rect 1081 43 1111 69
rect 1217 43 1247 69
rect 1289 43 1319 69
rect 1493 51 1523 113
rect 1565 51 1595 113
rect 1674 99 1704 125
rect 1746 99 1776 125
rect 1871 174 1934 188
rect 1968 174 1984 208
rect 1871 158 1984 174
rect 1871 51 1901 158
rect 2035 116 2065 419
rect 2175 366 2205 419
rect 2284 397 2334 419
rect 2453 397 2483 549
rect 2561 495 2591 521
rect 2284 367 2483 397
rect 2136 350 2205 366
rect 2136 316 2152 350
rect 2186 319 2205 350
rect 2453 345 2483 367
rect 2561 345 2591 367
rect 2186 316 2243 319
rect 2136 289 2243 316
rect 2213 262 2243 289
rect 2291 262 2321 288
rect 2363 262 2393 319
rect 2453 315 2591 345
rect 2670 329 2700 367
rect 2555 215 2585 315
rect 2633 313 2700 329
rect 2633 279 2649 313
rect 2683 279 2700 313
rect 2633 263 2700 279
rect 2670 225 2700 263
rect 2555 185 2591 215
rect 2213 152 2243 178
rect 1493 21 1901 51
rect 1961 100 2065 116
rect 1961 66 1977 100
rect 2011 66 2065 100
rect 1961 50 2065 66
rect 2291 130 2321 178
rect 2363 130 2393 178
rect 2561 141 2591 185
rect 2291 114 2393 130
rect 2291 80 2320 114
rect 2354 80 2393 114
rect 2291 64 2393 80
rect 2561 31 2591 57
rect 2670 31 2700 57
<< polycont >>
rect 735 497 769 531
rect 133 327 167 361
rect 88 213 122 247
rect 340 366 374 400
rect 448 366 482 400
rect 1074 448 1108 482
rect 1618 565 1652 599
rect 268 252 302 286
rect 376 252 410 286
rect 2469 565 2503 599
rect 1618 369 1652 403
rect 930 261 964 295
rect 1038 268 1072 302
rect 1206 235 1240 269
rect 1274 235 1308 269
rect 1726 301 1760 335
rect 1834 295 1868 329
rect 664 67 698 101
rect 1934 174 1968 208
rect 2152 316 2186 350
rect 2649 279 2683 313
rect 1977 66 2011 100
rect 2320 80 2354 114
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 17 593 77 609
rect 17 559 43 593
rect 17 523 77 559
rect 17 489 43 523
rect 17 416 77 489
rect 113 593 179 649
rect 113 559 129 593
rect 163 559 179 593
rect 113 523 179 559
rect 113 489 129 523
rect 163 489 179 523
rect 113 473 179 489
rect 277 593 343 609
rect 277 559 293 593
rect 327 559 343 593
rect 277 523 343 559
rect 480 587 530 649
rect 1099 627 1165 649
rect 480 553 496 587
rect 480 532 530 553
rect 564 587 885 615
rect 564 581 835 587
rect 277 489 293 523
rect 327 498 343 523
rect 564 498 598 581
rect 819 553 835 581
rect 869 553 885 587
rect 327 489 598 498
rect 277 464 598 489
rect 641 531 785 547
rect 675 497 735 531
rect 769 497 785 531
rect 641 481 785 497
rect 17 400 381 416
rect 17 382 340 400
rect 17 135 51 382
rect 117 366 340 382
rect 374 366 381 400
rect 117 361 381 366
rect 117 327 133 361
rect 167 350 381 361
rect 415 400 498 430
rect 415 366 448 400
rect 482 366 498 400
rect 415 350 498 366
rect 167 327 183 350
rect 117 311 183 327
rect 217 286 318 302
rect 85 247 151 263
rect 85 213 88 247
rect 122 213 151 247
rect 217 252 268 286
rect 302 252 318 286
rect 217 236 318 252
rect 359 286 455 302
rect 359 252 376 286
rect 410 252 455 286
rect 359 236 455 252
rect 532 236 566 464
rect 641 430 691 481
rect 819 447 885 553
rect 85 202 151 213
rect 359 202 393 236
rect 497 202 566 236
rect 600 396 691 430
rect 727 413 885 447
rect 919 587 985 615
rect 1099 593 1115 627
rect 1149 593 1165 627
rect 1199 599 1668 615
rect 919 553 935 587
rect 969 559 985 587
rect 1199 581 1618 599
rect 1199 559 1233 581
rect 969 553 1233 559
rect 919 525 1233 553
rect 1602 565 1618 581
rect 1652 565 1668 599
rect 1602 549 1668 565
rect 1747 599 1813 615
rect 1747 565 1763 599
rect 1797 565 1813 599
rect 85 197 393 202
rect 117 168 393 197
rect 427 168 531 202
rect 17 110 83 135
rect 427 134 461 168
rect 600 135 634 396
rect 727 227 761 413
rect 919 379 985 525
rect 1267 501 1333 547
rect 1267 491 1283 501
rect 1058 482 1283 491
rect 1058 448 1074 482
rect 1108 467 1283 482
rect 1317 467 1333 501
rect 1108 448 1333 467
rect 1058 421 1333 448
rect 1439 531 1505 547
rect 1439 497 1455 531
rect 1489 497 1505 531
rect 1439 487 1505 497
rect 1747 503 1813 565
rect 1945 592 2001 615
rect 1945 581 1967 592
rect 1945 547 1951 581
rect 1985 547 2001 558
rect 1945 536 2001 547
rect 2035 581 2205 615
rect 1747 487 1763 503
rect 1439 469 1763 487
rect 1797 502 1813 503
rect 2035 502 2069 581
rect 1797 469 2069 502
rect 1439 468 2069 469
rect 2103 498 2137 547
rect 1439 453 1813 468
rect 2171 502 2205 581
rect 2239 592 2273 615
rect 2239 536 2273 547
rect 2307 599 2519 615
rect 2307 565 2469 599
rect 2503 565 2519 599
rect 2307 549 2519 565
rect 2609 607 2659 649
rect 2609 573 2625 607
rect 2307 502 2341 549
rect 2171 468 2341 502
rect 2375 482 2425 515
rect 2609 510 2659 573
rect 1439 425 1505 453
rect 2103 434 2137 464
rect 2409 448 2425 482
rect 2375 434 2425 448
rect 695 206 761 227
rect 695 172 711 206
rect 745 172 761 206
rect 695 151 761 172
rect 797 345 1088 379
rect 797 198 847 345
rect 831 164 847 198
rect 914 295 980 311
rect 914 261 930 295
rect 964 261 980 295
rect 914 225 980 261
rect 1022 302 1088 345
rect 1022 268 1038 302
rect 1072 268 1088 302
rect 1022 259 1088 268
rect 1122 225 1156 421
rect 1439 391 1455 425
rect 1489 391 1505 425
rect 1847 419 2270 434
rect 1439 319 1505 391
rect 1602 403 2270 419
rect 1602 369 1618 403
rect 1652 400 2270 403
rect 1652 385 1881 400
rect 1652 369 1668 385
rect 1602 353 1668 369
rect 1710 335 1776 351
rect 1945 350 2202 366
rect 1710 319 1726 335
rect 1408 301 1726 319
rect 1760 301 1776 335
rect 1408 285 1776 301
rect 1818 329 1884 345
rect 1818 295 1834 329
rect 1868 295 1884 329
rect 1945 316 2152 350
rect 2186 316 2202 350
rect 1945 300 2202 316
rect 914 191 1156 225
rect 797 135 847 164
rect 1122 177 1156 191
rect 17 76 49 110
rect 17 51 83 76
rect 119 105 185 134
rect 119 71 135 105
rect 169 71 185 105
rect 119 17 185 71
rect 305 109 461 134
rect 305 75 321 109
rect 355 100 461 109
rect 495 105 529 134
rect 355 75 371 100
rect 305 51 371 75
rect 495 17 529 71
rect 565 117 634 135
rect 881 123 1088 157
rect 565 110 714 117
rect 565 76 581 110
rect 615 101 714 110
rect 615 76 664 101
rect 565 67 664 76
rect 698 85 714 101
rect 881 85 915 123
rect 698 67 915 85
rect 565 51 915 67
rect 961 73 1011 89
rect 961 39 977 73
rect 1054 85 1088 123
rect 1122 119 1156 143
rect 1190 269 1308 285
rect 1190 235 1206 269
rect 1240 235 1274 269
rect 1190 219 1308 235
rect 1190 85 1224 219
rect 1408 185 1442 285
rect 1818 251 1884 295
rect 2236 266 2270 400
rect 1376 169 1442 185
rect 1410 135 1442 169
rect 1376 119 1442 135
rect 1476 217 1884 251
rect 2129 243 2270 266
rect 1476 85 1556 217
rect 1918 208 1984 224
rect 1918 183 1934 208
rect 1054 51 1556 85
rect 1590 163 1656 183
rect 1590 129 1606 163
rect 1640 129 1656 163
rect 961 17 1011 39
rect 1590 17 1656 129
rect 1794 174 1934 183
rect 1968 183 1984 208
rect 2129 209 2145 243
rect 2179 232 2270 243
rect 2304 400 2425 434
rect 2500 483 2566 499
rect 2500 449 2516 483
rect 2550 449 2566 483
rect 2500 413 2566 449
rect 2179 209 2195 232
rect 2129 187 2195 209
rect 2304 198 2338 400
rect 2500 379 2516 413
rect 2550 379 2566 413
rect 2500 329 2566 379
rect 2609 476 2625 510
rect 2609 413 2659 476
rect 2609 379 2625 413
rect 2609 363 2659 379
rect 2695 599 2767 615
rect 2695 565 2711 599
rect 2745 565 2767 599
rect 2695 506 2767 565
rect 2695 472 2711 506
rect 2745 472 2767 506
rect 2695 413 2767 472
rect 2695 379 2711 413
rect 2745 379 2767 413
rect 2695 363 2767 379
rect 2500 313 2699 329
rect 2500 279 2649 313
rect 2683 279 2699 313
rect 1968 174 2095 183
rect 1794 167 2095 174
rect 1794 133 1810 167
rect 1844 153 2095 167
rect 2229 164 2338 198
rect 2404 237 2454 266
rect 2438 203 2454 237
rect 2229 153 2263 164
rect 1844 149 2263 153
rect 1844 133 1860 149
rect 1794 117 1860 133
rect 2061 119 2263 149
rect 1961 100 2027 115
rect 1961 66 1977 100
rect 2011 85 2027 100
rect 2304 114 2370 130
rect 2304 85 2320 114
rect 2011 80 2320 85
rect 2354 80 2370 114
rect 2011 66 2370 80
rect 1961 51 2370 66
rect 2404 17 2454 203
rect 2500 263 2699 279
rect 2500 116 2566 263
rect 2733 229 2767 363
rect 2500 82 2516 116
rect 2550 82 2566 116
rect 2500 53 2566 82
rect 2609 213 2659 229
rect 2609 179 2625 213
rect 2609 103 2659 179
rect 2609 69 2625 103
rect 2609 17 2659 69
rect 2695 213 2767 229
rect 2695 179 2711 213
rect 2745 179 2767 213
rect 2695 103 2767 179
rect 2695 69 2711 103
rect 2745 69 2767 103
rect 2695 53 2767 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 1951 558 1967 581
rect 1967 558 1985 581
rect 1951 547 1985 558
rect 2239 558 2273 581
rect 2239 547 2273 558
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 14 581 2770 589
rect 14 547 1951 581
rect 1985 547 2239 581
rect 2273 547 2770 581
rect 14 535 2770 547
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 srsdfxtp_1
flabel metal1 s 14 535 2770 589 0 FreeSans 340 0 0 0 KAPWR
port 6 nsew power bidirectional
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 2719 94 2753 128 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 2719 168 2753 202 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2143 316 2177 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2335 94 2369 128 0 FreeSans 340 0 0 0 SLEEP_B
port 5 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6342382
string GDS_START 6323742
<< end >>
