magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 1165 186 1589 263
rect 1 157 427 178
rect 1165 157 2015 186
rect 1 49 2015 157
rect 0 0 2016 49
<< scnmos >>
rect 84 68 114 152
rect 156 68 186 152
rect 242 68 272 152
rect 314 68 344 152
rect 1247 153 1277 237
rect 1319 153 1349 237
rect 1405 153 1435 237
rect 1477 153 1507 237
rect 512 47 542 131
rect 584 47 614 131
rect 728 47 758 131
rect 806 47 836 131
rect 920 47 950 131
rect 1028 47 1058 131
rect 1673 76 1703 160
rect 1745 76 1775 160
rect 1831 76 1861 160
rect 1903 76 1933 160
<< scpmoshvt >>
rect 96 396 146 596
rect 202 396 252 596
rect 508 419 558 619
rect 648 419 698 619
rect 746 419 796 619
rect 854 419 904 619
rect 952 419 1002 619
rect 1120 419 1170 619
rect 1226 419 1276 619
rect 1500 419 1550 619
rect 1725 374 1775 574
rect 1831 374 1881 574
<< ndiff >>
rect 27 127 84 152
rect 27 93 39 127
rect 73 93 84 127
rect 27 68 84 93
rect 114 68 156 152
rect 186 127 242 152
rect 186 93 197 127
rect 231 93 242 127
rect 186 68 242 93
rect 272 68 314 152
rect 344 127 401 152
rect 1191 225 1247 237
rect 1191 191 1202 225
rect 1236 191 1247 225
rect 1191 153 1247 191
rect 1277 153 1319 237
rect 1349 199 1405 237
rect 1349 165 1360 199
rect 1394 165 1405 199
rect 1349 153 1405 165
rect 1435 153 1477 237
rect 1507 212 1563 237
rect 1507 178 1518 212
rect 1552 178 1563 212
rect 1507 153 1563 178
rect 344 93 355 127
rect 389 93 401 127
rect 344 68 401 93
rect 455 111 512 131
rect 455 77 467 111
rect 501 77 512 111
rect 455 47 512 77
rect 542 47 584 131
rect 614 106 728 131
rect 614 72 625 106
rect 659 72 728 106
rect 614 47 728 72
rect 758 47 806 131
rect 836 111 920 131
rect 836 77 875 111
rect 909 77 920 111
rect 836 47 920 77
rect 950 47 1028 131
rect 1058 85 1130 131
rect 1058 51 1085 85
rect 1119 51 1130 85
rect 1617 135 1673 160
rect 1617 101 1628 135
rect 1662 101 1673 135
rect 1617 76 1673 101
rect 1703 76 1745 160
rect 1775 135 1831 160
rect 1775 101 1786 135
rect 1820 101 1831 135
rect 1775 76 1831 101
rect 1861 76 1903 160
rect 1933 135 1989 160
rect 1933 101 1944 135
rect 1978 101 1989 135
rect 1933 76 1989 101
rect 1058 47 1130 51
rect 1073 39 1130 47
<< pdiff >>
rect 39 584 96 596
rect 39 550 51 584
rect 85 550 96 584
rect 39 513 96 550
rect 39 479 51 513
rect 85 479 96 513
rect 39 442 96 479
rect 39 408 51 442
rect 85 408 96 442
rect 39 396 96 408
rect 146 583 202 596
rect 146 549 157 583
rect 191 549 202 583
rect 146 396 202 549
rect 252 442 308 596
rect 252 408 263 442
rect 297 408 308 442
rect 252 396 308 408
rect 451 496 508 619
rect 451 462 463 496
rect 497 462 508 496
rect 451 419 508 462
rect 558 607 648 619
rect 558 573 603 607
rect 637 573 648 607
rect 558 531 648 573
rect 558 497 603 531
rect 637 497 648 531
rect 558 419 648 497
rect 698 419 746 619
rect 796 597 854 619
rect 796 563 809 597
rect 843 563 854 597
rect 796 465 854 563
rect 796 431 809 465
rect 843 431 854 465
rect 796 419 854 431
rect 904 419 952 619
rect 1002 607 1120 619
rect 1002 573 1013 607
rect 1047 573 1120 607
rect 1002 527 1120 573
rect 1002 493 1013 527
rect 1047 493 1120 527
rect 1002 419 1120 493
rect 1170 597 1226 619
rect 1170 563 1181 597
rect 1215 563 1226 597
rect 1170 465 1226 563
rect 1170 431 1181 465
rect 1215 431 1226 465
rect 1170 419 1226 431
rect 1276 607 1500 619
rect 1276 573 1455 607
rect 1489 573 1500 607
rect 1276 536 1500 573
rect 1276 502 1455 536
rect 1489 502 1500 536
rect 1276 465 1500 502
rect 1276 431 1455 465
rect 1489 431 1500 465
rect 1276 419 1500 431
rect 1550 597 1607 619
rect 1550 563 1561 597
rect 1595 563 1607 597
rect 1550 465 1607 563
rect 1550 431 1561 465
rect 1595 431 1607 465
rect 1550 419 1607 431
rect 1668 562 1725 574
rect 1668 528 1680 562
rect 1714 528 1725 562
rect 1668 491 1725 528
rect 1668 457 1680 491
rect 1714 457 1725 491
rect 1668 420 1725 457
rect 1668 386 1680 420
rect 1714 386 1725 420
rect 1668 374 1725 386
rect 1775 562 1831 574
rect 1775 528 1786 562
rect 1820 528 1831 562
rect 1775 491 1831 528
rect 1775 457 1786 491
rect 1820 457 1831 491
rect 1775 420 1831 457
rect 1775 386 1786 420
rect 1820 386 1831 420
rect 1775 374 1831 386
rect 1881 562 1938 574
rect 1881 528 1892 562
rect 1926 528 1938 562
rect 1881 491 1938 528
rect 1881 457 1892 491
rect 1926 457 1938 491
rect 1881 420 1938 457
rect 1881 386 1892 420
rect 1926 386 1938 420
rect 1881 374 1938 386
<< ndiffc >>
rect 39 93 73 127
rect 197 93 231 127
rect 1202 191 1236 225
rect 1360 165 1394 199
rect 1518 178 1552 212
rect 355 93 389 127
rect 467 77 501 111
rect 625 72 659 106
rect 875 77 909 111
rect 1085 51 1119 85
rect 1628 101 1662 135
rect 1786 101 1820 135
rect 1944 101 1978 135
<< pdiffc >>
rect 51 550 85 584
rect 51 479 85 513
rect 51 408 85 442
rect 157 549 191 583
rect 263 408 297 442
rect 463 462 497 496
rect 603 573 637 607
rect 603 497 637 531
rect 809 563 843 597
rect 809 431 843 465
rect 1013 573 1047 607
rect 1013 493 1047 527
rect 1181 563 1215 597
rect 1181 431 1215 465
rect 1455 573 1489 607
rect 1455 502 1489 536
rect 1455 431 1489 465
rect 1561 563 1595 597
rect 1561 431 1595 465
rect 1680 528 1714 562
rect 1680 457 1714 491
rect 1680 386 1714 420
rect 1786 528 1820 562
rect 1786 457 1820 491
rect 1786 386 1820 420
rect 1892 528 1926 562
rect 1892 457 1926 491
rect 1892 386 1926 420
<< poly >>
rect 96 596 146 622
rect 202 596 252 622
rect 508 619 558 645
rect 648 619 698 645
rect 746 619 796 645
rect 854 619 904 645
rect 952 619 1002 645
rect 1120 619 1170 645
rect 1226 619 1276 645
rect 1500 619 1550 645
rect 340 510 406 526
rect 340 476 356 510
rect 390 476 406 510
rect 340 442 406 476
rect 340 408 356 442
rect 390 408 406 442
rect 1725 574 1775 600
rect 1831 574 1881 600
rect 340 404 406 408
rect 508 404 558 419
rect 96 352 146 396
rect 84 336 154 352
rect 84 302 104 336
rect 138 302 154 336
rect 84 268 154 302
rect 202 326 252 396
rect 340 374 558 404
rect 648 387 698 419
rect 202 310 300 326
rect 202 296 250 310
rect 84 234 104 268
rect 138 248 154 268
rect 234 276 250 296
rect 284 276 300 310
rect 528 305 558 374
rect 632 371 698 387
rect 632 337 648 371
rect 682 337 698 371
rect 746 351 796 419
rect 854 377 904 419
rect 632 321 698 337
rect 740 335 806 351
rect 874 335 904 377
rect 138 234 186 248
rect 84 218 186 234
rect 84 152 114 218
rect 156 152 186 218
rect 234 242 300 276
rect 234 208 250 242
rect 284 222 300 242
rect 486 289 558 305
rect 486 255 502 289
rect 536 255 558 289
rect 284 208 344 222
rect 234 192 344 208
rect 242 152 272 192
rect 314 152 344 192
rect 486 221 558 255
rect 486 187 502 221
rect 536 201 558 221
rect 536 187 614 201
rect 486 171 614 187
rect 512 131 542 171
rect 584 131 614 171
rect 662 176 692 321
rect 740 301 756 335
rect 790 301 806 335
rect 740 285 806 301
rect 848 305 904 335
rect 952 371 1002 419
rect 1120 379 1170 419
rect 1226 387 1276 419
rect 952 355 1064 371
rect 952 321 1009 355
rect 1043 321 1064 355
rect 952 305 1064 321
rect 1112 363 1178 379
rect 1112 329 1128 363
rect 1162 329 1178 363
rect 1112 313 1178 329
rect 1226 371 1349 387
rect 1226 337 1283 371
rect 1317 337 1349 371
rect 1226 321 1349 337
rect 1500 325 1550 419
rect 848 237 878 305
rect 806 221 878 237
rect 806 187 822 221
rect 856 207 878 221
rect 920 241 986 257
rect 920 207 936 241
rect 970 207 986 241
rect 856 187 872 207
rect 662 146 758 176
rect 728 131 758 146
rect 806 171 872 187
rect 920 191 986 207
rect 806 131 836 171
rect 920 131 950 191
rect 1028 131 1058 305
rect 1146 131 1176 313
rect 1247 237 1277 263
rect 1319 237 1349 321
rect 1400 309 1550 325
rect 1400 275 1416 309
rect 1450 289 1550 309
rect 1725 289 1775 374
rect 1450 275 1775 289
rect 1400 259 1775 275
rect 1405 237 1435 259
rect 1477 237 1507 259
rect 1673 160 1703 259
rect 1745 160 1775 259
rect 1831 334 1881 374
rect 1831 318 1897 334
rect 1831 284 1847 318
rect 1881 284 1897 318
rect 1831 250 1897 284
rect 1831 216 1847 250
rect 1881 230 1897 250
rect 1881 216 1933 230
rect 1831 200 1933 216
rect 1831 160 1861 200
rect 1903 160 1933 200
rect 1247 131 1277 153
rect 84 42 114 68
rect 156 42 186 68
rect 242 42 272 68
rect 314 42 344 68
rect 1146 115 1277 131
rect 1319 127 1349 153
rect 1405 127 1435 153
rect 1477 127 1507 153
rect 1146 81 1187 115
rect 1221 101 1277 115
rect 1221 81 1237 101
rect 1146 65 1237 81
rect 1673 50 1703 76
rect 1745 50 1775 76
rect 1831 50 1861 76
rect 1903 50 1933 76
rect 512 21 542 47
rect 584 21 614 47
rect 728 21 758 47
rect 806 21 836 47
rect 920 21 950 47
rect 1028 21 1058 47
<< polycont >>
rect 356 476 390 510
rect 356 408 390 442
rect 104 302 138 336
rect 104 234 138 268
rect 250 276 284 310
rect 648 337 682 371
rect 250 208 284 242
rect 502 255 536 289
rect 502 187 536 221
rect 756 301 790 335
rect 1009 321 1043 355
rect 1128 329 1162 363
rect 1283 337 1317 371
rect 822 187 856 221
rect 936 207 970 241
rect 1416 275 1450 309
rect 1847 284 1881 318
rect 1847 216 1881 250
rect 1187 81 1221 115
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 18 584 101 600
rect 18 550 51 584
rect 85 550 101 584
rect 18 513 101 550
rect 141 583 207 649
rect 141 549 157 583
rect 191 549 207 583
rect 141 548 207 549
rect 243 579 567 613
rect 18 479 51 513
rect 85 512 101 513
rect 243 512 277 579
rect 85 479 277 512
rect 18 478 277 479
rect 339 510 393 526
rect 18 442 101 478
rect 339 476 356 510
rect 390 476 393 510
rect 339 442 393 476
rect 18 408 51 442
rect 85 408 101 442
rect 18 392 101 408
rect 247 408 263 442
rect 297 408 356 442
rect 390 408 393 442
rect 247 392 393 408
rect 18 156 52 392
rect 88 336 167 356
rect 88 302 104 336
rect 138 302 167 336
rect 88 268 167 302
rect 88 234 104 268
rect 138 234 167 268
rect 88 218 167 234
rect 217 310 300 356
rect 217 276 250 310
rect 284 276 300 310
rect 217 242 300 276
rect 217 208 250 242
rect 284 208 300 242
rect 217 192 300 208
rect 18 127 89 156
rect 18 93 39 127
rect 73 93 89 127
rect 18 64 89 93
rect 181 127 247 156
rect 181 93 197 127
rect 231 93 247 127
rect 181 17 247 93
rect 339 127 393 392
rect 339 93 355 127
rect 389 93 393 127
rect 339 64 393 93
rect 429 496 497 543
rect 429 462 463 496
rect 429 375 497 462
rect 533 445 567 579
rect 603 607 653 649
rect 637 573 653 607
rect 603 531 653 573
rect 637 497 653 531
rect 603 481 653 497
rect 793 597 859 613
rect 793 563 809 597
rect 843 563 859 597
rect 793 465 859 563
rect 997 607 1063 649
rect 997 573 1013 607
rect 1047 573 1063 607
rect 997 527 1063 573
rect 997 493 1013 527
rect 1047 493 1063 527
rect 997 477 1063 493
rect 1165 597 1231 613
rect 1165 563 1181 597
rect 1215 574 1231 597
rect 1439 607 1505 649
rect 1215 563 1403 574
rect 1165 540 1403 563
rect 533 411 698 445
rect 429 341 609 375
rect 429 135 463 341
rect 499 289 539 305
rect 499 255 502 289
rect 536 255 539 289
rect 499 221 539 255
rect 575 285 609 341
rect 645 371 698 411
rect 793 431 809 465
rect 843 441 859 465
rect 1165 465 1231 540
rect 843 431 1129 441
rect 793 407 1129 431
rect 1165 431 1181 465
rect 1215 431 1231 465
rect 1165 415 1231 431
rect 1095 379 1129 407
rect 645 337 648 371
rect 682 337 698 371
rect 993 355 1059 371
rect 645 321 698 337
rect 736 335 806 351
rect 736 301 756 335
rect 790 319 806 335
rect 993 321 1009 355
rect 1043 321 1059 355
rect 790 301 954 319
rect 993 305 1059 321
rect 1095 363 1178 379
rect 1095 329 1128 363
rect 1162 329 1178 363
rect 1095 313 1178 329
rect 1267 371 1333 504
rect 1267 337 1283 371
rect 1317 337 1333 371
rect 1267 321 1333 337
rect 1369 325 1403 540
rect 1439 573 1455 607
rect 1489 573 1505 607
rect 1439 536 1505 573
rect 1439 502 1455 536
rect 1489 502 1505 536
rect 1439 465 1505 502
rect 1439 431 1455 465
rect 1489 431 1505 465
rect 1439 415 1505 431
rect 1541 597 1611 613
rect 1541 563 1561 597
rect 1595 563 1611 597
rect 1541 465 1611 563
rect 1541 431 1561 465
rect 1595 431 1611 465
rect 736 285 954 301
rect 575 251 770 285
rect 920 257 954 285
rect 920 241 986 257
rect 499 187 502 221
rect 536 205 539 221
rect 806 221 872 237
rect 806 205 822 221
rect 536 187 822 205
rect 856 187 872 221
rect 920 207 936 241
rect 970 207 986 241
rect 920 191 986 207
rect 1025 241 1059 305
rect 1369 309 1466 325
rect 1369 285 1416 309
rect 1218 275 1416 285
rect 1450 275 1466 309
rect 1218 251 1466 275
rect 1218 241 1252 251
rect 1541 241 1611 431
rect 1025 225 1252 241
rect 1025 191 1202 225
rect 1236 191 1252 225
rect 1502 236 1611 241
rect 1647 562 1730 578
rect 1647 528 1680 562
rect 1714 528 1730 562
rect 1647 491 1730 528
rect 1647 457 1680 491
rect 1714 457 1730 491
rect 1647 420 1730 457
rect 1647 386 1680 420
rect 1714 386 1730 420
rect 1344 199 1410 215
rect 499 171 872 187
rect 1344 165 1360 199
rect 1394 165 1410 199
rect 908 135 1237 155
rect 429 111 517 135
rect 429 77 467 111
rect 501 77 517 111
rect 429 53 517 77
rect 609 106 675 135
rect 609 72 625 106
rect 659 72 675 106
rect 609 17 675 72
rect 859 121 1237 135
rect 859 111 942 121
rect 859 77 875 111
rect 909 77 942 111
rect 1171 115 1237 121
rect 859 53 942 77
rect 1069 51 1085 85
rect 1119 51 1135 85
rect 1171 81 1187 115
rect 1221 81 1237 115
rect 1171 65 1237 81
rect 1069 17 1135 51
rect 1344 17 1410 165
rect 1502 212 1575 236
rect 1502 178 1518 212
rect 1552 178 1575 212
rect 1502 149 1575 178
rect 1647 234 1730 386
rect 1770 562 1836 649
rect 1770 528 1786 562
rect 1820 528 1836 562
rect 1770 491 1836 528
rect 1770 457 1786 491
rect 1820 457 1836 491
rect 1770 420 1836 457
rect 1770 386 1786 420
rect 1820 386 1836 420
rect 1770 370 1836 386
rect 1876 562 1994 578
rect 1876 528 1892 562
rect 1926 528 1994 562
rect 1876 491 1994 528
rect 1876 457 1892 491
rect 1926 457 1994 491
rect 1876 420 1994 457
rect 1876 386 1892 420
rect 1926 386 1994 420
rect 1876 370 1994 386
rect 1831 318 1897 334
rect 1831 284 1847 318
rect 1881 284 1897 318
rect 1831 250 1897 284
rect 1831 234 1847 250
rect 1647 216 1847 234
rect 1881 216 1897 250
rect 1647 200 1897 216
rect 1647 164 1681 200
rect 1960 164 1994 370
rect 1612 135 1681 164
rect 1612 101 1628 135
rect 1662 101 1681 135
rect 1612 72 1681 101
rect 1770 135 1836 164
rect 1770 101 1786 135
rect 1820 101 1836 135
rect 1770 17 1836 101
rect 1928 135 1994 164
rect 1928 101 1944 135
rect 1978 101 1994 135
rect 1928 72 1994 101
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrbn_lp
flabel comment s 1179 88 1179 88 0 FreeSans 300 180 0 0 no_jumper_check
flabel comment s 1179 340 1179 340 0 FreeSans 300 180 0 0 no_jumper_check
flabel comment s 526 271 526 271 0 FreeSans 200 270 0 0 no_jumper_check
flabel comment s 379 418 379 418 0 FreeSans 200 270 0 0 no_jumper_check
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1279 464 1313 498 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1951 390 1985 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1951 464 1985 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1951 538 1985 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6249008
string GDS_START 6234180
<< end >>
