magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 760 241
rect 0 0 768 49
<< scnmos >>
rect 80 47 110 215
rect 243 47 273 215
rect 333 47 363 215
rect 423 47 453 215
rect 543 47 573 215
rect 651 47 681 215
<< scpmoshvt >>
rect 129 367 159 619
rect 229 367 259 619
rect 315 367 345 619
rect 471 367 501 619
rect 579 367 609 619
rect 651 367 681 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 101 80 169
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 127 243 215
rect 110 93 121 127
rect 155 93 198 127
rect 232 93 243 127
rect 110 47 243 93
rect 273 47 333 215
rect 363 47 423 215
rect 453 203 543 215
rect 453 169 481 203
rect 515 169 543 203
rect 453 101 543 169
rect 453 67 481 101
rect 515 67 543 101
rect 453 47 543 67
rect 573 129 651 215
rect 573 95 592 129
rect 626 95 651 129
rect 573 47 651 95
rect 681 203 734 215
rect 681 169 692 203
rect 726 169 734 203
rect 681 93 734 169
rect 681 59 692 93
rect 726 59 734 93
rect 681 47 734 59
<< pdiff >>
rect 76 599 129 619
rect 76 565 84 599
rect 118 565 129 599
rect 76 519 129 565
rect 76 485 84 519
rect 118 485 129 519
rect 76 441 129 485
rect 76 407 84 441
rect 118 407 129 441
rect 76 367 129 407
rect 159 607 229 619
rect 159 573 178 607
rect 212 573 229 607
rect 159 532 229 573
rect 159 498 178 532
rect 212 498 229 532
rect 159 457 229 498
rect 159 423 178 457
rect 212 423 229 457
rect 159 367 229 423
rect 259 599 315 619
rect 259 565 270 599
rect 304 565 315 599
rect 259 522 315 565
rect 259 488 270 522
rect 304 488 315 522
rect 259 441 315 488
rect 259 407 270 441
rect 304 407 315 441
rect 259 367 315 407
rect 345 607 471 619
rect 345 573 356 607
rect 390 573 426 607
rect 460 573 471 607
rect 345 513 471 573
rect 345 479 356 513
rect 390 479 426 513
rect 460 479 471 513
rect 345 367 471 479
rect 501 607 579 619
rect 501 573 526 607
rect 560 573 579 607
rect 501 529 579 573
rect 501 495 526 529
rect 560 495 579 529
rect 501 441 579 495
rect 501 407 526 441
rect 560 407 579 441
rect 501 367 579 407
rect 609 367 651 619
rect 681 607 734 619
rect 681 573 692 607
rect 726 573 734 607
rect 681 508 734 573
rect 681 474 692 508
rect 726 474 734 508
rect 681 413 734 474
rect 681 379 692 413
rect 726 379 734 413
rect 681 367 734 379
<< ndiffc >>
rect 35 169 69 203
rect 35 67 69 101
rect 121 93 155 127
rect 198 93 232 127
rect 481 169 515 203
rect 481 67 515 101
rect 592 95 626 129
rect 692 169 726 203
rect 692 59 726 93
<< pdiffc >>
rect 84 565 118 599
rect 84 485 118 519
rect 84 407 118 441
rect 178 573 212 607
rect 178 498 212 532
rect 178 423 212 457
rect 270 565 304 599
rect 270 488 304 522
rect 270 407 304 441
rect 356 573 390 607
rect 426 573 460 607
rect 356 479 390 513
rect 426 479 460 513
rect 526 573 560 607
rect 526 495 560 529
rect 526 407 560 441
rect 692 573 726 607
rect 692 474 726 508
rect 692 379 726 413
<< poly >>
rect 129 619 159 645
rect 229 619 259 645
rect 315 619 345 645
rect 471 619 501 645
rect 579 619 609 645
rect 651 619 681 645
rect 129 303 159 367
rect 229 305 259 367
rect 80 287 159 303
rect 80 253 105 287
rect 139 253 159 287
rect 80 237 159 253
rect 207 289 273 305
rect 207 255 223 289
rect 257 255 273 289
rect 207 239 273 255
rect 80 215 110 237
rect 243 215 273 239
rect 315 303 345 367
rect 471 305 501 367
rect 315 287 381 303
rect 315 253 331 287
rect 365 253 381 287
rect 315 237 381 253
rect 423 289 501 305
rect 579 303 609 367
rect 423 255 439 289
rect 473 255 501 289
rect 423 239 501 255
rect 543 287 609 303
rect 543 253 559 287
rect 593 253 609 287
rect 333 215 363 237
rect 423 215 453 239
rect 543 237 609 253
rect 651 305 681 367
rect 651 289 747 305
rect 651 255 697 289
rect 731 255 747 289
rect 651 239 747 255
rect 543 215 573 237
rect 651 215 681 239
rect 80 21 110 47
rect 243 21 273 47
rect 333 21 363 47
rect 423 21 453 47
rect 543 21 573 47
rect 651 21 681 47
<< polycont >>
rect 105 253 139 287
rect 223 255 257 289
rect 331 253 365 287
rect 439 255 473 289
rect 559 253 593 287
rect 697 255 731 289
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 599 134 615
rect 17 565 84 599
rect 118 565 134 599
rect 17 519 134 565
rect 17 485 84 519
rect 118 485 134 519
rect 17 441 134 485
rect 17 407 84 441
rect 118 407 134 441
rect 168 607 220 649
rect 168 573 178 607
rect 212 573 220 607
rect 168 532 220 573
rect 168 498 178 532
rect 212 498 220 532
rect 168 457 220 498
rect 168 423 178 457
rect 212 423 220 457
rect 168 407 220 423
rect 254 599 306 615
rect 254 565 270 599
rect 304 565 306 599
rect 254 522 306 565
rect 254 488 270 522
rect 304 488 306 522
rect 254 441 306 488
rect 340 607 476 649
rect 340 573 356 607
rect 390 573 426 607
rect 460 573 476 607
rect 340 513 476 573
rect 340 479 356 513
rect 390 479 426 513
rect 460 479 476 513
rect 340 475 476 479
rect 510 607 576 615
rect 510 573 526 607
rect 560 573 576 607
rect 510 529 576 573
rect 510 495 526 529
rect 560 495 576 529
rect 510 441 576 495
rect 254 407 270 441
rect 304 407 526 441
rect 560 407 576 441
rect 676 607 742 615
rect 676 573 692 607
rect 726 573 742 607
rect 676 508 742 573
rect 676 474 692 508
rect 726 474 742 508
rect 676 413 742 474
rect 17 203 71 407
rect 676 379 692 413
rect 726 379 742 413
rect 676 373 742 379
rect 121 339 742 373
rect 121 303 168 339
rect 17 169 35 203
rect 69 169 71 203
rect 105 287 168 303
rect 139 253 168 287
rect 105 205 168 253
rect 202 289 273 305
rect 202 255 223 289
rect 257 255 273 289
rect 202 239 273 255
rect 307 287 381 305
rect 307 253 331 287
rect 365 253 381 287
rect 307 239 381 253
rect 415 289 473 305
rect 415 255 439 289
rect 415 239 473 255
rect 507 287 643 305
rect 507 253 559 287
rect 593 253 643 287
rect 507 239 643 253
rect 677 289 751 305
rect 677 255 697 289
rect 731 255 751 289
rect 677 239 751 255
rect 105 203 742 205
rect 105 171 481 203
rect 17 101 71 169
rect 465 169 481 171
rect 515 171 692 203
rect 515 169 531 171
rect 17 67 35 101
rect 69 67 71 101
rect 17 51 71 67
rect 105 127 248 137
rect 105 93 121 127
rect 155 93 198 127
rect 232 93 248 127
rect 105 17 248 93
rect 465 101 531 169
rect 676 169 692 171
rect 726 169 742 203
rect 465 67 481 101
rect 515 67 531 101
rect 465 51 531 67
rect 576 129 642 137
rect 576 95 592 129
rect 626 95 642 129
rect 576 17 642 95
rect 676 93 742 169
rect 676 59 692 93
rect 726 59 742 93
rect 676 51 742 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a311o_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3907544
string GDS_START 3899860
<< end >>
