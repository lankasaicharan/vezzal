magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 58 49 534 241
rect 0 0 576 49
<< scnmos >>
rect 137 131 167 215
rect 245 47 275 215
rect 336 47 366 215
rect 425 47 455 215
<< scpmoshvt >>
rect 137 367 167 451
rect 245 367 275 619
rect 331 367 361 619
rect 425 367 455 619
<< ndiff >>
rect 84 203 137 215
rect 84 169 92 203
rect 126 169 137 203
rect 84 131 137 169
rect 167 183 245 215
rect 167 149 180 183
rect 214 149 245 183
rect 167 131 245 149
rect 192 93 245 131
rect 192 59 200 93
rect 234 59 245 93
rect 192 47 245 59
rect 275 47 336 215
rect 366 47 425 215
rect 455 183 508 215
rect 455 149 466 183
rect 500 149 508 183
rect 455 93 508 149
rect 455 59 466 93
rect 500 59 508 93
rect 455 47 508 59
<< pdiff >>
rect 192 607 245 619
rect 192 573 200 607
rect 234 573 245 607
rect 192 521 245 573
rect 192 487 200 521
rect 234 487 245 521
rect 192 451 245 487
rect 84 426 137 451
rect 84 392 92 426
rect 126 392 137 426
rect 84 367 137 392
rect 167 434 245 451
rect 167 400 178 434
rect 212 400 245 434
rect 167 367 245 400
rect 275 599 331 619
rect 275 565 286 599
rect 320 565 331 599
rect 275 510 331 565
rect 275 476 286 510
rect 320 476 331 510
rect 275 418 331 476
rect 275 384 286 418
rect 320 384 331 418
rect 275 367 331 384
rect 361 611 425 619
rect 361 577 377 611
rect 411 577 425 611
rect 361 490 425 577
rect 361 456 377 490
rect 411 456 425 490
rect 361 367 425 456
rect 455 599 508 619
rect 455 565 466 599
rect 500 565 508 599
rect 455 510 508 565
rect 455 476 466 510
rect 500 476 508 510
rect 455 418 508 476
rect 455 384 466 418
rect 500 384 508 418
rect 455 367 508 384
<< ndiffc >>
rect 92 169 126 203
rect 180 149 214 183
rect 200 59 234 93
rect 466 149 500 183
rect 466 59 500 93
<< pdiffc >>
rect 200 573 234 607
rect 200 487 234 521
rect 92 392 126 426
rect 178 400 212 434
rect 286 565 320 599
rect 286 476 320 510
rect 286 384 320 418
rect 377 577 411 611
rect 377 456 411 490
rect 466 565 500 599
rect 466 476 500 510
rect 466 384 500 418
<< poly >>
rect 245 619 275 645
rect 331 619 361 645
rect 425 619 455 645
rect 137 451 167 477
rect 137 335 167 367
rect 245 335 275 367
rect 331 335 361 367
rect 101 319 167 335
rect 101 285 117 319
rect 151 285 167 319
rect 101 269 167 285
rect 209 319 275 335
rect 209 285 225 319
rect 259 285 275 319
rect 209 269 275 285
rect 317 319 383 335
rect 317 285 333 319
rect 367 285 383 319
rect 317 269 383 285
rect 425 303 455 367
rect 425 287 491 303
rect 137 215 167 269
rect 245 215 275 269
rect 336 215 366 269
rect 425 253 441 287
rect 475 253 491 287
rect 425 237 491 253
rect 425 215 455 237
rect 137 105 167 131
rect 245 21 275 47
rect 336 21 366 47
rect 425 21 455 47
<< polycont >>
rect 117 285 151 319
rect 225 285 259 319
rect 333 285 367 319
rect 441 253 475 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 176 607 236 649
rect 176 573 200 607
rect 234 573 236 607
rect 176 521 236 573
rect 176 487 200 521
rect 234 487 236 521
rect 31 426 142 442
rect 31 392 92 426
rect 126 392 142 426
rect 31 384 142 392
rect 176 434 236 487
rect 176 400 178 434
rect 212 400 236 434
rect 176 384 236 400
rect 270 599 327 615
rect 270 565 286 599
rect 320 565 327 599
rect 270 510 327 565
rect 270 476 286 510
rect 320 476 327 510
rect 270 418 327 476
rect 361 611 427 649
rect 361 577 377 611
rect 411 577 427 611
rect 361 490 427 577
rect 361 456 377 490
rect 411 456 427 490
rect 361 452 427 456
rect 462 599 559 615
rect 462 565 466 599
rect 500 565 559 599
rect 462 510 559 565
rect 462 476 466 510
rect 500 476 559 510
rect 462 418 559 476
rect 270 384 286 418
rect 320 384 466 418
rect 500 384 559 418
rect 31 251 65 384
rect 101 319 175 350
rect 101 285 117 319
rect 151 285 175 319
rect 209 319 275 350
rect 209 285 225 319
rect 259 285 275 319
rect 309 319 383 350
rect 309 285 333 319
rect 367 285 383 319
rect 425 287 475 303
rect 425 253 441 287
rect 425 251 475 253
rect 31 217 475 251
rect 31 203 130 217
rect 31 169 92 203
rect 126 169 130 203
rect 509 183 559 384
rect 31 153 130 169
rect 164 149 180 183
rect 214 149 238 183
rect 164 93 238 149
rect 164 59 200 93
rect 234 59 238 93
rect 164 17 238 59
rect 441 149 466 183
rect 500 149 559 183
rect 441 93 559 149
rect 441 59 466 93
rect 500 59 559 93
rect 441 55 559 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand3b_1
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3710078
string GDS_START 3704210
<< end >>
