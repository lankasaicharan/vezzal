magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3026 1975
<< nwell >>
rect -38 331 1766 704
<< pwell >>
rect 1 201 813 241
rect 1511 201 1721 241
rect 1 49 1721 201
rect 0 0 1728 49
<< scnmos >>
rect 84 47 114 215
rect 170 47 200 215
rect 256 47 286 215
rect 342 47 372 215
rect 428 47 458 215
rect 514 47 544 215
rect 614 47 644 215
rect 700 47 730 215
rect 809 47 839 175
rect 895 47 925 175
rect 995 47 1025 175
rect 1095 47 1125 175
rect 1213 47 1243 175
rect 1299 47 1329 175
rect 1385 47 1415 175
rect 1485 47 1515 175
rect 1608 47 1638 215
<< scpmoshvt >>
rect 84 367 114 619
rect 170 367 200 619
rect 256 367 286 619
rect 342 367 372 619
rect 428 367 458 619
rect 514 367 544 619
rect 600 367 630 619
rect 686 367 716 619
rect 813 419 843 619
rect 913 419 943 619
rect 999 419 1029 619
rect 1099 419 1129 619
rect 1213 419 1243 619
rect 1299 419 1329 619
rect 1399 419 1429 619
rect 1501 419 1531 619
rect 1610 367 1640 619
<< ndiff >>
rect 27 207 84 215
rect 27 173 39 207
rect 73 173 84 207
rect 27 89 84 173
rect 27 55 39 89
rect 73 55 84 89
rect 27 47 84 55
rect 114 203 170 215
rect 114 169 125 203
rect 159 169 170 203
rect 114 93 170 169
rect 114 59 125 93
rect 159 59 170 93
rect 114 47 170 59
rect 200 114 256 215
rect 200 80 211 114
rect 245 80 256 114
rect 200 47 256 80
rect 286 203 342 215
rect 286 169 297 203
rect 331 169 342 203
rect 286 93 342 169
rect 286 59 297 93
rect 331 59 342 93
rect 286 47 342 59
rect 372 114 428 215
rect 372 80 383 114
rect 417 80 428 114
rect 372 47 428 80
rect 458 203 514 215
rect 458 169 469 203
rect 503 169 514 203
rect 458 93 514 169
rect 458 59 469 93
rect 503 59 514 93
rect 458 47 514 59
rect 544 114 614 215
rect 544 80 555 114
rect 589 80 614 114
rect 544 47 614 80
rect 644 203 700 215
rect 644 169 655 203
rect 689 169 700 203
rect 644 93 700 169
rect 644 59 655 93
rect 689 59 700 93
rect 644 47 700 59
rect 730 203 787 215
rect 730 169 741 203
rect 775 175 787 203
rect 1537 175 1608 215
rect 775 169 809 175
rect 730 93 809 169
rect 730 59 741 93
rect 775 59 809 93
rect 730 47 809 59
rect 839 102 895 175
rect 839 68 850 102
rect 884 68 895 102
rect 839 47 895 68
rect 925 154 995 175
rect 925 120 950 154
rect 984 120 995 154
rect 925 47 995 120
rect 1025 102 1095 175
rect 1025 68 1050 102
rect 1084 68 1095 102
rect 1025 47 1095 68
rect 1125 87 1213 175
rect 1125 53 1152 87
rect 1186 53 1213 87
rect 1125 47 1213 53
rect 1243 93 1299 175
rect 1243 59 1254 93
rect 1288 59 1299 93
rect 1243 47 1299 59
rect 1329 162 1385 175
rect 1329 128 1340 162
rect 1374 128 1385 162
rect 1329 47 1385 128
rect 1415 122 1485 175
rect 1415 88 1440 122
rect 1474 88 1485 122
rect 1415 47 1485 88
rect 1515 122 1608 175
rect 1515 88 1549 122
rect 1583 88 1608 122
rect 1515 47 1608 88
rect 1638 203 1695 215
rect 1638 169 1649 203
rect 1683 169 1695 203
rect 1638 101 1695 169
rect 1638 67 1649 101
rect 1683 67 1695 101
rect 1638 47 1695 67
rect 1140 41 1198 47
<< pdiff >>
rect 27 607 84 619
rect 27 573 39 607
rect 73 573 84 607
rect 27 503 84 573
rect 27 469 39 503
rect 73 469 84 503
rect 27 409 84 469
rect 27 375 39 409
rect 73 375 84 409
rect 27 367 84 375
rect 114 599 170 619
rect 114 565 125 599
rect 159 565 170 599
rect 114 506 170 565
rect 114 472 125 506
rect 159 472 170 506
rect 114 413 170 472
rect 114 379 125 413
rect 159 379 170 413
rect 114 367 170 379
rect 200 607 256 619
rect 200 573 211 607
rect 245 573 256 607
rect 200 481 256 573
rect 200 447 211 481
rect 245 447 256 481
rect 200 367 256 447
rect 286 599 342 619
rect 286 565 297 599
rect 331 565 342 599
rect 286 506 342 565
rect 286 472 297 506
rect 331 472 342 506
rect 286 413 342 472
rect 286 379 297 413
rect 331 379 342 413
rect 286 367 342 379
rect 372 607 428 619
rect 372 573 383 607
rect 417 573 428 607
rect 372 481 428 573
rect 372 447 383 481
rect 417 447 428 481
rect 372 367 428 447
rect 458 599 514 619
rect 458 565 469 599
rect 503 565 514 599
rect 458 506 514 565
rect 458 472 469 506
rect 503 472 514 506
rect 458 413 514 472
rect 458 379 469 413
rect 503 379 514 413
rect 458 367 514 379
rect 544 607 600 619
rect 544 573 555 607
rect 589 573 600 607
rect 544 481 600 573
rect 544 447 555 481
rect 589 447 600 481
rect 544 367 600 447
rect 630 599 686 619
rect 630 565 641 599
rect 675 565 686 599
rect 630 506 686 565
rect 630 472 641 506
rect 675 472 686 506
rect 630 413 686 472
rect 630 379 641 413
rect 675 379 686 413
rect 630 367 686 379
rect 716 594 813 619
rect 716 560 727 594
rect 761 560 813 594
rect 716 419 813 560
rect 843 599 913 619
rect 843 565 854 599
rect 888 565 913 599
rect 843 419 913 565
rect 943 531 999 619
rect 943 497 954 531
rect 988 497 999 531
rect 943 419 999 497
rect 1029 599 1099 619
rect 1029 565 1054 599
rect 1088 565 1099 599
rect 1029 419 1099 565
rect 1129 606 1213 619
rect 1129 572 1154 606
rect 1188 572 1213 606
rect 1129 419 1213 572
rect 1243 594 1299 619
rect 1243 560 1254 594
rect 1288 560 1299 594
rect 1243 419 1299 560
rect 1329 534 1399 619
rect 1329 500 1354 534
rect 1388 500 1399 534
rect 1329 419 1399 500
rect 1429 590 1501 619
rect 1429 556 1454 590
rect 1488 556 1501 590
rect 1429 419 1501 556
rect 1531 594 1610 619
rect 1531 560 1565 594
rect 1599 560 1610 594
rect 1531 419 1610 560
rect 716 367 773 419
rect 1553 367 1610 419
rect 1640 599 1697 619
rect 1640 565 1651 599
rect 1685 565 1697 599
rect 1640 509 1697 565
rect 1640 475 1651 509
rect 1685 475 1697 509
rect 1640 419 1697 475
rect 1640 385 1651 419
rect 1685 385 1697 419
rect 1640 367 1697 385
<< ndiffc >>
rect 39 173 73 207
rect 39 55 73 89
rect 125 169 159 203
rect 125 59 159 93
rect 211 80 245 114
rect 297 169 331 203
rect 297 59 331 93
rect 383 80 417 114
rect 469 169 503 203
rect 469 59 503 93
rect 555 80 589 114
rect 655 169 689 203
rect 655 59 689 93
rect 741 169 775 203
rect 741 59 775 93
rect 850 68 884 102
rect 950 120 984 154
rect 1050 68 1084 102
rect 1152 53 1186 87
rect 1254 59 1288 93
rect 1340 128 1374 162
rect 1440 88 1474 122
rect 1549 88 1583 122
rect 1649 169 1683 203
rect 1649 67 1683 101
<< pdiffc >>
rect 39 573 73 607
rect 39 469 73 503
rect 39 375 73 409
rect 125 565 159 599
rect 125 472 159 506
rect 125 379 159 413
rect 211 573 245 607
rect 211 447 245 481
rect 297 565 331 599
rect 297 472 331 506
rect 297 379 331 413
rect 383 573 417 607
rect 383 447 417 481
rect 469 565 503 599
rect 469 472 503 506
rect 469 379 503 413
rect 555 573 589 607
rect 555 447 589 481
rect 641 565 675 599
rect 641 472 675 506
rect 641 379 675 413
rect 727 560 761 594
rect 854 565 888 599
rect 954 497 988 531
rect 1054 565 1088 599
rect 1154 572 1188 606
rect 1254 560 1288 594
rect 1354 500 1388 534
rect 1454 556 1488 590
rect 1565 560 1599 594
rect 1651 565 1685 599
rect 1651 475 1685 509
rect 1651 385 1685 419
<< poly >>
rect 84 619 114 645
rect 170 619 200 645
rect 256 619 286 645
rect 342 619 372 645
rect 428 619 458 645
rect 514 619 544 645
rect 600 619 630 645
rect 686 619 716 645
rect 813 619 843 645
rect 913 619 943 645
rect 999 619 1029 645
rect 1099 619 1129 645
rect 1213 619 1243 645
rect 1299 619 1329 645
rect 1399 619 1429 645
rect 1501 619 1531 645
rect 1610 619 1640 645
rect 813 387 843 419
rect 805 371 871 387
rect 84 319 114 367
rect 170 319 200 367
rect 256 319 286 367
rect 342 319 372 367
rect 428 319 458 367
rect 514 319 544 367
rect 600 319 630 367
rect 686 319 716 367
rect 805 337 821 371
rect 855 337 871 371
rect 913 379 943 419
rect 999 379 1029 419
rect 913 363 1029 379
rect 1099 377 1129 419
rect 1213 377 1243 419
rect 1299 385 1329 419
rect 1399 385 1429 419
rect 913 349 979 363
rect 805 321 871 337
rect 963 329 979 349
rect 1013 329 1029 363
rect 84 303 750 319
rect 84 269 224 303
rect 258 269 292 303
rect 326 269 360 303
rect 394 269 428 303
rect 462 269 496 303
rect 530 269 564 303
rect 598 269 632 303
rect 666 269 700 303
rect 734 269 750 303
rect 84 253 750 269
rect 84 215 114 253
rect 170 215 200 253
rect 256 215 286 253
rect 342 215 372 253
rect 428 215 458 253
rect 514 215 544 253
rect 614 215 644 253
rect 700 215 730 253
rect 809 175 839 321
rect 963 313 1029 329
rect 1071 361 1137 377
rect 1071 327 1087 361
rect 1121 327 1137 361
rect 1071 311 1137 327
rect 1179 361 1245 377
rect 1179 327 1195 361
rect 1229 327 1245 361
rect 1299 369 1429 385
rect 1299 355 1369 369
rect 1179 311 1245 327
rect 1353 335 1369 355
rect 1403 335 1429 369
rect 1353 319 1429 335
rect 895 255 961 271
rect 895 221 911 255
rect 945 235 961 255
rect 945 221 1025 235
rect 895 205 1025 221
rect 895 175 925 205
rect 995 175 1025 205
rect 1095 175 1125 311
rect 1213 175 1243 311
rect 1501 303 1531 419
rect 1610 335 1640 367
rect 1608 319 1674 335
rect 1473 287 1539 303
rect 1353 255 1419 271
rect 1353 235 1369 255
rect 1299 221 1369 235
rect 1403 221 1419 255
rect 1473 253 1489 287
rect 1523 253 1539 287
rect 1473 237 1539 253
rect 1608 285 1624 319
rect 1658 285 1674 319
rect 1608 269 1674 285
rect 1299 205 1419 221
rect 1299 175 1329 205
rect 1385 175 1415 205
rect 1485 175 1515 237
rect 1608 215 1638 269
rect 84 21 114 47
rect 170 21 200 47
rect 256 21 286 47
rect 342 21 372 47
rect 428 21 458 47
rect 514 21 544 47
rect 614 21 644 47
rect 700 21 730 47
rect 809 21 839 47
rect 895 21 925 47
rect 995 21 1025 47
rect 1095 21 1125 47
rect 1213 21 1243 47
rect 1299 21 1329 47
rect 1385 21 1415 47
rect 1485 21 1515 47
rect 1608 21 1638 47
<< polycont >>
rect 821 337 855 371
rect 979 329 1013 363
rect 224 269 258 303
rect 292 269 326 303
rect 360 269 394 303
rect 428 269 462 303
rect 496 269 530 303
rect 564 269 598 303
rect 632 269 666 303
rect 700 269 734 303
rect 1087 327 1121 361
rect 1195 327 1229 361
rect 1369 335 1403 369
rect 911 221 945 255
rect 1369 221 1403 255
rect 1489 253 1523 287
rect 1624 285 1658 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 23 607 73 649
rect 23 573 39 607
rect 23 503 73 573
rect 23 469 39 503
rect 23 409 73 469
rect 23 375 39 409
rect 23 359 73 375
rect 109 599 175 615
rect 109 565 125 599
rect 159 565 175 599
rect 109 506 175 565
rect 109 472 125 506
rect 159 472 175 506
rect 109 413 175 472
rect 211 607 245 649
rect 211 481 245 573
rect 211 431 245 447
rect 281 599 347 615
rect 281 565 297 599
rect 331 565 347 599
rect 281 506 347 565
rect 281 472 297 506
rect 331 472 347 506
rect 109 379 125 413
rect 159 397 175 413
rect 281 413 347 472
rect 383 607 417 649
rect 383 481 417 573
rect 383 431 417 447
rect 453 599 519 615
rect 453 565 469 599
rect 503 565 519 599
rect 453 506 519 565
rect 453 472 469 506
rect 503 472 519 506
rect 281 397 297 413
rect 159 379 297 397
rect 331 397 347 413
rect 453 413 519 472
rect 555 607 589 649
rect 555 481 589 573
rect 555 431 589 447
rect 625 599 675 615
rect 625 565 641 599
rect 625 506 675 565
rect 711 594 777 649
rect 711 560 727 594
rect 761 560 777 594
rect 711 532 777 560
rect 838 599 1104 615
rect 838 565 854 599
rect 888 581 1054 599
rect 888 565 904 581
rect 838 549 904 565
rect 1038 565 1054 581
rect 1088 565 1104 599
rect 1038 549 1104 565
rect 1138 606 1204 649
rect 1138 572 1154 606
rect 1188 572 1204 606
rect 1138 555 1204 572
rect 1238 594 1504 615
rect 1238 560 1254 594
rect 1288 590 1504 594
rect 1288 581 1454 590
rect 1288 560 1304 581
rect 1238 555 1304 560
rect 1438 556 1454 581
rect 1488 556 1504 590
rect 938 531 1004 547
rect 938 515 954 531
rect 625 472 641 506
rect 811 498 954 515
rect 453 397 469 413
rect 331 379 469 397
rect 503 397 519 413
rect 625 413 675 472
rect 625 397 641 413
rect 503 379 641 397
rect 109 363 675 379
rect 725 497 954 498
rect 988 515 1004 531
rect 1338 534 1404 547
rect 1338 521 1354 534
rect 1138 515 1354 521
rect 988 500 1354 515
rect 1388 500 1404 534
rect 1438 532 1504 556
rect 1549 594 1615 649
rect 1549 560 1565 594
rect 1599 560 1615 594
rect 1549 532 1615 560
rect 1651 599 1701 615
rect 1685 565 1701 599
rect 988 497 1404 500
rect 1651 509 1701 565
rect 725 487 1404 497
rect 725 481 1172 487
rect 725 464 845 481
rect 1473 475 1651 498
rect 1685 475 1701 509
rect 1473 464 1701 475
rect 23 207 75 223
rect 23 173 39 207
rect 73 173 75 207
rect 23 89 75 173
rect 23 55 39 89
rect 73 55 75 89
rect 109 219 175 363
rect 725 319 759 464
rect 1473 453 1507 464
rect 1206 447 1507 453
rect 879 430 1137 447
rect 793 424 1137 430
rect 793 413 1087 424
rect 793 396 913 413
rect 793 371 861 396
rect 1071 390 1087 413
rect 1121 390 1137 424
rect 793 337 821 371
rect 855 337 861 371
rect 963 363 1029 379
rect 793 321 861 337
rect 895 350 929 356
rect 224 303 759 319
rect 258 269 292 303
rect 326 269 360 303
rect 394 269 428 303
rect 462 269 496 303
rect 530 269 564 303
rect 598 269 632 303
rect 666 269 700 303
rect 734 287 759 303
rect 734 269 861 287
rect 224 253 861 269
rect 109 203 705 219
rect 109 169 125 203
rect 159 185 297 203
rect 159 169 175 185
rect 109 93 175 169
rect 281 169 297 185
rect 331 185 469 203
rect 331 169 347 185
rect 109 59 125 93
rect 159 59 175 93
rect 211 114 245 151
rect 23 17 75 55
rect 211 17 245 80
rect 281 93 347 169
rect 453 169 469 185
rect 503 185 655 203
rect 503 169 519 185
rect 281 59 297 93
rect 331 59 347 93
rect 383 114 417 151
rect 383 17 417 80
rect 453 93 519 169
rect 639 169 655 185
rect 689 169 705 203
rect 453 59 469 93
rect 503 59 519 93
rect 555 114 605 151
rect 589 80 605 114
rect 555 17 605 80
rect 639 93 705 169
rect 639 59 655 93
rect 689 59 705 93
rect 741 203 791 219
rect 775 169 791 203
rect 741 93 791 169
rect 827 171 861 253
rect 895 271 929 316
rect 963 329 979 363
rect 1013 329 1029 363
rect 963 313 1029 329
rect 895 255 961 271
rect 895 221 911 255
rect 945 221 961 255
rect 895 205 961 221
rect 995 239 1029 313
rect 1071 361 1137 390
rect 1071 327 1087 361
rect 1121 327 1137 361
rect 1071 311 1137 327
rect 1179 419 1507 447
rect 1179 361 1237 419
rect 1179 327 1195 361
rect 1229 327 1237 361
rect 1179 311 1237 327
rect 1271 369 1419 385
rect 1271 350 1369 369
rect 1271 316 1279 350
rect 1313 335 1369 350
rect 1403 335 1419 369
rect 1313 316 1419 335
rect 1271 313 1419 316
rect 1271 310 1319 313
rect 1473 303 1507 419
rect 1561 424 1607 430
rect 1561 390 1567 424
rect 1601 390 1607 424
rect 1561 384 1607 390
rect 1573 335 1607 384
rect 1651 419 1701 464
rect 1685 385 1701 419
rect 1651 369 1701 385
rect 1573 319 1674 335
rect 1473 287 1539 303
rect 1353 255 1419 279
rect 1353 239 1369 255
rect 995 221 1369 239
rect 1403 221 1419 255
rect 995 205 1419 221
rect 1473 253 1489 287
rect 1523 253 1539 287
rect 1573 285 1624 319
rect 1658 285 1674 319
rect 1573 269 1674 285
rect 1473 235 1539 253
rect 1473 203 1699 235
rect 1473 201 1649 203
rect 827 162 1390 171
rect 1633 169 1649 201
rect 1683 169 1699 203
rect 827 154 1340 162
rect 827 137 950 154
rect 934 120 950 137
rect 984 137 1340 154
rect 984 120 1000 137
rect 1324 128 1340 137
rect 1374 128 1390 162
rect 1324 127 1390 128
rect 934 119 1000 120
rect 1424 122 1490 167
rect 775 59 791 93
rect 741 17 791 59
rect 834 102 900 103
rect 834 68 850 102
rect 884 85 900 102
rect 1034 102 1100 103
rect 1034 85 1050 102
rect 884 68 1050 85
rect 1084 68 1100 102
rect 834 51 1100 68
rect 1136 87 1202 103
rect 1424 93 1440 122
rect 1136 53 1152 87
rect 1186 53 1202 87
rect 1238 59 1254 93
rect 1288 88 1440 93
rect 1474 88 1490 122
rect 1288 59 1490 88
rect 1533 122 1599 167
rect 1533 88 1549 122
rect 1583 88 1599 122
rect 1136 17 1202 53
rect 1533 17 1599 88
rect 1633 101 1699 169
rect 1633 67 1649 101
rect 1683 67 1699 101
rect 1633 51 1699 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1087 390 1121 424
rect 895 316 929 350
rect 1279 316 1313 350
rect 1567 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 1075 424 1133 430
rect 1075 390 1087 424
rect 1121 421 1133 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 1121 393 1567 421
rect 1121 390 1133 393
rect 1075 384 1133 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 883 350 941 356
rect 883 316 895 350
rect 929 347 941 350
rect 1267 350 1325 356
rect 1267 347 1279 350
rect 929 319 1279 347
rect 929 316 941 319
rect 883 310 941 316
rect 1267 316 1279 319
rect 1313 316 1325 350
rect 1267 310 1325 316
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2_8
flabel metal1 s 1087 390 1121 424 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel metal1 s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1732612
string GDS_START 1718754
<< end >>
