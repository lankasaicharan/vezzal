magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4178 1975
<< nwell >>
rect -38 331 2918 704
rect 2375 327 2695 331
<< pwell >>
rect 7 163 203 289
rect 1763 241 2662 251
rect 489 201 787 222
rect 1763 206 2879 241
rect 1371 201 2879 206
rect 489 163 2879 201
rect 7 49 2879 163
rect 0 0 2880 49
<< scnmos >>
rect 90 179 120 263
rect 288 53 318 137
rect 374 53 404 137
rect 572 112 602 196
rect 658 112 688 196
rect 880 91 910 175
rect 974 91 1004 175
rect 1067 91 1097 175
rect 1192 47 1222 175
rect 1477 96 1507 180
rect 1617 96 1647 180
rect 1846 141 1876 225
rect 1956 57 1986 225
rect 2038 57 2068 225
rect 2211 141 2241 225
rect 2433 141 2463 225
rect 2551 57 2581 225
rect 2768 47 2798 215
<< scpmoshvt >>
rect 90 481 120 609
rect 343 423 373 507
rect 429 423 459 507
rect 501 423 531 507
rect 587 423 617 507
rect 872 396 902 480
rect 958 396 988 480
rect 1150 457 1180 541
rect 1257 373 1287 541
rect 1449 396 1479 524
rect 1643 396 1673 524
rect 1835 367 1865 619
rect 1941 388 1971 472
rect 2133 367 2163 619
rect 2241 417 2271 501
rect 2465 363 2495 491
rect 2573 363 2603 615
rect 2769 367 2799 619
<< ndiff >>
rect 33 238 90 263
rect 33 204 45 238
rect 79 204 90 238
rect 33 179 90 204
rect 120 238 177 263
rect 120 204 131 238
rect 165 204 177 238
rect 120 179 177 204
rect 515 178 572 196
rect 515 144 527 178
rect 561 144 572 178
rect 231 114 288 137
rect 231 80 243 114
rect 277 80 288 114
rect 231 53 288 80
rect 318 112 374 137
rect 318 78 329 112
rect 363 78 374 112
rect 318 53 374 78
rect 404 108 461 137
rect 515 112 572 144
rect 602 178 658 196
rect 602 144 613 178
rect 647 144 658 178
rect 602 112 658 144
rect 688 163 761 196
rect 1789 200 1846 225
rect 688 129 715 163
rect 749 129 761 163
rect 688 112 761 129
rect 815 150 880 175
rect 815 116 827 150
rect 861 116 880 150
rect 404 74 415 108
rect 449 74 461 108
rect 815 91 880 116
rect 910 150 974 175
rect 910 116 929 150
rect 963 116 974 150
rect 910 91 974 116
rect 1004 91 1067 175
rect 1097 150 1192 175
rect 1097 116 1108 150
rect 1142 116 1192 150
rect 1097 91 1192 116
rect 404 53 461 74
rect 1142 47 1192 91
rect 1222 124 1279 175
rect 1222 90 1233 124
rect 1267 90 1279 124
rect 1397 155 1477 180
rect 1397 121 1409 155
rect 1443 121 1477 155
rect 1397 96 1477 121
rect 1507 155 1617 180
rect 1507 121 1556 155
rect 1590 121 1617 155
rect 1507 96 1617 121
rect 1647 155 1704 180
rect 1647 121 1658 155
rect 1692 121 1704 155
rect 1789 166 1801 200
rect 1835 166 1846 200
rect 1789 141 1846 166
rect 1876 141 1956 225
rect 1647 96 1704 121
rect 1898 115 1956 141
rect 1222 47 1279 90
rect 1898 81 1910 115
rect 1944 81 1956 115
rect 1898 57 1956 81
rect 1986 57 2038 225
rect 2068 141 2211 225
rect 2241 209 2318 225
rect 2241 175 2274 209
rect 2308 175 2318 209
rect 2241 141 2318 175
rect 2068 73 2148 141
rect 2378 213 2433 225
rect 2378 179 2388 213
rect 2422 179 2433 213
rect 2378 141 2433 179
rect 2463 141 2551 225
rect 2068 57 2102 73
rect 2090 39 2102 57
rect 2136 39 2148 73
rect 2478 73 2551 141
rect 2090 27 2148 39
rect 2478 39 2490 73
rect 2524 57 2551 73
rect 2581 213 2636 225
rect 2581 179 2592 213
rect 2626 179 2636 213
rect 2581 57 2636 179
rect 2690 73 2768 215
rect 2524 39 2536 57
rect 2478 27 2536 39
rect 2690 39 2700 73
rect 2734 47 2768 73
rect 2798 203 2853 215
rect 2798 169 2809 203
rect 2843 169 2853 203
rect 2798 103 2853 169
rect 2798 69 2809 103
rect 2843 69 2853 103
rect 2798 47 2853 69
rect 2734 39 2746 47
rect 2690 27 2746 39
<< pdiff >>
rect 33 597 90 609
rect 33 563 45 597
rect 79 563 90 597
rect 33 527 90 563
rect 33 493 45 527
rect 79 493 90 527
rect 33 481 90 493
rect 120 597 177 609
rect 120 563 131 597
rect 165 563 177 597
rect 120 527 177 563
rect 120 493 131 527
rect 165 493 177 527
rect 120 481 177 493
rect 286 482 343 507
rect 286 448 298 482
rect 332 448 343 482
rect 286 423 343 448
rect 373 482 429 507
rect 373 448 384 482
rect 418 448 429 482
rect 373 423 429 448
rect 459 423 501 507
rect 531 482 587 507
rect 531 448 542 482
rect 576 448 587 482
rect 531 423 587 448
rect 617 482 674 507
rect 617 448 628 482
rect 662 448 674 482
rect 1096 516 1150 541
rect 1096 482 1105 516
rect 1139 482 1150 516
rect 617 423 674 448
rect 761 455 872 480
rect 761 421 773 455
rect 807 421 872 455
rect 761 396 872 421
rect 902 449 958 480
rect 902 415 913 449
rect 947 415 958 449
rect 902 396 958 415
rect 988 455 1042 480
rect 1096 457 1150 482
rect 1180 496 1257 541
rect 1180 462 1212 496
rect 1246 462 1257 496
rect 1180 457 1257 462
rect 988 421 999 455
rect 1033 421 1042 455
rect 988 396 1042 421
rect 1202 373 1257 457
rect 1287 529 1341 541
rect 1287 495 1298 529
rect 1332 495 1341 529
rect 1781 607 1835 619
rect 1781 573 1790 607
rect 1824 573 1835 607
rect 1287 419 1341 495
rect 1287 385 1298 419
rect 1332 385 1341 419
rect 1395 512 1449 524
rect 1395 478 1404 512
rect 1438 478 1449 512
rect 1395 442 1449 478
rect 1395 408 1404 442
rect 1438 408 1449 442
rect 1395 396 1449 408
rect 1479 512 1643 524
rect 1479 478 1544 512
rect 1578 478 1643 512
rect 1479 396 1643 478
rect 1673 446 1727 524
rect 1673 412 1684 446
rect 1718 412 1727 446
rect 1673 396 1727 412
rect 1287 373 1341 385
rect 1781 367 1835 573
rect 1865 494 1919 619
rect 2079 594 2133 619
rect 2079 560 2088 594
rect 2122 560 2133 594
rect 1865 460 1876 494
rect 1910 472 1919 494
rect 1910 460 1941 472
rect 1865 388 1941 460
rect 1971 451 2025 472
rect 1971 417 1982 451
rect 2016 417 2025 451
rect 1971 388 2025 417
rect 1865 367 1919 388
rect 2079 367 2133 560
rect 2163 607 2219 619
rect 2163 573 2174 607
rect 2208 573 2219 607
rect 2163 501 2219 573
rect 2517 596 2573 615
rect 2517 562 2528 596
rect 2562 562 2573 596
rect 2163 417 2241 501
rect 2271 478 2357 501
rect 2517 491 2573 562
rect 2271 444 2314 478
rect 2348 444 2357 478
rect 2271 417 2357 444
rect 2163 367 2219 417
rect 2411 413 2465 491
rect 2411 379 2420 413
rect 2454 379 2465 413
rect 2411 363 2465 379
rect 2495 363 2573 491
rect 2603 417 2659 615
rect 2603 383 2614 417
rect 2648 383 2659 417
rect 2603 363 2659 383
rect 2713 598 2769 619
rect 2713 564 2724 598
rect 2758 564 2769 598
rect 2713 367 2769 564
rect 2799 597 2853 619
rect 2799 563 2810 597
rect 2844 563 2853 597
rect 2799 505 2853 563
rect 2799 471 2810 505
rect 2844 471 2853 505
rect 2799 413 2853 471
rect 2799 379 2810 413
rect 2844 379 2853 413
rect 2799 367 2853 379
<< ndiffc >>
rect 45 204 79 238
rect 131 204 165 238
rect 527 144 561 178
rect 243 80 277 114
rect 329 78 363 112
rect 613 144 647 178
rect 715 129 749 163
rect 827 116 861 150
rect 415 74 449 108
rect 929 116 963 150
rect 1108 116 1142 150
rect 1233 90 1267 124
rect 1409 121 1443 155
rect 1556 121 1590 155
rect 1658 121 1692 155
rect 1801 166 1835 200
rect 1910 81 1944 115
rect 2274 175 2308 209
rect 2388 179 2422 213
rect 2102 39 2136 73
rect 2490 39 2524 73
rect 2592 179 2626 213
rect 2700 39 2734 73
rect 2809 169 2843 203
rect 2809 69 2843 103
<< pdiffc >>
rect 45 563 79 597
rect 45 493 79 527
rect 131 563 165 597
rect 131 493 165 527
rect 298 448 332 482
rect 384 448 418 482
rect 542 448 576 482
rect 628 448 662 482
rect 1105 482 1139 516
rect 773 421 807 455
rect 913 415 947 449
rect 1212 462 1246 496
rect 999 421 1033 455
rect 1298 495 1332 529
rect 1790 573 1824 607
rect 1298 385 1332 419
rect 1404 478 1438 512
rect 1404 408 1438 442
rect 1544 478 1578 512
rect 1684 412 1718 446
rect 2088 560 2122 594
rect 1876 460 1910 494
rect 1982 417 2016 451
rect 2174 573 2208 607
rect 2528 562 2562 596
rect 2314 444 2348 478
rect 2420 379 2454 413
rect 2614 383 2648 417
rect 2724 564 2758 598
rect 2810 563 2844 597
rect 2810 471 2844 505
rect 2810 379 2844 413
<< poly >>
rect 90 609 120 635
rect 872 615 1673 645
rect 1835 619 1865 645
rect 2133 619 2163 645
rect 217 597 283 613
rect 217 563 233 597
rect 267 563 283 597
rect 217 547 283 563
rect 90 381 120 481
rect 217 401 247 547
rect 343 507 373 533
rect 429 507 459 533
rect 501 507 531 533
rect 587 507 617 533
rect 872 480 902 615
rect 1150 541 1180 567
rect 1257 541 1287 567
rect 958 480 988 506
rect 343 401 373 423
rect 217 381 373 401
rect 90 371 373 381
rect 90 351 318 371
rect 90 263 120 351
rect 90 153 120 179
rect 288 137 318 351
rect 429 313 459 423
rect 374 297 459 313
rect 374 263 390 297
rect 424 283 459 297
rect 501 302 531 423
rect 587 380 617 423
rect 587 350 764 380
rect 658 340 764 350
rect 658 306 714 340
rect 748 306 764 340
rect 872 354 902 396
rect 958 356 988 396
rect 1150 377 1180 457
rect 1097 361 1180 377
rect 1449 524 1479 550
rect 1643 524 1673 615
rect 872 324 910 354
rect 501 286 567 302
rect 424 263 440 283
rect 374 247 440 263
rect 501 252 517 286
rect 551 266 567 286
rect 658 290 764 306
rect 551 252 602 266
rect 374 137 404 247
rect 501 236 602 252
rect 572 196 602 236
rect 658 196 688 290
rect 880 175 910 324
rect 958 340 1049 356
rect 958 306 999 340
rect 1033 306 1049 340
rect 958 290 1049 306
rect 1097 327 1120 361
rect 1154 327 1180 361
rect 1097 311 1180 327
rect 974 175 1004 290
rect 1097 242 1127 311
rect 1257 263 1287 373
rect 1449 364 1479 396
rect 1449 334 1507 364
rect 1643 354 1673 396
rect 1941 472 1971 498
rect 1067 212 1127 242
rect 1192 247 1287 263
rect 1192 213 1210 247
rect 1244 213 1287 247
rect 1368 270 1434 286
rect 1368 236 1384 270
rect 1418 250 1434 270
rect 1477 250 1507 334
rect 1418 236 1507 250
rect 1368 220 1507 236
rect 1555 345 1673 354
rect 1835 345 1865 367
rect 1555 338 1876 345
rect 1555 304 1571 338
rect 1605 315 1876 338
rect 1941 315 1971 388
rect 2573 615 2603 641
rect 2769 619 2799 645
rect 2241 501 2271 527
rect 2465 491 2495 517
rect 2133 335 2163 367
rect 2241 349 2271 417
rect 2313 369 2379 385
rect 2313 349 2329 369
rect 2038 319 2163 335
rect 1605 304 1647 315
rect 1555 270 1647 304
rect 1555 236 1571 270
rect 1605 236 1647 270
rect 1555 220 1647 236
rect 1846 225 1876 315
rect 1924 299 1990 315
rect 1924 265 1940 299
rect 1974 265 1990 299
rect 1924 249 1990 265
rect 2038 285 2054 319
rect 2088 305 2163 319
rect 2211 335 2329 349
rect 2363 335 2379 369
rect 2211 319 2379 335
rect 2088 285 2104 305
rect 2038 269 2104 285
rect 1956 225 1986 249
rect 2038 225 2068 269
rect 2211 225 2241 319
rect 2465 277 2495 363
rect 2573 331 2603 363
rect 2333 247 2495 277
rect 2537 315 2603 331
rect 2537 281 2553 315
rect 2587 281 2603 315
rect 2769 303 2799 367
rect 2537 265 2603 281
rect 2708 287 2799 303
rect 1067 175 1097 212
rect 1192 197 1287 213
rect 1192 175 1222 197
rect 1477 180 1507 220
rect 1617 180 1647 220
rect 572 86 602 112
rect 658 86 688 112
rect 880 65 910 91
rect 974 65 1004 91
rect 1067 65 1097 91
rect 288 27 318 53
rect 374 27 404 53
rect 1846 115 1876 141
rect 1477 70 1507 96
rect 1617 70 1647 96
rect 2211 115 2241 141
rect 2333 119 2363 247
rect 2433 225 2463 247
rect 2551 225 2581 265
rect 2708 253 2724 287
rect 2758 253 2799 287
rect 2708 237 2799 253
rect 1192 21 1222 47
rect 1956 31 1986 57
rect 2038 31 2068 57
rect 2297 103 2363 119
rect 2433 115 2463 141
rect 2297 69 2313 103
rect 2347 69 2363 103
rect 2297 53 2363 69
rect 2768 215 2798 237
rect 2551 31 2581 57
rect 2768 21 2798 47
<< polycont >>
rect 233 563 267 597
rect 390 263 424 297
rect 714 306 748 340
rect 517 252 551 286
rect 999 306 1033 340
rect 1120 327 1154 361
rect 1210 213 1244 247
rect 1384 236 1418 270
rect 1571 304 1605 338
rect 1571 236 1605 270
rect 1940 265 1974 299
rect 2054 285 2088 319
rect 2329 335 2363 369
rect 2553 281 2587 315
rect 2724 253 2758 287
rect 2313 69 2347 103
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 29 597 79 649
rect 29 563 45 597
rect 29 527 79 563
rect 29 493 45 527
rect 29 477 79 493
rect 115 597 181 613
rect 115 563 131 597
rect 165 563 181 597
rect 115 527 181 563
rect 115 493 131 527
rect 165 493 181 527
rect 115 313 181 493
rect 217 597 283 613
rect 217 563 233 597
rect 267 563 283 597
rect 217 547 283 563
rect 217 384 262 547
rect 298 482 348 511
rect 332 448 348 482
rect 298 383 348 448
rect 384 482 418 649
rect 384 419 418 448
rect 454 547 662 581
rect 454 383 488 547
rect 298 349 488 383
rect 526 482 576 511
rect 526 448 542 482
rect 526 383 576 448
rect 612 482 662 547
rect 612 448 628 482
rect 612 419 662 448
rect 773 579 1155 613
rect 773 455 807 579
rect 698 424 737 430
rect 698 390 703 424
rect 773 392 807 421
rect 843 509 1049 543
rect 526 349 662 383
rect 115 297 440 313
rect 29 238 79 267
rect 29 204 45 238
rect 29 17 79 204
rect 115 263 390 297
rect 424 263 440 297
rect 115 247 440 263
rect 501 286 567 302
rect 501 252 517 286
rect 551 252 567 286
rect 115 238 181 247
rect 115 204 131 238
rect 165 204 181 238
rect 501 236 567 252
rect 628 254 662 349
rect 698 356 737 390
rect 698 340 764 356
rect 698 306 714 340
rect 748 306 764 340
rect 698 290 764 306
rect 843 254 877 509
rect 628 220 877 254
rect 115 175 181 204
rect 227 200 433 211
rect 628 200 663 220
rect 227 178 561 200
rect 227 177 527 178
rect 227 114 277 177
rect 399 166 527 177
rect 511 144 527 166
rect 227 80 243 114
rect 227 53 277 80
rect 313 112 363 141
rect 313 78 329 112
rect 313 17 363 78
rect 399 108 465 130
rect 511 123 561 144
rect 597 178 663 200
rect 597 144 613 178
rect 647 144 663 178
rect 597 123 663 144
rect 699 163 765 184
rect 699 129 715 163
rect 749 129 765 163
rect 399 74 415 108
rect 449 87 465 108
rect 699 87 765 129
rect 811 150 877 220
rect 811 116 827 150
rect 861 116 877 150
rect 811 87 877 116
rect 913 449 947 473
rect 913 249 947 415
rect 983 455 1049 509
rect 983 421 999 455
rect 1033 421 1049 455
rect 1089 516 1155 579
rect 1089 482 1105 516
rect 1139 482 1155 516
rect 1089 453 1155 482
rect 1196 496 1246 649
rect 1196 462 1212 496
rect 983 392 1049 421
rect 1196 413 1246 462
rect 1282 564 1508 598
rect 1282 529 1332 564
rect 1282 495 1298 529
rect 1282 419 1332 495
rect 1282 385 1298 419
rect 1282 377 1332 385
rect 1104 361 1332 377
rect 983 350 1049 356
rect 983 316 991 350
rect 1025 340 1049 350
rect 983 306 999 316
rect 1033 306 1049 340
rect 1104 327 1120 361
rect 1154 327 1332 361
rect 1104 311 1332 327
rect 1388 512 1438 528
rect 1388 478 1404 512
rect 1388 442 1438 478
rect 1388 408 1404 442
rect 1388 356 1438 408
rect 1474 426 1508 564
rect 1544 512 1578 649
rect 1774 607 2138 613
rect 1774 573 1790 607
rect 1824 594 2138 607
rect 1824 573 2088 594
rect 2072 560 2088 573
rect 2122 560 2138 594
rect 2072 557 2138 560
rect 2174 607 2208 649
rect 2512 596 2578 649
rect 2174 557 2208 573
rect 2244 541 2476 575
rect 1544 462 1578 478
rect 1614 503 1824 537
rect 1614 426 1648 503
rect 1474 392 1648 426
rect 1684 446 1734 467
rect 1718 412 1734 446
rect 1684 356 1734 412
rect 1388 322 1504 356
rect 983 290 1049 306
rect 1194 249 1260 263
rect 913 247 1260 249
rect 913 215 1210 247
rect 913 150 979 215
rect 1194 213 1210 215
rect 1244 213 1260 247
rect 1194 197 1260 213
rect 913 116 929 150
rect 963 116 979 150
rect 913 87 979 116
rect 1092 150 1158 179
rect 1298 161 1332 311
rect 1368 270 1434 286
rect 1368 236 1384 270
rect 1418 236 1434 270
rect 1368 220 1434 236
rect 1470 254 1504 322
rect 1555 338 1621 354
rect 1555 304 1571 338
rect 1605 304 1621 338
rect 1555 270 1621 304
rect 1555 254 1571 270
rect 1470 236 1571 254
rect 1605 236 1621 270
rect 1470 220 1621 236
rect 1657 350 1734 356
rect 1657 316 1663 350
rect 1697 316 1734 350
rect 1790 381 1824 503
rect 1860 521 1926 537
rect 2244 521 2278 541
rect 1860 494 2278 521
rect 1860 460 1876 494
rect 1910 487 2278 494
rect 1910 460 1926 487
rect 1860 417 1926 460
rect 2314 478 2364 505
rect 1966 417 1982 451
rect 2016 444 2314 451
rect 2348 444 2364 478
rect 2442 503 2476 541
rect 2512 562 2528 596
rect 2562 562 2578 596
rect 2512 539 2578 562
rect 2708 598 2774 649
rect 2708 564 2724 598
rect 2758 564 2774 598
rect 2708 539 2774 564
rect 2810 597 2860 613
rect 2844 563 2860 597
rect 2810 505 2860 563
rect 2442 469 2773 503
rect 2016 417 2364 444
rect 2404 424 2471 433
rect 2404 413 2431 424
rect 2404 381 2420 413
rect 2465 390 2471 424
rect 1790 347 2104 381
rect 1657 311 1734 316
rect 2038 319 2104 347
rect 2313 379 2420 381
rect 2454 379 2471 390
rect 2313 369 2471 379
rect 2313 335 2329 369
rect 2363 335 2471 369
rect 2521 417 2672 433
rect 2521 383 2614 417
rect 2648 383 2672 417
rect 2521 367 2672 383
rect 2313 331 2471 335
rect 2313 319 2602 331
rect 1657 299 1990 311
rect 1657 277 1940 299
rect 1470 184 1504 220
rect 1657 184 1708 277
rect 1924 265 1940 277
rect 1974 265 1990 299
rect 2038 285 2054 319
rect 2088 285 2104 319
rect 2038 269 2104 285
rect 2372 315 2602 319
rect 2372 281 2553 315
rect 2587 281 2602 315
rect 1924 249 1990 265
rect 2372 265 2602 281
rect 1092 116 1108 150
rect 1142 116 1158 150
rect 449 74 765 87
rect 399 53 765 74
rect 1092 17 1158 116
rect 1217 124 1332 161
rect 1217 90 1233 124
rect 1267 90 1332 124
rect 1393 155 1504 184
rect 1393 121 1409 155
rect 1443 150 1504 155
rect 1540 155 1606 184
rect 1443 121 1459 150
rect 1393 108 1459 121
rect 1540 121 1556 155
rect 1590 121 1606 155
rect 1217 53 1332 90
rect 1540 17 1606 121
rect 1642 155 1708 184
rect 1642 121 1658 155
rect 1692 121 1708 155
rect 1785 213 1851 229
rect 2258 213 2324 229
rect 1785 209 2324 213
rect 1785 200 2274 209
rect 1785 166 1801 200
rect 1835 179 2274 200
rect 1835 166 1851 179
rect 1785 137 1851 166
rect 2258 175 2274 179
rect 2308 175 2324 209
rect 2372 213 2438 265
rect 2638 229 2672 367
rect 2372 179 2388 213
rect 2422 179 2438 213
rect 2576 213 2672 229
rect 2576 179 2592 213
rect 2626 179 2672 213
rect 2708 287 2773 469
rect 2844 471 2860 505
rect 2810 430 2860 471
rect 2708 253 2724 287
rect 2758 253 2773 287
rect 2258 155 2324 175
rect 2708 143 2773 253
rect 1642 92 1708 121
rect 1894 119 2222 143
rect 2360 119 2773 143
rect 1894 115 2773 119
rect 1894 81 1910 115
rect 1944 109 2773 115
rect 2809 413 2860 430
rect 2809 379 2810 413
rect 2844 379 2860 413
rect 2809 203 2860 379
rect 2843 169 2860 203
rect 1944 81 1960 109
rect 1894 53 1960 81
rect 2188 103 2394 109
rect 2086 39 2102 73
rect 2136 39 2152 73
rect 2188 69 2313 103
rect 2347 69 2394 103
rect 2809 103 2860 169
rect 2188 53 2394 69
rect 2086 17 2152 39
rect 2474 39 2490 73
rect 2524 39 2540 73
rect 2474 17 2540 39
rect 2684 39 2700 73
rect 2734 39 2750 73
rect 2843 69 2860 103
rect 2809 53 2860 69
rect 2684 17 2750 39
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 703 390 737 424
rect 991 340 1025 350
rect 991 316 999 340
rect 999 316 1025 340
rect 1663 316 1697 350
rect 2431 413 2465 424
rect 2431 390 2454 413
rect 2454 390 2465 413
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
<< metal1 >>
rect 0 683 2880 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2880 683
rect 0 617 2880 649
rect 691 424 749 430
rect 691 390 703 424
rect 737 421 749 424
rect 2419 424 2477 430
rect 2419 421 2431 424
rect 737 393 2431 421
rect 737 390 749 393
rect 691 384 749 390
rect 2419 390 2431 393
rect 2465 390 2477 424
rect 2419 384 2477 390
rect 979 350 1037 356
rect 979 316 991 350
rect 1025 347 1037 350
rect 1651 350 1709 356
rect 1651 347 1663 350
rect 1025 319 1663 347
rect 1025 316 1037 319
rect 979 310 1037 316
rect 1651 316 1663 319
rect 1697 316 1709 350
rect 1651 310 1709 316
rect 0 17 2880 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2880 17
rect 0 -49 2880 -17
<< labels >>
flabel pwell s 0 0 2880 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2880 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 edfxbp_1
flabel metal1 s 0 617 2880 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2880 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2815 94 2849 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2815 168 2849 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2815 242 2849 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2815 316 2849 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2815 390 2849 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 DE
port 3 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 DE
port 3 nsew signal input
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 DE
port 3 nsew signal input
flabel locali s 2527 390 2561 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2623 390 2657 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2880 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3124154
string GDS_START 3104926
<< end >>
