magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 383 231 1049 241
rect 19 49 1049 231
rect 0 0 1056 49
<< scnmos >>
rect 98 121 128 205
rect 184 121 214 205
rect 270 121 300 205
rect 462 131 492 215
rect 534 131 564 215
rect 651 47 681 215
rect 737 47 767 215
rect 854 47 884 215
rect 940 47 970 215
<< scpmoshvt >>
rect 125 397 155 525
rect 197 397 227 525
rect 305 397 335 525
rect 460 397 490 525
rect 546 397 576 525
rect 651 367 681 619
rect 737 367 767 619
rect 823 367 853 619
rect 909 367 939 619
<< ndiff >>
rect 45 180 98 205
rect 45 146 53 180
rect 87 146 98 180
rect 45 121 98 146
rect 128 165 184 205
rect 128 131 139 165
rect 173 131 184 165
rect 128 121 184 131
rect 214 180 270 205
rect 214 146 225 180
rect 259 146 270 180
rect 214 121 270 146
rect 300 180 353 205
rect 300 146 311 180
rect 345 146 353 180
rect 300 121 353 146
rect 409 190 462 215
rect 409 156 417 190
rect 451 156 462 190
rect 409 131 462 156
rect 492 131 534 215
rect 564 194 651 215
rect 564 160 575 194
rect 609 160 651 194
rect 564 131 651 160
rect 598 97 651 131
rect 598 63 606 97
rect 640 63 651 97
rect 598 47 651 63
rect 681 187 737 215
rect 681 153 692 187
rect 726 153 737 187
rect 681 101 737 153
rect 681 67 692 101
rect 726 67 737 101
rect 681 47 737 67
rect 767 203 854 215
rect 767 169 795 203
rect 829 169 854 203
rect 767 93 854 169
rect 767 59 795 93
rect 829 59 854 93
rect 767 47 854 59
rect 884 207 940 215
rect 884 173 895 207
rect 929 173 940 207
rect 884 101 940 173
rect 884 67 895 101
rect 929 67 940 101
rect 884 47 940 67
rect 970 203 1023 215
rect 970 169 981 203
rect 1015 169 1023 203
rect 970 93 1023 169
rect 970 59 981 93
rect 1015 59 1023 93
rect 970 47 1023 59
<< pdiff >>
rect 598 601 651 619
rect 598 567 606 601
rect 640 567 651 601
rect 598 525 651 567
rect 72 513 125 525
rect 72 479 80 513
rect 114 479 125 513
rect 72 445 125 479
rect 72 411 80 445
rect 114 411 125 445
rect 72 397 125 411
rect 155 397 197 525
rect 227 511 305 525
rect 227 477 238 511
rect 272 477 305 511
rect 227 443 305 477
rect 227 409 238 443
rect 272 409 305 443
rect 227 397 305 409
rect 335 501 460 525
rect 335 467 361 501
rect 395 467 460 501
rect 335 397 460 467
rect 490 445 546 525
rect 490 411 501 445
rect 535 411 546 445
rect 490 397 546 411
rect 576 397 651 525
rect 598 367 651 397
rect 681 445 737 619
rect 681 411 692 445
rect 726 411 737 445
rect 681 367 737 411
rect 767 601 823 619
rect 767 567 778 601
rect 812 567 823 601
rect 767 367 823 567
rect 853 599 909 619
rect 853 565 864 599
rect 898 565 909 599
rect 853 499 909 565
rect 853 465 864 499
rect 898 465 909 499
rect 853 413 909 465
rect 853 379 864 413
rect 898 379 909 413
rect 853 367 909 379
rect 939 607 1007 619
rect 939 573 963 607
rect 997 573 1007 607
rect 939 505 1007 573
rect 939 471 963 505
rect 997 471 1007 505
rect 939 413 1007 471
rect 939 379 963 413
rect 997 379 1007 413
rect 939 367 1007 379
<< ndiffc >>
rect 53 146 87 180
rect 139 131 173 165
rect 225 146 259 180
rect 311 146 345 180
rect 417 156 451 190
rect 575 160 609 194
rect 606 63 640 97
rect 692 153 726 187
rect 692 67 726 101
rect 795 169 829 203
rect 795 59 829 93
rect 895 173 929 207
rect 895 67 929 101
rect 981 169 1015 203
rect 981 59 1015 93
<< pdiffc >>
rect 606 567 640 601
rect 80 479 114 513
rect 80 411 114 445
rect 238 477 272 511
rect 238 409 272 443
rect 361 467 395 501
rect 501 411 535 445
rect 692 411 726 445
rect 778 567 812 601
rect 864 565 898 599
rect 864 465 898 499
rect 864 379 898 413
rect 963 573 997 607
rect 963 471 997 505
rect 963 379 997 413
<< poly >>
rect 125 599 576 629
rect 651 619 681 645
rect 737 619 767 645
rect 823 619 853 645
rect 909 619 939 645
rect 125 525 155 599
rect 197 525 227 551
rect 305 525 335 551
rect 460 525 490 551
rect 546 525 576 599
rect 125 365 155 397
rect 70 349 155 365
rect 70 315 86 349
rect 120 335 155 349
rect 197 365 227 397
rect 197 349 263 365
rect 120 315 136 335
rect 70 299 136 315
rect 197 315 213 349
rect 247 315 263 349
rect 197 299 263 315
rect 305 303 335 397
rect 460 375 490 397
rect 546 375 576 397
rect 460 345 492 375
rect 98 205 128 299
rect 197 257 228 299
rect 305 287 420 303
rect 305 257 370 287
rect 184 227 228 257
rect 270 253 370 257
rect 404 253 420 287
rect 270 237 420 253
rect 270 227 336 237
rect 184 205 214 227
rect 270 205 300 227
rect 462 215 492 345
rect 534 345 576 375
rect 534 215 564 345
rect 651 303 681 367
rect 606 287 681 303
rect 606 253 622 287
rect 656 267 681 287
rect 737 267 767 367
rect 823 303 853 367
rect 909 303 939 367
rect 656 253 767 267
rect 606 237 767 253
rect 809 287 970 303
rect 809 253 825 287
rect 859 273 970 287
rect 859 253 884 273
rect 809 237 884 253
rect 651 215 681 237
rect 737 215 767 237
rect 854 215 884 237
rect 940 215 970 273
rect 98 95 128 121
rect 184 53 214 121
rect 270 95 300 121
rect 462 53 492 131
rect 534 105 564 131
rect 184 23 492 53
rect 651 21 681 47
rect 737 21 767 47
rect 854 21 884 47
rect 940 21 970 47
<< polycont >>
rect 86 315 120 349
rect 213 315 247 349
rect 370 253 404 287
rect 622 253 656 287
rect 825 253 859 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 64 513 130 649
rect 64 479 80 513
rect 114 479 130 513
rect 64 445 130 479
rect 64 411 80 445
rect 114 411 130 445
rect 64 395 130 411
rect 222 511 278 527
rect 222 477 238 511
rect 272 477 278 511
rect 222 443 278 477
rect 356 501 399 649
rect 590 601 656 649
rect 590 567 606 601
rect 640 567 656 601
rect 590 563 656 567
rect 762 601 828 649
rect 762 567 778 601
rect 812 567 828 601
rect 762 563 828 567
rect 862 599 929 615
rect 862 565 864 599
rect 898 565 929 599
rect 356 467 361 501
rect 395 467 399 501
rect 356 451 399 467
rect 433 495 828 529
rect 222 409 238 443
rect 272 427 278 443
rect 272 409 331 427
rect 222 393 331 409
rect 297 371 331 393
rect 433 371 467 495
rect 17 349 163 361
rect 17 315 86 349
rect 120 315 163 349
rect 17 299 163 315
rect 197 349 263 359
rect 197 315 213 349
rect 247 315 263 349
rect 197 299 263 315
rect 297 337 467 371
rect 501 445 539 461
rect 535 411 539 445
rect 37 215 263 249
rect 37 180 103 215
rect 37 146 53 180
rect 87 146 103 180
rect 37 130 103 146
rect 137 165 187 181
rect 137 131 139 165
rect 173 131 187 165
rect 137 17 187 131
rect 221 180 263 215
rect 221 146 225 180
rect 259 146 263 180
rect 221 130 263 146
rect 297 196 332 337
rect 501 303 539 411
rect 690 445 745 461
rect 690 411 692 445
rect 726 411 745 445
rect 368 287 656 303
rect 368 253 370 287
rect 404 253 622 287
rect 368 237 656 253
rect 368 230 467 237
rect 297 180 361 196
rect 297 146 311 180
rect 345 146 361 180
rect 297 130 361 146
rect 395 190 467 230
rect 690 203 745 411
rect 794 303 828 495
rect 862 499 929 565
rect 862 465 864 499
rect 898 465 929 499
rect 862 413 929 465
rect 862 379 864 413
rect 898 379 929 413
rect 862 339 929 379
rect 963 607 1003 649
rect 997 573 1003 607
rect 963 505 1003 573
rect 997 471 1003 505
rect 963 413 1003 471
rect 997 379 1003 413
rect 963 363 1003 379
rect 794 287 859 303
rect 794 253 825 287
rect 794 237 859 253
rect 893 207 929 339
rect 395 156 417 190
rect 451 156 467 190
rect 395 140 467 156
rect 559 194 644 203
rect 559 160 575 194
rect 609 160 644 194
rect 559 97 644 160
rect 559 63 606 97
rect 640 63 644 97
rect 559 17 644 63
rect 678 187 745 203
rect 678 153 692 187
rect 726 153 745 187
rect 678 101 745 153
rect 678 67 692 101
rect 726 67 745 101
rect 678 51 745 67
rect 779 169 795 203
rect 829 169 845 203
rect 779 93 845 169
rect 779 59 795 93
rect 829 59 845 93
rect 779 17 845 59
rect 893 173 895 207
rect 893 101 929 173
rect 893 67 895 101
rect 893 51 929 67
rect 965 203 1031 219
rect 965 169 981 203
rect 1015 169 1031 203
rect 965 93 1031 169
rect 965 59 981 93
rect 1015 59 1031 93
rect 965 17 1031 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ha_2
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 895 94 929 128 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 895 464 929 498 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 895 538 929 572 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6731474
string GDS_START 6722334
<< end >>
