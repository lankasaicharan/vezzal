magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 5 157 384 241
rect 5 49 767 157
rect 0 0 768 49
<< scnmos >>
rect 84 131 114 215
rect 189 47 219 215
rect 275 47 305 215
rect 380 47 410 131
rect 466 47 496 131
rect 572 47 602 131
rect 658 47 688 131
<< scpmoshvt >>
rect 84 367 114 451
rect 189 367 219 619
rect 275 367 305 619
rect 406 385 436 469
rect 478 385 508 469
rect 586 385 616 469
rect 658 385 688 469
<< ndiff >>
rect 31 190 84 215
rect 31 156 39 190
rect 73 156 84 190
rect 31 131 84 156
rect 114 163 189 215
rect 114 131 144 163
rect 136 129 144 131
rect 178 129 189 163
rect 136 93 189 129
rect 136 59 144 93
rect 178 59 189 93
rect 136 47 189 59
rect 219 203 275 215
rect 219 169 230 203
rect 264 169 275 203
rect 219 101 275 169
rect 219 67 230 101
rect 264 67 275 101
rect 219 47 275 67
rect 305 167 358 215
rect 305 133 316 167
rect 350 133 358 167
rect 305 131 358 133
rect 305 93 380 131
rect 305 59 335 93
rect 369 59 380 93
rect 305 47 380 59
rect 410 106 466 131
rect 410 72 421 106
rect 455 72 466 106
rect 410 47 466 72
rect 496 106 572 131
rect 496 72 513 106
rect 547 72 572 106
rect 496 47 572 72
rect 602 106 658 131
rect 602 72 613 106
rect 647 72 658 106
rect 602 47 658 72
rect 688 95 741 131
rect 688 61 699 95
rect 733 61 741 95
rect 688 47 741 61
<< pdiff >>
rect 136 577 189 619
rect 136 543 144 577
rect 178 543 189 577
rect 136 451 189 543
rect 31 426 84 451
rect 31 392 39 426
rect 73 392 84 426
rect 31 367 84 392
rect 114 367 189 451
rect 219 419 275 619
rect 219 385 230 419
rect 264 385 275 419
rect 219 367 275 385
rect 305 577 358 619
rect 305 543 316 577
rect 350 543 358 577
rect 305 469 358 543
rect 305 385 406 469
rect 436 385 478 469
rect 508 385 586 469
rect 616 385 658 469
rect 688 431 741 469
rect 688 397 699 431
rect 733 397 741 431
rect 688 385 741 397
rect 305 367 358 385
<< ndiffc >>
rect 39 156 73 190
rect 144 129 178 163
rect 144 59 178 93
rect 230 169 264 203
rect 230 67 264 101
rect 316 133 350 167
rect 335 59 369 93
rect 421 72 455 106
rect 513 72 547 106
rect 613 72 647 106
rect 699 61 733 95
<< pdiffc >>
rect 144 543 178 577
rect 39 392 73 426
rect 230 385 264 419
rect 316 543 350 577
rect 699 397 733 431
<< poly >>
rect 189 619 219 645
rect 275 619 305 645
rect 84 451 114 477
rect 620 593 688 609
rect 620 559 636 593
rect 670 559 688 593
rect 620 543 688 559
rect 406 469 436 495
rect 478 469 508 495
rect 586 469 616 495
rect 658 469 688 543
rect 84 325 114 367
rect 30 309 114 325
rect 30 275 46 309
rect 80 275 114 309
rect 30 259 114 275
rect 84 215 114 259
rect 189 333 219 367
rect 275 333 305 367
rect 406 335 436 385
rect 189 317 322 333
rect 189 283 272 317
rect 306 283 322 317
rect 189 267 322 283
rect 370 319 436 335
rect 370 285 386 319
rect 420 285 436 319
rect 370 269 436 285
rect 478 297 508 385
rect 478 281 544 297
rect 189 215 219 267
rect 275 215 305 267
rect 84 105 114 131
rect 380 131 410 269
rect 478 247 494 281
rect 528 247 544 281
rect 478 231 544 247
rect 586 291 616 385
rect 658 363 688 385
rect 658 333 730 363
rect 586 275 652 291
rect 586 241 602 275
rect 636 241 652 275
rect 478 221 508 231
rect 466 191 508 221
rect 586 225 652 241
rect 466 131 496 191
rect 586 183 616 225
rect 700 183 730 333
rect 572 153 616 183
rect 658 153 730 183
rect 572 131 602 153
rect 658 131 688 153
rect 189 21 219 47
rect 275 21 305 47
rect 380 21 410 47
rect 466 21 496 47
rect 572 21 602 47
rect 658 21 688 47
<< polycont >>
rect 636 559 670 593
rect 46 275 80 309
rect 272 283 306 317
rect 386 285 420 319
rect 494 247 528 281
rect 602 241 636 275
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 128 577 194 649
rect 128 543 144 577
rect 178 543 194 577
rect 128 539 194 543
rect 300 577 366 649
rect 300 543 316 577
rect 350 543 366 577
rect 300 539 366 543
rect 620 593 688 609
rect 620 559 636 593
rect 670 559 688 593
rect 620 505 688 559
rect 132 471 688 505
rect 132 452 166 471
rect 23 426 166 452
rect 23 392 39 426
rect 73 392 166 426
rect 23 384 166 392
rect 17 309 96 350
rect 17 275 46 309
rect 80 275 96 309
rect 130 231 166 384
rect 23 197 166 231
rect 202 419 264 437
rect 202 385 230 419
rect 202 369 264 385
rect 300 431 749 437
rect 300 401 699 431
rect 202 231 236 369
rect 300 333 334 401
rect 683 397 699 401
rect 733 397 749 431
rect 270 317 334 333
rect 270 283 272 317
rect 306 283 334 317
rect 270 267 334 283
rect 370 319 455 367
rect 370 285 386 319
rect 420 285 455 319
rect 370 269 455 285
rect 489 281 553 367
rect 300 235 334 267
rect 489 247 494 281
rect 528 247 553 281
rect 202 203 266 231
rect 202 197 230 203
rect 23 190 89 197
rect 23 156 39 190
rect 73 156 89 190
rect 228 169 230 197
rect 264 169 266 203
rect 300 201 455 235
rect 23 140 89 156
rect 128 129 144 163
rect 178 129 194 163
rect 128 93 194 129
rect 128 59 144 93
rect 178 59 194 93
rect 128 17 194 59
rect 228 101 266 169
rect 228 67 230 101
rect 264 67 266 101
rect 228 51 266 67
rect 300 133 316 167
rect 350 133 378 167
rect 300 93 378 133
rect 300 59 335 93
rect 369 59 378 93
rect 300 17 378 59
rect 412 106 455 201
rect 489 168 553 247
rect 587 275 649 367
rect 587 241 602 275
rect 636 241 649 275
rect 587 225 649 241
rect 683 179 749 397
rect 597 145 749 179
rect 412 72 421 106
rect 412 56 455 72
rect 491 106 563 122
rect 491 72 513 106
rect 547 72 563 106
rect 491 17 563 72
rect 597 106 663 145
rect 597 72 613 106
rect 647 72 663 106
rect 597 51 663 72
rect 697 95 749 111
rect 697 61 699 95
rect 733 61 749 95
rect 697 17 749 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or4b_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2932782
string GDS_START 2925920
<< end >>
