magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 1109 157 1535 167
rect 1 49 1535 157
rect 0 0 1536 49
<< scnmos >>
rect 84 47 114 131
rect 156 47 186 131
rect 242 47 272 131
rect 320 47 350 131
rect 524 47 554 131
rect 596 47 626 131
rect 682 47 712 131
rect 760 47 790 131
rect 868 47 898 131
rect 982 47 1012 131
rect 1192 57 1222 141
rect 1264 57 1294 141
rect 1350 57 1380 141
rect 1422 57 1452 141
<< scpmoshvt >>
rect 108 415 158 615
rect 214 415 264 615
rect 456 415 506 615
rect 596 415 646 615
rect 694 415 744 615
rect 851 415 901 615
rect 949 415 999 615
rect 1128 415 1178 615
rect 1234 415 1284 615
rect 1361 415 1411 615
<< ndiff >>
rect 27 111 84 131
rect 27 77 39 111
rect 73 77 84 111
rect 27 47 84 77
rect 114 47 156 131
rect 186 106 242 131
rect 186 72 197 106
rect 231 72 242 106
rect 186 47 242 72
rect 272 47 320 131
rect 350 95 407 131
rect 350 61 361 95
rect 395 61 407 95
rect 350 47 407 61
rect 467 111 524 131
rect 467 77 479 111
rect 513 77 524 111
rect 467 47 524 77
rect 554 47 596 131
rect 626 95 682 131
rect 626 61 637 95
rect 671 61 682 95
rect 626 47 682 61
rect 712 47 760 131
rect 790 95 868 131
rect 790 61 823 95
rect 857 61 868 95
rect 790 47 868 61
rect 898 47 982 131
rect 1012 106 1081 131
rect 1012 72 1035 106
rect 1069 72 1081 106
rect 1012 47 1081 72
rect 1135 116 1192 141
rect 1135 82 1147 116
rect 1181 82 1192 116
rect 1135 57 1192 82
rect 1222 57 1264 141
rect 1294 111 1350 141
rect 1294 77 1305 111
rect 1339 77 1350 111
rect 1294 57 1350 77
rect 1380 57 1422 141
rect 1452 116 1509 141
rect 1452 82 1463 116
rect 1497 82 1509 116
rect 1452 57 1509 82
<< pdiff >>
rect 51 597 108 615
rect 51 563 63 597
rect 97 563 108 597
rect 51 529 108 563
rect 51 495 63 529
rect 97 495 108 529
rect 51 461 108 495
rect 51 427 63 461
rect 97 427 108 461
rect 51 415 108 427
rect 158 603 214 615
rect 158 569 169 603
rect 203 569 214 603
rect 158 415 214 569
rect 264 462 321 615
rect 264 428 275 462
rect 309 428 321 462
rect 264 415 321 428
rect 399 471 456 615
rect 399 437 411 471
rect 445 437 456 471
rect 399 415 456 437
rect 506 603 596 615
rect 506 569 551 603
rect 585 569 596 603
rect 506 469 596 569
rect 506 435 551 469
rect 585 435 596 469
rect 506 415 596 435
rect 646 415 694 615
rect 744 597 851 615
rect 744 563 806 597
rect 840 563 851 597
rect 744 529 851 563
rect 744 495 806 529
rect 840 495 851 529
rect 744 461 851 495
rect 744 427 806 461
rect 840 427 851 461
rect 744 415 851 427
rect 901 415 949 615
rect 999 603 1128 615
rect 999 569 1051 603
rect 1085 569 1128 603
rect 999 532 1128 569
rect 999 498 1051 532
rect 1085 498 1128 532
rect 999 461 1128 498
rect 999 427 1051 461
rect 1085 427 1128 461
rect 999 415 1128 427
rect 1178 597 1234 615
rect 1178 563 1189 597
rect 1223 563 1234 597
rect 1178 529 1234 563
rect 1178 495 1189 529
rect 1223 495 1234 529
rect 1178 461 1234 495
rect 1178 427 1189 461
rect 1223 427 1234 461
rect 1178 415 1234 427
rect 1284 603 1361 615
rect 1284 569 1295 603
rect 1329 569 1361 603
rect 1284 531 1361 569
rect 1284 497 1295 531
rect 1329 497 1361 531
rect 1284 415 1361 497
rect 1411 597 1468 615
rect 1411 563 1422 597
rect 1456 563 1468 597
rect 1411 529 1468 563
rect 1411 495 1422 529
rect 1456 495 1468 529
rect 1411 461 1468 495
rect 1411 427 1422 461
rect 1456 427 1468 461
rect 1411 415 1468 427
<< ndiffc >>
rect 39 77 73 111
rect 197 72 231 106
rect 361 61 395 95
rect 479 77 513 111
rect 637 61 671 95
rect 823 61 857 95
rect 1035 72 1069 106
rect 1147 82 1181 116
rect 1305 77 1339 111
rect 1463 82 1497 116
<< pdiffc >>
rect 63 563 97 597
rect 63 495 97 529
rect 63 427 97 461
rect 169 569 203 603
rect 275 428 309 462
rect 411 437 445 471
rect 551 569 585 603
rect 551 435 585 469
rect 806 563 840 597
rect 806 495 840 529
rect 806 427 840 461
rect 1051 569 1085 603
rect 1051 498 1085 532
rect 1051 427 1085 461
rect 1189 563 1223 597
rect 1189 495 1223 529
rect 1189 427 1223 461
rect 1295 569 1329 603
rect 1295 497 1329 531
rect 1422 563 1456 597
rect 1422 495 1456 529
rect 1422 427 1456 461
<< poly >>
rect 108 615 158 641
rect 214 615 264 641
rect 456 615 506 641
rect 596 615 646 641
rect 694 615 744 641
rect 851 615 901 641
rect 949 615 999 641
rect 1128 615 1178 641
rect 1234 615 1284 641
rect 1361 615 1411 641
rect 108 356 158 415
rect 214 358 264 415
rect 314 367 380 383
rect 84 340 158 356
rect 84 306 108 340
rect 142 306 158 340
rect 84 272 158 306
rect 84 238 108 272
rect 142 238 158 272
rect 84 222 158 238
rect 206 342 272 358
rect 206 308 222 342
rect 256 308 272 342
rect 314 333 330 367
rect 364 347 380 367
rect 456 347 506 415
rect 596 383 646 415
rect 694 383 744 415
rect 364 333 506 347
rect 314 317 506 333
rect 580 367 646 383
rect 580 333 596 367
rect 630 333 646 367
rect 580 317 646 333
rect 688 367 754 383
rect 688 333 704 367
rect 738 333 754 367
rect 851 365 901 415
rect 688 317 754 333
rect 796 335 901 365
rect 949 365 999 415
rect 949 335 1012 365
rect 1128 351 1178 415
rect 1234 375 1284 415
rect 1234 359 1300 375
rect 206 274 272 308
rect 206 240 222 274
rect 256 254 272 274
rect 476 269 506 317
rect 616 269 646 317
rect 796 269 826 335
rect 256 240 350 254
rect 206 224 350 240
rect 84 176 114 222
rect 84 146 186 176
rect 84 131 114 146
rect 156 131 186 146
rect 242 131 272 224
rect 320 131 350 224
rect 476 253 554 269
rect 476 219 504 253
rect 538 219 554 253
rect 616 239 712 269
rect 476 203 554 219
rect 524 191 554 203
rect 524 161 626 191
rect 524 131 554 161
rect 596 131 626 161
rect 682 131 712 239
rect 760 253 826 269
rect 760 219 776 253
rect 810 219 826 253
rect 760 203 826 219
rect 868 271 934 287
rect 868 237 884 271
rect 918 237 934 271
rect 868 203 934 237
rect 760 131 790 203
rect 868 169 884 203
rect 918 169 934 203
rect 868 153 934 169
rect 982 237 1012 335
rect 1075 335 1192 351
rect 1075 301 1091 335
rect 1125 301 1192 335
rect 1075 285 1192 301
rect 982 221 1101 237
rect 982 187 1051 221
rect 1085 187 1101 221
rect 982 171 1101 187
rect 1162 193 1192 285
rect 1234 325 1250 359
rect 1284 325 1300 359
rect 1234 291 1300 325
rect 1361 305 1411 415
rect 1234 257 1250 291
rect 1284 257 1300 291
rect 1234 241 1300 257
rect 1342 289 1411 305
rect 1342 255 1358 289
rect 1392 255 1411 289
rect 868 131 898 153
rect 982 131 1012 171
rect 1162 163 1222 193
rect 1192 141 1222 163
rect 1264 141 1294 241
rect 1342 221 1411 255
rect 1342 187 1358 221
rect 1392 201 1411 221
rect 1392 187 1452 201
rect 1342 171 1452 187
rect 1350 141 1380 171
rect 1422 141 1452 171
rect 84 21 114 47
rect 156 21 186 47
rect 242 21 272 47
rect 320 21 350 47
rect 524 21 554 47
rect 596 21 626 47
rect 682 21 712 47
rect 760 21 790 47
rect 868 21 898 47
rect 982 21 1012 47
rect 1192 31 1222 57
rect 1264 31 1294 57
rect 1350 31 1380 57
rect 1422 31 1452 57
<< polycont >>
rect 108 306 142 340
rect 108 238 142 272
rect 222 308 256 342
rect 330 333 364 367
rect 596 333 630 367
rect 704 333 738 367
rect 222 240 256 274
rect 504 219 538 253
rect 776 219 810 253
rect 884 237 918 271
rect 884 169 918 203
rect 1091 301 1125 335
rect 1051 187 1085 221
rect 1250 325 1284 359
rect 1250 257 1284 291
rect 1358 255 1392 289
rect 1358 187 1392 221
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 22 597 113 613
rect 22 563 63 597
rect 97 563 113 597
rect 153 603 219 649
rect 153 569 169 603
rect 203 569 219 603
rect 551 603 601 649
rect 585 569 601 603
rect 22 533 113 563
rect 255 533 515 567
rect 22 529 289 533
rect 22 495 63 529
rect 97 499 289 529
rect 97 495 113 499
rect 22 461 113 495
rect 411 471 445 497
rect 22 427 63 461
rect 97 427 113 461
rect 22 411 113 427
rect 259 462 375 463
rect 259 428 275 462
rect 309 428 375 462
rect 259 411 375 428
rect 22 135 56 411
rect 314 367 375 411
rect 92 340 167 356
rect 92 306 108 340
rect 142 306 167 340
rect 92 272 167 306
rect 92 238 108 272
rect 142 238 167 272
rect 92 222 167 238
rect 206 342 272 358
rect 206 308 222 342
rect 256 308 272 342
rect 206 274 272 308
rect 206 240 222 274
rect 256 240 272 274
rect 206 224 272 240
rect 314 333 330 367
rect 364 333 375 367
rect 22 111 89 135
rect 22 77 39 111
rect 73 77 89 111
rect 22 53 89 77
rect 181 106 247 135
rect 181 72 197 106
rect 231 72 247 106
rect 181 17 247 72
rect 314 97 375 333
rect 411 167 445 437
rect 481 383 515 533
rect 551 469 601 569
rect 585 435 601 469
rect 551 419 601 435
rect 790 597 856 613
rect 790 563 806 597
rect 840 563 856 597
rect 790 529 856 563
rect 790 495 806 529
rect 840 495 856 529
rect 790 461 856 495
rect 790 427 806 461
rect 840 445 856 461
rect 1035 603 1101 649
rect 1035 569 1051 603
rect 1085 569 1101 603
rect 1035 532 1101 569
rect 1035 498 1051 532
rect 1085 498 1101 532
rect 1035 461 1101 498
rect 840 427 999 445
rect 790 411 999 427
rect 1035 427 1051 461
rect 1085 427 1101 461
rect 1035 411 1101 427
rect 1173 597 1239 613
rect 1173 563 1189 597
rect 1223 563 1239 597
rect 1173 529 1239 563
rect 1173 495 1189 529
rect 1223 495 1239 529
rect 1173 461 1239 495
rect 1279 603 1345 649
rect 1279 569 1295 603
rect 1329 569 1345 603
rect 1279 531 1345 569
rect 1279 497 1295 531
rect 1329 497 1345 531
rect 1279 481 1345 497
rect 1406 597 1513 613
rect 1406 563 1422 597
rect 1456 563 1513 597
rect 1406 529 1513 563
rect 1406 495 1422 529
rect 1456 495 1513 529
rect 1173 427 1189 461
rect 1223 445 1239 461
rect 1406 461 1513 495
rect 1223 427 1370 445
rect 1173 411 1370 427
rect 1406 427 1422 461
rect 1456 427 1513 461
rect 1406 411 1513 427
rect 481 367 646 383
rect 481 333 596 367
rect 630 333 646 367
rect 481 317 646 333
rect 688 367 754 383
rect 688 333 704 367
rect 738 351 754 367
rect 965 351 999 411
rect 1177 359 1300 375
rect 738 333 896 351
rect 688 317 896 333
rect 862 287 896 317
rect 965 335 1141 351
rect 965 301 1091 335
rect 1125 301 1141 335
rect 862 271 929 287
rect 488 253 826 269
rect 488 219 504 253
rect 538 219 776 253
rect 810 219 826 253
rect 488 203 826 219
rect 862 237 884 271
rect 918 237 929 271
rect 862 203 929 237
rect 862 169 884 203
rect 918 169 929 203
rect 862 167 929 169
rect 411 133 929 167
rect 965 285 1141 301
rect 1177 325 1250 359
rect 1284 325 1300 359
rect 1177 291 1300 325
rect 463 111 529 133
rect 314 95 411 97
rect 314 61 361 95
rect 395 61 411 95
rect 314 59 411 61
rect 463 77 479 111
rect 513 77 529 111
rect 965 97 999 285
rect 1177 257 1250 291
rect 1284 257 1300 291
rect 1177 241 1300 257
rect 1336 305 1370 411
rect 1336 289 1408 305
rect 1336 255 1358 289
rect 1392 255 1408 289
rect 1035 221 1101 237
rect 1035 187 1051 221
rect 1085 205 1101 221
rect 1336 221 1408 255
rect 1336 205 1358 221
rect 1085 187 1358 205
rect 1392 187 1408 221
rect 1035 171 1408 187
rect 463 53 529 77
rect 621 95 687 97
rect 621 61 637 95
rect 671 61 687 95
rect 621 17 687 61
rect 807 95 999 97
rect 807 61 823 95
rect 857 61 999 95
rect 807 59 999 61
rect 1035 106 1085 135
rect 1069 72 1085 106
rect 1035 17 1085 72
rect 1131 116 1197 171
rect 1131 82 1147 116
rect 1181 82 1197 116
rect 1131 53 1197 82
rect 1289 111 1355 135
rect 1289 77 1305 111
rect 1339 77 1355 111
rect 1289 17 1355 77
rect 1447 116 1513 411
rect 1447 82 1463 116
rect 1497 82 1513 116
rect 1447 53 1513 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrtn_lp
flabel comment s 544 242 544 242 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1471 94 1505 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 168 1505 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 390 1505 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 464 1505 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 538 1505 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2678076
string GDS_START 2666284
<< end >>
