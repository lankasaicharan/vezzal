magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1778 1975
<< nwell >>
rect -38 331 518 704
<< pwell >>
rect 199 157 473 241
rect 8 49 473 157
rect 0 0 480 49
<< scnmos >>
rect 87 47 117 131
rect 173 47 203 131
rect 278 47 308 215
rect 364 47 394 215
<< scpmoshvt >>
rect 101 390 131 474
rect 173 390 203 474
rect 278 367 308 619
rect 364 367 394 619
<< ndiff >>
rect 225 131 278 215
rect 34 106 87 131
rect 34 72 42 106
rect 76 72 87 106
rect 34 47 87 72
rect 117 101 173 131
rect 117 67 128 101
rect 162 67 173 101
rect 117 47 173 67
rect 203 103 278 131
rect 203 69 224 103
rect 258 69 278 103
rect 203 47 278 69
rect 308 203 364 215
rect 308 169 319 203
rect 353 169 364 203
rect 308 101 364 169
rect 308 67 319 101
rect 353 67 364 101
rect 308 47 364 67
rect 394 203 447 215
rect 394 169 405 203
rect 439 169 447 203
rect 394 93 447 169
rect 394 59 405 93
rect 439 59 447 93
rect 394 47 447 59
<< pdiff >>
rect 225 607 278 619
rect 225 573 233 607
rect 267 573 278 607
rect 225 522 278 573
rect 225 488 233 522
rect 267 488 278 522
rect 225 474 278 488
rect 48 436 101 474
rect 48 402 56 436
rect 90 402 101 436
rect 48 390 101 402
rect 131 390 173 474
rect 203 444 278 474
rect 203 410 214 444
rect 248 410 278 444
rect 203 390 278 410
rect 225 367 278 390
rect 308 599 364 619
rect 308 565 319 599
rect 353 565 364 599
rect 308 506 364 565
rect 308 472 319 506
rect 353 472 364 506
rect 308 413 364 472
rect 308 379 319 413
rect 353 379 364 413
rect 308 367 364 379
rect 394 607 447 619
rect 394 573 405 607
rect 439 573 447 607
rect 394 513 447 573
rect 394 479 405 513
rect 439 479 447 513
rect 394 413 447 479
rect 394 379 405 413
rect 439 379 447 413
rect 394 367 447 379
<< ndiffc >>
rect 42 72 76 106
rect 128 67 162 101
rect 224 69 258 103
rect 319 169 353 203
rect 319 67 353 101
rect 405 169 439 203
rect 405 59 439 93
<< pdiffc >>
rect 233 573 267 607
rect 233 488 267 522
rect 56 402 90 436
rect 214 410 248 444
rect 319 565 353 599
rect 319 472 353 506
rect 319 379 353 413
rect 405 573 439 607
rect 405 479 439 513
rect 405 379 439 413
<< poly >>
rect 278 619 308 645
rect 364 619 394 645
rect 101 474 131 500
rect 173 474 203 500
rect 101 368 131 390
rect 57 338 131 368
rect 57 292 87 338
rect 173 296 203 390
rect 278 321 308 367
rect 364 321 394 367
rect 21 276 87 292
rect 21 242 37 276
rect 71 242 87 276
rect 21 208 87 242
rect 129 280 203 296
rect 129 246 145 280
rect 179 246 203 280
rect 245 305 394 321
rect 245 271 261 305
rect 295 271 394 305
rect 245 255 394 271
rect 129 230 203 246
rect 21 174 37 208
rect 71 188 87 208
rect 71 174 117 188
rect 21 158 117 174
rect 87 131 117 158
rect 173 131 203 230
rect 278 215 308 255
rect 364 215 394 255
rect 87 21 117 47
rect 173 21 203 47
rect 278 21 308 47
rect 364 21 394 47
<< polycont >>
rect 37 242 71 276
rect 145 246 179 280
rect 261 271 295 305
rect 37 174 71 208
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 192 607 275 649
rect 192 573 233 607
rect 267 573 275 607
rect 192 522 275 573
rect 192 488 233 522
rect 267 488 275 522
rect 52 436 94 452
rect 52 402 56 436
rect 90 402 94 436
rect 52 360 94 402
rect 192 444 275 488
rect 192 410 214 444
rect 248 410 275 444
rect 192 394 275 410
rect 309 599 355 615
rect 309 565 319 599
rect 353 565 355 599
rect 309 506 355 565
rect 309 472 319 506
rect 353 472 355 506
rect 309 413 355 472
rect 389 607 455 649
rect 389 573 405 607
rect 439 573 455 607
rect 389 513 455 573
rect 389 479 405 513
rect 439 479 455 513
rect 389 419 455 479
rect 309 379 319 413
rect 353 385 355 413
rect 397 413 455 419
rect 353 379 363 385
rect 52 326 275 360
rect 309 353 363 379
rect 397 379 405 413
rect 439 379 455 413
rect 397 363 455 379
rect 237 321 275 326
rect 237 305 295 321
rect 17 276 81 292
rect 17 242 37 276
rect 71 242 81 276
rect 17 208 81 242
rect 115 280 195 292
rect 115 246 145 280
rect 179 246 195 280
rect 115 230 195 246
rect 237 271 261 305
rect 237 255 295 271
rect 17 174 37 208
rect 71 174 81 208
rect 237 179 283 255
rect 329 228 363 353
rect 17 158 81 174
rect 118 145 283 179
rect 317 203 363 228
rect 317 169 319 203
rect 353 201 363 203
rect 397 203 455 219
rect 353 169 355 201
rect 26 106 84 122
rect 26 72 42 106
rect 76 72 84 106
rect 26 17 84 72
rect 118 101 174 145
rect 118 67 128 101
rect 162 67 174 101
rect 118 51 174 67
rect 208 103 274 111
rect 208 69 224 103
rect 258 69 274 103
rect 208 17 274 69
rect 317 101 355 169
rect 397 169 405 203
rect 439 169 455 203
rect 397 167 455 169
rect 317 67 319 101
rect 353 67 355 101
rect 317 51 355 67
rect 389 93 455 167
rect 389 59 405 93
rect 439 59 455 93
rect 389 17 455 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or2_2
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6096006
string GDS_START 6090726
<< end >>
