magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
<< pwell >>
rect 16 49 1245 241
rect 0 0 1248 49
<< scnmos >>
rect 95 47 125 215
rect 249 47 279 215
rect 335 47 365 215
rect 421 47 451 215
rect 509 47 539 215
rect 690 47 720 215
rect 776 47 806 215
rect 878 47 908 215
rect 964 47 994 215
rect 1050 47 1080 215
rect 1136 47 1166 215
<< scpmoshvt >>
rect 102 367 132 619
rect 188 367 218 619
rect 274 367 304 619
rect 360 367 390 619
rect 446 367 476 619
rect 698 367 728 619
rect 784 367 814 619
rect 870 367 900 619
rect 964 367 994 619
rect 1050 367 1080 619
rect 1136 367 1166 619
<< ndiff >>
rect 42 190 95 215
rect 42 156 50 190
rect 84 156 95 190
rect 42 101 95 156
rect 42 67 50 101
rect 84 67 95 101
rect 42 47 95 67
rect 125 167 249 215
rect 125 133 136 167
rect 170 133 204 167
rect 238 133 249 167
rect 125 93 249 133
rect 125 59 136 93
rect 170 59 204 93
rect 238 59 249 93
rect 125 47 249 59
rect 279 203 335 215
rect 279 169 290 203
rect 324 169 335 203
rect 279 101 335 169
rect 279 67 290 101
rect 324 67 335 101
rect 279 47 335 67
rect 365 165 421 215
rect 365 131 376 165
rect 410 131 421 165
rect 365 93 421 131
rect 365 59 376 93
rect 410 59 421 93
rect 365 47 421 59
rect 451 203 509 215
rect 451 169 462 203
rect 496 169 509 203
rect 451 101 509 169
rect 451 67 462 101
rect 496 67 509 101
rect 451 47 509 67
rect 539 165 690 215
rect 539 131 550 165
rect 584 131 645 165
rect 679 131 690 165
rect 539 89 690 131
rect 539 55 550 89
rect 584 55 645 89
rect 679 55 690 89
rect 539 47 690 55
rect 720 207 776 215
rect 720 173 731 207
rect 765 173 776 207
rect 720 101 776 173
rect 720 67 731 101
rect 765 67 776 101
rect 720 47 776 67
rect 806 165 878 215
rect 806 131 817 165
rect 851 131 878 165
rect 806 89 878 131
rect 806 55 817 89
rect 851 55 878 89
rect 806 47 878 55
rect 908 165 964 215
rect 908 131 919 165
rect 953 131 964 165
rect 908 91 964 131
rect 908 57 919 91
rect 953 57 964 91
rect 908 47 964 57
rect 994 169 1050 215
rect 994 135 1005 169
rect 1039 135 1050 169
rect 994 47 1050 135
rect 1080 203 1136 215
rect 1080 169 1091 203
rect 1125 169 1136 203
rect 1080 101 1136 169
rect 1080 67 1091 101
rect 1125 67 1136 101
rect 1080 47 1136 67
rect 1166 203 1219 215
rect 1166 169 1177 203
rect 1211 169 1219 203
rect 1166 93 1219 169
rect 1166 59 1177 93
rect 1211 59 1219 93
rect 1166 47 1219 59
<< pdiff >>
rect 49 599 102 619
rect 49 565 57 599
rect 91 565 102 599
rect 49 516 102 565
rect 49 482 57 516
rect 91 482 102 516
rect 49 436 102 482
rect 49 402 57 436
rect 91 402 102 436
rect 49 367 102 402
rect 132 592 188 619
rect 132 558 143 592
rect 177 558 188 592
rect 132 367 188 558
rect 218 424 274 619
rect 218 390 229 424
rect 263 390 274 424
rect 218 367 274 390
rect 304 592 360 619
rect 304 558 315 592
rect 349 558 360 592
rect 304 367 360 558
rect 390 424 446 619
rect 390 390 401 424
rect 435 390 446 424
rect 390 367 446 390
rect 476 592 529 619
rect 476 558 487 592
rect 521 558 529 592
rect 476 367 529 558
rect 645 599 698 619
rect 645 565 653 599
rect 687 565 698 599
rect 645 529 698 565
rect 645 495 653 529
rect 687 495 698 529
rect 645 459 698 495
rect 645 425 653 459
rect 687 425 698 459
rect 645 367 698 425
rect 728 547 784 619
rect 728 513 739 547
rect 773 513 784 547
rect 728 479 784 513
rect 728 445 739 479
rect 773 445 784 479
rect 728 411 784 445
rect 728 377 739 411
rect 773 377 784 411
rect 728 367 784 377
rect 814 599 870 619
rect 814 565 825 599
rect 859 565 870 599
rect 814 498 870 565
rect 814 464 825 498
rect 859 464 870 498
rect 814 409 870 464
rect 814 375 825 409
rect 859 375 870 409
rect 814 367 870 375
rect 900 567 964 619
rect 900 533 911 567
rect 945 533 964 567
rect 900 367 964 533
rect 994 599 1050 619
rect 994 565 1005 599
rect 1039 565 1050 599
rect 994 508 1050 565
rect 994 474 1005 508
rect 1039 474 1050 508
rect 994 367 1050 474
rect 1080 567 1136 619
rect 1080 533 1091 567
rect 1125 533 1136 567
rect 1080 367 1136 533
rect 1166 599 1219 619
rect 1166 565 1177 599
rect 1211 565 1219 599
rect 1166 498 1219 565
rect 1166 464 1177 498
rect 1211 464 1219 498
rect 1166 413 1219 464
rect 1166 379 1177 413
rect 1211 379 1219 413
rect 1166 367 1219 379
<< ndiffc >>
rect 50 156 84 190
rect 50 67 84 101
rect 136 133 170 167
rect 204 133 238 167
rect 136 59 170 93
rect 204 59 238 93
rect 290 169 324 203
rect 290 67 324 101
rect 376 131 410 165
rect 376 59 410 93
rect 462 169 496 203
rect 462 67 496 101
rect 550 131 584 165
rect 645 131 679 165
rect 550 55 584 89
rect 645 55 679 89
rect 731 173 765 207
rect 731 67 765 101
rect 817 131 851 165
rect 817 55 851 89
rect 919 131 953 165
rect 919 57 953 91
rect 1005 135 1039 169
rect 1091 169 1125 203
rect 1091 67 1125 101
rect 1177 169 1211 203
rect 1177 59 1211 93
<< pdiffc >>
rect 57 565 91 599
rect 57 482 91 516
rect 57 402 91 436
rect 143 558 177 592
rect 229 390 263 424
rect 315 558 349 592
rect 401 390 435 424
rect 487 558 521 592
rect 653 565 687 599
rect 653 495 687 529
rect 653 425 687 459
rect 739 513 773 547
rect 739 445 773 479
rect 739 377 773 411
rect 825 565 859 599
rect 825 464 859 498
rect 825 375 859 409
rect 911 533 945 567
rect 1005 565 1039 599
rect 1005 474 1039 508
rect 1091 533 1125 567
rect 1177 565 1211 599
rect 1177 464 1211 498
rect 1177 379 1211 413
<< poly >>
rect 102 619 132 645
rect 188 619 218 645
rect 274 619 304 645
rect 360 619 390 645
rect 446 619 476 645
rect 698 619 728 645
rect 784 619 814 645
rect 870 619 900 645
rect 964 619 994 645
rect 1050 619 1080 645
rect 1136 619 1166 645
rect 102 308 132 367
rect 188 345 218 367
rect 274 345 304 367
rect 188 321 304 345
rect 360 321 390 367
rect 446 321 476 367
rect 698 335 728 367
rect 784 335 814 367
rect 188 315 539 321
rect 74 292 140 308
rect 74 258 90 292
rect 124 258 140 292
rect 74 242 140 258
rect 249 305 539 315
rect 249 271 285 305
rect 319 271 353 305
rect 387 271 421 305
rect 455 271 489 305
rect 523 271 539 305
rect 249 255 539 271
rect 582 319 814 335
rect 870 325 900 367
rect 964 335 994 367
rect 1050 335 1080 367
rect 582 285 614 319
rect 648 285 814 319
rect 582 269 814 285
rect 856 309 922 325
rect 856 275 872 309
rect 906 275 922 309
rect 95 215 125 242
rect 249 215 279 255
rect 335 215 365 255
rect 421 215 451 255
rect 509 215 539 255
rect 690 215 720 269
rect 776 215 806 269
rect 856 259 922 275
rect 964 319 1080 335
rect 964 285 1003 319
rect 1037 285 1080 319
rect 964 269 1080 285
rect 878 215 908 259
rect 964 215 994 269
rect 1050 215 1080 269
rect 1136 335 1166 367
rect 1136 319 1202 335
rect 1136 285 1152 319
rect 1186 285 1202 319
rect 1136 269 1202 285
rect 1136 215 1166 269
rect 95 21 125 47
rect 249 21 279 47
rect 335 21 365 47
rect 421 21 451 47
rect 509 21 539 47
rect 690 21 720 47
rect 776 21 806 47
rect 878 21 908 47
rect 964 21 994 47
rect 1050 21 1080 47
rect 1136 21 1166 47
<< polycont >>
rect 90 258 124 292
rect 285 271 319 305
rect 353 271 387 305
rect 421 271 455 305
rect 489 271 523 305
rect 614 285 648 319
rect 872 275 906 309
rect 1003 285 1037 319
rect 1152 285 1186 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 18 599 91 615
rect 18 565 57 599
rect 18 516 91 565
rect 127 592 193 649
rect 127 558 143 592
rect 177 558 193 592
rect 127 542 193 558
rect 299 592 365 649
rect 299 558 315 592
rect 349 558 365 592
rect 299 542 365 558
rect 471 592 537 649
rect 471 558 487 592
rect 521 558 537 592
rect 471 542 537 558
rect 649 599 861 615
rect 649 565 653 599
rect 687 581 825 599
rect 687 565 689 581
rect 18 482 57 516
rect 649 529 689 565
rect 823 565 825 581
rect 859 565 861 599
rect 91 482 615 508
rect 18 474 615 482
rect 18 436 91 474
rect 18 402 57 436
rect 18 386 91 402
rect 127 424 545 440
rect 127 390 229 424
rect 263 390 401 424
rect 435 390 545 424
rect 127 386 545 390
rect 18 206 54 386
rect 199 360 545 386
rect 581 375 615 474
rect 649 495 653 529
rect 687 495 689 529
rect 649 459 689 495
rect 649 425 653 459
rect 687 425 689 459
rect 649 409 689 425
rect 723 513 739 547
rect 773 513 789 547
rect 723 479 789 513
rect 723 445 739 479
rect 773 445 789 479
rect 723 411 789 445
rect 723 377 739 411
rect 773 377 789 411
rect 88 292 161 352
rect 88 258 90 292
rect 124 258 161 292
rect 88 240 161 258
rect 199 235 233 360
rect 581 341 664 375
rect 598 319 664 341
rect 269 305 564 307
rect 269 271 285 305
rect 319 271 353 305
rect 387 271 421 305
rect 455 271 489 305
rect 523 271 564 305
rect 18 190 86 206
rect 199 203 496 235
rect 199 201 290 203
rect 18 156 50 190
rect 84 156 86 190
rect 288 169 290 201
rect 324 201 462 203
rect 324 169 326 201
rect 18 101 86 156
rect 18 67 50 101
rect 84 67 86 101
rect 18 51 86 67
rect 120 133 136 167
rect 170 133 204 167
rect 238 133 254 167
rect 120 93 254 133
rect 120 59 136 93
rect 170 59 204 93
rect 238 59 254 93
rect 120 17 254 59
rect 288 101 326 169
rect 460 169 462 201
rect 530 233 564 271
rect 598 285 614 319
rect 648 285 664 319
rect 598 269 664 285
rect 723 233 789 377
rect 823 498 861 565
rect 895 567 961 649
rect 895 533 911 567
rect 945 533 961 567
rect 895 526 961 533
rect 995 599 1041 615
rect 995 565 1005 599
rect 1039 565 1041 599
rect 823 464 825 498
rect 859 492 861 498
rect 995 508 1041 565
rect 1075 567 1141 649
rect 1075 533 1091 567
rect 1125 533 1141 567
rect 1075 526 1141 533
rect 1175 599 1227 615
rect 1175 565 1177 599
rect 1211 565 1227 599
rect 995 492 1005 508
rect 859 474 1005 492
rect 1039 492 1041 508
rect 1175 498 1227 565
rect 1175 492 1177 498
rect 1039 474 1177 492
rect 859 464 1177 474
rect 1211 464 1227 498
rect 823 458 1227 464
rect 823 409 861 458
rect 823 375 825 409
rect 859 375 861 409
rect 823 359 861 375
rect 895 388 1133 424
rect 895 325 929 388
rect 856 309 929 325
rect 856 275 872 309
rect 906 275 929 309
rect 856 267 929 275
rect 980 319 1053 354
rect 980 285 1003 319
rect 1037 285 1053 319
rect 980 269 1053 285
rect 1087 329 1133 388
rect 1167 413 1227 458
rect 1167 379 1177 413
rect 1211 379 1227 413
rect 1167 363 1227 379
rect 1087 319 1202 329
rect 1087 285 1152 319
rect 1186 285 1202 319
rect 1087 268 1202 285
rect 530 207 1043 233
rect 530 199 731 207
rect 288 67 290 101
rect 324 67 326 101
rect 288 51 326 67
rect 360 131 376 165
rect 410 131 426 165
rect 360 93 426 131
rect 360 59 376 93
rect 410 59 426 93
rect 360 17 426 59
rect 460 101 496 169
rect 729 173 731 199
rect 765 199 1043 207
rect 765 173 767 199
rect 460 67 462 101
rect 460 51 496 67
rect 534 131 550 165
rect 584 131 645 165
rect 679 131 695 165
rect 534 89 695 131
rect 534 55 550 89
rect 584 55 645 89
rect 679 55 695 89
rect 534 17 695 55
rect 729 101 767 173
rect 1003 169 1043 199
rect 729 67 731 101
rect 765 67 767 101
rect 729 51 767 67
rect 801 131 817 165
rect 851 131 867 165
rect 801 89 867 131
rect 801 55 817 89
rect 851 55 867 89
rect 801 17 867 55
rect 903 131 919 165
rect 953 131 969 165
rect 903 91 969 131
rect 1003 135 1005 169
rect 1039 135 1043 169
rect 1003 119 1043 135
rect 1087 203 1137 219
rect 1087 169 1091 203
rect 1125 169 1137 203
rect 903 57 919 91
rect 953 85 969 91
rect 1087 101 1137 169
rect 1087 85 1091 101
rect 953 67 1091 85
rect 1125 67 1137 101
rect 953 57 1137 67
rect 903 51 1137 57
rect 1171 203 1227 219
rect 1171 169 1177 203
rect 1211 169 1227 203
rect 1171 93 1227 169
rect 1171 59 1177 93
rect 1211 59 1227 93
rect 1171 17 1227 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21bo_4
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1087 390 1121 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3763162
string GDS_START 3752382
<< end >>
