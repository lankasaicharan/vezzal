magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
rect 616 309 1090 331
<< pwell >>
rect 4 241 450 243
rect 4 49 1518 241
rect 0 0 1536 49
<< scnmos >>
rect 83 49 113 217
rect 169 49 199 217
rect 255 49 285 217
rect 341 49 371 217
rect 533 47 563 215
rect 619 47 649 215
rect 705 47 735 215
rect 791 47 821 215
rect 877 47 907 215
rect 963 47 993 215
rect 1049 47 1079 215
rect 1233 47 1263 215
rect 1319 47 1349 215
rect 1405 47 1435 215
<< scpmoshvt >>
rect 83 367 113 619
rect 169 367 199 619
rect 255 367 285 619
rect 341 367 371 619
rect 427 367 457 619
rect 513 367 543 619
rect 705 345 735 597
rect 791 345 821 597
rect 877 345 907 597
rect 963 345 993 597
rect 1161 367 1191 619
rect 1247 367 1277 619
rect 1333 367 1363 619
rect 1419 367 1449 619
<< ndiff >>
rect 30 174 83 217
rect 30 140 38 174
rect 72 140 83 174
rect 30 95 83 140
rect 30 61 38 95
rect 72 61 83 95
rect 30 49 83 61
rect 113 205 169 217
rect 113 171 124 205
rect 158 171 169 205
rect 113 101 169 171
rect 113 67 124 101
rect 158 67 169 101
rect 113 49 169 67
rect 199 175 255 217
rect 199 141 210 175
rect 244 141 255 175
rect 199 91 255 141
rect 199 57 210 91
rect 244 57 255 91
rect 199 49 255 57
rect 285 205 341 217
rect 285 171 296 205
rect 330 171 341 205
rect 285 101 341 171
rect 285 67 296 101
rect 330 67 341 101
rect 285 49 341 67
rect 371 205 424 217
rect 371 171 382 205
rect 416 171 424 205
rect 371 95 424 171
rect 371 61 382 95
rect 416 61 424 95
rect 371 49 424 61
rect 480 122 533 215
rect 480 88 488 122
rect 522 88 533 122
rect 480 47 533 88
rect 563 164 619 215
rect 563 130 574 164
rect 608 130 619 164
rect 563 47 619 130
rect 649 192 705 215
rect 649 158 660 192
rect 694 158 705 192
rect 649 103 705 158
rect 649 69 660 103
rect 694 69 705 103
rect 649 47 705 69
rect 735 124 791 215
rect 735 90 746 124
rect 780 90 791 124
rect 735 47 791 90
rect 821 192 877 215
rect 821 158 832 192
rect 866 158 877 192
rect 821 101 877 158
rect 821 67 832 101
rect 866 67 877 101
rect 821 47 877 67
rect 907 124 963 215
rect 907 90 918 124
rect 952 90 963 124
rect 907 47 963 90
rect 993 192 1049 215
rect 993 158 1004 192
rect 1038 158 1049 192
rect 993 101 1049 158
rect 993 67 1004 101
rect 1038 67 1049 101
rect 993 47 1049 67
rect 1079 124 1233 215
rect 1079 90 1090 124
rect 1124 90 1188 124
rect 1222 90 1233 124
rect 1079 47 1233 90
rect 1263 192 1319 215
rect 1263 158 1274 192
rect 1308 158 1319 192
rect 1263 101 1319 158
rect 1263 67 1274 101
rect 1308 67 1319 101
rect 1263 47 1319 67
rect 1349 124 1405 215
rect 1349 90 1360 124
rect 1394 90 1405 124
rect 1349 47 1405 90
rect 1435 192 1492 215
rect 1435 158 1450 192
rect 1484 158 1492 192
rect 1435 103 1492 158
rect 1435 69 1450 103
rect 1484 69 1492 103
rect 1435 47 1492 69
<< pdiff >>
rect 30 607 83 619
rect 30 573 38 607
rect 72 573 83 607
rect 30 532 83 573
rect 30 498 38 532
rect 72 498 83 532
rect 30 453 83 498
rect 30 419 38 453
rect 72 419 83 453
rect 30 367 83 419
rect 113 599 169 619
rect 113 565 124 599
rect 158 565 169 599
rect 113 506 169 565
rect 113 472 124 506
rect 158 472 169 506
rect 113 413 169 472
rect 113 379 124 413
rect 158 379 169 413
rect 113 367 169 379
rect 199 607 255 619
rect 199 573 210 607
rect 244 573 255 607
rect 199 532 255 573
rect 199 498 210 532
rect 244 498 255 532
rect 199 455 255 498
rect 199 421 210 455
rect 244 421 255 455
rect 199 367 255 421
rect 285 599 341 619
rect 285 565 296 599
rect 330 565 341 599
rect 285 506 341 565
rect 285 472 296 506
rect 330 472 341 506
rect 285 413 341 472
rect 285 379 296 413
rect 330 379 341 413
rect 285 367 341 379
rect 371 607 427 619
rect 371 573 382 607
rect 416 573 427 607
rect 371 506 427 573
rect 371 472 382 506
rect 416 472 427 506
rect 371 413 427 472
rect 371 379 382 413
rect 416 379 427 413
rect 371 367 427 379
rect 457 599 513 619
rect 457 565 468 599
rect 502 565 513 599
rect 457 506 513 565
rect 457 472 468 506
rect 502 472 513 506
rect 457 413 513 472
rect 457 379 468 413
rect 502 379 513 413
rect 457 367 513 379
rect 543 607 596 619
rect 543 573 554 607
rect 588 573 596 607
rect 543 517 596 573
rect 543 483 554 517
rect 588 483 596 517
rect 543 431 596 483
rect 543 397 554 431
rect 588 397 596 431
rect 543 367 596 397
rect 652 585 705 597
rect 652 551 660 585
rect 694 551 705 585
rect 652 510 705 551
rect 652 476 660 510
rect 694 476 705 510
rect 652 431 705 476
rect 652 397 660 431
rect 694 397 705 431
rect 652 345 705 397
rect 735 531 791 597
rect 735 497 746 531
rect 780 497 791 531
rect 735 463 791 497
rect 735 429 746 463
rect 780 429 791 463
rect 735 387 791 429
rect 735 353 746 387
rect 780 353 791 387
rect 735 345 791 353
rect 821 585 877 597
rect 821 551 832 585
rect 866 551 877 585
rect 821 489 877 551
rect 821 455 832 489
rect 866 455 877 489
rect 821 391 877 455
rect 821 357 832 391
rect 866 357 877 391
rect 821 345 877 357
rect 907 585 963 597
rect 907 551 918 585
rect 952 551 963 585
rect 907 517 963 551
rect 907 483 918 517
rect 952 483 963 517
rect 907 439 963 483
rect 907 405 918 439
rect 952 405 963 439
rect 907 345 963 405
rect 993 545 1054 597
rect 993 511 1004 545
rect 1038 511 1054 545
rect 993 471 1054 511
rect 993 437 1004 471
rect 1038 437 1054 471
rect 993 391 1054 437
rect 993 357 1004 391
rect 1038 357 1054 391
rect 1108 529 1161 619
rect 1108 495 1116 529
rect 1150 495 1161 529
rect 1108 413 1161 495
rect 1108 379 1116 413
rect 1150 379 1161 413
rect 1108 367 1161 379
rect 1191 597 1247 619
rect 1191 563 1202 597
rect 1236 563 1247 597
rect 1191 521 1247 563
rect 1191 487 1202 521
rect 1236 487 1247 521
rect 1191 445 1247 487
rect 1191 411 1202 445
rect 1236 411 1247 445
rect 1191 367 1247 411
rect 1277 599 1333 619
rect 1277 565 1288 599
rect 1322 565 1333 599
rect 1277 506 1333 565
rect 1277 472 1288 506
rect 1322 472 1333 506
rect 1277 409 1333 472
rect 1277 375 1288 409
rect 1322 375 1333 409
rect 1277 367 1333 375
rect 1363 607 1419 619
rect 1363 573 1374 607
rect 1408 573 1419 607
rect 1363 531 1419 573
rect 1363 497 1374 531
rect 1408 497 1419 531
rect 1363 455 1419 497
rect 1363 421 1374 455
rect 1408 421 1419 455
rect 1363 367 1419 421
rect 1449 599 1502 619
rect 1449 565 1460 599
rect 1494 565 1502 599
rect 1449 506 1502 565
rect 1449 472 1460 506
rect 1494 472 1502 506
rect 1449 413 1502 472
rect 1449 379 1460 413
rect 1494 379 1502 413
rect 1449 367 1502 379
rect 993 345 1054 357
<< ndiffc >>
rect 38 140 72 174
rect 38 61 72 95
rect 124 171 158 205
rect 124 67 158 101
rect 210 141 244 175
rect 210 57 244 91
rect 296 171 330 205
rect 296 67 330 101
rect 382 171 416 205
rect 382 61 416 95
rect 488 88 522 122
rect 574 130 608 164
rect 660 158 694 192
rect 660 69 694 103
rect 746 90 780 124
rect 832 158 866 192
rect 832 67 866 101
rect 918 90 952 124
rect 1004 158 1038 192
rect 1004 67 1038 101
rect 1090 90 1124 124
rect 1188 90 1222 124
rect 1274 158 1308 192
rect 1274 67 1308 101
rect 1360 90 1394 124
rect 1450 158 1484 192
rect 1450 69 1484 103
<< pdiffc >>
rect 38 573 72 607
rect 38 498 72 532
rect 38 419 72 453
rect 124 565 158 599
rect 124 472 158 506
rect 124 379 158 413
rect 210 573 244 607
rect 210 498 244 532
rect 210 421 244 455
rect 296 565 330 599
rect 296 472 330 506
rect 296 379 330 413
rect 382 573 416 607
rect 382 472 416 506
rect 382 379 416 413
rect 468 565 502 599
rect 468 472 502 506
rect 468 379 502 413
rect 554 573 588 607
rect 554 483 588 517
rect 554 397 588 431
rect 660 551 694 585
rect 660 476 694 510
rect 660 397 694 431
rect 746 497 780 531
rect 746 429 780 463
rect 746 353 780 387
rect 832 551 866 585
rect 832 455 866 489
rect 832 357 866 391
rect 918 551 952 585
rect 918 483 952 517
rect 918 405 952 439
rect 1004 511 1038 545
rect 1004 437 1038 471
rect 1004 357 1038 391
rect 1116 495 1150 529
rect 1116 379 1150 413
rect 1202 563 1236 597
rect 1202 487 1236 521
rect 1202 411 1236 445
rect 1288 565 1322 599
rect 1288 472 1322 506
rect 1288 375 1322 409
rect 1374 573 1408 607
rect 1374 497 1408 531
rect 1374 421 1408 455
rect 1460 565 1494 599
rect 1460 472 1494 506
rect 1460 379 1494 413
<< poly >>
rect 83 619 113 645
rect 169 619 199 645
rect 255 619 285 645
rect 341 619 371 645
rect 427 619 457 645
rect 513 619 543 645
rect 705 597 735 623
rect 791 597 821 623
rect 877 597 907 623
rect 963 597 993 623
rect 1161 619 1191 645
rect 1247 619 1277 645
rect 1333 619 1363 645
rect 1419 619 1449 645
rect 83 331 113 367
rect 169 331 199 367
rect 255 331 285 367
rect 341 331 371 367
rect 83 315 371 331
rect 83 281 117 315
rect 151 281 185 315
rect 219 281 253 315
rect 287 281 321 315
rect 355 281 371 315
rect 83 265 371 281
rect 83 217 113 265
rect 169 217 199 265
rect 255 217 285 265
rect 341 217 371 265
rect 427 303 457 367
rect 513 303 543 367
rect 705 303 735 345
rect 791 303 821 345
rect 877 303 907 345
rect 963 303 993 345
rect 1161 303 1191 367
rect 1247 303 1277 367
rect 1333 305 1363 367
rect 427 287 649 303
rect 427 253 554 287
rect 588 253 649 287
rect 427 237 649 253
rect 697 287 821 303
rect 697 253 713 287
rect 747 253 821 287
rect 697 237 821 253
rect 863 287 1007 303
rect 863 253 879 287
rect 913 253 957 287
rect 991 253 1007 287
rect 863 237 1007 253
rect 1049 287 1277 303
rect 1049 253 1103 287
rect 1137 253 1195 287
rect 1229 253 1277 287
rect 1049 237 1277 253
rect 1319 303 1363 305
rect 1419 303 1449 367
rect 1319 287 1453 303
rect 1319 253 1335 287
rect 1369 253 1403 287
rect 1437 253 1453 287
rect 1319 237 1453 253
rect 533 215 563 237
rect 619 215 649 237
rect 705 215 735 237
rect 791 215 821 237
rect 877 215 907 237
rect 963 215 993 237
rect 1049 215 1079 237
rect 1233 215 1263 237
rect 1319 215 1349 237
rect 1405 215 1435 237
rect 83 23 113 49
rect 169 23 199 49
rect 255 23 285 49
rect 341 23 371 49
rect 533 21 563 47
rect 619 21 649 47
rect 705 21 735 47
rect 791 21 821 47
rect 877 21 907 47
rect 963 21 993 47
rect 1049 21 1079 47
rect 1233 21 1263 47
rect 1319 21 1349 47
rect 1405 21 1435 47
<< polycont >>
rect 117 281 151 315
rect 185 281 219 315
rect 253 281 287 315
rect 321 281 355 315
rect 554 253 588 287
rect 713 253 747 287
rect 879 253 913 287
rect 957 253 991 287
rect 1103 253 1137 287
rect 1195 253 1229 287
rect 1335 253 1369 287
rect 1403 253 1437 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 22 607 88 649
rect 22 573 38 607
rect 72 573 88 607
rect 22 532 88 573
rect 22 498 38 532
rect 72 498 88 532
rect 22 453 88 498
rect 22 419 38 453
rect 72 419 88 453
rect 122 599 160 615
rect 122 565 124 599
rect 158 565 160 599
rect 122 506 160 565
rect 122 472 124 506
rect 158 472 160 506
rect 122 413 160 472
rect 194 607 260 649
rect 194 573 210 607
rect 244 573 260 607
rect 194 532 260 573
rect 194 498 210 532
rect 244 498 260 532
rect 194 455 260 498
rect 194 421 210 455
rect 244 421 260 455
rect 294 599 332 615
rect 294 565 296 599
rect 330 565 332 599
rect 294 506 332 565
rect 294 472 296 506
rect 330 472 332 506
rect 122 385 124 413
rect 17 379 124 385
rect 158 385 160 413
rect 294 413 332 472
rect 294 385 296 413
rect 158 379 296 385
rect 330 379 332 413
rect 17 351 332 379
rect 366 607 432 649
rect 366 573 382 607
rect 416 573 432 607
rect 366 506 432 573
rect 366 472 382 506
rect 416 472 432 506
rect 366 413 432 472
rect 366 379 382 413
rect 416 379 432 413
rect 366 363 432 379
rect 466 599 504 615
rect 466 565 468 599
rect 502 565 504 599
rect 466 506 504 565
rect 466 472 468 506
rect 502 472 504 506
rect 466 413 504 472
rect 466 379 468 413
rect 502 379 504 413
rect 538 607 604 649
rect 538 573 554 607
rect 588 573 604 607
rect 538 517 604 573
rect 538 483 554 517
rect 588 483 604 517
rect 538 431 604 483
rect 538 397 554 431
rect 588 397 604 431
rect 644 585 882 615
rect 644 551 660 585
rect 694 581 832 585
rect 694 551 710 581
rect 644 510 710 551
rect 816 551 832 581
rect 866 551 882 585
rect 644 476 660 510
rect 694 476 710 510
rect 644 431 710 476
rect 644 397 660 431
rect 694 397 710 431
rect 744 531 782 547
rect 744 497 746 531
rect 780 497 782 531
rect 744 463 782 497
rect 744 429 746 463
rect 780 429 782 463
rect 466 363 504 379
rect 744 387 782 429
rect 744 363 746 387
rect 466 353 746 363
rect 780 353 782 387
rect 17 245 67 351
rect 466 321 782 353
rect 816 489 882 551
rect 816 455 832 489
rect 866 455 882 489
rect 816 391 882 455
rect 816 357 832 391
rect 866 357 882 391
rect 916 597 1252 615
rect 916 585 1202 597
rect 916 551 918 585
rect 952 579 1202 585
rect 952 551 954 579
rect 916 517 954 551
rect 1186 563 1202 579
rect 1236 563 1252 597
rect 916 483 918 517
rect 952 483 954 517
rect 916 439 954 483
rect 916 405 918 439
rect 952 405 954 439
rect 916 389 954 405
rect 988 511 1004 545
rect 1038 511 1054 545
rect 988 471 1054 511
rect 988 437 1004 471
rect 1038 437 1054 471
rect 988 391 1054 437
rect 816 355 882 357
rect 988 357 1004 391
rect 1038 357 1054 391
rect 988 355 1054 357
rect 816 321 1054 355
rect 1100 529 1152 545
rect 1100 495 1116 529
rect 1150 495 1152 529
rect 1100 413 1152 495
rect 1100 379 1116 413
rect 1150 379 1152 413
rect 1186 521 1252 563
rect 1186 487 1202 521
rect 1236 487 1252 521
rect 1186 445 1252 487
rect 1186 411 1202 445
rect 1236 411 1252 445
rect 1286 599 1324 615
rect 1286 565 1288 599
rect 1322 565 1324 599
rect 1286 506 1324 565
rect 1286 472 1288 506
rect 1322 472 1324 506
rect 1100 375 1152 379
rect 1286 409 1324 472
rect 1358 607 1424 649
rect 1358 573 1374 607
rect 1408 573 1424 607
rect 1358 531 1424 573
rect 1358 497 1374 531
rect 1408 497 1424 531
rect 1358 455 1424 497
rect 1358 421 1374 455
rect 1408 421 1424 455
rect 1458 599 1498 615
rect 1458 565 1460 599
rect 1494 565 1498 599
rect 1458 506 1498 565
rect 1458 472 1460 506
rect 1494 472 1498 506
rect 1286 375 1288 409
rect 1322 375 1324 409
rect 1458 413 1498 472
rect 1458 379 1460 413
rect 1494 379 1498 413
rect 1458 375 1498 379
rect 1100 341 1498 375
rect 466 317 502 321
rect 101 315 502 317
rect 101 281 117 315
rect 151 281 185 315
rect 219 281 253 315
rect 287 281 321 315
rect 355 281 502 315
rect 101 279 502 281
rect 17 211 332 245
rect 122 205 160 211
rect 22 174 88 177
rect 22 140 38 174
rect 72 140 88 174
rect 22 95 88 140
rect 22 61 38 95
rect 72 61 88 95
rect 22 17 88 61
rect 122 171 124 205
rect 158 171 160 205
rect 294 205 332 211
rect 122 101 160 171
rect 122 67 124 101
rect 158 67 160 101
rect 122 51 160 67
rect 194 175 260 177
rect 194 141 210 175
rect 244 141 260 175
rect 194 91 260 141
rect 194 57 210 91
rect 244 57 260 91
rect 194 17 260 57
rect 294 171 296 205
rect 330 171 332 205
rect 294 101 332 171
rect 294 67 296 101
rect 330 67 332 101
rect 294 51 332 67
rect 366 205 430 221
rect 366 171 382 205
rect 416 171 430 205
rect 464 208 502 279
rect 538 253 554 287
rect 588 253 657 287
rect 538 242 657 253
rect 691 253 713 287
rect 747 253 763 287
rect 691 242 763 253
rect 797 253 879 287
rect 913 253 957 287
rect 991 253 1035 287
rect 797 242 1035 253
rect 1069 253 1103 287
rect 1137 253 1195 287
rect 1229 253 1245 287
rect 1069 242 1245 253
rect 1279 253 1335 287
rect 1369 253 1403 287
rect 1437 253 1519 287
rect 1279 242 1519 253
rect 464 172 624 208
rect 366 95 430 171
rect 558 164 624 172
rect 366 61 382 95
rect 416 61 430 95
rect 366 17 430 61
rect 472 122 524 138
rect 472 88 488 122
rect 522 88 524 122
rect 558 130 574 164
rect 608 130 624 164
rect 558 119 624 130
rect 658 192 1500 208
rect 658 158 660 192
rect 694 174 832 192
rect 694 158 703 174
rect 472 85 524 88
rect 658 103 703 158
rect 823 158 832 174
rect 866 174 1004 192
rect 866 158 875 174
rect 658 85 660 103
rect 472 69 660 85
rect 694 69 703 103
rect 472 51 703 69
rect 737 124 789 140
rect 737 90 746 124
rect 780 90 789 124
rect 737 17 789 90
rect 823 101 875 158
rect 994 158 1004 174
rect 1038 174 1274 192
rect 1038 158 1047 174
rect 823 67 832 101
rect 866 67 875 101
rect 823 51 875 67
rect 909 124 960 140
rect 909 90 918 124
rect 952 90 960 124
rect 909 17 960 90
rect 994 101 1047 158
rect 1264 158 1274 174
rect 1308 174 1450 192
rect 1308 158 1317 174
rect 994 67 1004 101
rect 1038 67 1047 101
rect 994 51 1047 67
rect 1081 124 1230 140
rect 1081 90 1090 124
rect 1124 90 1188 124
rect 1222 90 1230 124
rect 1081 17 1230 90
rect 1264 101 1317 158
rect 1437 158 1450 174
rect 1484 158 1500 192
rect 1264 67 1274 101
rect 1308 67 1317 101
rect 1264 51 1317 67
rect 1351 124 1403 140
rect 1351 90 1360 124
rect 1394 90 1403 124
rect 1351 17 1403 90
rect 1437 103 1500 158
rect 1437 69 1450 103
rect 1484 69 1500 103
rect 1437 53 1500 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o41a_4
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 525976
string GDS_START 512132
<< end >>
