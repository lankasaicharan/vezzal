magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 1 157 427 167
rect 1364 157 1631 193
rect 1 49 1631 157
rect 0 0 1632 49
<< scnmos >>
rect 84 57 114 141
rect 156 57 186 141
rect 242 57 272 141
rect 314 57 344 141
rect 512 47 542 131
rect 584 47 614 131
rect 670 47 700 131
rect 748 47 778 131
rect 850 47 880 131
rect 928 47 958 131
rect 1177 47 1207 131
rect 1249 47 1279 131
rect 1447 83 1477 167
rect 1519 83 1549 167
<< scpmoshvt >>
rect 84 409 134 609
rect 190 409 240 609
rect 509 419 559 619
rect 716 419 766 619
rect 814 419 864 619
rect 922 419 972 619
rect 1036 419 1086 619
rect 1183 419 1233 619
rect 1447 381 1497 581
<< ndiff >>
rect 27 116 84 141
rect 27 82 39 116
rect 73 82 84 116
rect 27 57 84 82
rect 114 57 156 141
rect 186 116 242 141
rect 186 82 197 116
rect 231 82 242 116
rect 186 57 242 82
rect 272 57 314 141
rect 344 116 401 141
rect 1390 142 1447 167
rect 344 82 355 116
rect 389 82 401 116
rect 344 57 401 82
rect 455 111 512 131
rect 455 77 467 111
rect 501 77 512 111
rect 455 47 512 77
rect 542 47 584 131
rect 614 106 670 131
rect 614 72 625 106
rect 659 72 670 106
rect 614 47 670 72
rect 700 47 748 131
rect 778 97 850 131
rect 778 63 805 97
rect 839 63 850 97
rect 778 47 850 63
rect 880 47 928 131
rect 958 106 1177 131
rect 958 72 1098 106
rect 1132 72 1177 106
rect 958 47 1177 72
rect 1207 47 1249 131
rect 1279 111 1336 131
rect 1279 77 1290 111
rect 1324 77 1336 111
rect 1390 108 1402 142
rect 1436 108 1447 142
rect 1390 83 1447 108
rect 1477 83 1519 167
rect 1549 142 1605 167
rect 1549 108 1560 142
rect 1594 108 1605 142
rect 1549 83 1605 108
rect 1279 47 1336 77
<< pdiff >>
rect 574 621 632 633
rect 574 619 586 621
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 596 190 609
rect 134 562 145 596
rect 179 562 190 596
rect 134 409 190 562
rect 240 455 297 609
rect 452 465 509 619
rect 240 421 251 455
rect 285 421 297 455
rect 240 409 297 421
rect 452 431 464 465
rect 498 431 509 465
rect 452 419 509 431
rect 559 587 586 619
rect 620 619 632 621
rect 620 587 716 619
rect 559 419 716 587
rect 766 419 814 619
rect 864 597 922 619
rect 864 563 877 597
rect 911 563 922 597
rect 864 465 922 563
rect 864 431 877 465
rect 911 431 922 465
rect 864 419 922 431
rect 972 419 1036 619
rect 1086 607 1183 619
rect 1086 573 1098 607
rect 1132 573 1183 607
rect 1086 536 1183 573
rect 1086 502 1098 536
rect 1132 502 1183 536
rect 1086 465 1183 502
rect 1086 431 1098 465
rect 1132 431 1183 465
rect 1086 419 1183 431
rect 1233 597 1290 619
rect 1233 563 1244 597
rect 1278 563 1290 597
rect 1233 465 1290 563
rect 1233 431 1244 465
rect 1278 431 1290 465
rect 1233 419 1290 431
rect 1390 569 1447 581
rect 1390 535 1402 569
rect 1436 535 1447 569
rect 1390 498 1447 535
rect 1390 464 1402 498
rect 1436 464 1447 498
rect 1390 427 1447 464
rect 1390 393 1402 427
rect 1436 393 1447 427
rect 1390 381 1447 393
rect 1497 569 1554 581
rect 1497 535 1508 569
rect 1542 535 1554 569
rect 1497 498 1554 535
rect 1497 464 1508 498
rect 1542 464 1554 498
rect 1497 427 1554 464
rect 1497 393 1508 427
rect 1542 393 1554 427
rect 1497 381 1554 393
<< ndiffc >>
rect 39 82 73 116
rect 197 82 231 116
rect 355 82 389 116
rect 467 77 501 111
rect 625 72 659 106
rect 805 63 839 97
rect 1098 72 1132 106
rect 1290 77 1324 111
rect 1402 108 1436 142
rect 1560 108 1594 142
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 562 179 596
rect 251 421 285 455
rect 464 431 498 465
rect 586 587 620 621
rect 877 563 911 597
rect 877 431 911 465
rect 1098 573 1132 607
rect 1098 502 1132 536
rect 1098 431 1132 465
rect 1244 563 1278 597
rect 1244 431 1278 465
rect 1402 535 1436 569
rect 1402 464 1436 498
rect 1402 393 1436 427
rect 1508 535 1542 569
rect 1508 464 1542 498
rect 1508 393 1542 427
<< poly >>
rect 84 609 134 635
rect 190 609 240 635
rect 509 619 559 645
rect 339 439 405 455
rect 84 315 134 409
rect 190 369 240 409
rect 339 405 355 439
rect 389 405 405 439
rect 716 619 766 645
rect 814 619 864 645
rect 922 619 972 645
rect 1036 619 1086 645
rect 1183 619 1233 645
rect 1447 581 1497 607
rect 339 371 405 405
rect 210 353 276 369
rect 210 319 226 353
rect 260 319 276 353
rect 339 337 355 371
rect 389 351 405 371
rect 509 387 559 419
rect 716 387 766 419
rect 509 371 616 387
rect 509 351 566 371
rect 389 337 566 351
rect 600 337 616 371
rect 339 321 616 337
rect 664 371 766 387
rect 664 337 680 371
rect 714 337 766 371
rect 664 321 766 337
rect 814 333 864 419
rect 922 379 972 419
rect 922 363 988 379
rect 84 299 159 315
rect 84 265 109 299
rect 143 265 159 299
rect 84 231 159 265
rect 210 285 276 319
rect 210 251 226 285
rect 260 265 276 285
rect 512 303 616 321
rect 512 269 566 303
rect 600 269 616 303
rect 260 251 344 265
rect 210 235 344 251
rect 84 197 109 231
rect 143 197 159 231
rect 84 187 159 197
rect 84 157 186 187
rect 84 141 114 157
rect 156 141 186 157
rect 242 141 272 235
rect 314 141 344 235
rect 512 253 616 269
rect 512 131 542 253
rect 584 131 614 253
rect 670 131 700 321
rect 814 317 880 333
rect 814 283 830 317
rect 864 283 880 317
rect 814 267 880 283
rect 742 203 808 219
rect 742 169 758 203
rect 792 169 808 203
rect 742 153 808 169
rect 748 131 778 153
rect 850 131 880 267
rect 922 329 938 363
rect 972 329 988 363
rect 922 295 988 329
rect 922 261 938 295
rect 972 261 988 295
rect 922 245 988 261
rect 1036 375 1086 419
rect 1036 359 1135 375
rect 1036 325 1085 359
rect 1119 325 1135 359
rect 1036 291 1135 325
rect 1183 305 1233 419
rect 1327 325 1393 341
rect 1036 257 1085 291
rect 1119 257 1135 291
rect 1036 241 1135 257
rect 1177 289 1243 305
rect 1177 255 1193 289
rect 1227 255 1243 289
rect 1036 176 1066 241
rect 928 146 1066 176
rect 1177 221 1243 255
rect 1177 187 1193 221
rect 1227 201 1243 221
rect 1327 291 1343 325
rect 1377 291 1393 325
rect 1327 257 1393 291
rect 1327 223 1343 257
rect 1377 237 1393 257
rect 1447 237 1497 381
rect 1377 223 1549 237
rect 1327 207 1549 223
rect 1227 187 1279 201
rect 1177 171 1279 187
rect 928 131 958 146
rect 1177 131 1207 171
rect 1249 131 1279 171
rect 1447 167 1477 207
rect 1519 167 1549 207
rect 84 31 114 57
rect 156 31 186 57
rect 242 31 272 57
rect 314 31 344 57
rect 1447 57 1477 83
rect 1519 57 1549 83
rect 512 21 542 47
rect 584 21 614 47
rect 670 21 700 47
rect 748 21 778 47
rect 850 21 880 47
rect 928 21 958 47
rect 1177 21 1207 47
rect 1249 21 1279 47
<< polycont >>
rect 355 405 389 439
rect 226 319 260 353
rect 355 337 389 371
rect 566 337 600 371
rect 680 337 714 371
rect 109 265 143 299
rect 226 251 260 285
rect 566 269 600 303
rect 109 197 143 231
rect 830 283 864 317
rect 758 169 792 203
rect 938 329 972 363
rect 938 261 972 295
rect 1085 325 1119 359
rect 1085 257 1119 291
rect 1193 255 1227 289
rect 1193 187 1227 221
rect 1343 291 1377 325
rect 1343 223 1377 257
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 526 89 563
rect 129 596 195 649
rect 129 562 145 596
rect 179 562 195 596
rect 570 621 636 649
rect 570 587 586 621
rect 620 587 636 621
rect 861 597 927 613
rect 129 561 195 562
rect 861 563 877 597
rect 911 563 927 597
rect 23 492 39 526
rect 73 525 89 526
rect 231 525 730 551
rect 73 517 730 525
rect 73 492 265 517
rect 23 491 265 492
rect 23 455 89 491
rect 448 465 514 481
rect 23 421 39 455
rect 73 421 89 455
rect 23 405 89 421
rect 235 421 251 455
rect 285 439 405 455
rect 285 421 355 439
rect 235 405 355 421
rect 389 405 405 439
rect 23 145 57 405
rect 339 371 405 405
rect 93 299 167 356
rect 93 265 109 299
rect 143 265 167 299
rect 93 231 167 265
rect 210 353 276 369
rect 210 319 226 353
rect 260 319 276 353
rect 210 285 276 319
rect 210 251 226 285
rect 260 251 276 285
rect 210 235 276 251
rect 339 337 355 371
rect 389 337 405 371
rect 93 197 109 231
rect 143 197 167 231
rect 93 181 167 197
rect 23 116 89 145
rect 23 82 39 116
rect 73 82 89 116
rect 23 53 89 82
rect 181 116 247 145
rect 181 82 197 116
rect 231 82 247 116
rect 181 17 247 82
rect 339 116 405 337
rect 339 82 355 116
rect 389 82 405 116
rect 339 53 405 82
rect 448 431 464 465
rect 498 431 514 465
rect 448 217 514 431
rect 550 371 616 387
rect 550 337 566 371
rect 600 337 616 371
rect 550 303 616 337
rect 664 371 730 517
rect 861 465 927 563
rect 861 431 877 465
rect 911 449 927 465
rect 1082 607 1148 649
rect 1082 573 1098 607
rect 1132 573 1148 607
rect 1082 536 1148 573
rect 1082 502 1098 536
rect 1132 502 1148 536
rect 1082 465 1148 502
rect 911 431 1046 449
rect 861 415 1046 431
rect 1082 431 1098 465
rect 1132 431 1148 465
rect 1082 415 1148 431
rect 1228 597 1313 613
rect 1228 563 1244 597
rect 1278 563 1313 597
rect 1228 465 1313 563
rect 1228 431 1244 465
rect 1278 431 1313 465
rect 1228 415 1313 431
rect 664 337 680 371
rect 714 337 730 371
rect 664 323 730 337
rect 922 363 976 379
rect 550 269 566 303
rect 600 287 616 303
rect 814 317 880 333
rect 814 287 830 317
rect 600 283 830 287
rect 864 283 880 317
rect 600 269 880 283
rect 550 253 880 269
rect 922 329 938 363
rect 972 329 976 363
rect 922 295 976 329
rect 922 261 938 295
rect 972 261 976 295
rect 922 217 976 261
rect 448 203 976 217
rect 448 183 758 203
rect 448 111 517 183
rect 742 169 758 183
rect 792 169 976 203
rect 742 153 976 169
rect 1012 205 1046 415
rect 1279 375 1313 415
rect 1386 569 1452 649
rect 1386 535 1402 569
rect 1436 535 1452 569
rect 1386 498 1452 535
rect 1386 464 1402 498
rect 1436 464 1452 498
rect 1386 427 1452 464
rect 1386 393 1402 427
rect 1436 393 1452 427
rect 1386 377 1452 393
rect 1492 569 1610 585
rect 1492 535 1508 569
rect 1542 535 1610 569
rect 1492 498 1610 535
rect 1492 464 1508 498
rect 1542 464 1610 498
rect 1492 427 1610 464
rect 1492 393 1508 427
rect 1542 393 1610 427
rect 1082 359 1313 375
rect 1082 325 1085 359
rect 1119 341 1313 359
rect 1119 325 1135 341
rect 1082 291 1135 325
rect 1279 325 1393 341
rect 1082 257 1085 291
rect 1119 257 1135 291
rect 1082 241 1135 257
rect 1177 289 1243 305
rect 1177 255 1193 289
rect 1227 255 1243 289
rect 1177 221 1243 255
rect 1177 205 1193 221
rect 1012 187 1193 205
rect 1227 187 1243 221
rect 1012 171 1243 187
rect 1279 291 1343 325
rect 1377 291 1393 325
rect 1279 257 1393 291
rect 1279 223 1343 257
rect 1377 223 1393 257
rect 1279 207 1393 223
rect 448 77 467 111
rect 501 77 517 111
rect 448 53 517 77
rect 609 106 675 135
rect 1012 117 1046 171
rect 1279 135 1340 207
rect 609 72 625 106
rect 659 72 675 106
rect 609 17 675 72
rect 789 97 1046 117
rect 789 63 805 97
rect 839 63 1046 97
rect 789 59 1046 63
rect 1082 106 1148 135
rect 1082 72 1098 106
rect 1132 72 1148 106
rect 1082 17 1148 72
rect 1274 111 1340 135
rect 1274 77 1290 111
rect 1324 77 1340 111
rect 1274 53 1340 77
rect 1386 142 1452 171
rect 1386 108 1402 142
rect 1436 108 1452 142
rect 1386 17 1452 108
rect 1492 142 1610 393
rect 1492 108 1560 142
rect 1594 108 1610 142
rect 1492 88 1610 108
rect 1544 79 1610 88
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlxtp_lp2
flabel comment s 469 329 469 329 0 FreeSans 200 180 0 0 no_jumper_check
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 234706
string GDS_START 223020
<< end >>
