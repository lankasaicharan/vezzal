magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 48 49 846 241
rect 0 0 864 49
<< scnmos >>
rect 131 47 161 215
rect 217 47 247 215
rect 303 47 333 215
rect 389 47 419 215
rect 475 47 505 215
rect 561 47 591 215
rect 647 47 677 215
rect 733 47 763 215
<< scpmoshvt >>
rect 131 367 161 619
rect 217 367 247 619
rect 303 367 333 619
rect 389 367 419 619
rect 475 367 505 619
rect 561 367 591 619
rect 647 367 677 619
rect 733 367 763 619
<< ndiff >>
rect 74 159 131 215
rect 74 125 86 159
rect 120 125 131 159
rect 74 91 131 125
rect 74 57 86 91
rect 120 57 131 91
rect 74 47 131 57
rect 161 185 217 215
rect 161 151 172 185
rect 206 151 217 185
rect 161 110 217 151
rect 161 76 172 110
rect 206 76 217 110
rect 161 47 217 76
rect 247 159 303 215
rect 247 125 258 159
rect 292 125 303 159
rect 247 91 303 125
rect 247 57 258 91
rect 292 57 303 91
rect 247 47 303 57
rect 333 185 389 215
rect 333 151 344 185
rect 378 151 389 185
rect 333 110 389 151
rect 333 76 344 110
rect 378 76 389 110
rect 333 47 389 76
rect 419 114 475 215
rect 419 80 430 114
rect 464 80 475 114
rect 419 47 475 80
rect 505 185 561 215
rect 505 151 516 185
rect 550 151 561 185
rect 505 110 561 151
rect 505 76 516 110
rect 550 76 561 110
rect 505 47 561 76
rect 591 159 647 215
rect 591 125 602 159
rect 636 125 647 159
rect 591 91 647 125
rect 591 57 602 91
rect 636 57 647 91
rect 591 47 647 57
rect 677 185 733 215
rect 677 151 688 185
rect 722 151 733 185
rect 677 110 733 151
rect 677 76 688 110
rect 722 76 733 110
rect 677 47 733 76
rect 763 159 820 215
rect 763 125 774 159
rect 808 125 820 159
rect 763 91 820 125
rect 763 57 774 91
rect 808 57 820 91
rect 763 47 820 57
<< pdiff >>
rect 74 607 131 619
rect 74 573 86 607
rect 120 573 131 607
rect 74 539 131 573
rect 74 505 86 539
rect 120 505 131 539
rect 74 471 131 505
rect 74 437 86 471
rect 120 437 131 471
rect 74 367 131 437
rect 161 589 217 619
rect 161 555 172 589
rect 206 555 217 589
rect 161 510 217 555
rect 161 476 172 510
rect 206 476 217 510
rect 161 431 217 476
rect 161 397 172 431
rect 206 397 217 431
rect 161 367 217 397
rect 247 605 303 619
rect 247 571 258 605
rect 292 571 303 605
rect 247 537 303 571
rect 247 503 258 537
rect 292 503 303 537
rect 247 469 303 503
rect 247 435 258 469
rect 292 435 303 469
rect 247 367 303 435
rect 333 589 389 619
rect 333 555 344 589
rect 378 555 389 589
rect 333 510 389 555
rect 333 476 344 510
rect 378 476 389 510
rect 333 431 389 476
rect 333 397 344 431
rect 378 397 389 431
rect 333 367 389 397
rect 419 605 475 619
rect 419 571 430 605
rect 464 571 475 605
rect 419 537 475 571
rect 419 503 430 537
rect 464 503 475 537
rect 419 469 475 503
rect 419 435 430 469
rect 464 435 475 469
rect 419 367 475 435
rect 505 589 561 619
rect 505 555 516 589
rect 550 555 561 589
rect 505 510 561 555
rect 505 476 516 510
rect 550 476 561 510
rect 505 431 561 476
rect 505 397 516 431
rect 550 397 561 431
rect 505 367 561 397
rect 591 605 647 619
rect 591 571 602 605
rect 636 571 647 605
rect 591 537 647 571
rect 591 503 602 537
rect 636 503 647 537
rect 591 469 647 503
rect 591 435 602 469
rect 636 435 647 469
rect 591 367 647 435
rect 677 589 733 619
rect 677 555 688 589
rect 722 555 733 589
rect 677 510 733 555
rect 677 476 688 510
rect 722 476 733 510
rect 677 431 733 476
rect 677 397 688 431
rect 722 397 733 431
rect 677 367 733 397
rect 763 605 820 619
rect 763 571 774 605
rect 808 571 820 605
rect 763 537 820 571
rect 763 503 774 537
rect 808 503 820 537
rect 763 469 820 503
rect 763 435 774 469
rect 808 435 820 469
rect 763 367 820 435
<< ndiffc >>
rect 86 125 120 159
rect 86 57 120 91
rect 172 151 206 185
rect 172 76 206 110
rect 258 125 292 159
rect 258 57 292 91
rect 344 151 378 185
rect 344 76 378 110
rect 430 80 464 114
rect 516 151 550 185
rect 516 76 550 110
rect 602 125 636 159
rect 602 57 636 91
rect 688 151 722 185
rect 688 76 722 110
rect 774 125 808 159
rect 774 57 808 91
<< pdiffc >>
rect 86 573 120 607
rect 86 505 120 539
rect 86 437 120 471
rect 172 555 206 589
rect 172 476 206 510
rect 172 397 206 431
rect 258 571 292 605
rect 258 503 292 537
rect 258 435 292 469
rect 344 555 378 589
rect 344 476 378 510
rect 344 397 378 431
rect 430 571 464 605
rect 430 503 464 537
rect 430 435 464 469
rect 516 555 550 589
rect 516 476 550 510
rect 516 397 550 431
rect 602 571 636 605
rect 602 503 636 537
rect 602 435 636 469
rect 688 555 722 589
rect 688 476 722 510
rect 688 397 722 431
rect 774 571 808 605
rect 774 503 808 537
rect 774 435 808 469
<< poly >>
rect 131 619 161 645
rect 217 619 247 645
rect 303 619 333 645
rect 389 619 419 645
rect 475 619 505 645
rect 561 619 591 645
rect 647 619 677 645
rect 733 619 763 645
rect 131 329 161 367
rect 217 329 247 367
rect 303 329 333 367
rect 389 329 419 367
rect 475 329 505 367
rect 561 329 591 367
rect 647 329 677 367
rect 733 329 763 367
rect 85 313 763 329
rect 85 279 101 313
rect 135 279 169 313
rect 203 279 237 313
rect 271 279 305 313
rect 339 279 373 313
rect 407 279 441 313
rect 475 279 509 313
rect 543 279 577 313
rect 611 279 645 313
rect 679 279 713 313
rect 747 279 763 313
rect 85 263 763 279
rect 131 215 161 263
rect 217 215 247 263
rect 303 215 333 263
rect 389 215 419 263
rect 475 215 505 263
rect 561 215 591 263
rect 647 215 677 263
rect 733 215 763 263
rect 131 21 161 47
rect 217 21 247 47
rect 303 21 333 47
rect 389 21 419 47
rect 475 21 505 47
rect 561 21 591 47
rect 647 21 677 47
rect 733 21 763 47
<< polycont >>
rect 101 279 135 313
rect 169 279 203 313
rect 237 279 271 313
rect 305 279 339 313
rect 373 279 407 313
rect 441 279 475 313
rect 509 279 543 313
rect 577 279 611 313
rect 645 279 679 313
rect 713 279 747 313
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 70 607 129 649
rect 70 573 86 607
rect 120 573 129 607
rect 70 539 129 573
rect 70 505 86 539
rect 120 505 129 539
rect 70 471 129 505
rect 70 437 86 471
rect 120 437 129 471
rect 70 421 129 437
rect 163 589 215 615
rect 163 555 172 589
rect 206 555 215 589
rect 163 510 215 555
rect 163 476 172 510
rect 206 476 215 510
rect 163 431 215 476
rect 163 397 172 431
rect 206 397 215 431
rect 249 605 301 649
rect 249 571 258 605
rect 292 571 301 605
rect 249 537 301 571
rect 249 503 258 537
rect 292 503 301 537
rect 249 469 301 503
rect 249 435 258 469
rect 292 435 301 469
rect 249 419 301 435
rect 335 589 387 615
rect 335 555 344 589
rect 378 555 387 589
rect 335 510 387 555
rect 335 476 344 510
rect 378 476 387 510
rect 335 431 387 476
rect 163 385 215 397
rect 335 397 344 431
rect 378 397 387 431
rect 421 605 473 649
rect 421 571 430 605
rect 464 571 473 605
rect 421 537 473 571
rect 421 503 430 537
rect 464 503 473 537
rect 421 469 473 503
rect 421 435 430 469
rect 464 435 473 469
rect 421 419 473 435
rect 507 589 559 615
rect 507 555 516 589
rect 550 555 559 589
rect 507 510 559 555
rect 507 476 516 510
rect 550 476 559 510
rect 507 431 559 476
rect 335 385 387 397
rect 507 397 516 431
rect 550 397 559 431
rect 593 605 645 649
rect 593 571 602 605
rect 636 571 645 605
rect 593 537 645 571
rect 593 503 602 537
rect 636 503 645 537
rect 593 469 645 503
rect 593 435 602 469
rect 636 435 645 469
rect 593 419 645 435
rect 679 589 731 615
rect 679 555 688 589
rect 722 555 731 589
rect 679 510 731 555
rect 679 476 688 510
rect 722 476 731 510
rect 679 431 731 476
rect 507 385 559 397
rect 679 397 688 431
rect 722 397 731 431
rect 765 605 824 649
rect 765 571 774 605
rect 808 571 824 605
rect 765 537 824 571
rect 765 503 774 537
rect 808 503 824 537
rect 765 469 824 503
rect 765 435 774 469
rect 808 435 824 469
rect 765 419 824 435
rect 679 385 731 397
rect 17 351 845 385
rect 17 243 51 351
rect 85 313 763 317
rect 85 279 101 313
rect 135 279 169 313
rect 203 279 237 313
rect 271 279 305 313
rect 339 279 373 313
rect 407 279 441 313
rect 475 279 509 313
rect 543 279 577 313
rect 611 279 645 313
rect 679 279 713 313
rect 747 279 763 313
rect 412 277 763 279
rect 17 209 378 243
rect 412 232 473 277
rect 797 243 845 351
rect 163 185 215 209
rect 70 159 129 175
rect 70 125 86 159
rect 120 125 129 159
rect 70 91 129 125
rect 70 57 86 91
rect 120 57 129 91
rect 70 17 129 57
rect 163 151 172 185
rect 206 151 215 185
rect 335 198 378 209
rect 507 209 845 243
rect 507 198 559 209
rect 335 185 559 198
rect 163 110 215 151
rect 163 76 172 110
rect 206 76 215 110
rect 163 51 215 76
rect 249 159 301 175
rect 249 125 258 159
rect 292 125 301 159
rect 249 91 301 125
rect 249 57 258 91
rect 292 57 301 91
rect 249 17 301 57
rect 335 151 344 185
rect 378 164 516 185
rect 378 151 387 164
rect 335 110 387 151
rect 507 151 516 164
rect 550 151 559 185
rect 679 185 731 209
rect 335 76 344 110
rect 378 76 387 110
rect 335 51 387 76
rect 421 114 473 130
rect 421 80 430 114
rect 464 80 473 114
rect 421 17 473 80
rect 507 110 559 151
rect 507 76 516 110
rect 550 76 559 110
rect 507 51 559 76
rect 593 159 645 175
rect 593 125 602 159
rect 636 125 645 159
rect 593 91 645 125
rect 593 57 602 91
rect 636 57 645 91
rect 593 17 645 57
rect 679 151 688 185
rect 722 151 731 185
rect 679 110 731 151
rect 679 76 688 110
rect 722 76 731 110
rect 679 51 731 76
rect 765 159 824 175
rect 765 125 774 159
rect 808 125 824 159
rect 765 91 824 125
rect 765 57 774 91
rect 808 57 824 91
rect 765 17 824 57
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 inv_8
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4486962
string GDS_START 4479180
<< end >>
