magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 352 2150 704
rect -38 332 1382 352
rect 1655 332 2150 352
<< pwell >>
rect 1424 275 1613 294
rect 1424 274 1728 275
rect 1424 248 2104 274
rect 5 49 2104 248
rect 0 0 2112 49
<< scpmos >>
rect 111 392 147 592
rect 231 392 267 592
rect 441 392 477 592
rect 585 392 621 592
rect 669 392 705 592
rect 807 392 843 592
rect 981 392 1017 592
rect 1119 392 1155 592
rect 1203 392 1239 592
rect 1410 392 1446 592
rect 1500 392 1536 592
rect 1727 388 1763 588
rect 1904 368 1940 592
rect 1994 368 2030 592
<< nmoslvt >>
rect 88 94 118 222
rect 225 74 255 222
rect 303 74 333 222
rect 477 74 507 222
rect 663 74 693 222
rect 801 74 831 222
rect 879 74 909 222
rect 1017 74 1047 222
rect 1203 74 1233 222
rect 1399 74 1429 222
rect 1500 120 1530 268
rect 1727 120 1757 248
rect 1905 100 1935 248
rect 1991 100 2021 248
<< ndiff >>
rect 1450 222 1500 268
rect 31 167 88 222
rect 31 133 43 167
rect 77 133 88 167
rect 31 94 88 133
rect 118 188 225 222
rect 118 154 180 188
rect 214 154 225 188
rect 118 120 225 154
rect 118 94 180 120
rect 168 86 180 94
rect 214 86 225 120
rect 168 74 225 86
rect 255 74 303 222
rect 333 202 477 222
rect 333 168 399 202
rect 433 168 477 202
rect 333 74 477 168
rect 507 74 663 222
rect 693 188 801 222
rect 693 154 713 188
rect 747 154 801 188
rect 693 120 801 154
rect 693 86 713 120
rect 747 86 801 120
rect 693 74 801 86
rect 831 74 879 222
rect 909 188 1017 222
rect 909 154 954 188
rect 988 154 1017 188
rect 909 120 1017 154
rect 909 86 954 120
rect 988 86 1017 120
rect 909 74 1017 86
rect 1047 74 1203 222
rect 1233 120 1289 222
rect 1233 86 1244 120
rect 1278 86 1289 120
rect 1233 74 1289 86
rect 1343 188 1399 222
rect 1343 154 1354 188
rect 1388 154 1399 188
rect 1343 120 1399 154
rect 1343 86 1354 120
rect 1388 86 1399 120
rect 1343 74 1399 86
rect 1429 120 1500 222
rect 1530 256 1587 268
rect 1530 222 1541 256
rect 1575 222 1587 256
rect 1530 120 1587 222
rect 1641 248 1702 249
rect 1641 237 1727 248
rect 1641 203 1654 237
rect 1688 203 1727 237
rect 1641 120 1727 203
rect 1757 220 1905 248
rect 1757 186 1860 220
rect 1894 186 1905 220
rect 1757 152 1905 186
rect 1757 120 1860 152
rect 1429 86 1440 120
rect 1474 86 1485 120
rect 1429 74 1485 86
rect 1848 118 1860 120
rect 1894 118 1905 152
rect 1848 100 1905 118
rect 1935 236 1991 248
rect 1935 202 1946 236
rect 1980 202 1991 236
rect 1935 146 1991 202
rect 1935 112 1946 146
rect 1980 112 1991 146
rect 1935 100 1991 112
rect 2021 236 2078 248
rect 2021 202 2032 236
rect 2066 202 2078 236
rect 2021 146 2078 202
rect 2021 112 2032 146
rect 2066 112 2078 146
rect 2021 100 2078 112
<< pdiff >>
rect 55 580 111 592
rect 55 546 67 580
rect 101 546 111 580
rect 55 509 111 546
rect 55 475 67 509
rect 101 475 111 509
rect 55 438 111 475
rect 55 404 67 438
rect 101 404 111 438
rect 55 392 111 404
rect 147 580 231 592
rect 147 546 167 580
rect 201 546 231 580
rect 147 510 231 546
rect 147 476 167 510
rect 201 476 231 510
rect 147 440 231 476
rect 147 406 167 440
rect 201 406 231 440
rect 147 392 231 406
rect 267 392 441 592
rect 477 580 585 592
rect 477 546 515 580
rect 549 546 585 580
rect 477 510 585 546
rect 477 476 515 510
rect 549 476 585 510
rect 477 440 585 476
rect 477 406 515 440
rect 549 406 585 440
rect 477 392 585 406
rect 621 392 669 592
rect 705 580 807 592
rect 705 546 739 580
rect 773 546 807 580
rect 705 508 807 546
rect 705 474 739 508
rect 773 474 807 508
rect 705 392 807 474
rect 843 392 981 592
rect 1017 566 1119 592
rect 1017 532 1051 566
rect 1085 532 1119 566
rect 1017 392 1119 532
rect 1155 392 1203 592
rect 1239 578 1295 592
rect 1239 544 1249 578
rect 1283 544 1295 578
rect 1239 392 1295 544
rect 1349 440 1410 592
rect 1349 406 1363 440
rect 1397 406 1410 440
rect 1349 392 1410 406
rect 1446 578 1500 592
rect 1446 544 1456 578
rect 1490 544 1500 578
rect 1446 392 1500 544
rect 1536 508 1591 592
rect 1854 588 1904 592
rect 1536 474 1546 508
rect 1580 474 1591 508
rect 1536 440 1591 474
rect 1536 406 1546 440
rect 1580 406 1591 440
rect 1536 392 1591 406
rect 1645 448 1727 588
rect 1645 414 1656 448
rect 1690 414 1727 448
rect 1645 388 1727 414
rect 1763 576 1904 588
rect 1763 542 1860 576
rect 1894 542 1904 576
rect 1763 498 1904 542
rect 1763 464 1860 498
rect 1894 464 1904 498
rect 1763 420 1904 464
rect 1763 388 1860 420
rect 1848 386 1860 388
rect 1894 386 1904 420
rect 1848 368 1904 386
rect 1940 580 1994 592
rect 1940 546 1950 580
rect 1984 546 1994 580
rect 1940 497 1994 546
rect 1940 463 1950 497
rect 1984 463 1994 497
rect 1940 414 1994 463
rect 1940 380 1950 414
rect 1984 380 1994 414
rect 1940 368 1994 380
rect 2030 580 2085 592
rect 2030 546 2040 580
rect 2074 546 2085 580
rect 2030 497 2085 546
rect 2030 463 2040 497
rect 2074 463 2085 497
rect 2030 414 2085 463
rect 2030 380 2040 414
rect 2074 380 2085 414
rect 2030 368 2085 380
<< ndiffc >>
rect 43 133 77 167
rect 180 154 214 188
rect 180 86 214 120
rect 399 168 433 202
rect 713 154 747 188
rect 713 86 747 120
rect 954 154 988 188
rect 954 86 988 120
rect 1244 86 1278 120
rect 1354 154 1388 188
rect 1354 86 1388 120
rect 1541 222 1575 256
rect 1654 203 1688 237
rect 1860 186 1894 220
rect 1440 86 1474 120
rect 1860 118 1894 152
rect 1946 202 1980 236
rect 1946 112 1980 146
rect 2032 202 2066 236
rect 2032 112 2066 146
<< pdiffc >>
rect 67 546 101 580
rect 67 475 101 509
rect 67 404 101 438
rect 167 546 201 580
rect 167 476 201 510
rect 167 406 201 440
rect 515 546 549 580
rect 515 476 549 510
rect 515 406 549 440
rect 739 546 773 580
rect 739 474 773 508
rect 1051 532 1085 566
rect 1249 544 1283 578
rect 1363 406 1397 440
rect 1456 544 1490 578
rect 1546 474 1580 508
rect 1546 406 1580 440
rect 1656 414 1690 448
rect 1860 542 1894 576
rect 1860 464 1894 498
rect 1860 386 1894 420
rect 1950 546 1984 580
rect 1950 463 1984 497
rect 1950 380 1984 414
rect 2040 546 2074 580
rect 2040 463 2074 497
rect 2040 380 2074 414
<< poly >>
rect 111 592 147 618
rect 231 592 267 618
rect 441 592 477 618
rect 585 592 621 618
rect 669 592 705 618
rect 807 592 843 618
rect 981 592 1017 618
rect 1119 592 1155 618
rect 1203 592 1239 618
rect 1410 592 1446 618
rect 1500 592 1536 618
rect 1727 588 1763 614
rect 1904 592 1940 618
rect 1994 592 2030 618
rect 111 310 147 392
rect 231 356 267 392
rect 441 356 477 392
rect 585 356 621 392
rect 669 356 705 392
rect 807 358 843 392
rect 981 358 1017 392
rect 807 356 837 358
rect 195 346 267 356
rect 195 340 261 346
rect 87 294 153 310
rect 87 260 103 294
rect 137 260 153 294
rect 195 306 211 340
rect 245 306 261 340
rect 411 340 477 356
rect 195 290 261 306
rect 303 302 369 318
rect 87 244 153 260
rect 88 222 118 244
rect 225 222 255 290
rect 303 268 319 302
rect 353 268 369 302
rect 411 306 427 340
rect 461 320 477 340
rect 555 340 621 356
rect 461 306 507 320
rect 411 290 507 306
rect 555 306 571 340
rect 605 306 621 340
rect 555 290 621 306
rect 663 340 729 356
rect 663 306 679 340
rect 713 306 729 340
rect 303 252 369 268
rect 303 222 333 252
rect 477 222 507 290
rect 663 248 729 306
rect 771 340 837 356
rect 771 306 787 340
rect 821 306 837 340
rect 987 342 1053 358
rect 1119 350 1155 392
rect 771 290 837 306
rect 879 294 945 310
rect 663 222 693 248
rect 801 222 831 290
rect 879 260 895 294
rect 929 260 945 294
rect 987 308 1003 342
rect 1037 308 1053 342
rect 987 292 1053 308
rect 1095 334 1161 350
rect 1095 300 1111 334
rect 1145 300 1161 334
rect 879 244 945 260
rect 879 222 909 244
rect 1017 222 1047 292
rect 1095 284 1161 300
rect 1203 310 1239 392
rect 1410 356 1446 392
rect 1380 340 1446 356
rect 1203 294 1269 310
rect 1203 260 1219 294
rect 1253 260 1269 294
rect 1380 306 1396 340
rect 1430 306 1446 340
rect 1380 290 1446 306
rect 1500 356 1536 392
rect 1500 340 1679 356
rect 1500 306 1561 340
rect 1595 306 1629 340
rect 1663 306 1679 340
rect 1500 290 1679 306
rect 1203 244 1269 260
rect 1203 222 1233 244
rect 1399 222 1429 290
rect 1500 268 1530 290
rect 88 68 118 94
rect 1727 263 1763 388
rect 1904 336 1940 368
rect 1811 330 1940 336
rect 1994 330 2030 368
rect 1811 320 2030 330
rect 1811 286 1827 320
rect 1861 300 2030 320
rect 1861 286 2021 300
rect 1811 270 2021 286
rect 1727 248 1757 263
rect 1905 248 1935 270
rect 1991 248 2021 270
rect 1500 94 1530 120
rect 225 48 255 74
rect 303 48 333 74
rect 477 48 507 74
rect 663 48 693 74
rect 801 48 831 74
rect 879 48 909 74
rect 1017 48 1047 74
rect 1203 48 1233 74
rect 1399 52 1429 74
rect 1727 52 1757 120
rect 1905 74 1935 100
rect 1991 74 2021 100
rect 1399 22 1757 52
<< polycont >>
rect 103 260 137 294
rect 211 306 245 340
rect 319 268 353 302
rect 427 306 461 340
rect 571 306 605 340
rect 679 306 713 340
rect 787 306 821 340
rect 895 260 929 294
rect 1003 308 1037 342
rect 1111 300 1145 334
rect 1219 260 1253 294
rect 1396 306 1430 340
rect 1561 306 1595 340
rect 1629 306 1663 340
rect 1827 286 1861 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 51 580 117 596
rect 51 546 67 580
rect 101 546 117 580
rect 51 509 117 546
rect 51 475 67 509
rect 101 475 117 509
rect 51 438 117 475
rect 51 430 67 438
rect 19 424 67 430
rect 19 390 31 424
rect 65 404 67 424
rect 101 404 117 438
rect 65 390 117 404
rect 151 580 217 649
rect 151 546 167 580
rect 201 546 217 580
rect 151 510 217 546
rect 151 476 167 510
rect 201 476 217 510
rect 151 440 217 476
rect 151 406 167 440
rect 201 406 217 440
rect 499 580 689 596
rect 499 546 515 580
rect 549 546 689 580
rect 499 510 689 546
rect 499 476 515 510
rect 549 476 689 510
rect 499 440 689 476
rect 723 580 789 649
rect 723 546 739 580
rect 773 546 789 580
rect 723 508 789 546
rect 1011 566 1189 582
rect 1011 532 1051 566
rect 1085 532 1189 566
rect 1233 578 1299 649
rect 1233 544 1249 578
rect 1283 544 1299 578
rect 1233 542 1299 544
rect 1440 581 1826 615
rect 1440 578 1506 581
rect 1440 544 1456 578
rect 1490 544 1506 578
rect 1440 542 1506 544
rect 723 474 739 508
rect 773 474 789 508
rect 1155 508 1189 532
rect 1562 513 1758 547
rect 1562 508 1596 513
rect 723 458 789 474
rect 823 464 1121 498
rect 1155 474 1546 508
rect 1580 474 1596 508
rect 151 390 217 406
rect 409 424 465 430
rect 409 390 415 424
rect 449 390 465 424
rect 19 384 117 390
rect 19 202 53 384
rect 195 340 263 356
rect 87 294 161 310
rect 87 260 103 294
rect 137 260 161 294
rect 195 306 211 340
rect 245 306 263 340
rect 409 340 465 390
rect 195 290 263 306
rect 297 302 369 318
rect 87 256 161 260
rect 297 268 319 302
rect 353 268 369 302
rect 409 306 427 340
rect 461 306 465 340
rect 409 290 465 306
rect 499 406 515 440
rect 549 424 689 440
rect 823 424 857 464
rect 1087 440 1121 464
rect 1530 440 1596 474
rect 549 406 857 424
rect 499 390 857 406
rect 985 424 1053 430
rect 985 390 991 424
rect 1025 390 1053 424
rect 1087 406 1363 440
rect 1397 406 1416 440
rect 1087 392 1416 406
rect 297 256 369 268
rect 87 252 369 256
rect 87 236 331 252
rect 127 222 331 236
rect 19 167 93 202
rect 19 133 43 167
rect 77 133 93 167
rect 19 100 93 133
rect 164 154 180 188
rect 214 154 230 188
rect 164 120 230 154
rect 164 86 180 120
rect 214 86 230 120
rect 164 17 230 86
rect 297 118 331 222
rect 499 218 533 390
rect 370 202 533 218
rect 370 168 399 202
rect 433 168 533 202
rect 370 152 533 168
rect 567 340 621 356
rect 567 306 571 340
rect 605 306 621 340
rect 567 256 621 306
rect 663 340 737 356
rect 663 306 679 340
rect 713 306 737 340
rect 663 290 737 306
rect 771 340 839 356
rect 771 306 787 340
rect 821 306 839 340
rect 985 342 1053 390
rect 1312 390 1416 392
rect 1530 406 1546 440
rect 1580 406 1596 440
rect 1530 390 1596 406
rect 1640 448 1690 479
rect 1640 414 1656 448
rect 771 290 839 306
rect 879 294 945 310
rect 879 260 895 294
rect 929 260 945 294
rect 985 308 1003 342
rect 1037 308 1053 342
rect 985 292 1053 308
rect 1095 334 1149 350
rect 1095 300 1111 334
rect 1145 300 1149 334
rect 879 256 945 260
rect 1095 256 1149 300
rect 567 222 1149 256
rect 1183 294 1269 356
rect 1183 260 1219 294
rect 1253 260 1269 294
rect 1183 236 1269 260
rect 1312 256 1346 390
rect 1640 356 1690 414
rect 1380 340 1511 356
rect 1380 306 1396 340
rect 1430 306 1511 340
rect 1380 290 1511 306
rect 1545 340 1690 356
rect 1545 306 1561 340
rect 1595 306 1629 340
rect 1663 306 1690 340
rect 1545 290 1690 306
rect 1312 222 1541 256
rect 1575 222 1591 256
rect 1637 237 1690 290
rect 567 118 621 222
rect 1637 203 1654 237
rect 1688 203 1690 237
rect 297 84 621 118
rect 689 154 713 188
rect 747 154 785 188
rect 689 120 785 154
rect 689 86 713 120
rect 747 86 785 120
rect 689 17 785 86
rect 906 154 954 188
rect 988 154 1354 188
rect 1388 154 1603 188
rect 1637 187 1690 203
rect 906 120 1021 154
rect 1338 120 1388 154
rect 1569 153 1603 154
rect 1724 153 1758 513
rect 906 86 954 120
rect 988 86 1021 120
rect 906 70 1021 86
rect 1228 86 1244 120
rect 1278 86 1294 120
rect 1228 17 1294 86
rect 1338 86 1354 120
rect 1338 70 1388 86
rect 1424 86 1440 120
rect 1474 86 1490 120
rect 1569 119 1758 153
rect 1792 336 1826 581
rect 1860 576 1894 649
rect 1860 498 1894 542
rect 1860 420 1894 464
rect 1860 370 1894 386
rect 1930 580 2000 596
rect 1930 546 1950 580
rect 1984 546 2000 580
rect 1930 497 2000 546
rect 1930 463 1950 497
rect 1984 463 2000 497
rect 1930 414 2000 463
rect 1930 380 1950 414
rect 1984 380 2000 414
rect 1930 364 2000 380
rect 2040 580 2090 649
rect 2074 546 2090 580
rect 2040 497 2090 546
rect 2074 463 2090 497
rect 2040 414 2090 463
rect 2074 380 2090 414
rect 2040 364 2090 380
rect 1792 320 1877 336
rect 1792 286 1827 320
rect 1861 286 1877 320
rect 1792 270 1877 286
rect 1424 85 1490 86
rect 1792 85 1826 270
rect 1930 236 1996 364
rect 1424 51 1826 85
rect 1860 220 1894 236
rect 1860 152 1894 186
rect 1860 17 1894 118
rect 1930 202 1946 236
rect 1980 202 1996 236
rect 1930 146 1996 202
rect 1930 112 1946 146
rect 1980 112 1996 146
rect 1930 88 1996 112
rect 2032 236 2082 252
rect 2066 202 2082 236
rect 2032 146 2082 202
rect 2066 112 2082 146
rect 2032 17 2082 112
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 390 65 424
rect 415 390 449 424
rect 991 390 1025 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 19 424 77 430
rect 19 390 31 424
rect 65 421 77 424
rect 403 424 461 430
rect 403 421 415 424
rect 65 393 415 421
rect 65 390 77 393
rect 19 384 77 390
rect 403 390 415 393
rect 449 421 461 424
rect 979 424 1037 430
rect 979 421 991 424
rect 449 393 991 421
rect 449 390 461 393
rect 403 384 461 390
rect 979 390 991 393
rect 1025 390 1037 424
rect 979 384 1037 390
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux4_2
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 1951 94 1985 128 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 168 1985 202 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 390 1985 424 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 464 1985 498 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 538 1985 572 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 482396
string GDS_START 467340
<< end >>
