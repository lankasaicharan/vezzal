magic
tech sky130A
timestamp 1627202621
<< checkpaint >>
rect -649 -654 23189 1198
use sky130_fd_sc_hdll__muxb4to1_1  sky130_fd_sc_hdll__muxb4to1_1_0
timestamp 1627202621
transform 1 0 1564 0 1 0
box -19 -24 893 296
use sky130_fd_sc_hdll__muxb4to1_2  sky130_fd_sc_hdll__muxb4to1_2_0
timestamp 1627202621
transform 1 0 2438 0 1 0
box -19 -24 1307 296
use sky130_fd_sc_hdll__muxb4to1_4  sky130_fd_sc_hdll__muxb4to1_4_0
timestamp 1627202621
transform 1 0 3726 0 1 0
box -19 -24 2595 296
use sky130_fd_sc_hdll__muxb8to1_1  sky130_fd_sc_hdll__muxb8to1_1_0
timestamp 1627202621
transform 1 0 6302 0 1 0
box -19 -24 1721 296
use sky130_fd_sc_hdll__muxb16to1_1  sky130_fd_sc_hdll__muxb16to1_1_0
timestamp 1627202621
transform 1 0 13064 0 1 0
box -19 -24 1721 568
use sky130_fd_sc_hdll__muxb8to1_2  sky130_fd_sc_hdll__muxb8to1_2_0
timestamp 1627202621
transform 1 0 8004 0 1 0
box -19 -24 2595 296
use sky130_fd_sc_hdll__muxb8to1_4  sky130_fd_sc_hdll__muxb8to1_4_0
timestamp 1627202621
transform 1 0 10580 0 1 0
box -19 -24 2503 568
use sky130_fd_sc_hdll__muxb16to1_2  sky130_fd_sc_hdll__muxb16to1_2_0
timestamp 1627202621
transform 1 0 14766 0 1 0
box -19 -24 2595 568
use sky130_fd_sc_hdll__muxb16to1_4  sky130_fd_sc_hdll__muxb16to1_4_0
timestamp 1627202621
transform 1 0 17342 0 1 0
box -19 -24 5217 568
use sky130_fd_sc_hdll__clkmux2_1  sky130_fd_sc_hdll__clkmux2_1_0
timestamp 1627202621
transform 1 0 0 0 1 0
box -19 -24 479 296
use sky130_fd_sc_hdll__clkmux2_2  sky130_fd_sc_hdll__clkmux2_2_0
timestamp 1627202621
transform 1 0 460 0 1 0
box -19 -24 525 296
use sky130_fd_sc_hdll__clkmux2_4  sky130_fd_sc_hdll__clkmux2_4_0
timestamp 1627202621
transform 1 0 966 0 1 0
box -19 -24 617 296
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX -19 -24 22559 568
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string GDS_END 3646992
string GDS_START 3646346
<< end >>
