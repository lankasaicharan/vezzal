magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4850 1975
<< nwell >>
rect -38 331 3590 704
<< pwell >>
rect 964 241 1068 271
rect 559 211 1194 241
rect 377 195 1194 211
rect 88 157 1194 195
rect 1425 201 1916 241
rect 1425 157 3292 201
rect 88 49 3292 157
rect 0 0 3552 49
<< scnmos >>
rect 171 85 201 169
rect 273 85 303 169
rect 351 85 381 169
rect 696 47 726 215
rect 782 47 812 215
rect 938 47 968 215
rect 1064 47 1094 215
rect 1208 47 1238 131
rect 1308 47 1338 131
rect 1508 47 1538 215
rect 1594 47 1624 215
rect 1696 47 1726 215
rect 1798 47 1828 215
rect 2061 47 2091 175
rect 2147 47 2177 175
rect 2233 47 2263 175
rect 2319 47 2349 175
rect 2405 47 2435 175
rect 2491 47 2521 175
rect 2577 47 2607 175
rect 2663 47 2693 175
rect 2749 47 2779 175
rect 2835 47 2865 175
rect 2921 47 2951 175
rect 3007 47 3037 175
rect 3093 47 3123 175
rect 3179 47 3209 175
<< scpmos >>
rect 81 367 111 535
rect 187 367 217 619
rect 273 367 303 619
rect 375 451 405 619
rect 461 451 491 619
rect 720 367 750 619
rect 806 367 836 619
rect 908 367 938 619
rect 994 367 1024 619
rect 1230 373 1260 541
rect 1308 373 1338 541
rect 1514 367 1544 619
rect 1600 367 1630 619
rect 1803 367 1833 619
rect 1889 367 1919 619
rect 1975 367 2005 619
rect 2061 367 2091 619
rect 2147 367 2177 619
rect 2233 367 2263 619
rect 2319 367 2349 619
rect 2405 367 2435 619
rect 2491 367 2521 619
rect 2577 367 2607 619
rect 2663 367 2693 619
rect 2749 367 2779 619
rect 2835 367 2865 619
rect 2921 367 2951 619
rect 3007 367 3037 619
rect 3093 367 3123 619
rect 3179 367 3209 619
rect 3265 367 3295 619
rect 3351 367 3381 619
rect 3437 367 3467 619
<< ndiff >>
rect 990 233 1042 245
rect 990 215 999 233
rect 403 173 461 185
rect 403 169 415 173
rect 114 139 171 169
rect 114 105 126 139
rect 160 105 171 139
rect 114 85 171 105
rect 201 139 273 169
rect 201 105 228 139
rect 262 105 273 139
rect 201 85 273 105
rect 303 85 351 169
rect 381 139 415 169
rect 449 139 461 173
rect 381 85 461 139
rect 585 105 696 215
rect 585 71 597 105
rect 631 71 696 105
rect 585 47 696 71
rect 726 188 782 215
rect 726 154 737 188
rect 771 154 782 188
rect 726 47 782 154
rect 812 93 938 215
rect 812 59 893 93
rect 927 59 938 93
rect 812 47 938 59
rect 968 199 999 215
rect 1033 215 1042 233
rect 1033 199 1064 215
rect 968 47 1064 199
rect 1094 131 1168 215
rect 1094 77 1208 131
rect 1094 47 1125 77
rect 1116 43 1125 47
rect 1159 47 1208 77
rect 1238 111 1308 131
rect 1238 77 1249 111
rect 1283 77 1308 111
rect 1238 47 1308 77
rect 1338 93 1397 131
rect 1338 59 1351 93
rect 1385 59 1397 93
rect 1338 47 1397 59
rect 1451 93 1508 215
rect 1451 59 1463 93
rect 1497 59 1508 93
rect 1451 47 1508 59
rect 1538 113 1594 215
rect 1538 79 1549 113
rect 1583 79 1594 113
rect 1538 47 1594 79
rect 1624 203 1696 215
rect 1624 169 1651 203
rect 1685 169 1696 203
rect 1624 103 1696 169
rect 1624 69 1651 103
rect 1685 69 1696 103
rect 1624 47 1696 69
rect 1726 180 1798 215
rect 1726 146 1753 180
rect 1787 146 1798 180
rect 1726 47 1798 146
rect 1828 203 1890 215
rect 1828 169 1844 203
rect 1878 169 1890 203
rect 1828 103 1890 169
rect 1828 69 1844 103
rect 1878 69 1890 103
rect 1828 47 1890 69
rect 2004 157 2061 175
rect 2004 123 2016 157
rect 2050 123 2061 157
rect 2004 89 2061 123
rect 2004 55 2016 89
rect 2050 55 2061 89
rect 2004 47 2061 55
rect 2091 157 2147 175
rect 2091 123 2102 157
rect 2136 123 2147 157
rect 2091 89 2147 123
rect 2091 55 2102 89
rect 2136 55 2147 89
rect 2091 47 2147 55
rect 2177 157 2233 175
rect 2177 123 2188 157
rect 2222 123 2233 157
rect 2177 89 2233 123
rect 2177 55 2188 89
rect 2222 55 2233 89
rect 2177 47 2233 55
rect 2263 157 2319 175
rect 2263 123 2274 157
rect 2308 123 2319 157
rect 2263 89 2319 123
rect 2263 55 2274 89
rect 2308 55 2319 89
rect 2263 47 2319 55
rect 2349 157 2405 175
rect 2349 123 2360 157
rect 2394 123 2405 157
rect 2349 89 2405 123
rect 2349 55 2360 89
rect 2394 55 2405 89
rect 2349 47 2405 55
rect 2435 157 2491 175
rect 2435 123 2446 157
rect 2480 123 2491 157
rect 2435 89 2491 123
rect 2435 55 2446 89
rect 2480 55 2491 89
rect 2435 47 2491 55
rect 2521 157 2577 175
rect 2521 123 2532 157
rect 2566 123 2577 157
rect 2521 89 2577 123
rect 2521 55 2532 89
rect 2566 55 2577 89
rect 2521 47 2577 55
rect 2607 157 2663 175
rect 2607 123 2618 157
rect 2652 123 2663 157
rect 2607 89 2663 123
rect 2607 55 2618 89
rect 2652 55 2663 89
rect 2607 47 2663 55
rect 2693 157 2749 175
rect 2693 123 2704 157
rect 2738 123 2749 157
rect 2693 89 2749 123
rect 2693 55 2704 89
rect 2738 55 2749 89
rect 2693 47 2749 55
rect 2779 157 2835 175
rect 2779 123 2790 157
rect 2824 123 2835 157
rect 2779 89 2835 123
rect 2779 55 2790 89
rect 2824 55 2835 89
rect 2779 47 2835 55
rect 2865 157 2921 175
rect 2865 123 2876 157
rect 2910 123 2921 157
rect 2865 89 2921 123
rect 2865 55 2876 89
rect 2910 55 2921 89
rect 2865 47 2921 55
rect 2951 157 3007 175
rect 2951 123 2962 157
rect 2996 123 3007 157
rect 2951 89 3007 123
rect 2951 55 2962 89
rect 2996 55 3007 89
rect 2951 47 3007 55
rect 3037 157 3093 175
rect 3037 123 3048 157
rect 3082 123 3093 157
rect 3037 89 3093 123
rect 3037 55 3048 89
rect 3082 55 3093 89
rect 3037 47 3093 55
rect 3123 157 3179 175
rect 3123 123 3134 157
rect 3168 123 3179 157
rect 3123 89 3179 123
rect 3123 55 3134 89
rect 3168 55 3179 89
rect 3123 47 3179 55
rect 3209 157 3266 175
rect 3209 123 3220 157
rect 3254 123 3266 157
rect 3209 89 3266 123
rect 3209 55 3220 89
rect 3254 55 3266 89
rect 3209 47 3266 55
rect 1159 43 1168 47
rect 1116 31 1168 43
<< pdiff >>
rect 133 607 187 619
rect 133 573 142 607
rect 176 573 187 607
rect 133 535 187 573
rect 27 523 81 535
rect 27 489 36 523
rect 70 489 81 523
rect 27 413 81 489
rect 27 379 36 413
rect 70 379 81 413
rect 27 367 81 379
rect 111 522 187 535
rect 111 488 142 522
rect 176 488 187 522
rect 111 438 187 488
rect 111 404 142 438
rect 176 404 187 438
rect 111 367 187 404
rect 217 597 273 619
rect 217 563 228 597
rect 262 563 273 597
rect 217 517 273 563
rect 217 483 228 517
rect 262 483 273 517
rect 217 438 273 483
rect 217 404 228 438
rect 262 404 273 438
rect 217 367 273 404
rect 303 607 375 619
rect 303 573 314 607
rect 348 573 375 607
rect 303 508 375 573
rect 303 474 314 508
rect 348 474 375 508
rect 303 451 375 474
rect 405 597 461 619
rect 405 563 416 597
rect 450 563 461 597
rect 405 497 461 563
rect 405 463 416 497
rect 450 463 461 497
rect 405 451 461 463
rect 491 607 545 619
rect 491 573 502 607
rect 536 573 545 607
rect 491 537 545 573
rect 491 503 502 537
rect 536 503 545 537
rect 491 451 545 503
rect 658 597 720 619
rect 658 563 667 597
rect 701 563 720 597
rect 658 505 720 563
rect 658 471 667 505
rect 701 471 720 505
rect 303 367 353 451
rect 658 413 720 471
rect 658 379 667 413
rect 701 379 720 413
rect 658 367 720 379
rect 750 527 806 619
rect 750 493 761 527
rect 795 493 806 527
rect 750 413 806 493
rect 750 379 761 413
rect 795 379 806 413
rect 750 367 806 379
rect 836 597 908 619
rect 836 563 847 597
rect 881 563 908 597
rect 836 505 908 563
rect 836 471 847 505
rect 881 471 908 505
rect 836 413 908 471
rect 836 379 847 413
rect 881 379 908 413
rect 836 367 908 379
rect 938 596 994 619
rect 938 562 949 596
rect 983 562 994 596
rect 938 367 994 562
rect 1024 597 1113 619
rect 1024 563 1067 597
rect 1101 563 1113 597
rect 1024 509 1113 563
rect 1024 475 1067 509
rect 1101 475 1113 509
rect 1024 421 1113 475
rect 1024 387 1067 421
rect 1101 387 1113 421
rect 1024 367 1113 387
rect 1173 529 1230 541
rect 1173 495 1185 529
rect 1219 495 1230 529
rect 1173 419 1230 495
rect 1173 385 1185 419
rect 1219 385 1230 419
rect 1173 373 1230 385
rect 1260 373 1308 541
rect 1338 529 1395 541
rect 1338 495 1349 529
rect 1383 495 1395 529
rect 1338 419 1395 495
rect 1338 385 1349 419
rect 1383 385 1395 419
rect 1338 373 1395 385
rect 1457 607 1514 619
rect 1457 573 1469 607
rect 1503 573 1514 607
rect 1457 487 1514 573
rect 1457 453 1469 487
rect 1503 453 1514 487
rect 1457 367 1514 453
rect 1544 597 1600 619
rect 1544 563 1555 597
rect 1589 563 1600 597
rect 1544 505 1600 563
rect 1544 471 1555 505
rect 1589 471 1600 505
rect 1544 413 1600 471
rect 1544 379 1555 413
rect 1589 379 1600 413
rect 1544 367 1600 379
rect 1630 607 1803 619
rect 1630 437 1657 607
rect 1759 437 1803 607
rect 1630 367 1803 437
rect 1833 597 1889 619
rect 1833 563 1844 597
rect 1878 563 1889 597
rect 1833 519 1889 563
rect 1833 485 1844 519
rect 1878 485 1889 519
rect 1833 442 1889 485
rect 1833 408 1844 442
rect 1878 408 1889 442
rect 1833 367 1889 408
rect 1919 607 1975 619
rect 1919 573 1930 607
rect 1964 573 1975 607
rect 1919 512 1975 573
rect 1919 478 1930 512
rect 1964 478 1975 512
rect 1919 367 1975 478
rect 2005 597 2061 619
rect 2005 563 2016 597
rect 2050 563 2061 597
rect 2005 517 2061 563
rect 2005 483 2016 517
rect 2050 483 2061 517
rect 2005 438 2061 483
rect 2005 404 2016 438
rect 2050 404 2061 438
rect 2005 367 2061 404
rect 2091 607 2147 619
rect 2091 573 2102 607
rect 2136 573 2147 607
rect 2091 508 2147 573
rect 2091 474 2102 508
rect 2136 474 2147 508
rect 2091 367 2147 474
rect 2177 597 2233 619
rect 2177 563 2188 597
rect 2222 563 2233 597
rect 2177 517 2233 563
rect 2177 483 2188 517
rect 2222 483 2233 517
rect 2177 438 2233 483
rect 2177 404 2188 438
rect 2222 404 2233 438
rect 2177 367 2233 404
rect 2263 607 2319 619
rect 2263 573 2274 607
rect 2308 573 2319 607
rect 2263 508 2319 573
rect 2263 474 2274 508
rect 2308 474 2319 508
rect 2263 367 2319 474
rect 2349 597 2405 619
rect 2349 563 2360 597
rect 2394 563 2405 597
rect 2349 517 2405 563
rect 2349 483 2360 517
rect 2394 483 2405 517
rect 2349 438 2405 483
rect 2349 404 2360 438
rect 2394 404 2405 438
rect 2349 367 2405 404
rect 2435 607 2491 619
rect 2435 573 2446 607
rect 2480 573 2491 607
rect 2435 508 2491 573
rect 2435 474 2446 508
rect 2480 474 2491 508
rect 2435 367 2491 474
rect 2521 597 2577 619
rect 2521 563 2532 597
rect 2566 563 2577 597
rect 2521 517 2577 563
rect 2521 483 2532 517
rect 2566 483 2577 517
rect 2521 438 2577 483
rect 2521 404 2532 438
rect 2566 404 2577 438
rect 2521 367 2577 404
rect 2607 607 2663 619
rect 2607 573 2618 607
rect 2652 573 2663 607
rect 2607 508 2663 573
rect 2607 474 2618 508
rect 2652 474 2663 508
rect 2607 367 2663 474
rect 2693 597 2749 619
rect 2693 563 2704 597
rect 2738 563 2749 597
rect 2693 517 2749 563
rect 2693 483 2704 517
rect 2738 483 2749 517
rect 2693 438 2749 483
rect 2693 404 2704 438
rect 2738 404 2749 438
rect 2693 367 2749 404
rect 2779 607 2835 619
rect 2779 573 2790 607
rect 2824 573 2835 607
rect 2779 508 2835 573
rect 2779 474 2790 508
rect 2824 474 2835 508
rect 2779 367 2835 474
rect 2865 597 2921 619
rect 2865 563 2876 597
rect 2910 563 2921 597
rect 2865 517 2921 563
rect 2865 483 2876 517
rect 2910 483 2921 517
rect 2865 438 2921 483
rect 2865 404 2876 438
rect 2910 404 2921 438
rect 2865 367 2921 404
rect 2951 607 3007 619
rect 2951 573 2962 607
rect 2996 573 3007 607
rect 2951 508 3007 573
rect 2951 474 2962 508
rect 2996 474 3007 508
rect 2951 367 3007 474
rect 3037 597 3093 619
rect 3037 563 3048 597
rect 3082 563 3093 597
rect 3037 517 3093 563
rect 3037 483 3048 517
rect 3082 483 3093 517
rect 3037 438 3093 483
rect 3037 404 3048 438
rect 3082 404 3093 438
rect 3037 367 3093 404
rect 3123 607 3179 619
rect 3123 573 3134 607
rect 3168 573 3179 607
rect 3123 508 3179 573
rect 3123 474 3134 508
rect 3168 474 3179 508
rect 3123 367 3179 474
rect 3209 597 3265 619
rect 3209 563 3220 597
rect 3254 563 3265 597
rect 3209 517 3265 563
rect 3209 483 3220 517
rect 3254 483 3265 517
rect 3209 438 3265 483
rect 3209 404 3220 438
rect 3254 404 3265 438
rect 3209 367 3265 404
rect 3295 607 3351 619
rect 3295 573 3306 607
rect 3340 573 3351 607
rect 3295 508 3351 573
rect 3295 474 3306 508
rect 3340 474 3351 508
rect 3295 367 3351 474
rect 3381 597 3437 619
rect 3381 563 3392 597
rect 3426 563 3437 597
rect 3381 517 3437 563
rect 3381 483 3392 517
rect 3426 483 3437 517
rect 3381 438 3437 483
rect 3381 404 3392 438
rect 3426 404 3437 438
rect 3381 367 3437 404
rect 3467 607 3524 619
rect 3467 573 3478 607
rect 3512 573 3524 607
rect 3467 508 3524 573
rect 3467 474 3478 508
rect 3512 474 3524 508
rect 3467 367 3524 474
<< ndiffc >>
rect 126 105 160 139
rect 228 105 262 139
rect 415 139 449 173
rect 597 71 631 105
rect 737 154 771 188
rect 893 59 927 93
rect 999 199 1033 233
rect 1125 43 1159 77
rect 1249 77 1283 111
rect 1351 59 1385 93
rect 1463 59 1497 93
rect 1549 79 1583 113
rect 1651 169 1685 203
rect 1651 69 1685 103
rect 1753 146 1787 180
rect 1844 169 1878 203
rect 1844 69 1878 103
rect 2016 123 2050 157
rect 2016 55 2050 89
rect 2102 123 2136 157
rect 2102 55 2136 89
rect 2188 123 2222 157
rect 2188 55 2222 89
rect 2274 123 2308 157
rect 2274 55 2308 89
rect 2360 123 2394 157
rect 2360 55 2394 89
rect 2446 123 2480 157
rect 2446 55 2480 89
rect 2532 123 2566 157
rect 2532 55 2566 89
rect 2618 123 2652 157
rect 2618 55 2652 89
rect 2704 123 2738 157
rect 2704 55 2738 89
rect 2790 123 2824 157
rect 2790 55 2824 89
rect 2876 123 2910 157
rect 2876 55 2910 89
rect 2962 123 2996 157
rect 2962 55 2996 89
rect 3048 123 3082 157
rect 3048 55 3082 89
rect 3134 123 3168 157
rect 3134 55 3168 89
rect 3220 123 3254 157
rect 3220 55 3254 89
<< pdiffc >>
rect 142 573 176 607
rect 36 489 70 523
rect 36 379 70 413
rect 142 488 176 522
rect 142 404 176 438
rect 228 563 262 597
rect 228 483 262 517
rect 228 404 262 438
rect 314 573 348 607
rect 314 474 348 508
rect 416 563 450 597
rect 416 463 450 497
rect 502 573 536 607
rect 502 503 536 537
rect 667 563 701 597
rect 667 471 701 505
rect 667 379 701 413
rect 761 493 795 527
rect 761 379 795 413
rect 847 563 881 597
rect 847 471 881 505
rect 847 379 881 413
rect 949 562 983 596
rect 1067 563 1101 597
rect 1067 475 1101 509
rect 1067 387 1101 421
rect 1185 495 1219 529
rect 1185 385 1219 419
rect 1349 495 1383 529
rect 1349 385 1383 419
rect 1469 573 1503 607
rect 1469 453 1503 487
rect 1555 563 1589 597
rect 1555 471 1589 505
rect 1555 379 1589 413
rect 1657 437 1759 607
rect 1844 563 1878 597
rect 1844 485 1878 519
rect 1844 408 1878 442
rect 1930 573 1964 607
rect 1930 478 1964 512
rect 2016 563 2050 597
rect 2016 483 2050 517
rect 2016 404 2050 438
rect 2102 573 2136 607
rect 2102 474 2136 508
rect 2188 563 2222 597
rect 2188 483 2222 517
rect 2188 404 2222 438
rect 2274 573 2308 607
rect 2274 474 2308 508
rect 2360 563 2394 597
rect 2360 483 2394 517
rect 2360 404 2394 438
rect 2446 573 2480 607
rect 2446 474 2480 508
rect 2532 563 2566 597
rect 2532 483 2566 517
rect 2532 404 2566 438
rect 2618 573 2652 607
rect 2618 474 2652 508
rect 2704 563 2738 597
rect 2704 483 2738 517
rect 2704 404 2738 438
rect 2790 573 2824 607
rect 2790 474 2824 508
rect 2876 563 2910 597
rect 2876 483 2910 517
rect 2876 404 2910 438
rect 2962 573 2996 607
rect 2962 474 2996 508
rect 3048 563 3082 597
rect 3048 483 3082 517
rect 3048 404 3082 438
rect 3134 573 3168 607
rect 3134 474 3168 508
rect 3220 563 3254 597
rect 3220 483 3254 517
rect 3220 404 3254 438
rect 3306 573 3340 607
rect 3306 474 3340 508
rect 3392 563 3426 597
rect 3392 483 3426 517
rect 3392 404 3426 438
rect 3478 573 3512 607
rect 3478 474 3512 508
<< poly >>
rect 187 619 217 645
rect 273 619 303 645
rect 375 619 405 645
rect 461 619 491 645
rect 720 619 750 645
rect 806 619 836 645
rect 908 619 938 645
rect 994 619 1024 645
rect 81 535 111 561
rect 81 265 111 367
rect 187 343 217 367
rect 273 343 303 367
rect 375 343 405 451
rect 461 381 491 451
rect 187 319 405 343
rect 187 313 233 319
rect 217 285 233 313
rect 267 313 405 319
rect 447 365 513 381
rect 447 331 463 365
rect 497 331 513 365
rect 447 315 513 331
rect 560 365 626 381
rect 1128 615 1440 645
rect 1514 619 1544 645
rect 1600 619 1630 645
rect 1803 619 1833 645
rect 1889 619 1919 645
rect 1975 619 2005 645
rect 2061 619 2091 645
rect 2147 619 2177 645
rect 2233 619 2263 645
rect 2319 619 2349 645
rect 2405 619 2435 645
rect 2491 619 2521 645
rect 2577 619 2607 645
rect 2663 619 2693 645
rect 2749 619 2779 645
rect 2835 619 2865 645
rect 2921 619 2951 645
rect 3007 619 3037 645
rect 3093 619 3123 645
rect 3179 619 3209 645
rect 3265 619 3295 645
rect 3351 619 3381 645
rect 3437 619 3467 645
rect 560 331 576 365
rect 610 345 626 365
rect 720 345 750 367
rect 806 345 836 367
rect 610 331 836 345
rect 560 315 836 331
rect 267 285 303 313
rect 217 269 303 285
rect 81 249 167 265
rect 81 215 117 249
rect 151 221 167 249
rect 151 215 201 221
rect 81 191 201 215
rect 171 169 201 191
rect 273 169 303 269
rect 453 265 483 315
rect 908 299 938 367
rect 994 343 1024 367
rect 1128 343 1158 615
rect 1230 541 1260 567
rect 1308 541 1338 567
rect 994 319 1158 343
rect 994 299 1010 319
rect 908 285 1010 299
rect 1044 313 1158 319
rect 1044 285 1094 313
rect 908 269 1094 285
rect 351 235 483 265
rect 531 237 812 267
rect 351 169 381 235
rect 531 187 561 237
rect 696 215 726 237
rect 782 215 812 237
rect 938 215 968 269
rect 495 171 561 187
rect 495 137 511 171
rect 545 137 561 171
rect 495 103 561 137
rect 171 59 201 85
rect 273 59 303 85
rect 351 59 381 85
rect 495 69 511 103
rect 545 69 561 103
rect 495 53 561 69
rect 1064 215 1094 269
rect 1230 265 1260 373
rect 1308 333 1338 373
rect 1410 345 1440 615
rect 1514 345 1544 367
rect 1600 345 1630 367
rect 1190 249 1260 265
rect 1190 215 1206 249
rect 1240 215 1260 249
rect 1190 199 1260 215
rect 1302 317 1368 333
rect 1302 283 1318 317
rect 1352 283 1368 317
rect 1410 315 1630 345
rect 1803 345 1833 367
rect 1889 345 1919 367
rect 1975 345 2005 367
rect 2061 345 2091 367
rect 2147 345 2177 367
rect 2233 345 2263 367
rect 2319 345 2349 367
rect 2405 345 2435 367
rect 2491 345 2521 367
rect 2577 345 2607 367
rect 2663 345 2693 367
rect 2749 345 2779 367
rect 2835 345 2865 367
rect 2921 345 2951 367
rect 3007 345 3037 367
rect 3093 345 3123 367
rect 3179 345 3209 367
rect 3265 345 3295 367
rect 3351 345 3381 367
rect 3437 345 3467 367
rect 1302 249 1368 283
rect 1302 215 1318 249
rect 1352 215 1368 249
rect 1508 215 1538 315
rect 1594 215 1624 315
rect 1672 305 1738 321
rect 1803 319 3467 345
rect 1803 315 2788 319
rect 1672 271 1688 305
rect 1722 271 1738 305
rect 2772 285 2788 315
rect 2822 285 2960 319
rect 2994 285 3132 319
rect 3166 285 3304 319
rect 3338 285 3372 319
rect 3406 285 3467 319
rect 1672 267 1738 271
rect 1672 237 1828 267
rect 1696 215 1726 237
rect 1798 215 1828 237
rect 1905 257 2670 273
rect 2772 269 3467 285
rect 1905 223 1932 257
rect 1966 223 2104 257
rect 2138 223 2272 257
rect 2306 223 2448 257
rect 2482 223 2620 257
rect 2654 227 2670 257
rect 2654 223 3209 227
rect 1302 199 1368 215
rect 1208 131 1238 199
rect 1308 131 1338 199
rect 696 21 726 47
rect 782 21 812 47
rect 938 21 968 47
rect 1064 21 1094 47
rect 1905 207 3209 223
rect 2061 175 2091 207
rect 2147 175 2177 207
rect 2233 175 2263 207
rect 2319 175 2349 207
rect 2405 197 3209 207
rect 2405 175 2435 197
rect 2491 175 2521 197
rect 2577 175 2607 197
rect 2663 175 2693 197
rect 2749 175 2779 197
rect 2835 175 2865 197
rect 2921 175 2951 197
rect 3007 175 3037 197
rect 3093 175 3123 197
rect 3179 175 3209 197
rect 1208 21 1238 47
rect 1308 21 1338 47
rect 1508 21 1538 47
rect 1594 21 1624 47
rect 1696 21 1726 47
rect 1798 21 1828 47
rect 2061 21 2091 47
rect 2147 21 2177 47
rect 2233 21 2263 47
rect 2319 21 2349 47
rect 2405 21 2435 47
rect 2491 21 2521 47
rect 2577 21 2607 47
rect 2663 21 2693 47
rect 2749 21 2779 47
rect 2835 21 2865 47
rect 2921 21 2951 47
rect 3007 21 3037 47
rect 3093 21 3123 47
rect 3179 21 3209 47
<< polycont >>
rect 233 285 267 319
rect 463 331 497 365
rect 576 331 610 365
rect 117 215 151 249
rect 1010 285 1044 319
rect 511 137 545 171
rect 511 69 545 103
rect 1206 215 1240 249
rect 1318 283 1352 317
rect 1318 215 1352 249
rect 1688 271 1722 305
rect 2788 285 2822 319
rect 2960 285 2994 319
rect 3132 285 3166 319
rect 3304 285 3338 319
rect 3372 285 3406 319
rect 1932 223 1966 257
rect 2104 223 2138 257
rect 2272 223 2306 257
rect 2448 223 2482 257
rect 2620 223 2654 257
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3552 683
rect 126 607 176 649
rect 126 573 142 607
rect 20 523 86 539
rect 20 489 36 523
rect 70 489 86 523
rect 20 413 86 489
rect 20 379 36 413
rect 70 379 86 413
rect 126 522 176 573
rect 126 488 142 522
rect 126 438 176 488
rect 126 404 142 438
rect 126 388 176 404
rect 212 597 278 613
rect 212 563 228 597
rect 262 563 278 597
rect 212 517 278 563
rect 212 483 228 517
rect 262 483 278 517
rect 212 438 278 483
rect 314 607 364 649
rect 348 573 364 607
rect 314 508 364 573
rect 348 474 364 508
rect 314 458 364 474
rect 400 597 466 613
rect 400 563 416 597
rect 450 563 466 597
rect 400 497 466 563
rect 400 463 416 497
rect 450 463 466 497
rect 502 607 552 649
rect 536 573 552 607
rect 502 537 552 573
rect 536 503 552 537
rect 502 487 552 503
rect 667 597 897 613
rect 701 579 847 597
rect 667 505 701 563
rect 831 563 847 579
rect 881 563 897 597
rect 212 404 228 438
rect 262 422 278 438
rect 400 451 466 463
rect 262 404 353 422
rect 400 417 626 451
rect 212 388 353 404
rect 20 352 86 379
rect 20 319 283 352
rect 20 318 233 319
rect 20 163 54 318
rect 217 285 233 318
rect 267 285 283 319
rect 319 344 353 388
rect 409 365 513 381
rect 409 350 463 365
rect 409 344 415 350
rect 319 316 415 344
rect 449 331 463 350
rect 497 331 513 365
rect 449 316 513 331
rect 319 310 513 316
rect 560 365 626 417
rect 560 331 576 365
rect 610 331 626 365
rect 667 413 701 471
rect 667 363 701 379
rect 737 527 795 543
rect 737 493 761 527
rect 737 413 795 493
rect 737 379 761 413
rect 737 363 795 379
rect 831 505 897 563
rect 933 596 999 649
rect 933 562 949 596
rect 983 562 999 596
rect 933 536 999 562
rect 1067 597 1117 613
rect 1101 563 1117 597
rect 831 471 847 505
rect 881 500 897 505
rect 1067 509 1117 563
rect 881 475 1067 500
rect 1101 475 1117 509
rect 881 471 1117 475
rect 831 466 1117 471
rect 831 413 897 466
rect 831 379 847 413
rect 881 379 897 413
rect 831 363 897 379
rect 560 315 626 331
rect 101 249 167 282
rect 217 269 283 285
rect 560 274 594 315
rect 101 215 117 249
rect 151 233 167 249
rect 399 240 594 274
rect 151 215 348 233
rect 101 199 348 215
rect 20 139 176 163
rect 20 129 126 139
rect 110 105 126 129
rect 160 105 176 139
rect 110 81 176 105
rect 212 139 278 163
rect 212 105 228 139
rect 262 105 278 139
rect 212 17 278 105
rect 314 87 348 199
rect 399 173 449 240
rect 737 233 771 363
rect 985 335 1031 430
rect 1067 421 1117 466
rect 1101 387 1117 421
rect 1067 371 1117 387
rect 1169 529 1235 649
rect 1453 607 1503 649
rect 1453 573 1469 607
rect 1169 495 1185 529
rect 1219 495 1235 529
rect 1169 419 1235 495
rect 1169 385 1185 419
rect 1219 385 1235 419
rect 1169 369 1235 385
rect 1333 529 1399 545
rect 1333 495 1349 529
rect 1383 495 1399 529
rect 1333 419 1399 495
rect 1453 487 1503 573
rect 1453 453 1469 487
rect 1453 437 1503 453
rect 1539 597 1605 613
rect 1539 563 1555 597
rect 1589 563 1605 597
rect 1539 505 1605 563
rect 1539 471 1555 505
rect 1589 471 1605 505
rect 1333 385 1349 419
rect 1383 403 1399 419
rect 1539 413 1605 471
rect 1641 607 1775 649
rect 1641 437 1657 607
rect 1759 437 1775 607
rect 1641 427 1775 437
rect 1844 597 1878 613
rect 1844 519 1878 563
rect 1844 442 1878 485
rect 1914 607 1964 649
rect 1914 573 1930 607
rect 1914 512 1964 573
rect 1914 478 1930 512
rect 1914 462 1964 478
rect 2000 597 2066 613
rect 2000 563 2016 597
rect 2050 563 2066 597
rect 2000 517 2066 563
rect 2000 483 2016 517
rect 2050 483 2066 517
rect 1383 385 1438 403
rect 1333 369 1438 385
rect 985 319 1051 335
rect 985 285 1010 319
rect 1044 285 1051 319
rect 985 269 1051 285
rect 1279 317 1368 333
rect 1279 283 1318 317
rect 1352 283 1368 317
rect 1087 276 1127 282
rect 1121 242 1127 276
rect 1279 276 1368 283
rect 1087 233 1127 242
rect 399 139 415 173
rect 399 123 449 139
rect 495 171 701 204
rect 495 137 511 171
rect 545 170 701 171
rect 545 137 561 170
rect 495 103 561 137
rect 495 87 511 103
rect 314 69 511 87
rect 545 69 561 103
rect 314 53 561 69
rect 597 105 631 134
rect 597 17 631 71
rect 667 87 701 170
rect 737 199 999 233
rect 1033 199 1127 233
rect 1163 249 1243 265
rect 1163 215 1206 249
rect 1240 215 1243 249
rect 1163 199 1243 215
rect 1313 249 1368 276
rect 1313 242 1318 249
rect 1279 215 1318 242
rect 1352 215 1368 249
rect 1279 199 1368 215
rect 1404 321 1438 369
rect 1539 379 1555 413
rect 1589 391 1605 413
rect 2000 438 2066 483
rect 2102 607 2136 649
rect 2102 508 2136 573
rect 2102 458 2136 474
rect 2172 597 2238 613
rect 2172 563 2188 597
rect 2222 563 2238 597
rect 2172 517 2238 563
rect 2172 483 2188 517
rect 2222 483 2238 517
rect 2000 426 2016 438
rect 1589 379 1808 391
rect 1878 390 2016 426
rect 2050 390 2066 438
rect 1539 357 1808 379
rect 1774 356 1808 357
rect 1774 350 1895 356
rect 1404 305 1738 321
rect 1404 271 1688 305
rect 1722 271 1738 305
rect 1404 255 1738 271
rect 1774 316 1855 350
rect 1889 316 1895 350
rect 1774 310 1895 316
rect 737 188 771 199
rect 1163 163 1197 199
rect 1404 163 1438 255
rect 1774 219 1808 310
rect 1928 276 1966 282
rect 1928 223 1932 276
rect 737 123 771 154
rect 807 129 1197 163
rect 1233 129 1438 163
rect 1472 203 1701 219
rect 1472 185 1651 203
rect 807 87 841 129
rect 1233 111 1299 129
rect 667 53 841 87
rect 877 59 893 93
rect 927 59 943 93
rect 877 17 943 59
rect 1109 77 1175 93
rect 1109 43 1125 77
rect 1159 43 1175 77
rect 1233 77 1249 111
rect 1283 77 1299 111
rect 1472 93 1513 185
rect 1635 169 1651 185
rect 1685 169 1701 203
rect 1233 53 1299 77
rect 1335 59 1351 93
rect 1385 59 1401 93
rect 1447 59 1463 93
rect 1497 59 1513 93
rect 1549 113 1599 149
rect 1583 79 1599 113
rect 1109 17 1175 43
rect 1335 17 1401 59
rect 1549 17 1599 79
rect 1635 103 1701 169
rect 1737 180 1808 219
rect 1737 146 1753 180
rect 1787 146 1808 180
rect 1737 123 1808 146
rect 1844 203 1894 219
rect 1928 207 1966 223
rect 1878 169 1894 203
rect 1635 69 1651 103
rect 1685 87 1701 103
rect 1844 103 1894 169
rect 1685 69 1844 87
rect 1878 69 1894 103
rect 1635 53 1894 69
rect 2000 157 2066 390
rect 2172 438 2238 483
rect 2274 607 2308 649
rect 2274 508 2308 573
rect 2274 458 2308 474
rect 2344 597 2410 613
rect 2344 563 2360 597
rect 2394 563 2410 597
rect 2344 517 2410 563
rect 2344 483 2360 517
rect 2394 483 2410 517
rect 2172 390 2188 438
rect 2222 390 2238 438
rect 2100 276 2138 282
rect 2100 223 2104 276
rect 2100 207 2138 223
rect 2000 123 2016 157
rect 2050 123 2066 157
rect 2000 89 2066 123
rect 2000 55 2016 89
rect 2050 55 2066 89
rect 2000 51 2066 55
rect 2102 157 2136 173
rect 2102 89 2136 123
rect 2102 17 2136 55
rect 2172 157 2238 390
rect 2344 438 2410 483
rect 2446 607 2480 649
rect 2446 508 2480 573
rect 2446 458 2480 474
rect 2516 597 2582 613
rect 2516 563 2532 597
rect 2566 563 2582 597
rect 2516 517 2582 563
rect 2516 483 2532 517
rect 2566 483 2582 517
rect 2344 390 2360 438
rect 2394 390 2410 438
rect 2272 276 2310 282
rect 2272 257 2276 276
rect 2306 223 2310 242
rect 2272 207 2310 223
rect 2172 123 2188 157
rect 2222 123 2238 157
rect 2172 89 2238 123
rect 2172 55 2188 89
rect 2222 55 2238 89
rect 2172 51 2238 55
rect 2274 157 2308 173
rect 2274 89 2308 123
rect 2274 17 2308 55
rect 2344 157 2410 390
rect 2516 438 2582 483
rect 2618 607 2652 649
rect 2618 508 2652 573
rect 2618 458 2652 474
rect 2688 597 2754 613
rect 2688 563 2704 597
rect 2738 563 2754 597
rect 2688 517 2754 563
rect 2688 483 2704 517
rect 2738 483 2754 517
rect 2516 390 2532 438
rect 2566 390 2582 438
rect 2444 276 2482 282
rect 2444 223 2448 276
rect 2444 207 2482 223
rect 2344 123 2360 157
rect 2394 123 2410 157
rect 2344 89 2410 123
rect 2344 55 2360 89
rect 2394 55 2410 89
rect 2344 51 2410 55
rect 2446 157 2480 173
rect 2446 89 2480 123
rect 2446 17 2480 55
rect 2516 157 2582 390
rect 2688 438 2754 483
rect 2790 607 2824 649
rect 2790 508 2824 573
rect 2790 458 2824 474
rect 2860 597 2926 613
rect 2860 563 2876 597
rect 2910 563 2926 597
rect 2860 517 2926 563
rect 2860 483 2876 517
rect 2910 483 2926 517
rect 2688 390 2704 438
rect 2738 390 2754 438
rect 2616 276 2654 282
rect 2616 223 2620 276
rect 2616 207 2654 223
rect 2516 123 2532 157
rect 2566 123 2582 157
rect 2516 89 2582 123
rect 2516 55 2532 89
rect 2566 55 2582 89
rect 2516 51 2582 55
rect 2618 157 2652 173
rect 2618 89 2652 123
rect 2618 17 2652 55
rect 2688 157 2754 390
rect 2860 438 2926 483
rect 2962 607 2996 649
rect 2962 508 2996 573
rect 2962 458 2996 474
rect 3032 597 3098 613
rect 3032 563 3048 597
rect 3082 563 3098 597
rect 3032 517 3098 563
rect 3032 483 3048 517
rect 3082 483 3098 517
rect 2860 390 2876 438
rect 2910 390 2926 438
rect 2788 350 2826 352
rect 2822 285 2826 350
rect 2788 269 2826 285
rect 2688 123 2704 157
rect 2738 123 2754 157
rect 2688 89 2754 123
rect 2688 55 2704 89
rect 2738 55 2754 89
rect 2688 51 2754 55
rect 2790 157 2824 173
rect 2790 89 2824 123
rect 2790 17 2824 55
rect 2860 157 2926 390
rect 3032 438 3098 483
rect 3134 607 3168 649
rect 3134 508 3168 573
rect 3134 458 3168 474
rect 3204 597 3270 613
rect 3204 563 3220 597
rect 3254 563 3270 597
rect 3204 517 3270 563
rect 3204 483 3220 517
rect 3254 483 3270 517
rect 3032 390 3048 438
rect 3082 390 3098 438
rect 2960 350 2998 352
rect 2994 285 2998 350
rect 2960 269 2998 285
rect 2860 123 2876 157
rect 2910 123 2926 157
rect 2860 89 2926 123
rect 2860 55 2876 89
rect 2910 55 2926 89
rect 2860 51 2926 55
rect 2962 157 2996 173
rect 2962 89 2996 123
rect 2962 17 2996 55
rect 3032 157 3098 390
rect 3204 438 3270 483
rect 3306 607 3340 649
rect 3306 508 3340 573
rect 3306 458 3340 474
rect 3376 597 3442 613
rect 3376 563 3392 597
rect 3426 563 3442 597
rect 3376 517 3442 563
rect 3376 483 3392 517
rect 3426 483 3442 517
rect 3204 390 3220 438
rect 3254 390 3270 438
rect 3132 350 3170 352
rect 3166 285 3170 350
rect 3132 269 3170 285
rect 3032 123 3048 157
rect 3082 123 3098 157
rect 3032 89 3098 123
rect 3032 55 3048 89
rect 3082 55 3098 89
rect 3032 52 3098 55
rect 3134 157 3168 173
rect 3134 89 3168 123
rect 3134 17 3168 55
rect 3204 157 3270 390
rect 3376 438 3442 483
rect 3478 607 3528 649
rect 3512 573 3528 607
rect 3478 508 3528 573
rect 3512 474 3528 508
rect 3478 458 3528 474
rect 3376 390 3392 438
rect 3426 390 3442 438
rect 3376 388 3442 390
rect 3304 350 3422 352
rect 3338 319 3376 350
rect 3338 285 3372 319
rect 3410 316 3422 350
rect 3406 285 3422 316
rect 3304 269 3422 285
rect 3204 123 3220 157
rect 3254 123 3270 157
rect 3204 89 3270 123
rect 3204 55 3220 89
rect 3254 55 3270 89
rect 3204 51 3270 55
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 415 316 449 350
rect 1087 242 1121 276
rect 1279 242 1313 276
rect 1844 408 1878 424
rect 1844 390 1878 408
rect 2016 404 2050 424
rect 2016 390 2050 404
rect 1855 316 1889 350
rect 1932 257 1966 276
rect 1932 242 1966 257
rect 2188 404 2222 424
rect 2188 390 2222 404
rect 2104 257 2138 276
rect 2104 242 2138 257
rect 2360 404 2394 424
rect 2360 390 2394 404
rect 2276 257 2310 276
rect 2276 242 2306 257
rect 2306 242 2310 257
rect 2532 404 2566 424
rect 2532 390 2566 404
rect 2448 257 2482 276
rect 2448 242 2482 257
rect 2704 404 2738 424
rect 2704 390 2738 404
rect 2620 257 2654 276
rect 2620 242 2654 257
rect 2876 404 2910 424
rect 2876 390 2910 404
rect 2788 319 2822 350
rect 2788 316 2822 319
rect 3048 404 3082 424
rect 3048 390 3082 404
rect 2960 319 2994 350
rect 2960 316 2994 319
rect 3220 404 3254 424
rect 3220 390 3254 404
rect 3132 319 3166 350
rect 3132 316 3166 319
rect 3392 404 3426 424
rect 3392 390 3426 404
rect 3304 319 3338 350
rect 3376 319 3410 350
rect 3304 316 3338 319
rect 3376 316 3406 319
rect 3406 316 3410 319
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
<< metal1 >>
rect 0 683 3552 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3552 683
rect 0 617 3552 649
rect 1832 424 3438 430
rect 1832 390 1844 424
rect 1878 390 2016 424
rect 2050 390 2188 424
rect 2222 390 2360 424
rect 2394 390 2532 424
rect 2566 390 2704 424
rect 2738 390 2876 424
rect 2910 390 3048 424
rect 3082 390 3220 424
rect 3254 390 3392 424
rect 3426 390 3438 424
rect 1832 384 3438 390
rect 403 350 461 356
rect 403 316 415 350
rect 449 347 461 350
rect 1843 350 3422 356
rect 1843 347 1855 350
rect 449 319 1855 347
rect 449 316 461 319
rect 403 310 461 316
rect 1843 316 1855 319
rect 1889 316 2788 350
rect 2822 316 2960 350
rect 2994 316 3132 350
rect 3166 316 3304 350
rect 3338 316 3376 350
rect 3410 316 3422 350
rect 1843 310 3422 316
rect 1075 276 1133 282
rect 1075 242 1087 276
rect 1121 273 1133 276
rect 1267 276 1325 282
rect 1267 273 1279 276
rect 1121 245 1279 273
rect 1121 242 1133 245
rect 1075 236 1133 242
rect 1267 242 1279 245
rect 1313 273 1325 276
rect 1920 276 2666 282
rect 1920 273 1932 276
rect 1313 245 1932 273
rect 1313 242 1325 245
rect 1267 236 1325 242
rect 1920 242 1932 245
rect 1966 242 2104 276
rect 2138 242 2276 276
rect 2310 242 2448 276
rect 2482 242 2620 276
rect 2654 242 2666 276
rect 1920 236 2666 242
rect 0 17 3552 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
rect 0 -49 3552 -17
<< labels >>
flabel pwell s 0 0 3552 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 3552 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 busdrivernovlp_20
flabel metal1 s 1832 384 3438 430 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel metal1 s 0 617 3552 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 3552 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3552 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y
string GDS_END 721358
string GDS_START 694268
<< end >>
