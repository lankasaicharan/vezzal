magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 1 49 671 157
rect 0 0 672 49
<< scnmos >>
rect 80 47 110 131
rect 310 47 340 131
rect 398 47 428 131
rect 490 47 520 131
rect 562 47 592 131
<< scpmoshvt >>
rect 208 485 238 613
rect 310 485 340 613
rect 382 485 412 613
rect 476 485 506 613
rect 562 485 592 613
<< ndiff >>
rect 27 106 80 131
rect 27 72 35 106
rect 69 72 80 106
rect 27 47 80 72
rect 110 106 163 131
rect 110 72 121 106
rect 155 72 163 106
rect 110 47 163 72
rect 257 106 310 131
rect 257 72 265 106
rect 299 72 310 106
rect 257 47 310 72
rect 340 106 398 131
rect 340 72 353 106
rect 387 72 398 106
rect 340 47 398 72
rect 428 106 490 131
rect 428 72 445 106
rect 479 72 490 106
rect 428 47 490 72
rect 520 47 562 131
rect 592 106 645 131
rect 592 72 603 106
rect 637 72 645 106
rect 592 47 645 72
<< pdiff >>
rect 87 601 208 613
rect 87 567 95 601
rect 129 567 163 601
rect 197 567 208 601
rect 87 531 208 567
rect 87 497 95 531
rect 129 497 163 531
rect 197 497 208 531
rect 87 485 208 497
rect 238 601 310 613
rect 238 567 265 601
rect 299 567 310 601
rect 238 531 310 567
rect 238 497 265 531
rect 299 497 310 531
rect 238 485 310 497
rect 340 485 382 613
rect 412 599 476 613
rect 412 565 423 599
rect 457 565 476 599
rect 412 527 476 565
rect 412 493 423 527
rect 457 493 476 527
rect 412 485 476 493
rect 506 601 562 613
rect 506 567 517 601
rect 551 567 562 601
rect 506 531 562 567
rect 506 497 517 531
rect 551 497 562 531
rect 506 485 562 497
rect 592 601 645 613
rect 592 567 603 601
rect 637 567 645 601
rect 592 531 645 567
rect 592 497 603 531
rect 637 497 645 531
rect 592 485 645 497
<< ndiffc >>
rect 35 72 69 106
rect 121 72 155 106
rect 265 72 299 106
rect 353 72 387 106
rect 445 72 479 106
rect 603 72 637 106
<< pdiffc >>
rect 95 567 129 601
rect 163 567 197 601
rect 95 497 129 531
rect 163 497 197 531
rect 265 567 299 601
rect 265 497 299 531
rect 423 565 457 599
rect 423 493 457 527
rect 517 567 551 601
rect 517 497 551 531
rect 603 567 637 601
rect 603 497 637 531
<< poly >>
rect 208 613 238 639
rect 310 613 340 639
rect 382 613 412 639
rect 476 613 506 639
rect 562 613 592 639
rect 208 453 238 485
rect 80 437 243 453
rect 80 403 125 437
rect 159 403 193 437
rect 227 403 243 437
rect 80 387 243 403
rect 80 131 110 387
rect 310 313 340 485
rect 206 297 340 313
rect 206 263 222 297
rect 256 263 290 297
rect 324 263 340 297
rect 206 247 340 263
rect 310 131 340 247
rect 382 367 412 485
rect 476 445 506 485
rect 476 415 520 445
rect 490 372 520 415
rect 562 444 592 485
rect 562 414 649 444
rect 382 351 448 367
rect 382 317 398 351
rect 432 317 448 351
rect 382 283 448 317
rect 382 249 398 283
rect 432 249 448 283
rect 382 233 448 249
rect 490 356 577 372
rect 490 322 506 356
rect 540 322 577 356
rect 490 300 577 322
rect 398 131 428 233
rect 490 131 520 300
rect 619 219 649 414
rect 562 203 649 219
rect 562 169 599 203
rect 633 169 649 203
rect 562 153 649 169
rect 562 131 592 153
rect 80 21 110 47
rect 310 21 340 47
rect 398 21 428 47
rect 490 21 520 47
rect 562 21 592 47
<< polycont >>
rect 125 403 159 437
rect 193 403 227 437
rect 222 263 256 297
rect 290 263 324 297
rect 398 317 432 351
rect 398 249 432 283
rect 506 322 540 356
rect 599 169 633 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 17 601 213 615
rect 17 567 95 601
rect 129 567 163 601
rect 197 567 213 601
rect 17 531 213 567
rect 17 497 95 531
rect 129 497 163 531
rect 197 497 213 531
rect 17 481 213 497
rect 249 601 315 649
rect 249 567 265 601
rect 299 567 315 601
rect 249 531 315 567
rect 249 497 265 531
rect 299 497 315 531
rect 249 481 315 497
rect 413 599 467 615
rect 413 565 423 599
rect 457 565 467 599
rect 413 527 467 565
rect 413 493 423 527
rect 457 493 467 527
rect 17 106 73 481
rect 413 447 467 493
rect 501 601 553 649
rect 501 567 517 601
rect 551 567 553 601
rect 501 531 553 567
rect 501 497 517 531
rect 551 497 553 531
rect 501 481 553 497
rect 587 601 653 615
rect 587 567 603 601
rect 637 567 653 601
rect 587 531 653 567
rect 587 497 603 531
rect 637 497 653 531
rect 587 447 653 497
rect 109 437 653 447
rect 109 403 125 437
rect 159 403 193 437
rect 227 410 653 437
rect 227 403 358 410
rect 109 387 358 403
rect 392 351 456 367
rect 392 317 398 351
rect 432 317 456 351
rect 206 297 340 313
rect 206 263 222 297
rect 256 263 290 297
rect 324 263 340 297
rect 206 224 340 263
rect 392 283 456 317
rect 490 356 553 372
rect 490 322 506 356
rect 540 322 553 356
rect 490 306 553 322
rect 392 249 398 283
rect 432 249 456 283
rect 587 272 653 410
rect 392 233 456 249
rect 515 238 653 272
rect 251 156 481 190
rect 17 72 35 106
rect 69 72 73 106
rect 17 53 73 72
rect 109 106 175 123
rect 109 72 121 106
rect 155 72 175 106
rect 109 17 175 72
rect 251 106 315 156
rect 251 72 265 106
rect 299 72 315 106
rect 251 56 315 72
rect 349 106 401 122
rect 349 72 353 106
rect 387 72 401 106
rect 349 17 401 72
rect 435 106 481 156
rect 435 72 445 106
rect 479 72 481 106
rect 435 56 481 72
rect 515 121 549 238
rect 583 203 649 204
rect 583 169 599 203
rect 633 169 649 203
rect 583 155 649 169
rect 515 106 653 121
rect 515 72 603 106
rect 637 72 653 106
rect 515 56 653 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o211a_0
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2802084
string GDS_START 2794990
<< end >>
