magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4370 1975
<< nwell >>
rect -38 331 3110 704
<< pwell >>
rect 1606 229 1903 273
rect 2206 241 2598 243
rect 2206 229 3061 241
rect 1054 183 3061 229
rect 811 157 3061 183
rect 51 49 3061 157
rect 0 0 3072 49
<< scnmos >>
rect 130 47 160 131
rect 238 47 268 131
rect 310 47 340 131
rect 441 47 471 131
rect 513 47 543 131
rect 599 47 629 131
rect 890 73 920 157
rect 1133 119 1163 203
rect 1219 119 1249 203
rect 1291 119 1321 203
rect 1500 119 1530 203
rect 1572 119 1602 203
rect 1705 119 1735 247
rect 1794 119 1824 247
rect 1899 119 1929 203
rect 1971 119 2001 203
rect 2043 119 2073 203
rect 2285 133 2315 217
rect 2403 49 2433 217
rect 2489 49 2519 217
rect 2594 49 2624 133
rect 2792 47 2822 215
rect 2952 47 2982 215
<< scpmoshvt >>
rect 80 467 110 595
rect 166 467 196 595
rect 238 467 268 595
rect 346 467 376 595
rect 448 467 478 595
rect 641 467 671 595
rect 890 389 920 517
rect 1159 463 1189 547
rect 1245 463 1275 547
rect 1317 463 1347 547
rect 1435 463 1465 547
rect 1521 463 1551 547
rect 1667 379 1697 547
rect 1769 408 1799 576
rect 1874 492 1904 576
rect 1946 492 1976 576
rect 2064 492 2094 576
rect 2328 367 2358 451
rect 2433 367 2463 619
rect 2519 367 2549 619
rect 2624 367 2654 495
rect 2866 367 2896 619
rect 2952 367 2982 619
<< ndiff >>
rect 1632 203 1705 247
rect 1080 178 1133 203
rect 77 105 130 131
rect 77 71 85 105
rect 119 71 130 105
rect 77 47 130 71
rect 160 105 238 131
rect 160 71 182 105
rect 216 71 238 105
rect 160 47 238 71
rect 268 47 310 131
rect 340 106 441 131
rect 340 72 394 106
rect 428 72 441 106
rect 340 47 441 72
rect 471 47 513 131
rect 543 99 599 131
rect 543 65 554 99
rect 588 65 599 99
rect 543 47 599 65
rect 629 105 682 131
rect 629 71 640 105
rect 674 71 682 105
rect 837 129 890 157
rect 837 95 845 129
rect 879 95 890 129
rect 837 73 890 95
rect 920 130 973 157
rect 920 96 931 130
rect 965 96 973 130
rect 1080 144 1088 178
rect 1122 144 1133 178
rect 1080 119 1133 144
rect 1163 178 1219 203
rect 1163 144 1174 178
rect 1208 144 1219 178
rect 1163 119 1219 144
rect 1249 119 1291 203
rect 1321 178 1374 203
rect 1321 144 1332 178
rect 1366 144 1374 178
rect 1321 119 1374 144
rect 1447 178 1500 203
rect 1447 144 1455 178
rect 1489 144 1500 178
rect 1447 119 1500 144
rect 1530 119 1572 203
rect 1602 135 1705 203
rect 1602 119 1644 135
rect 920 73 973 96
rect 629 47 682 71
rect 1632 101 1644 119
rect 1678 119 1705 135
rect 1735 119 1794 247
rect 1824 203 1877 247
rect 1824 168 1899 203
rect 1824 134 1843 168
rect 1877 134 1899 168
rect 1824 119 1899 134
rect 1929 119 1971 203
rect 2001 119 2043 203
rect 2073 175 2126 203
rect 2073 141 2084 175
rect 2118 141 2126 175
rect 2073 119 2126 141
rect 2232 192 2285 217
rect 2232 158 2240 192
rect 2274 158 2285 192
rect 2232 133 2285 158
rect 2315 183 2403 217
rect 2315 149 2326 183
rect 2360 149 2403 183
rect 2315 133 2403 149
rect 1678 101 1690 119
rect 1632 93 1690 101
rect 2337 95 2403 133
rect 2337 61 2358 95
rect 2392 61 2403 95
rect 2337 49 2403 61
rect 2433 205 2489 217
rect 2433 171 2444 205
rect 2478 171 2489 205
rect 2433 103 2489 171
rect 2433 69 2444 103
rect 2478 69 2489 103
rect 2433 49 2489 69
rect 2519 205 2572 217
rect 2519 171 2530 205
rect 2564 171 2572 205
rect 2519 133 2572 171
rect 2739 203 2792 215
rect 2739 169 2747 203
rect 2781 169 2792 203
rect 2519 95 2594 133
rect 2519 61 2549 95
rect 2583 61 2594 95
rect 2519 49 2594 61
rect 2624 108 2677 133
rect 2624 74 2635 108
rect 2669 74 2677 108
rect 2624 49 2677 74
rect 2739 93 2792 169
rect 2739 59 2747 93
rect 2781 59 2792 93
rect 2739 47 2792 59
rect 2822 203 2952 215
rect 2822 169 2833 203
rect 2867 169 2907 203
rect 2941 169 2952 203
rect 2822 101 2952 169
rect 2822 67 2833 101
rect 2867 67 2907 101
rect 2941 67 2952 101
rect 2822 47 2952 67
rect 2982 203 3035 215
rect 2982 169 2993 203
rect 3027 169 3035 203
rect 2982 93 3035 169
rect 2982 59 2993 93
rect 3027 59 3035 93
rect 2982 47 3035 59
<< pdiff >>
rect 493 631 551 639
rect 493 597 505 631
rect 539 597 551 631
rect 493 595 551 597
rect 27 581 80 595
rect 27 547 35 581
rect 69 547 80 581
rect 27 513 80 547
rect 27 479 35 513
rect 69 479 80 513
rect 27 467 80 479
rect 110 587 166 595
rect 110 553 121 587
rect 155 553 166 587
rect 110 467 166 553
rect 196 467 238 595
rect 268 557 346 595
rect 268 523 301 557
rect 335 523 346 557
rect 268 467 346 523
rect 376 467 448 595
rect 478 467 641 595
rect 671 509 728 595
rect 671 475 682 509
rect 716 475 728 509
rect 671 467 728 475
rect 810 585 868 595
rect 810 551 822 585
rect 856 551 868 585
rect 810 517 868 551
rect 2380 607 2433 619
rect 1991 576 2049 605
rect 1362 564 1420 572
rect 1362 547 1374 564
rect 1106 522 1159 547
rect 810 389 890 517
rect 920 431 977 517
rect 1106 488 1114 522
rect 1148 488 1159 522
rect 1106 463 1159 488
rect 1189 522 1245 547
rect 1189 488 1200 522
rect 1234 488 1245 522
rect 1189 463 1245 488
rect 1275 463 1317 547
rect 1347 530 1374 547
rect 1408 547 1420 564
rect 1594 564 1652 572
rect 1594 547 1606 564
rect 1408 530 1435 547
rect 1347 463 1435 530
rect 1465 522 1521 547
rect 1465 488 1476 522
rect 1510 488 1521 522
rect 1465 463 1521 488
rect 1551 530 1606 547
rect 1640 547 1652 564
rect 1719 547 1769 576
rect 1640 530 1667 547
rect 1551 463 1667 530
rect 920 397 931 431
rect 965 397 977 431
rect 920 389 977 397
rect 1617 379 1667 463
rect 1697 408 1769 547
rect 1799 561 1874 576
rect 1799 527 1810 561
rect 1844 527 1874 561
rect 1799 492 1874 527
rect 1904 492 1946 576
rect 1976 551 2064 576
rect 1976 517 2003 551
rect 2037 517 2064 551
rect 1976 492 2064 517
rect 2094 551 2151 576
rect 2094 517 2105 551
rect 2139 517 2151 551
rect 2094 492 2151 517
rect 2380 573 2388 607
rect 2422 573 2433 607
rect 2380 513 2433 573
rect 1799 408 1852 492
rect 1697 379 1747 408
rect 2380 479 2388 513
rect 2422 479 2433 513
rect 2380 451 2433 479
rect 2275 413 2328 451
rect 2275 379 2283 413
rect 2317 379 2328 413
rect 2275 367 2328 379
rect 2358 367 2433 451
rect 2463 599 2519 619
rect 2463 565 2474 599
rect 2508 565 2519 599
rect 2463 507 2519 565
rect 2463 473 2474 507
rect 2508 473 2519 507
rect 2463 413 2519 473
rect 2463 379 2474 413
rect 2508 379 2519 413
rect 2463 367 2519 379
rect 2549 607 2602 619
rect 2549 573 2560 607
rect 2594 573 2602 607
rect 2549 506 2602 573
rect 2813 607 2866 619
rect 2813 573 2821 607
rect 2855 573 2866 607
rect 2549 472 2560 506
rect 2594 495 2602 506
rect 2813 508 2866 573
rect 2594 472 2624 495
rect 2549 413 2624 472
rect 2549 379 2569 413
rect 2603 379 2624 413
rect 2549 367 2624 379
rect 2654 483 2707 495
rect 2654 449 2665 483
rect 2699 449 2707 483
rect 2654 413 2707 449
rect 2654 379 2665 413
rect 2699 379 2707 413
rect 2654 367 2707 379
rect 2813 474 2821 508
rect 2855 474 2866 508
rect 2813 414 2866 474
rect 2813 380 2821 414
rect 2855 380 2866 414
rect 2813 367 2866 380
rect 2896 599 2952 619
rect 2896 565 2907 599
rect 2941 565 2952 599
rect 2896 498 2952 565
rect 2896 464 2907 498
rect 2941 464 2952 498
rect 2896 409 2952 464
rect 2896 375 2907 409
rect 2941 375 2952 409
rect 2896 367 2952 375
rect 2982 607 3035 619
rect 2982 573 2993 607
rect 3027 573 3035 607
rect 2982 508 3035 573
rect 2982 474 2993 508
rect 3027 474 3035 508
rect 2982 414 3035 474
rect 2982 380 2993 414
rect 3027 380 3035 414
rect 2982 367 3035 380
<< ndiffc >>
rect 85 71 119 105
rect 182 71 216 105
rect 394 72 428 106
rect 554 65 588 99
rect 640 71 674 105
rect 845 95 879 129
rect 931 96 965 130
rect 1088 144 1122 178
rect 1174 144 1208 178
rect 1332 144 1366 178
rect 1455 144 1489 178
rect 1644 101 1678 135
rect 1843 134 1877 168
rect 2084 141 2118 175
rect 2240 158 2274 192
rect 2326 149 2360 183
rect 2358 61 2392 95
rect 2444 171 2478 205
rect 2444 69 2478 103
rect 2530 171 2564 205
rect 2747 169 2781 203
rect 2549 61 2583 95
rect 2635 74 2669 108
rect 2747 59 2781 93
rect 2833 169 2867 203
rect 2907 169 2941 203
rect 2833 67 2867 101
rect 2907 67 2941 101
rect 2993 169 3027 203
rect 2993 59 3027 93
<< pdiffc >>
rect 505 597 539 631
rect 35 547 69 581
rect 35 479 69 513
rect 121 553 155 587
rect 301 523 335 557
rect 682 475 716 509
rect 822 551 856 585
rect 1114 488 1148 522
rect 1200 488 1234 522
rect 1374 530 1408 564
rect 1476 488 1510 522
rect 1606 530 1640 564
rect 931 397 965 431
rect 1810 527 1844 561
rect 2003 517 2037 551
rect 2105 517 2139 551
rect 2388 573 2422 607
rect 2388 479 2422 513
rect 2283 379 2317 413
rect 2474 565 2508 599
rect 2474 473 2508 507
rect 2474 379 2508 413
rect 2560 573 2594 607
rect 2821 573 2855 607
rect 2560 472 2594 506
rect 2569 379 2603 413
rect 2665 449 2699 483
rect 2665 379 2699 413
rect 2821 474 2855 508
rect 2821 380 2855 414
rect 2907 565 2941 599
rect 2907 464 2941 498
rect 2907 375 2941 409
rect 2993 573 3027 607
rect 2993 474 3027 508
rect 2993 380 3027 414
<< poly >>
rect 80 595 110 621
rect 166 595 196 621
rect 238 595 268 621
rect 346 595 376 621
rect 448 595 478 621
rect 641 595 671 621
rect 890 615 1799 645
rect 2433 619 2463 645
rect 2519 619 2549 645
rect 2866 619 2896 645
rect 2952 619 2982 645
rect 890 517 920 615
rect 1159 547 1189 573
rect 1245 547 1275 615
rect 1769 576 1799 615
rect 1874 576 1904 602
rect 1946 576 1976 602
rect 2064 576 2094 602
rect 1317 547 1347 573
rect 80 435 110 467
rect 166 435 196 467
rect 80 419 196 435
rect 80 385 127 419
rect 161 385 196 419
rect 80 369 196 385
rect 238 429 268 467
rect 238 413 304 429
rect 238 379 254 413
rect 288 379 304 413
rect 80 321 110 369
rect 238 363 304 379
rect 80 291 160 321
rect 346 297 376 467
rect 448 445 478 467
rect 448 415 592 445
rect 130 131 160 291
rect 202 281 376 297
rect 202 247 218 281
rect 252 267 376 281
rect 418 351 484 367
rect 418 317 434 351
rect 468 317 484 351
rect 418 283 484 317
rect 252 247 268 267
rect 202 213 268 247
rect 418 249 434 283
rect 468 249 484 283
rect 418 233 484 249
rect 526 366 592 415
rect 526 332 542 366
rect 576 332 592 366
rect 526 316 592 332
rect 202 179 218 213
rect 252 179 268 213
rect 202 163 268 179
rect 238 131 268 163
rect 310 203 376 219
rect 310 169 326 203
rect 360 169 376 203
rect 310 153 376 169
rect 310 131 340 153
rect 441 131 471 233
rect 526 185 556 316
rect 641 219 671 467
rect 1435 547 1465 573
rect 1521 547 1551 573
rect 1667 547 1697 573
rect 1009 415 1075 431
rect 890 313 920 389
rect 513 155 556 185
rect 599 203 671 219
rect 599 169 615 203
rect 649 169 671 203
rect 815 297 920 313
rect 1009 381 1025 415
rect 1059 381 1075 415
rect 1009 369 1075 381
rect 1159 369 1189 463
rect 1245 437 1275 463
rect 1317 441 1347 463
rect 1317 415 1393 441
rect 1317 411 1343 415
rect 1327 381 1343 411
rect 1377 381 1393 415
rect 1009 353 1285 369
rect 1327 365 1393 381
rect 1009 347 1235 353
rect 1009 313 1025 347
rect 1059 339 1235 347
rect 1059 313 1075 339
rect 1009 297 1075 313
rect 1219 319 1235 339
rect 1269 319 1285 353
rect 1219 303 1285 319
rect 815 263 831 297
rect 865 263 920 297
rect 815 229 920 263
rect 815 195 831 229
rect 865 195 920 229
rect 1133 203 1163 229
rect 1219 203 1249 303
rect 1333 255 1363 365
rect 1291 225 1363 255
rect 1435 291 1465 463
rect 1521 431 1551 463
rect 1507 415 1602 431
rect 1507 381 1523 415
rect 1557 381 1602 415
rect 1507 365 1602 381
rect 1769 382 1799 408
rect 1435 275 1501 291
rect 1435 241 1451 275
rect 1485 255 1501 275
rect 1485 241 1530 255
rect 1435 225 1530 241
rect 1291 203 1321 225
rect 1500 203 1530 225
rect 1572 203 1602 365
rect 1667 335 1697 379
rect 1874 340 1904 492
rect 1946 399 1976 492
rect 2064 460 2094 492
rect 2064 444 2193 460
rect 2328 451 2358 477
rect 2064 430 2143 444
rect 2127 410 2143 430
rect 2177 410 2193 444
rect 1946 369 2001 399
rect 2127 376 2193 410
rect 1663 319 1729 335
rect 1663 285 1679 319
rect 1713 299 1729 319
rect 1777 324 1904 340
rect 1713 285 1735 299
rect 1663 269 1735 285
rect 1777 290 1793 324
rect 1827 310 1904 324
rect 1971 353 2069 369
rect 1971 319 2019 353
rect 2053 319 2069 353
rect 1827 290 1843 310
rect 1777 274 1843 290
rect 1971 303 2069 319
rect 2127 342 2143 376
rect 2177 342 2193 376
rect 2624 495 2654 521
rect 2127 326 2193 342
rect 2328 335 2358 367
rect 1705 247 1735 269
rect 1794 247 1824 274
rect 815 179 920 195
rect 513 131 543 155
rect 599 153 671 169
rect 890 157 920 179
rect 599 131 629 153
rect 890 51 920 73
rect 1133 51 1163 119
rect 1219 93 1249 119
rect 1291 93 1321 119
rect 1500 93 1530 119
rect 1572 93 1602 119
rect 1899 203 1929 229
rect 1971 203 2001 303
rect 2127 255 2157 326
rect 2249 319 2358 335
rect 2249 285 2265 319
rect 2299 299 2358 319
rect 2433 299 2463 367
rect 2519 299 2549 367
rect 2624 299 2654 367
rect 2866 321 2896 367
rect 2952 321 2982 367
rect 2299 285 2654 299
rect 2249 269 2654 285
rect 2743 305 2982 321
rect 2743 271 2759 305
rect 2793 271 2837 305
rect 2871 271 2982 305
rect 2043 225 2157 255
rect 2043 203 2073 225
rect 2285 217 2315 269
rect 2403 217 2433 269
rect 2489 217 2519 269
rect 1705 93 1735 119
rect 1794 93 1824 119
rect 1899 51 1929 119
rect 1971 93 2001 119
rect 2043 93 2073 119
rect 2285 107 2315 133
rect 130 21 160 47
rect 238 21 268 47
rect 310 21 340 47
rect 441 21 471 47
rect 513 21 543 47
rect 599 21 629 47
rect 890 21 1929 51
rect 2594 133 2624 269
rect 2743 255 2982 271
rect 2792 215 2822 255
rect 2952 215 2982 255
rect 2403 23 2433 49
rect 2489 23 2519 49
rect 2594 23 2624 49
rect 2792 21 2822 47
rect 2952 21 2982 47
<< polycont >>
rect 127 385 161 419
rect 254 379 288 413
rect 218 247 252 281
rect 434 317 468 351
rect 434 249 468 283
rect 542 332 576 366
rect 218 179 252 213
rect 326 169 360 203
rect 615 169 649 203
rect 1025 381 1059 415
rect 1343 381 1377 415
rect 1025 313 1059 347
rect 1235 319 1269 353
rect 831 263 865 297
rect 831 195 865 229
rect 1523 381 1557 415
rect 1451 241 1485 275
rect 2143 410 2177 444
rect 1679 285 1713 319
rect 1793 290 1827 324
rect 2019 319 2053 353
rect 2143 342 2177 376
rect 2265 285 2299 319
rect 2759 271 2793 305
rect 2837 271 2871 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 19 581 71 597
rect 19 547 35 581
rect 69 547 71 581
rect 19 513 71 547
rect 105 587 171 649
rect 489 631 555 649
rect 489 597 505 631
rect 539 597 555 631
rect 489 595 555 597
rect 105 553 121 587
rect 155 553 171 587
rect 612 561 786 599
rect 105 532 171 553
rect 285 557 646 561
rect 285 523 301 557
rect 335 523 646 557
rect 285 517 646 523
rect 19 479 35 513
rect 69 479 71 513
rect 19 197 71 479
rect 111 483 197 498
rect 111 449 468 483
rect 111 419 177 449
rect 111 385 127 419
rect 161 385 177 419
rect 111 231 177 385
rect 238 413 360 415
rect 238 379 254 413
rect 288 379 360 413
rect 238 363 360 379
rect 211 281 269 297
rect 211 247 218 281
rect 252 247 269 281
rect 211 213 269 247
rect 211 197 218 213
rect 19 179 218 197
rect 252 179 269 213
rect 19 163 269 179
rect 303 203 360 363
rect 418 351 468 449
rect 418 317 434 351
rect 418 283 468 317
rect 502 366 578 450
rect 502 332 542 366
rect 576 332 578 366
rect 502 307 578 332
rect 418 249 434 283
rect 612 273 646 517
rect 418 233 468 249
rect 504 239 646 273
rect 680 509 718 527
rect 680 475 682 509
rect 716 475 718 509
rect 680 313 718 475
rect 752 501 786 561
rect 820 585 872 649
rect 820 551 822 585
rect 856 551 872 585
rect 820 535 872 551
rect 1358 564 1424 649
rect 1095 522 1156 541
rect 1095 501 1114 522
rect 752 488 1114 501
rect 1148 488 1156 522
rect 752 472 1156 488
rect 1190 522 1250 538
rect 1358 530 1374 564
rect 1408 530 1424 564
rect 1590 564 1656 649
rect 1358 528 1424 530
rect 1190 488 1200 522
rect 1234 488 1250 522
rect 1460 522 1526 538
rect 1590 530 1606 564
rect 1640 530 1656 564
rect 1590 528 1656 530
rect 1794 561 1967 577
rect 1460 494 1476 522
rect 752 467 1131 472
rect 915 431 1059 433
rect 915 397 931 431
rect 965 415 1059 431
rect 965 397 1025 415
rect 915 381 1025 397
rect 915 347 1059 381
rect 915 313 1025 347
rect 680 297 881 313
rect 680 263 831 297
rect 865 263 881 297
rect 680 239 881 263
rect 303 169 326 203
rect 504 175 538 239
rect 710 229 881 239
rect 19 105 132 163
rect 19 71 85 105
rect 119 71 132 105
rect 19 55 132 71
rect 166 105 232 121
rect 166 71 182 105
rect 216 71 232 105
rect 303 77 360 169
rect 394 141 538 175
rect 599 203 676 205
rect 599 169 615 203
rect 649 169 676 203
rect 599 155 676 169
rect 710 195 831 229
rect 865 195 881 229
rect 710 179 881 195
rect 915 297 1059 313
rect 394 106 444 141
rect 710 121 788 179
rect 166 17 232 71
rect 428 72 444 106
rect 394 56 444 72
rect 538 99 604 107
rect 538 65 554 99
rect 588 65 604 99
rect 538 17 604 65
rect 638 105 788 121
rect 638 71 640 105
rect 674 71 788 105
rect 638 55 788 71
rect 829 129 881 145
rect 829 95 845 129
rect 879 95 881 129
rect 829 17 881 95
rect 915 130 981 297
rect 1095 247 1131 467
rect 1190 438 1250 488
rect 915 96 931 130
rect 965 96 981 130
rect 1072 178 1131 247
rect 1072 144 1088 178
rect 1122 144 1131 178
rect 1072 128 1131 144
rect 1165 404 1250 438
rect 1327 488 1476 494
rect 1510 494 1526 522
rect 1794 527 1810 561
rect 1844 527 1967 561
rect 1794 511 1967 527
rect 1510 488 1643 494
rect 1327 475 1643 488
rect 1327 460 1897 475
rect 1327 415 1393 460
rect 1609 441 1897 460
rect 1165 269 1199 404
rect 1327 381 1343 415
rect 1377 381 1393 415
rect 1453 424 1573 426
rect 1453 390 1471 424
rect 1505 415 1573 424
rect 1505 390 1523 415
rect 1453 381 1523 390
rect 1557 381 1573 415
rect 1453 379 1573 381
rect 1609 371 1829 405
rect 1233 353 1285 369
rect 1233 319 1235 353
rect 1269 345 1285 353
rect 1609 345 1643 371
rect 1269 319 1643 345
rect 1233 309 1643 319
rect 1677 319 1715 335
rect 1233 303 1286 309
rect 1677 285 1679 319
rect 1713 285 1715 319
rect 1677 275 1715 285
rect 1435 269 1451 275
rect 1165 241 1451 269
rect 1485 241 1715 275
rect 1777 324 1829 371
rect 1777 290 1793 324
rect 1827 290 1829 324
rect 1777 274 1829 290
rect 1165 228 1501 241
rect 1863 240 1897 441
rect 1165 178 1224 228
rect 1749 207 1897 240
rect 1558 206 1897 207
rect 1933 467 1967 511
rect 2001 551 2039 649
rect 2372 607 2424 649
rect 2372 573 2388 607
rect 2422 573 2424 607
rect 2001 517 2003 551
rect 2037 517 2039 551
rect 2001 501 2039 517
rect 2073 551 2247 567
rect 2073 517 2105 551
rect 2139 517 2247 551
rect 2073 501 2247 517
rect 2073 467 2107 501
rect 1933 431 2107 467
rect 2141 444 2179 460
rect 1558 194 1783 206
rect 1165 144 1174 178
rect 1208 144 1224 178
rect 1165 128 1224 144
rect 1316 178 1382 194
rect 1316 144 1332 178
rect 1366 144 1382 178
rect 915 82 981 96
rect 1316 17 1382 144
rect 1451 178 1783 194
rect 1451 144 1455 178
rect 1489 173 1783 178
rect 1489 144 1592 173
rect 1933 172 1967 431
rect 2141 390 2143 444
rect 2177 390 2179 444
rect 2141 376 2179 390
rect 2003 353 2069 369
rect 2003 319 2019 353
rect 2053 319 2069 353
rect 2141 342 2143 376
rect 2177 342 2179 376
rect 2141 326 2179 342
rect 2213 329 2247 501
rect 2372 513 2424 573
rect 2372 479 2388 513
rect 2422 479 2424 513
rect 2372 463 2424 479
rect 2458 599 2517 615
rect 2458 565 2474 599
rect 2508 565 2517 599
rect 2458 507 2517 565
rect 2458 473 2474 507
rect 2508 473 2517 507
rect 2283 413 2385 429
rect 2458 424 2517 473
rect 2317 379 2385 413
rect 2283 363 2385 379
rect 2003 251 2069 319
rect 2213 319 2315 329
rect 2213 285 2265 319
rect 2299 285 2315 319
rect 2351 251 2385 363
rect 2003 217 2385 251
rect 2431 413 2517 424
rect 2431 379 2474 413
rect 2508 379 2517 413
rect 2431 363 2517 379
rect 2551 607 2619 649
rect 2551 573 2560 607
rect 2594 573 2619 607
rect 2551 506 2619 573
rect 2551 472 2560 506
rect 2594 472 2619 506
rect 2805 607 2871 649
rect 2805 573 2821 607
rect 2855 573 2871 607
rect 2805 508 2871 573
rect 2551 413 2619 472
rect 2551 379 2569 413
rect 2603 379 2619 413
rect 2551 363 2619 379
rect 2653 483 2715 499
rect 2653 449 2665 483
rect 2699 449 2715 483
rect 2653 413 2715 449
rect 2653 379 2665 413
rect 2699 379 2715 413
rect 2224 192 2276 217
rect 1451 128 1592 144
rect 1827 168 1967 172
rect 1628 135 1694 139
rect 1628 101 1644 135
rect 1678 101 1694 135
rect 1827 134 1843 168
rect 1877 134 1967 168
rect 1827 118 1967 134
rect 2068 175 2134 183
rect 2068 141 2084 175
rect 2118 141 2134 175
rect 2224 158 2240 192
rect 2274 158 2276 192
rect 2431 205 2492 363
rect 2653 321 2715 379
rect 2805 474 2821 508
rect 2855 474 2871 508
rect 2805 414 2871 474
rect 2805 380 2821 414
rect 2855 380 2871 414
rect 2805 364 2871 380
rect 2905 599 2955 615
rect 2905 565 2907 599
rect 2941 565 2955 599
rect 2905 498 2955 565
rect 2905 464 2907 498
rect 2941 464 2955 498
rect 2905 409 2955 464
rect 2905 375 2907 409
rect 2941 375 2955 409
rect 2653 305 2871 321
rect 2653 271 2759 305
rect 2793 271 2837 305
rect 2653 255 2871 271
rect 2224 142 2276 158
rect 2310 149 2326 183
rect 2360 149 2397 183
rect 1628 17 1694 101
rect 2068 17 2134 141
rect 2310 95 2397 149
rect 2310 61 2358 95
rect 2392 61 2397 95
rect 2310 17 2397 61
rect 2431 171 2444 205
rect 2478 171 2492 205
rect 2431 103 2492 171
rect 2431 69 2444 103
rect 2478 69 2492 103
rect 2431 53 2492 69
rect 2526 205 2593 221
rect 2526 171 2530 205
rect 2564 171 2593 205
rect 2526 95 2593 171
rect 2653 124 2695 255
rect 2905 219 2955 375
rect 2989 607 3043 649
rect 2989 573 2993 607
rect 3027 573 3043 607
rect 2989 508 3043 573
rect 2989 474 2993 508
rect 3027 474 3043 508
rect 2989 414 3043 474
rect 2989 380 2993 414
rect 3027 380 3043 414
rect 2989 364 3043 380
rect 2526 61 2549 95
rect 2583 61 2593 95
rect 2526 17 2593 61
rect 2627 108 2695 124
rect 2627 74 2635 108
rect 2669 74 2695 108
rect 2627 58 2695 74
rect 2731 203 2788 219
rect 2731 169 2747 203
rect 2781 169 2788 203
rect 2731 93 2788 169
rect 2731 59 2747 93
rect 2781 59 2788 93
rect 2731 17 2788 59
rect 2822 203 2955 219
rect 2822 169 2833 203
rect 2867 169 2907 203
rect 2941 169 2955 203
rect 2822 101 2955 169
rect 2822 67 2833 101
rect 2867 67 2907 101
rect 2941 67 2955 101
rect 2822 51 2955 67
rect 2989 203 3043 219
rect 2989 169 2993 203
rect 3027 169 3043 203
rect 2989 93 3043 169
rect 2989 59 2993 93
rect 3027 59 3043 93
rect 2989 17 3043 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 1471 390 1505 424
rect 2143 410 2177 424
rect 2143 390 2177 410
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 683 3072 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 0 617 3072 649
rect 1459 424 1517 430
rect 1459 390 1471 424
rect 1505 421 1517 424
rect 2131 424 2189 430
rect 2131 421 2143 424
rect 1505 393 2143 421
rect 1505 390 1517 393
rect 1459 384 1517 390
rect 2131 390 2143 393
rect 2177 390 2189 424
rect 2131 384 2189 390
rect 0 17 3072 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
rect 0 -49 3072 -17
<< labels >>
flabel pwell s 0 0 3072 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 3072 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfsbp_2
flabel comment s 1154 355 1154 355 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 2143 390 2177 424 0 FreeSans 200 0 0 0 SET_B
port 5 nsew signal input
flabel metal1 s 0 617 3072 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 3072 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 2911 94 2945 128 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2911 168 2945 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2911 242 2945 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2911 316 2945 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2911 390 2945 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2911 464 2945 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2911 538 2945 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2431 94 2465 128 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2431 168 2465 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2431 242 2465 276 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2431 316 2465 350 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2431 390 2465 424 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3072 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5615834
string GDS_START 5593972
<< end >>
