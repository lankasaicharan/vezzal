magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2494 1852
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1127 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 267 47 297 177
rect 371 47 401 177
rect 455 47 485 177
rect 559 47 589 177
rect 643 47 673 177
rect 747 47 777 177
rect 831 47 861 177
rect 935 47 965 177
rect 1019 47 1049 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
<< ndiff >>
rect 27 169 89 177
rect 27 135 45 169
rect 79 135 89 169
rect 27 101 89 135
rect 27 67 45 101
rect 79 67 89 101
rect 27 47 89 67
rect 119 97 183 177
rect 119 63 135 97
rect 169 63 183 97
rect 119 47 183 63
rect 213 169 267 177
rect 213 135 223 169
rect 257 135 267 169
rect 213 101 267 135
rect 213 67 223 101
rect 257 67 267 101
rect 213 47 267 67
rect 297 97 371 177
rect 297 63 317 97
rect 351 63 371 97
rect 297 47 371 63
rect 401 169 455 177
rect 401 135 411 169
rect 445 135 455 169
rect 401 101 455 135
rect 401 67 411 101
rect 445 67 455 101
rect 401 47 455 67
rect 485 97 559 177
rect 485 63 505 97
rect 539 63 559 97
rect 485 47 559 63
rect 589 169 643 177
rect 589 135 599 169
rect 633 135 643 169
rect 589 101 643 135
rect 589 67 599 101
rect 633 67 643 101
rect 589 47 643 67
rect 673 97 747 177
rect 673 63 693 97
rect 727 63 747 97
rect 673 47 747 63
rect 777 169 831 177
rect 777 135 787 169
rect 821 135 831 169
rect 777 101 831 135
rect 777 67 787 101
rect 821 67 831 101
rect 777 47 831 67
rect 861 97 935 177
rect 861 63 881 97
rect 915 63 935 97
rect 861 47 935 63
rect 965 169 1019 177
rect 965 135 975 169
rect 1009 135 1019 169
rect 965 101 1019 135
rect 965 67 975 101
rect 1009 67 1019 101
rect 965 47 1019 67
rect 1049 161 1101 177
rect 1049 127 1059 161
rect 1093 127 1101 161
rect 1049 93 1101 127
rect 1049 59 1059 93
rect 1093 59 1101 93
rect 1049 47 1101 59
<< pdiff >>
rect 27 479 81 497
rect 27 445 35 479
rect 69 445 81 479
rect 27 411 81 445
rect 27 377 35 411
rect 69 377 81 411
rect 27 343 81 377
rect 27 309 35 343
rect 69 309 81 343
rect 27 297 81 309
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 297 175 383
rect 211 479 269 497
rect 211 445 223 479
rect 257 445 269 479
rect 211 411 269 445
rect 211 377 223 411
rect 257 377 269 411
rect 211 343 269 377
rect 211 309 223 343
rect 257 309 269 343
rect 211 297 269 309
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 297 363 383
rect 399 463 457 497
rect 399 429 411 463
rect 445 429 457 463
rect 399 368 457 429
rect 399 334 411 368
rect 445 334 457 368
rect 399 297 457 334
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 297 551 383
rect 587 463 645 497
rect 587 429 599 463
rect 633 429 645 463
rect 587 368 645 429
rect 587 334 599 368
rect 633 334 645 368
rect 587 297 645 334
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 297 739 383
rect 775 463 833 497
rect 775 429 787 463
rect 821 429 833 463
rect 775 368 833 429
rect 775 334 787 368
rect 821 334 833 368
rect 775 297 833 334
rect 869 485 927 497
rect 869 451 881 485
rect 915 451 927 485
rect 869 417 927 451
rect 869 383 881 417
rect 915 383 927 417
rect 869 297 927 383
rect 963 463 1021 497
rect 963 429 975 463
rect 1009 429 1021 463
rect 963 368 1021 429
rect 963 334 975 368
rect 1009 334 1021 368
rect 963 297 1021 334
rect 1057 485 1111 497
rect 1057 451 1069 485
rect 1103 451 1111 485
rect 1057 417 1111 451
rect 1057 383 1069 417
rect 1103 383 1111 417
rect 1057 349 1111 383
rect 1057 315 1069 349
rect 1103 315 1111 349
rect 1057 297 1111 315
<< ndiffc >>
rect 45 135 79 169
rect 45 67 79 101
rect 135 63 169 97
rect 223 135 257 169
rect 223 67 257 101
rect 317 63 351 97
rect 411 135 445 169
rect 411 67 445 101
rect 505 63 539 97
rect 599 135 633 169
rect 599 67 633 101
rect 693 63 727 97
rect 787 135 821 169
rect 787 67 821 101
rect 881 63 915 97
rect 975 135 1009 169
rect 975 67 1009 101
rect 1059 127 1093 161
rect 1059 59 1093 93
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 129 451 163 485
rect 129 383 163 417
rect 223 445 257 479
rect 223 377 257 411
rect 223 309 257 343
rect 317 451 351 485
rect 317 383 351 417
rect 411 429 445 463
rect 411 334 445 368
rect 505 451 539 485
rect 505 383 539 417
rect 599 429 633 463
rect 599 334 633 368
rect 693 451 727 485
rect 693 383 727 417
rect 787 429 821 463
rect 787 334 821 368
rect 881 451 915 485
rect 881 383 915 417
rect 975 429 1009 463
rect 975 334 1009 368
rect 1069 451 1103 485
rect 1069 383 1103 417
rect 1069 315 1103 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 79 261 119 282
rect 28 259 119 261
rect 173 259 213 282
rect 267 259 307 282
rect 28 249 307 259
rect 28 215 44 249
rect 78 215 112 249
rect 146 215 180 249
rect 214 215 307 249
rect 28 205 307 215
rect 361 259 401 282
rect 455 259 495 282
rect 549 259 589 282
rect 643 259 683 282
rect 737 259 777 282
rect 831 259 871 282
rect 925 259 965 282
rect 1019 259 1059 282
rect 361 249 1059 259
rect 361 215 419 249
rect 453 215 487 249
rect 521 215 555 249
rect 589 215 623 249
rect 657 215 691 249
rect 725 215 759 249
rect 793 215 1059 249
rect 361 205 1059 215
rect 28 203 119 205
rect 89 177 119 203
rect 183 177 213 205
rect 267 177 297 205
rect 371 177 401 205
rect 455 177 485 205
rect 559 177 589 205
rect 643 177 673 205
rect 747 177 777 205
rect 831 177 861 205
rect 935 177 965 205
rect 1019 177 1049 205
rect 89 21 119 47
rect 183 21 213 47
rect 267 21 297 47
rect 371 21 401 47
rect 455 21 485 47
rect 559 21 589 47
rect 643 21 673 47
rect 747 21 777 47
rect 831 21 861 47
rect 935 21 965 47
rect 1019 21 1049 47
<< polycont >>
rect 44 215 78 249
rect 112 215 146 249
rect 180 215 214 249
rect 419 215 453 249
rect 487 215 521 249
rect 555 215 589 249
rect 623 215 657 249
rect 691 215 725 249
rect 759 215 793 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 19 479 85 493
rect 19 445 35 479
rect 69 445 85 479
rect 19 411 85 445
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 119 485 173 527
rect 119 451 129 485
rect 163 451 173 485
rect 119 417 173 451
rect 119 383 129 417
rect 163 383 173 417
rect 119 367 173 383
rect 207 479 273 493
rect 207 445 223 479
rect 257 445 273 479
rect 207 411 273 445
rect 207 377 223 411
rect 257 377 273 411
rect 19 309 35 343
rect 69 323 85 343
rect 207 343 273 377
rect 307 485 361 527
rect 307 451 317 485
rect 351 451 361 485
rect 307 417 361 451
rect 307 383 317 417
rect 351 383 361 417
rect 307 367 361 383
rect 395 463 461 493
rect 395 429 411 463
rect 445 429 461 463
rect 395 368 461 429
rect 207 323 223 343
rect 69 309 223 323
rect 257 323 273 343
rect 395 334 411 368
rect 445 334 461 368
rect 495 485 549 527
rect 495 451 505 485
rect 539 451 549 485
rect 495 417 549 451
rect 495 383 505 417
rect 539 383 549 417
rect 495 367 549 383
rect 583 463 649 493
rect 583 429 599 463
rect 633 429 649 463
rect 583 368 649 429
rect 395 323 461 334
rect 583 334 599 368
rect 633 334 649 368
rect 683 485 737 527
rect 683 451 693 485
rect 727 451 737 485
rect 683 417 737 451
rect 683 383 693 417
rect 727 383 737 417
rect 683 367 737 383
rect 771 463 837 493
rect 771 429 787 463
rect 821 429 837 463
rect 771 368 837 429
rect 583 323 649 334
rect 771 334 787 368
rect 821 334 837 368
rect 871 485 925 527
rect 871 451 881 485
rect 915 451 925 485
rect 871 417 925 451
rect 871 383 881 417
rect 915 383 925 417
rect 871 367 925 383
rect 959 463 1025 493
rect 959 429 975 463
rect 1009 429 1025 463
rect 959 368 1025 429
rect 771 323 837 334
rect 959 334 975 368
rect 1009 334 1025 368
rect 959 323 1025 334
rect 257 309 319 323
rect 19 289 319 309
rect 395 289 1025 323
rect 1059 485 1119 527
rect 1059 451 1069 485
rect 1103 451 1119 485
rect 1059 417 1119 451
rect 1059 383 1069 417
rect 1103 383 1119 417
rect 1059 349 1119 383
rect 1059 315 1069 349
rect 1103 315 1119 349
rect 1059 297 1119 315
rect 28 249 248 255
rect 28 215 44 249
rect 78 215 112 249
rect 146 215 180 249
rect 214 215 248 249
rect 284 249 319 289
rect 858 255 1025 289
rect 284 215 419 249
rect 453 215 487 249
rect 521 215 555 249
rect 589 215 623 249
rect 657 215 691 249
rect 725 215 759 249
rect 793 215 809 249
rect 858 221 912 255
rect 946 221 984 255
rect 1018 221 1025 255
rect 284 181 319 215
rect 858 181 1025 221
rect 29 169 319 181
rect 29 135 45 169
rect 79 147 223 169
rect 79 135 89 147
rect 29 101 89 135
rect 213 135 223 147
rect 257 147 319 169
rect 395 169 1025 181
rect 257 135 267 147
rect 29 67 45 101
rect 79 67 89 101
rect 29 51 89 67
rect 123 97 179 113
rect 123 63 135 97
rect 169 63 179 97
rect 123 17 179 63
rect 213 101 267 135
rect 395 135 411 169
rect 445 147 599 169
rect 445 135 461 147
rect 213 67 223 101
rect 257 67 267 101
rect 213 51 267 67
rect 301 97 361 113
rect 301 63 317 97
rect 351 63 361 97
rect 301 17 361 63
rect 395 101 461 135
rect 583 135 599 147
rect 633 147 787 169
rect 633 135 649 147
rect 395 67 411 101
rect 445 67 461 101
rect 395 51 461 67
rect 495 97 549 113
rect 495 63 505 97
rect 539 63 549 97
rect 495 17 549 63
rect 583 101 649 135
rect 771 135 787 147
rect 821 147 975 169
rect 821 135 837 147
rect 583 67 599 101
rect 633 67 649 101
rect 583 51 649 67
rect 683 97 737 113
rect 683 63 693 97
rect 727 63 737 97
rect 683 17 737 63
rect 771 101 837 135
rect 959 135 975 147
rect 1009 135 1025 169
rect 771 67 787 101
rect 821 67 837 101
rect 771 51 837 67
rect 871 97 925 113
rect 871 63 881 97
rect 915 63 925 97
rect 871 17 925 63
rect 959 101 1025 135
rect 959 67 975 101
rect 1009 67 1025 101
rect 959 51 1025 67
rect 1059 161 1109 177
rect 1093 127 1109 161
rect 1059 93 1109 127
rect 1093 59 1109 93
rect 1059 17 1109 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 912 221 946 255
rect 984 221 1018 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 693 212 699 264
rect 751 212 763 264
rect 815 261 821 264
rect 815 255 1030 261
rect 815 221 912 255
rect 946 221 984 255
rect 1018 221 1030 255
rect 815 215 1030 221
rect 815 212 821 215
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< via1 >>
rect 699 212 751 264
rect 763 212 815 264
<< metal2 >>
rect 689 266 825 275
rect 745 264 769 266
rect 751 212 763 264
rect 745 210 769 212
rect 689 201 825 210
<< via2 >>
rect 689 264 745 266
rect 769 264 825 266
rect 689 212 699 264
rect 699 212 745 264
rect 769 212 815 264
rect 815 212 825 264
rect 689 210 745 212
rect 769 210 825 212
<< metal3 >>
rect 679 270 835 271
rect 679 206 685 270
rect 749 206 765 270
rect 829 206 835 270
rect 679 205 835 206
<< via3 >>
rect 685 266 749 270
rect 685 210 689 266
rect 689 210 745 266
rect 745 210 749 266
rect 685 206 749 210
rect 765 266 829 270
rect 765 210 769 266
rect 769 210 825 266
rect 825 210 829 266
rect 765 206 829 210
<< metal4 >>
rect 510 136 594 372
<< via4 >>
rect 274 136 510 372
rect 594 270 830 372
rect 594 206 685 270
rect 685 206 749 270
rect 749 206 765 270
rect 765 206 829 270
rect 829 206 830 270
rect 594 136 830 206
<< metal5 >>
rect 250 390 854 432
rect 250 372 854 389
rect 250 136 274 372
rect 510 136 594 372
rect 830 136 854 372
rect 250 112 854 136
<< rm5 >>
rect 250 389 854 390
<< labels >>
flabel metal5 s 250 391 854 432 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground input
flabel locali s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground input
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power input
rlabel comment s 0 0 0 0 4 probe_p_8
rlabel metal1 s 0 -48 1196 48 1 VGND
port 2 nsew ground input
rlabel metal1 s 0 496 1196 592 1 VPWR
port 5 nsew power input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 3591032
string GDS_START 3580508
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
string path 17.325 5.950 20.525 5.950 
<< end >>
