magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3046 1852
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 5 21 1728 203
rect 29 -17 63 21
<< scnmos >>
rect 83 47 113 177
rect 177 47 207 177
rect 271 47 301 177
rect 375 47 405 177
rect 459 47 489 177
rect 553 47 583 177
rect 647 47 677 177
rect 751 47 781 177
rect 835 47 865 177
rect 1022 47 1052 177
rect 1116 47 1146 177
rect 1244 47 1274 177
rect 1328 47 1358 177
rect 1422 47 1452 177
rect 1516 47 1546 177
rect 1610 47 1640 177
<< scpmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 273 297 309 497
rect 367 297 403 497
rect 461 297 497 497
rect 555 297 591 497
rect 649 297 685 497
rect 743 297 779 497
rect 954 297 990 497
rect 1048 297 1084 497
rect 1142 297 1178 497
rect 1236 297 1272 497
rect 1330 297 1366 497
rect 1424 297 1460 497
rect 1518 297 1554 497
rect 1612 297 1648 497
<< ndiff >>
rect 31 161 83 177
rect 31 127 39 161
rect 73 127 83 161
rect 31 93 83 127
rect 31 59 39 93
rect 73 59 83 93
rect 31 47 83 59
rect 113 93 177 177
rect 113 59 133 93
rect 167 59 177 93
rect 113 47 177 59
rect 207 157 271 177
rect 207 123 227 157
rect 261 123 271 157
rect 207 89 271 123
rect 207 55 227 89
rect 261 55 271 89
rect 207 47 271 55
rect 301 93 375 177
rect 301 59 321 93
rect 355 59 375 93
rect 301 47 375 59
rect 405 157 459 177
rect 405 123 415 157
rect 449 123 459 157
rect 405 89 459 123
rect 405 55 415 89
rect 449 55 459 89
rect 405 47 459 55
rect 489 93 553 177
rect 489 59 509 93
rect 543 59 553 93
rect 489 47 553 59
rect 583 157 647 177
rect 583 123 603 157
rect 637 123 647 157
rect 583 89 647 123
rect 583 55 603 89
rect 637 55 647 89
rect 583 47 647 55
rect 677 93 751 177
rect 677 59 697 93
rect 731 59 751 93
rect 677 47 751 59
rect 781 157 835 177
rect 781 123 791 157
rect 825 123 835 157
rect 781 89 835 123
rect 781 55 791 89
rect 825 55 835 89
rect 781 47 835 55
rect 865 89 1022 177
rect 865 55 900 89
rect 934 55 968 89
rect 1002 55 1022 89
rect 865 47 1022 55
rect 1052 129 1116 177
rect 1052 95 1072 129
rect 1106 95 1116 129
rect 1052 47 1116 95
rect 1146 89 1244 177
rect 1146 55 1178 89
rect 1212 55 1244 89
rect 1146 47 1244 55
rect 1274 129 1328 177
rect 1274 95 1284 129
rect 1318 95 1328 129
rect 1274 47 1328 95
rect 1358 169 1422 177
rect 1358 135 1378 169
rect 1412 135 1422 169
rect 1358 47 1422 135
rect 1452 89 1516 177
rect 1452 55 1472 89
rect 1506 55 1516 89
rect 1452 47 1516 55
rect 1546 169 1610 177
rect 1546 135 1566 169
rect 1600 135 1610 169
rect 1546 47 1610 135
rect 1640 161 1702 177
rect 1640 127 1660 161
rect 1694 127 1702 161
rect 1640 93 1702 127
rect 1640 59 1660 93
rect 1694 59 1702 93
rect 1640 47 1702 59
<< pdiff >>
rect 27 489 85 497
rect 27 455 39 489
rect 73 455 85 489
rect 27 421 85 455
rect 27 387 39 421
rect 73 387 85 421
rect 27 353 85 387
rect 27 319 39 353
rect 73 319 85 353
rect 27 297 85 319
rect 121 485 179 497
rect 121 451 133 485
rect 167 451 179 485
rect 121 297 179 451
rect 215 489 273 497
rect 215 455 227 489
rect 261 455 273 489
rect 215 421 273 455
rect 215 387 227 421
rect 261 387 273 421
rect 215 353 273 387
rect 215 319 227 353
rect 261 319 273 353
rect 215 297 273 319
rect 309 485 367 497
rect 309 451 321 485
rect 355 451 367 485
rect 309 297 367 451
rect 403 489 461 497
rect 403 455 415 489
rect 449 455 461 489
rect 403 421 461 455
rect 403 387 415 421
rect 449 387 461 421
rect 403 353 461 387
rect 403 319 415 353
rect 449 319 461 353
rect 403 297 461 319
rect 497 369 555 497
rect 497 335 509 369
rect 543 335 555 369
rect 497 297 555 335
rect 591 489 649 497
rect 591 455 603 489
rect 637 455 649 489
rect 591 421 649 455
rect 591 387 603 421
rect 637 387 649 421
rect 591 297 649 387
rect 685 369 743 497
rect 685 335 697 369
rect 731 335 743 369
rect 685 297 743 335
rect 779 489 837 497
rect 779 455 791 489
rect 825 455 837 489
rect 779 297 837 455
rect 895 339 954 497
rect 895 305 908 339
rect 942 305 954 339
rect 895 297 954 305
rect 990 475 1048 497
rect 990 441 1002 475
rect 1036 441 1048 475
rect 990 407 1048 441
rect 990 373 1002 407
rect 1036 373 1048 407
rect 990 297 1048 373
rect 1084 339 1142 497
rect 1084 305 1096 339
rect 1130 305 1142 339
rect 1084 297 1142 305
rect 1178 475 1236 497
rect 1178 441 1190 475
rect 1224 441 1236 475
rect 1178 407 1236 441
rect 1178 373 1190 407
rect 1224 373 1236 407
rect 1178 297 1236 373
rect 1272 475 1330 497
rect 1272 441 1284 475
rect 1318 441 1330 475
rect 1272 407 1330 441
rect 1272 373 1284 407
rect 1318 373 1330 407
rect 1272 339 1330 373
rect 1272 305 1284 339
rect 1318 305 1330 339
rect 1272 297 1330 305
rect 1366 489 1424 497
rect 1366 455 1378 489
rect 1412 455 1424 489
rect 1366 421 1424 455
rect 1366 387 1378 421
rect 1412 387 1424 421
rect 1366 297 1424 387
rect 1460 475 1518 497
rect 1460 441 1472 475
rect 1506 441 1518 475
rect 1460 407 1518 441
rect 1460 373 1472 407
rect 1506 373 1518 407
rect 1460 339 1518 373
rect 1460 305 1472 339
rect 1506 305 1518 339
rect 1460 297 1518 305
rect 1554 489 1612 497
rect 1554 455 1566 489
rect 1600 455 1612 489
rect 1554 421 1612 455
rect 1554 387 1566 421
rect 1600 387 1612 421
rect 1554 297 1612 387
rect 1648 423 1702 497
rect 1648 389 1660 423
rect 1694 389 1702 423
rect 1648 355 1702 389
rect 1648 321 1660 355
rect 1694 321 1702 355
rect 1648 297 1702 321
<< ndiffc >>
rect 39 127 73 161
rect 39 59 73 93
rect 133 59 167 93
rect 227 123 261 157
rect 227 55 261 89
rect 321 59 355 93
rect 415 123 449 157
rect 415 55 449 89
rect 509 59 543 93
rect 603 123 637 157
rect 603 55 637 89
rect 697 59 731 93
rect 791 123 825 157
rect 791 55 825 89
rect 900 55 934 89
rect 968 55 1002 89
rect 1072 95 1106 129
rect 1178 55 1212 89
rect 1284 95 1318 129
rect 1378 135 1412 169
rect 1472 55 1506 89
rect 1566 135 1600 169
rect 1660 127 1694 161
rect 1660 59 1694 93
<< pdiffc >>
rect 39 455 73 489
rect 39 387 73 421
rect 39 319 73 353
rect 133 451 167 485
rect 227 455 261 489
rect 227 387 261 421
rect 227 319 261 353
rect 321 451 355 485
rect 415 455 449 489
rect 415 387 449 421
rect 415 319 449 353
rect 509 335 543 369
rect 603 455 637 489
rect 603 387 637 421
rect 697 335 731 369
rect 791 455 825 489
rect 908 305 942 339
rect 1002 441 1036 475
rect 1002 373 1036 407
rect 1096 305 1130 339
rect 1190 441 1224 475
rect 1190 373 1224 407
rect 1284 441 1318 475
rect 1284 373 1318 407
rect 1284 305 1318 339
rect 1378 455 1412 489
rect 1378 387 1412 421
rect 1472 441 1506 475
rect 1472 373 1506 407
rect 1472 305 1506 339
rect 1566 455 1600 489
rect 1566 387 1600 421
rect 1660 389 1694 423
rect 1660 321 1694 355
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 273 497 309 523
rect 367 497 403 523
rect 461 497 497 523
rect 555 497 591 523
rect 649 497 685 523
rect 743 497 779 523
rect 954 497 990 523
rect 1048 497 1084 523
rect 1142 497 1178 523
rect 1236 497 1272 523
rect 1330 497 1366 523
rect 1424 497 1460 523
rect 1518 497 1554 523
rect 1612 497 1648 523
rect 85 282 121 297
rect 179 282 215 297
rect 273 282 309 297
rect 367 282 403 297
rect 461 282 497 297
rect 555 282 591 297
rect 649 282 685 297
rect 743 282 779 297
rect 954 282 990 297
rect 1048 282 1084 297
rect 1142 282 1178 297
rect 1236 282 1272 297
rect 1330 282 1366 297
rect 1424 282 1460 297
rect 1518 282 1554 297
rect 1612 282 1648 297
rect 83 259 123 282
rect 177 259 217 282
rect 271 259 311 282
rect 365 259 405 282
rect 83 249 405 259
rect 83 215 102 249
rect 136 215 180 249
rect 214 215 258 249
rect 292 215 336 249
rect 370 215 405 249
rect 83 205 405 215
rect 83 177 113 205
rect 177 177 207 205
rect 271 177 301 205
rect 375 177 405 205
rect 459 259 499 282
rect 553 259 593 282
rect 647 259 687 282
rect 741 259 781 282
rect 952 259 992 282
rect 1046 259 1086 282
rect 1140 259 1180 282
rect 1234 259 1274 282
rect 459 249 781 259
rect 459 215 475 249
rect 509 215 553 249
rect 587 215 631 249
rect 665 215 709 249
rect 743 215 781 249
rect 459 205 781 215
rect 459 177 489 205
rect 553 177 583 205
rect 647 177 677 205
rect 751 177 781 205
rect 835 249 1274 259
rect 835 215 851 249
rect 885 215 929 249
rect 963 215 1007 249
rect 1041 215 1085 249
rect 1119 215 1163 249
rect 1197 215 1274 249
rect 835 205 1274 215
rect 835 177 865 205
rect 1022 177 1052 205
rect 1116 177 1146 205
rect 1244 177 1274 205
rect 1328 259 1368 282
rect 1422 259 1462 282
rect 1516 259 1556 282
rect 1610 259 1650 282
rect 1328 249 1665 259
rect 1328 215 1449 249
rect 1483 215 1527 249
rect 1561 215 1605 249
rect 1639 215 1665 249
rect 1328 205 1665 215
rect 1328 177 1358 205
rect 1422 177 1452 205
rect 1516 177 1546 205
rect 1610 177 1640 205
rect 83 21 113 47
rect 177 21 207 47
rect 271 21 301 47
rect 375 21 405 47
rect 459 21 489 47
rect 553 21 583 47
rect 647 21 677 47
rect 751 21 781 47
rect 835 21 865 47
rect 1022 21 1052 47
rect 1116 21 1146 47
rect 1244 21 1274 47
rect 1328 21 1358 47
rect 1422 21 1452 47
rect 1516 21 1546 47
rect 1610 21 1640 47
<< polycont >>
rect 102 215 136 249
rect 180 215 214 249
rect 258 215 292 249
rect 336 215 370 249
rect 475 215 509 249
rect 553 215 587 249
rect 631 215 665 249
rect 709 215 743 249
rect 851 215 885 249
rect 929 215 963 249
rect 1007 215 1041 249
rect 1085 215 1119 249
rect 1163 215 1197 249
rect 1449 215 1483 249
rect 1527 215 1561 249
rect 1605 215 1639 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 18 489 89 493
rect 18 455 39 489
rect 73 455 89 489
rect 18 421 89 455
rect 18 387 39 421
rect 73 387 89 421
rect 133 485 167 527
rect 133 413 167 451
rect 201 489 277 493
rect 201 455 227 489
rect 261 455 277 489
rect 201 421 277 455
rect 18 379 89 387
rect 201 387 227 421
rect 261 387 277 421
rect 321 485 355 527
rect 321 413 355 451
rect 389 489 857 493
rect 389 455 415 489
rect 449 455 603 489
rect 637 455 791 489
rect 825 455 857 489
rect 389 441 857 455
rect 906 475 1240 493
rect 906 441 1002 475
rect 1036 441 1190 475
rect 1224 441 1240 475
rect 389 421 465 441
rect 201 379 277 387
rect 389 387 415 421
rect 449 387 465 421
rect 577 421 653 441
rect 389 379 465 387
rect 18 353 465 379
rect 18 319 39 353
rect 73 319 227 353
rect 261 319 415 353
rect 449 319 465 353
rect 509 369 543 407
rect 577 387 603 421
rect 637 387 653 421
rect 906 407 1240 441
rect 697 373 1002 407
rect 1036 373 1190 407
rect 1224 373 1240 407
rect 1284 475 1318 493
rect 1284 407 1318 441
rect 1352 489 1428 527
rect 1352 455 1378 489
rect 1412 455 1428 489
rect 1352 421 1428 455
rect 1352 387 1378 421
rect 1412 387 1428 421
rect 1352 378 1428 387
rect 1472 475 1506 493
rect 1472 407 1506 441
rect 697 369 801 373
rect 543 335 697 353
rect 731 335 801 369
rect 1284 339 1318 373
rect 1540 489 1616 527
rect 1540 455 1566 489
rect 1600 455 1616 489
rect 1540 421 1616 455
rect 1540 387 1566 421
rect 1600 387 1616 421
rect 1540 378 1616 387
rect 1660 423 1725 493
rect 1694 389 1725 423
rect 1472 339 1506 373
rect 1660 355 1725 389
rect 509 319 801 335
rect 835 305 908 339
rect 942 305 1096 339
rect 1130 305 1284 339
rect 1318 305 1472 339
rect 1506 321 1660 339
rect 1694 321 1725 355
rect 1506 305 1725 321
rect 835 289 1725 305
rect 18 249 386 285
rect 18 215 102 249
rect 136 215 180 249
rect 214 215 258 249
rect 292 215 336 249
rect 370 215 386 249
rect 18 211 386 215
rect 430 249 801 285
rect 430 215 475 249
rect 509 215 553 249
rect 587 215 631 249
rect 665 215 709 249
rect 743 215 801 249
rect 430 211 801 215
rect 835 249 1318 255
rect 835 215 851 249
rect 885 215 929 249
rect 963 215 1007 249
rect 1041 215 1085 249
rect 1119 215 1163 249
rect 1197 215 1318 249
rect 835 211 1318 215
rect 1352 177 1399 289
rect 1433 249 1717 255
rect 1433 215 1449 249
rect 1483 215 1527 249
rect 1561 215 1605 249
rect 1639 215 1717 249
rect 1433 211 1717 215
rect 18 161 1318 177
rect 18 127 39 161
rect 73 157 1318 161
rect 73 143 227 157
rect 73 127 89 143
rect 18 93 89 127
rect 201 123 227 143
rect 261 143 415 157
rect 261 123 277 143
rect 18 59 39 93
rect 73 59 89 93
rect 18 51 89 59
rect 133 93 167 109
rect 133 17 167 59
rect 201 89 277 123
rect 389 123 415 143
rect 449 143 603 157
rect 449 123 465 143
rect 201 55 227 89
rect 261 55 277 89
rect 201 51 277 55
rect 321 93 355 109
rect 321 17 355 59
rect 389 89 465 123
rect 577 123 603 143
rect 637 143 791 157
rect 637 123 653 143
rect 389 55 415 89
rect 449 55 465 89
rect 389 51 465 55
rect 509 93 543 109
rect 509 17 543 59
rect 577 89 653 123
rect 765 123 791 143
rect 825 143 1318 157
rect 825 123 841 143
rect 577 55 603 89
rect 637 55 653 89
rect 577 51 653 55
rect 697 93 731 109
rect 697 17 731 59
rect 765 89 841 123
rect 1072 129 1106 143
rect 765 55 791 89
rect 825 55 841 89
rect 765 51 841 55
rect 889 89 1028 109
rect 889 55 900 89
rect 934 55 968 89
rect 1002 55 1028 89
rect 1284 129 1318 143
rect 1352 169 1616 177
rect 1352 135 1378 169
rect 1412 135 1566 169
rect 1600 135 1616 169
rect 1352 129 1616 135
rect 1660 161 1717 177
rect 1072 79 1106 95
rect 1158 89 1232 109
rect 889 17 1028 55
rect 1158 55 1178 89
rect 1212 55 1232 89
rect 1158 17 1232 55
rect 1694 127 1717 161
rect 1660 95 1717 127
rect 1284 93 1717 95
rect 1284 89 1660 93
rect 1284 55 1472 89
rect 1506 59 1660 89
rect 1694 59 1717 93
rect 1506 55 1717 59
rect 1284 51 1717 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel locali s 1049 221 1083 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 947 221 981 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 856 221 890 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1253 221 1287 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 744 221 778 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 642 221 676 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 540 221 574 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 438 221 472 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 336 221 370 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 234 221 268 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 132 221 166 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 853 289 887 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 947 289 981 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1047 289 1081 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1161 289 1195 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1362 289 1396 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1467 289 1501 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1569 289 1603 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1671 425 1705 459 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1671 357 1705 391 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1467 221 1501 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1569 221 1603 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1671 289 1705 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1671 221 1705 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1161 221 1195 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1258 289 1292 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 o31ai_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1748 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 621458
string GDS_START 606458
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
