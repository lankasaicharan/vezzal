magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 8 49 850 243
rect 0 0 864 49
<< scnmos >>
rect 155 49 185 217
rect 345 49 375 217
rect 431 49 461 217
rect 547 49 577 217
rect 633 49 663 217
rect 741 49 771 217
<< scpmoshvt >>
rect 192 367 222 619
rect 306 367 336 619
rect 417 367 447 619
rect 543 367 573 619
rect 633 367 663 619
rect 741 367 771 619
<< ndiff >>
rect 34 205 155 217
rect 34 171 42 205
rect 76 171 155 205
rect 34 169 155 171
rect 34 135 110 169
rect 144 135 155 169
rect 34 101 155 135
rect 34 97 110 101
rect 34 63 42 97
rect 76 67 110 97
rect 144 67 155 101
rect 76 63 155 67
rect 34 49 155 63
rect 185 163 238 217
rect 185 129 196 163
rect 230 129 238 163
rect 185 95 238 129
rect 185 61 196 95
rect 230 61 238 95
rect 185 49 238 61
rect 292 205 345 217
rect 292 171 300 205
rect 334 171 345 205
rect 292 101 345 171
rect 292 67 300 101
rect 334 67 345 101
rect 292 49 345 67
rect 375 205 431 217
rect 375 171 386 205
rect 420 171 431 205
rect 375 101 431 171
rect 375 67 386 101
rect 420 67 431 101
rect 375 49 431 67
rect 461 167 547 217
rect 461 133 486 167
rect 520 133 547 167
rect 461 91 547 133
rect 461 57 486 91
rect 520 57 547 91
rect 461 49 547 57
rect 577 205 633 217
rect 577 171 588 205
rect 622 171 633 205
rect 577 101 633 171
rect 577 67 588 101
rect 622 67 633 101
rect 577 49 633 67
rect 663 167 741 217
rect 663 133 688 167
rect 722 133 741 167
rect 663 91 741 133
rect 663 57 688 91
rect 722 57 741 91
rect 663 49 741 57
rect 771 205 824 217
rect 771 171 782 205
rect 816 171 824 205
rect 771 101 824 171
rect 771 67 782 101
rect 816 67 824 101
rect 771 49 824 67
<< pdiff >>
rect 71 599 192 619
rect 71 565 79 599
rect 113 565 147 599
rect 181 565 192 599
rect 71 511 192 565
rect 71 477 79 511
rect 113 477 147 511
rect 181 477 192 511
rect 71 413 192 477
rect 71 379 79 413
rect 113 379 147 413
rect 181 379 192 413
rect 71 367 192 379
rect 222 607 306 619
rect 222 573 247 607
rect 281 573 306 607
rect 222 495 306 573
rect 222 461 247 495
rect 281 461 306 495
rect 222 367 306 461
rect 336 599 417 619
rect 336 565 347 599
rect 381 565 417 599
rect 336 521 417 565
rect 336 487 347 521
rect 381 487 417 521
rect 336 435 417 487
rect 336 401 347 435
rect 381 401 417 435
rect 336 367 417 401
rect 447 367 543 619
rect 573 367 633 619
rect 663 367 741 619
rect 771 607 824 619
rect 771 573 782 607
rect 816 573 824 607
rect 771 518 824 573
rect 771 484 782 518
rect 816 484 824 518
rect 771 434 824 484
rect 771 400 782 434
rect 816 400 824 434
rect 771 367 824 400
<< ndiffc >>
rect 42 171 76 205
rect 110 135 144 169
rect 42 63 76 97
rect 110 67 144 101
rect 196 129 230 163
rect 196 61 230 95
rect 300 171 334 205
rect 300 67 334 101
rect 386 171 420 205
rect 386 67 420 101
rect 486 133 520 167
rect 486 57 520 91
rect 588 171 622 205
rect 588 67 622 101
rect 688 133 722 167
rect 688 57 722 91
rect 782 171 816 205
rect 782 67 816 101
<< pdiffc >>
rect 79 565 113 599
rect 147 565 181 599
rect 79 477 113 511
rect 147 477 181 511
rect 79 379 113 413
rect 147 379 181 413
rect 247 573 281 607
rect 247 461 281 495
rect 347 565 381 599
rect 347 487 381 521
rect 347 401 381 435
rect 782 573 816 607
rect 782 484 816 518
rect 782 400 816 434
<< poly >>
rect 192 619 222 645
rect 306 619 336 645
rect 417 619 447 645
rect 543 619 573 645
rect 633 619 663 645
rect 741 619 771 645
rect 192 305 222 367
rect 155 289 222 305
rect 155 255 172 289
rect 206 255 222 289
rect 306 335 336 367
rect 417 335 447 367
rect 543 335 573 367
rect 633 335 663 367
rect 306 319 375 335
rect 306 285 325 319
rect 359 285 375 319
rect 306 269 375 285
rect 417 319 483 335
rect 417 285 433 319
rect 467 285 483 319
rect 417 269 483 285
rect 525 319 591 335
rect 525 285 541 319
rect 575 285 591 319
rect 525 269 591 285
rect 633 319 699 335
rect 633 285 649 319
rect 683 285 699 319
rect 633 269 699 285
rect 741 325 771 367
rect 741 309 839 325
rect 741 275 789 309
rect 823 275 839 309
rect 155 239 222 255
rect 155 217 185 239
rect 345 217 375 269
rect 431 217 461 269
rect 547 217 577 269
rect 633 217 663 269
rect 741 259 839 275
rect 741 217 771 259
rect 155 23 185 49
rect 345 23 375 49
rect 431 23 461 49
rect 547 23 577 49
rect 633 23 663 49
rect 741 23 771 49
<< polycont >>
rect 172 255 206 289
rect 325 285 359 319
rect 433 285 467 319
rect 541 285 575 319
rect 649 285 683 319
rect 789 275 823 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 17 599 185 615
rect 17 565 79 599
rect 113 565 147 599
rect 181 565 185 599
rect 17 511 185 565
rect 17 477 79 511
rect 113 477 147 511
rect 181 477 185 511
rect 17 413 185 477
rect 231 607 297 649
rect 231 573 247 607
rect 281 573 297 607
rect 231 495 297 573
rect 231 461 247 495
rect 281 461 297 495
rect 231 454 297 461
rect 331 599 381 615
rect 331 565 347 599
rect 773 607 832 649
rect 331 521 381 565
rect 331 487 347 521
rect 331 435 381 487
rect 331 420 347 435
rect 17 379 79 413
rect 113 379 147 413
rect 181 379 185 413
rect 17 363 185 379
rect 251 401 347 420
rect 251 385 381 401
rect 17 285 115 363
rect 251 305 285 385
rect 156 289 285 305
rect 17 205 99 285
rect 156 255 172 289
rect 206 255 285 289
rect 319 319 381 350
rect 319 285 325 319
rect 359 285 381 319
rect 319 269 381 285
rect 415 319 467 596
rect 415 285 433 319
rect 415 269 467 285
rect 501 319 591 596
rect 655 335 739 596
rect 773 573 782 607
rect 816 573 832 607
rect 773 518 832 573
rect 773 484 782 518
rect 816 484 832 518
rect 773 434 832 484
rect 773 400 782 434
rect 816 400 832 434
rect 773 384 832 400
rect 501 285 541 319
rect 575 285 591 319
rect 633 319 739 335
rect 633 285 649 319
rect 683 285 739 319
rect 773 309 847 350
rect 501 269 591 285
rect 773 275 789 309
rect 823 275 847 309
rect 156 233 285 255
rect 156 219 342 233
rect 17 171 42 205
rect 76 185 99 205
rect 180 205 342 219
rect 180 199 300 205
rect 76 171 146 185
rect 17 169 146 171
rect 17 135 110 169
rect 144 135 146 169
rect 284 171 300 199
rect 334 171 342 205
rect 17 101 146 135
rect 17 97 110 101
rect 17 63 42 97
rect 76 67 110 97
rect 144 67 146 101
rect 76 63 146 67
rect 17 51 146 63
rect 180 129 196 163
rect 230 129 246 163
rect 180 95 246 129
rect 180 61 196 95
rect 230 61 246 95
rect 180 17 246 61
rect 284 101 342 171
rect 284 67 300 101
rect 334 67 342 101
rect 284 51 342 67
rect 376 205 832 235
rect 376 171 386 205
rect 420 201 588 205
rect 420 171 430 201
rect 376 101 430 171
rect 572 171 588 201
rect 622 201 782 205
rect 622 171 638 201
rect 376 67 386 101
rect 420 67 430 101
rect 376 51 430 67
rect 470 133 486 167
rect 520 133 536 167
rect 470 91 536 133
rect 470 57 486 91
rect 520 57 536 91
rect 470 17 536 57
rect 572 101 638 171
rect 772 171 782 201
rect 816 171 832 205
rect 572 67 588 101
rect 622 67 638 101
rect 572 51 638 67
rect 672 133 688 167
rect 722 133 738 167
rect 672 91 738 133
rect 672 57 688 91
rect 722 57 738 91
rect 672 17 738 57
rect 772 101 832 171
rect 772 67 782 101
rect 816 67 832 101
rect 772 51 832 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o41a_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 492572
string GDS_START 483194
<< end >>
