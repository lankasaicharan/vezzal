magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
rect 420 303 656 331
<< pwell >>
rect 57 49 807 157
rect 0 0 864 49
<< scnmos >>
rect 140 47 170 131
rect 218 47 248 131
rect 304 47 334 131
rect 376 47 406 131
rect 464 47 494 131
rect 536 47 566 131
rect 622 47 652 131
rect 694 47 724 131
<< scpmoshvt >>
rect 84 409 134 609
rect 190 409 240 609
rect 296 409 346 609
rect 513 339 563 539
rect 731 409 781 609
<< ndiff >>
rect 83 101 140 131
rect 83 67 95 101
rect 129 67 140 101
rect 83 47 140 67
rect 170 47 218 131
rect 248 111 304 131
rect 248 77 259 111
rect 293 77 304 111
rect 248 47 304 77
rect 334 47 376 131
rect 406 106 464 131
rect 406 72 417 106
rect 451 72 464 106
rect 406 47 464 72
rect 494 47 536 131
rect 566 103 622 131
rect 566 69 577 103
rect 611 69 622 103
rect 566 47 622 69
rect 652 47 694 131
rect 724 106 781 131
rect 724 72 735 106
rect 769 72 781 106
rect 724 47 781 72
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 190 609
rect 134 563 145 597
rect 179 563 190 597
rect 134 517 190 563
rect 134 483 145 517
rect 179 483 190 517
rect 134 409 190 483
rect 240 597 296 609
rect 240 563 251 597
rect 285 563 296 597
rect 240 526 296 563
rect 240 492 251 526
rect 285 492 296 526
rect 240 455 296 492
rect 240 421 251 455
rect 285 421 296 455
rect 240 409 296 421
rect 346 597 402 609
rect 346 563 357 597
rect 391 563 402 597
rect 674 597 731 609
rect 346 526 402 563
rect 674 563 686 597
rect 720 563 731 597
rect 346 492 357 526
rect 391 492 402 526
rect 346 455 402 492
rect 346 421 357 455
rect 391 421 402 455
rect 346 409 402 421
rect 456 527 513 539
rect 456 493 468 527
rect 502 493 513 527
rect 456 456 513 493
rect 456 422 468 456
rect 502 422 513 456
rect 456 385 513 422
rect 456 351 468 385
rect 502 351 513 385
rect 456 339 513 351
rect 563 527 620 539
rect 563 493 574 527
rect 608 493 620 527
rect 563 456 620 493
rect 563 422 574 456
rect 608 422 620 456
rect 563 385 620 422
rect 674 526 731 563
rect 674 492 686 526
rect 720 492 731 526
rect 674 455 731 492
rect 674 421 686 455
rect 720 421 731 455
rect 674 409 731 421
rect 781 597 837 609
rect 781 563 792 597
rect 826 563 837 597
rect 781 526 837 563
rect 781 492 792 526
rect 826 492 837 526
rect 781 455 837 492
rect 781 421 792 455
rect 826 421 837 455
rect 781 409 837 421
rect 563 351 574 385
rect 608 351 620 385
rect 563 339 620 351
<< ndiffc >>
rect 95 67 129 101
rect 259 77 293 111
rect 417 72 451 106
rect 577 69 611 103
rect 735 72 769 106
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 483 179 517
rect 251 563 285 597
rect 251 492 285 526
rect 251 421 285 455
rect 357 563 391 597
rect 686 563 720 597
rect 357 492 391 526
rect 357 421 391 455
rect 468 493 502 527
rect 468 422 502 456
rect 468 351 502 385
rect 574 493 608 527
rect 574 422 608 456
rect 686 492 720 526
rect 686 421 720 455
rect 792 563 826 597
rect 792 492 826 526
rect 792 421 826 455
rect 574 351 608 385
<< poly >>
rect 84 609 134 635
rect 190 609 240 635
rect 296 609 346 635
rect 731 609 781 635
rect 513 539 563 565
rect 84 228 134 409
rect 190 356 240 409
rect 182 340 248 356
rect 182 306 198 340
rect 232 306 248 340
rect 182 290 248 306
rect 68 212 134 228
rect 68 178 84 212
rect 118 192 134 212
rect 118 178 170 192
rect 68 162 170 178
rect 140 131 170 162
rect 218 131 248 290
rect 296 339 346 409
rect 731 356 781 409
rect 694 340 761 356
rect 296 255 326 339
rect 369 275 435 291
rect 369 255 385 275
rect 296 241 385 255
rect 419 241 435 275
rect 296 225 435 241
rect 296 176 326 225
rect 513 221 563 339
rect 694 306 711 340
rect 745 306 761 340
rect 694 272 761 306
rect 694 252 711 272
rect 622 238 711 252
rect 745 238 761 272
rect 622 222 761 238
rect 503 205 569 221
rect 503 177 519 205
rect 296 146 406 176
rect 304 131 334 146
rect 376 131 406 146
rect 464 171 519 177
rect 553 171 569 205
rect 464 147 569 171
rect 464 131 494 147
rect 536 131 566 147
rect 622 131 652 222
rect 694 131 724 222
rect 140 21 170 47
rect 218 21 248 47
rect 304 21 334 47
rect 376 21 406 47
rect 464 21 494 47
rect 536 21 566 47
rect 622 21 652 47
rect 694 21 724 47
<< polycont >>
rect 198 306 232 340
rect 84 178 118 212
rect 385 241 419 275
rect 711 306 745 340
rect 711 238 745 272
rect 519 171 553 205
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 526 89 563
rect 23 492 39 526
rect 73 492 89 526
rect 23 455 89 492
rect 129 597 195 649
rect 129 563 145 597
rect 179 563 195 597
rect 129 517 195 563
rect 129 483 145 517
rect 179 483 195 517
rect 129 467 195 483
rect 235 597 301 613
rect 235 563 251 597
rect 285 563 301 597
rect 235 526 301 563
rect 235 492 251 526
rect 285 492 301 526
rect 23 421 39 455
rect 73 431 89 455
rect 235 455 301 492
rect 235 431 251 455
rect 73 421 251 431
rect 285 421 301 455
rect 23 397 301 421
rect 341 597 407 613
rect 341 563 357 597
rect 391 563 407 597
rect 341 526 407 563
rect 341 492 357 526
rect 391 492 407 526
rect 341 455 407 492
rect 341 421 357 455
rect 391 421 407 455
rect 341 361 407 421
rect 25 340 263 356
rect 25 306 198 340
rect 232 306 263 340
rect 25 290 263 306
rect 299 327 407 361
rect 452 597 736 613
rect 452 579 686 597
rect 452 527 518 579
rect 670 563 686 579
rect 720 563 736 597
rect 452 493 468 527
rect 502 493 518 527
rect 452 456 518 493
rect 452 422 468 456
rect 502 422 518 456
rect 452 385 518 422
rect 452 351 468 385
rect 502 351 518 385
rect 452 335 518 351
rect 558 527 624 543
rect 558 493 574 527
rect 608 493 624 527
rect 558 456 624 493
rect 558 422 574 456
rect 608 422 624 456
rect 558 385 624 422
rect 670 526 736 563
rect 670 492 686 526
rect 720 492 736 526
rect 670 455 736 492
rect 670 421 686 455
rect 720 421 736 455
rect 670 405 736 421
rect 776 597 842 649
rect 776 563 792 597
rect 826 563 842 597
rect 776 526 842 563
rect 776 492 792 526
rect 826 492 842 526
rect 776 455 842 492
rect 776 421 792 455
rect 826 421 842 455
rect 776 405 842 421
rect 558 351 574 385
rect 608 351 624 385
rect 25 212 167 228
rect 25 178 84 212
rect 118 178 167 212
rect 25 162 167 178
rect 299 135 333 327
rect 558 291 624 351
rect 695 340 839 356
rect 695 306 711 340
rect 745 306 839 340
rect 369 275 639 291
rect 369 241 385 275
rect 419 257 639 275
rect 419 241 435 257
rect 369 225 435 241
rect 503 205 569 221
rect 503 171 519 205
rect 553 171 569 205
rect 503 155 569 171
rect 79 101 145 126
rect 79 67 95 101
rect 129 67 145 101
rect 79 17 145 67
rect 217 111 359 135
rect 217 77 259 111
rect 293 77 359 111
rect 217 53 359 77
rect 401 106 467 135
rect 605 119 639 257
rect 695 272 839 306
rect 695 238 711 272
rect 745 238 839 272
rect 695 222 839 238
rect 401 72 417 106
rect 451 72 467 106
rect 401 17 467 72
rect 561 103 639 119
rect 561 69 577 103
rect 611 69 639 103
rect 561 53 639 69
rect 719 106 785 135
rect 719 72 735 106
rect 769 72 785 106
rect 719 17 785 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2bb2oi_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3077816
string GDS_START 3069366
<< end >>
