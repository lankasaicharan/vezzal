magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 332 2054 704
<< pwell >>
rect 186 49 984 248
rect 1202 49 2000 248
rect 0 0 2016 49
<< scnmos >>
rect 265 74 295 222
rect 351 74 381 222
rect 437 74 467 222
rect 523 74 553 222
rect 789 74 819 222
rect 875 74 905 222
rect 1285 74 1315 222
rect 1371 74 1401 222
rect 1457 74 1487 222
rect 1543 74 1573 222
rect 1629 74 1659 222
rect 1715 74 1745 222
rect 1801 74 1831 222
rect 1887 74 1917 222
<< scpmoshvt >>
rect 84 368 114 592
rect 174 368 204 592
rect 264 368 294 592
rect 354 368 384 592
rect 444 368 474 592
rect 534 368 564 592
rect 624 368 654 592
rect 714 368 744 592
rect 912 368 942 592
rect 1002 368 1032 592
rect 1092 368 1122 592
rect 1182 368 1212 592
rect 1272 368 1302 592
rect 1362 368 1392 592
rect 1452 368 1482 592
rect 1542 368 1572 592
rect 1632 368 1662 592
rect 1722 368 1752 592
rect 1812 368 1842 592
rect 1902 368 1932 592
<< ndiff >>
rect 212 127 265 222
rect 212 93 220 127
rect 254 93 265 127
rect 212 74 265 93
rect 295 202 351 222
rect 295 168 306 202
rect 340 168 351 202
rect 295 116 351 168
rect 295 82 306 116
rect 340 82 351 116
rect 295 74 351 82
rect 381 127 437 222
rect 381 93 392 127
rect 426 93 437 127
rect 381 74 437 93
rect 467 210 523 222
rect 467 176 478 210
rect 512 176 523 210
rect 467 120 523 176
rect 467 86 478 120
rect 512 86 523 120
rect 467 74 523 86
rect 553 152 789 222
rect 553 118 564 152
rect 598 118 654 152
rect 688 118 744 152
rect 778 118 789 152
rect 553 74 789 118
rect 819 210 875 222
rect 819 176 830 210
rect 864 176 875 210
rect 819 120 875 176
rect 819 86 830 120
rect 864 86 875 120
rect 819 74 875 86
rect 905 145 958 222
rect 905 111 916 145
rect 950 111 958 145
rect 905 74 958 111
rect 1228 120 1285 222
rect 1228 86 1240 120
rect 1274 86 1285 120
rect 1228 74 1285 86
rect 1315 207 1371 222
rect 1315 173 1326 207
rect 1360 173 1371 207
rect 1315 74 1371 173
rect 1401 120 1457 222
rect 1401 86 1412 120
rect 1446 86 1457 120
rect 1401 74 1457 86
rect 1487 207 1543 222
rect 1487 173 1498 207
rect 1532 173 1543 207
rect 1487 74 1543 173
rect 1573 210 1629 222
rect 1573 176 1584 210
rect 1618 176 1629 210
rect 1573 120 1629 176
rect 1573 86 1584 120
rect 1618 86 1629 120
rect 1573 74 1629 86
rect 1659 152 1715 222
rect 1659 118 1670 152
rect 1704 118 1715 152
rect 1659 74 1715 118
rect 1745 210 1801 222
rect 1745 176 1756 210
rect 1790 176 1801 210
rect 1745 120 1801 176
rect 1745 86 1756 120
rect 1790 86 1801 120
rect 1745 74 1801 86
rect 1831 152 1887 222
rect 1831 118 1842 152
rect 1876 118 1887 152
rect 1831 74 1887 118
rect 1917 210 1974 222
rect 1917 176 1928 210
rect 1962 176 1974 210
rect 1917 120 1974 176
rect 1917 86 1928 120
rect 1962 86 1974 120
rect 1917 74 1974 86
<< pdiff >>
rect 29 580 84 592
rect 29 546 37 580
rect 71 546 84 580
rect 29 462 84 546
rect 29 428 37 462
rect 71 428 84 462
rect 29 368 84 428
rect 114 531 174 592
rect 114 497 127 531
rect 161 497 174 531
rect 114 414 174 497
rect 114 380 127 414
rect 161 380 174 414
rect 114 368 174 380
rect 204 580 264 592
rect 204 546 217 580
rect 251 546 264 580
rect 204 462 264 546
rect 204 428 217 462
rect 251 428 264 462
rect 204 368 264 428
rect 294 531 354 592
rect 294 497 307 531
rect 341 497 354 531
rect 294 414 354 497
rect 294 380 307 414
rect 341 380 354 414
rect 294 368 354 380
rect 384 580 444 592
rect 384 546 397 580
rect 431 546 444 580
rect 384 510 444 546
rect 384 476 397 510
rect 431 476 444 510
rect 384 424 444 476
rect 384 390 397 424
rect 431 390 444 424
rect 384 368 444 390
rect 474 584 534 592
rect 474 550 487 584
rect 521 550 534 584
rect 474 508 534 550
rect 474 474 487 508
rect 521 474 534 508
rect 474 368 534 474
rect 564 531 624 592
rect 564 497 577 531
rect 611 497 624 531
rect 564 424 624 497
rect 564 390 577 424
rect 611 390 624 424
rect 564 368 624 390
rect 654 584 714 592
rect 654 550 667 584
rect 701 550 714 584
rect 654 501 714 550
rect 654 467 667 501
rect 701 467 714 501
rect 654 368 714 467
rect 744 531 799 592
rect 744 497 757 531
rect 791 497 799 531
rect 744 427 799 497
rect 744 393 757 427
rect 791 393 799 427
rect 744 368 799 393
rect 853 531 912 592
rect 853 497 865 531
rect 899 497 912 531
rect 853 424 912 497
rect 853 390 865 424
rect 899 390 912 424
rect 853 368 912 390
rect 942 584 1002 592
rect 942 550 955 584
rect 989 550 1002 584
rect 942 498 1002 550
rect 942 464 955 498
rect 989 464 1002 498
rect 942 368 1002 464
rect 1032 531 1092 592
rect 1032 497 1045 531
rect 1079 497 1092 531
rect 1032 424 1092 497
rect 1032 390 1045 424
rect 1079 390 1092 424
rect 1032 368 1092 390
rect 1122 584 1182 592
rect 1122 550 1135 584
rect 1169 550 1182 584
rect 1122 498 1182 550
rect 1122 464 1135 498
rect 1169 464 1182 498
rect 1122 368 1182 464
rect 1212 580 1272 592
rect 1212 546 1225 580
rect 1259 546 1272 580
rect 1212 503 1272 546
rect 1212 469 1225 503
rect 1259 469 1272 503
rect 1212 424 1272 469
rect 1212 390 1225 424
rect 1259 390 1272 424
rect 1212 368 1272 390
rect 1302 580 1362 592
rect 1302 546 1315 580
rect 1349 546 1362 580
rect 1302 492 1362 546
rect 1302 458 1315 492
rect 1349 458 1362 492
rect 1302 368 1362 458
rect 1392 580 1452 592
rect 1392 546 1405 580
rect 1439 546 1452 580
rect 1392 503 1452 546
rect 1392 469 1405 503
rect 1439 469 1452 503
rect 1392 424 1452 469
rect 1392 390 1405 424
rect 1439 390 1452 424
rect 1392 368 1452 390
rect 1482 580 1542 592
rect 1482 546 1495 580
rect 1529 546 1542 580
rect 1482 492 1542 546
rect 1482 458 1495 492
rect 1529 458 1542 492
rect 1482 368 1542 458
rect 1572 580 1632 592
rect 1572 546 1585 580
rect 1619 546 1632 580
rect 1572 503 1632 546
rect 1572 469 1585 503
rect 1619 469 1632 503
rect 1572 424 1632 469
rect 1572 390 1585 424
rect 1619 390 1632 424
rect 1572 368 1632 390
rect 1662 580 1722 592
rect 1662 546 1675 580
rect 1709 546 1722 580
rect 1662 508 1722 546
rect 1662 474 1675 508
rect 1709 474 1722 508
rect 1662 368 1722 474
rect 1752 580 1812 592
rect 1752 546 1765 580
rect 1799 546 1812 580
rect 1752 503 1812 546
rect 1752 469 1765 503
rect 1799 469 1812 503
rect 1752 424 1812 469
rect 1752 390 1765 424
rect 1799 390 1812 424
rect 1752 368 1812 390
rect 1842 580 1902 592
rect 1842 546 1855 580
rect 1889 546 1902 580
rect 1842 508 1902 546
rect 1842 474 1855 508
rect 1889 474 1902 508
rect 1842 368 1902 474
rect 1932 580 1987 592
rect 1932 546 1945 580
rect 1979 546 1987 580
rect 1932 497 1987 546
rect 1932 463 1945 497
rect 1979 463 1987 497
rect 1932 414 1987 463
rect 1932 380 1945 414
rect 1979 380 1987 414
rect 1932 368 1987 380
<< ndiffc >>
rect 220 93 254 127
rect 306 168 340 202
rect 306 82 340 116
rect 392 93 426 127
rect 478 176 512 210
rect 478 86 512 120
rect 564 118 598 152
rect 654 118 688 152
rect 744 118 778 152
rect 830 176 864 210
rect 830 86 864 120
rect 916 111 950 145
rect 1240 86 1274 120
rect 1326 173 1360 207
rect 1412 86 1446 120
rect 1498 173 1532 207
rect 1584 176 1618 210
rect 1584 86 1618 120
rect 1670 118 1704 152
rect 1756 176 1790 210
rect 1756 86 1790 120
rect 1842 118 1876 152
rect 1928 176 1962 210
rect 1928 86 1962 120
<< pdiffc >>
rect 37 546 71 580
rect 37 428 71 462
rect 127 497 161 531
rect 127 380 161 414
rect 217 546 251 580
rect 217 428 251 462
rect 307 497 341 531
rect 307 380 341 414
rect 397 546 431 580
rect 397 476 431 510
rect 397 390 431 424
rect 487 550 521 584
rect 487 474 521 508
rect 577 497 611 531
rect 577 390 611 424
rect 667 550 701 584
rect 667 467 701 501
rect 757 497 791 531
rect 757 393 791 427
rect 865 497 899 531
rect 865 390 899 424
rect 955 550 989 584
rect 955 464 989 498
rect 1045 497 1079 531
rect 1045 390 1079 424
rect 1135 550 1169 584
rect 1135 464 1169 498
rect 1225 546 1259 580
rect 1225 469 1259 503
rect 1225 390 1259 424
rect 1315 546 1349 580
rect 1315 458 1349 492
rect 1405 546 1439 580
rect 1405 469 1439 503
rect 1405 390 1439 424
rect 1495 546 1529 580
rect 1495 458 1529 492
rect 1585 546 1619 580
rect 1585 469 1619 503
rect 1585 390 1619 424
rect 1675 546 1709 580
rect 1675 474 1709 508
rect 1765 546 1799 580
rect 1765 469 1799 503
rect 1765 390 1799 424
rect 1855 546 1889 580
rect 1855 474 1889 508
rect 1945 546 1979 580
rect 1945 463 1979 497
rect 1945 380 1979 414
<< poly >>
rect 84 592 114 618
rect 174 592 204 618
rect 264 592 294 618
rect 354 592 384 618
rect 444 592 474 618
rect 534 592 564 618
rect 624 592 654 618
rect 714 592 744 618
rect 912 592 942 618
rect 1002 592 1032 618
rect 1092 592 1122 618
rect 1182 592 1212 618
rect 1272 592 1302 618
rect 1362 592 1392 618
rect 1452 592 1482 618
rect 1542 592 1572 618
rect 1632 592 1662 618
rect 1722 592 1752 618
rect 1812 592 1842 618
rect 1902 592 1932 618
rect 84 353 114 368
rect 174 353 204 368
rect 264 353 294 368
rect 354 353 384 368
rect 444 353 474 368
rect 534 353 564 368
rect 624 353 654 368
rect 714 353 744 368
rect 912 353 942 368
rect 1002 353 1032 368
rect 1092 353 1122 368
rect 1182 353 1212 368
rect 1272 353 1302 368
rect 1362 353 1392 368
rect 1452 353 1482 368
rect 1542 353 1572 368
rect 1632 353 1662 368
rect 1722 353 1752 368
rect 1812 353 1842 368
rect 1902 353 1932 368
rect 81 310 117 353
rect 171 310 207 353
rect 261 310 297 353
rect 351 310 387 353
rect 444 336 477 353
rect 531 336 567 353
rect 621 342 657 353
rect 711 342 747 353
rect 621 336 747 342
rect 909 336 945 353
rect 999 336 1035 353
rect 1089 336 1125 353
rect 1179 336 1215 353
rect 81 294 387 310
rect 447 320 747 336
rect 447 294 463 320
rect 81 260 127 294
rect 161 260 195 294
rect 229 260 263 294
rect 297 260 331 294
rect 365 280 387 294
rect 437 286 463 294
rect 497 286 531 320
rect 565 286 599 320
rect 633 286 667 320
rect 701 286 747 320
rect 814 320 1215 336
rect 814 300 871 320
rect 365 260 381 280
rect 81 244 381 260
rect 265 222 295 244
rect 351 222 381 244
rect 437 264 747 286
rect 789 286 871 300
rect 905 286 939 320
rect 973 286 1013 320
rect 1047 286 1090 320
rect 1124 286 1165 320
rect 1199 286 1215 320
rect 789 270 1215 286
rect 1269 336 1305 353
rect 1359 336 1395 353
rect 1449 336 1485 353
rect 1539 336 1575 353
rect 1269 320 1575 336
rect 1269 286 1321 320
rect 1355 286 1389 320
rect 1423 286 1457 320
rect 1491 286 1525 320
rect 1559 286 1575 320
rect 1269 270 1575 286
rect 1629 336 1665 353
rect 1719 336 1755 353
rect 1809 336 1845 353
rect 1899 336 1935 353
rect 1629 320 1935 336
rect 1629 286 1657 320
rect 1691 286 1725 320
rect 1759 286 1793 320
rect 1827 286 1861 320
rect 1895 286 1935 320
rect 1629 270 1935 286
rect 437 222 467 264
rect 523 222 553 264
rect 789 222 819 270
rect 875 222 905 270
rect 1285 222 1315 270
rect 1371 222 1401 270
rect 1457 222 1487 270
rect 1543 222 1573 270
rect 1629 222 1659 270
rect 1715 222 1745 270
rect 1801 222 1831 270
rect 1887 222 1917 270
rect 265 48 295 74
rect 351 48 381 74
rect 437 48 467 74
rect 523 48 553 74
rect 789 48 819 74
rect 875 48 905 74
rect 1285 48 1315 74
rect 1371 48 1401 74
rect 1457 48 1487 74
rect 1543 48 1573 74
rect 1629 48 1659 74
rect 1715 48 1745 74
rect 1801 48 1831 74
rect 1887 48 1917 74
<< polycont >>
rect 127 260 161 294
rect 195 260 229 294
rect 263 260 297 294
rect 331 260 365 294
rect 463 286 497 320
rect 531 286 565 320
rect 599 286 633 320
rect 667 286 701 320
rect 871 286 905 320
rect 939 286 973 320
rect 1013 286 1047 320
rect 1090 286 1124 320
rect 1165 286 1199 320
rect 1321 286 1355 320
rect 1389 286 1423 320
rect 1457 286 1491 320
rect 1525 286 1559 320
rect 1657 286 1691 320
rect 1725 286 1759 320
rect 1793 286 1827 320
rect 1861 286 1895 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 21 581 447 615
rect 21 580 71 581
rect 21 546 37 580
rect 217 580 251 581
rect 21 462 71 546
rect 21 428 37 462
rect 21 412 71 428
rect 111 531 177 547
rect 111 497 127 531
rect 161 497 177 531
rect 111 414 177 497
rect 111 380 127 414
rect 161 380 177 414
rect 381 580 447 581
rect 217 462 251 546
rect 217 412 251 428
rect 291 531 341 547
rect 291 497 307 531
rect 291 414 341 497
rect 111 378 177 380
rect 291 380 307 414
rect 381 546 397 580
rect 431 546 447 580
rect 381 510 447 546
rect 381 476 397 510
rect 431 476 447 510
rect 381 424 447 476
rect 487 584 1185 615
rect 521 581 667 584
rect 521 550 537 581
rect 487 508 537 550
rect 651 550 667 581
rect 701 581 955 584
rect 701 550 717 581
rect 521 474 537 508
rect 487 458 537 474
rect 571 531 617 547
rect 571 497 577 531
rect 611 497 617 531
rect 571 424 617 497
rect 651 501 717 550
rect 939 550 955 581
rect 989 581 1135 584
rect 989 550 1005 581
rect 651 467 667 501
rect 701 467 717 501
rect 651 458 717 467
rect 751 531 807 547
rect 751 497 757 531
rect 791 497 807 531
rect 751 427 807 497
rect 751 424 757 427
rect 381 390 397 424
rect 431 390 577 424
rect 611 393 757 424
rect 791 393 807 427
rect 611 390 807 393
rect 849 531 905 547
rect 849 497 865 531
rect 899 497 905 531
rect 849 424 905 497
rect 939 498 1005 550
rect 1119 550 1135 581
rect 1169 550 1185 584
rect 939 464 955 498
rect 989 464 1005 498
rect 939 458 1005 464
rect 1039 531 1085 547
rect 1039 497 1045 531
rect 1079 497 1085 531
rect 1039 424 1085 497
rect 1119 498 1185 550
rect 1119 464 1135 498
rect 1169 464 1185 498
rect 1119 458 1185 464
rect 1225 580 1259 596
rect 1225 503 1259 546
rect 1225 424 1259 469
rect 1299 580 1365 649
rect 1299 546 1315 580
rect 1349 546 1365 580
rect 1299 492 1365 546
rect 1299 458 1315 492
rect 1349 458 1365 492
rect 1405 580 1439 596
rect 1405 503 1439 546
rect 1405 424 1439 469
rect 1479 580 1545 649
rect 1479 546 1495 580
rect 1529 546 1545 580
rect 1479 492 1545 546
rect 1479 458 1495 492
rect 1529 458 1545 492
rect 1585 580 1619 596
rect 1585 503 1619 546
rect 1585 424 1619 469
rect 1659 580 1709 649
rect 1659 546 1675 580
rect 1659 508 1709 546
rect 1659 474 1675 508
rect 1659 458 1709 474
rect 1749 580 1815 596
rect 1749 546 1765 580
rect 1799 546 1815 580
rect 1749 503 1815 546
rect 1749 469 1765 503
rect 1799 469 1815 503
rect 1749 424 1815 469
rect 1855 580 1905 649
rect 1889 546 1905 580
rect 1855 508 1905 546
rect 1889 474 1905 508
rect 1855 458 1905 474
rect 1945 580 1995 596
rect 1979 546 1995 580
rect 1945 497 1995 546
rect 1979 463 1995 497
rect 1945 424 1995 463
rect 849 390 865 424
rect 899 390 1045 424
rect 1079 390 1225 424
rect 1259 390 1405 424
rect 1439 390 1585 424
rect 1619 390 1765 424
rect 1799 414 1995 424
rect 1799 390 1945 414
rect 291 378 341 380
rect 25 344 341 378
rect 741 364 807 390
rect 1979 380 1995 414
rect 1945 364 1995 380
rect 25 202 71 344
rect 447 320 702 356
rect 111 294 381 310
rect 111 260 127 294
rect 161 260 195 294
rect 229 260 263 294
rect 297 260 331 294
rect 365 260 381 294
rect 447 286 463 320
rect 497 286 531 320
rect 565 286 599 320
rect 633 286 667 320
rect 701 286 702 320
rect 447 270 702 286
rect 855 320 1215 356
rect 855 286 871 320
rect 905 286 939 320
rect 973 286 1013 320
rect 1047 286 1090 320
rect 1124 286 1165 320
rect 1199 286 1215 320
rect 855 270 1215 286
rect 1290 320 1607 356
rect 1290 286 1321 320
rect 1355 286 1389 320
rect 1423 286 1457 320
rect 1491 286 1525 320
rect 1559 286 1607 320
rect 1290 270 1607 286
rect 1641 320 1911 356
rect 1641 286 1657 320
rect 1691 286 1725 320
rect 1759 286 1793 320
rect 1827 286 1861 320
rect 1895 286 1911 320
rect 1641 270 1911 286
rect 111 236 381 260
rect 478 226 1376 236
rect 478 210 1548 226
rect 25 168 306 202
rect 340 176 478 202
rect 512 202 830 210
rect 512 176 528 202
rect 340 168 528 176
rect 814 176 830 202
rect 864 207 1548 210
rect 864 195 1326 207
rect 204 127 270 134
rect 204 93 220 127
rect 254 93 270 127
rect 204 17 270 93
rect 306 116 340 168
rect 306 66 340 82
rect 376 127 442 134
rect 376 93 392 127
rect 426 93 442 127
rect 376 17 442 93
rect 478 120 528 168
rect 512 86 528 120
rect 478 70 528 86
rect 562 152 780 168
rect 562 118 564 152
rect 598 118 654 152
rect 688 118 744 152
rect 778 118 780 152
rect 562 17 780 118
rect 814 120 864 176
rect 1310 173 1326 195
rect 1360 183 1498 207
rect 1360 173 1376 183
rect 814 86 830 120
rect 814 70 864 86
rect 900 145 966 161
rect 1310 154 1376 173
rect 1482 173 1498 183
rect 1532 173 1548 207
rect 1482 154 1548 173
rect 1584 210 1978 236
rect 1618 202 1756 210
rect 900 111 916 145
rect 950 111 966 145
rect 900 17 966 111
rect 1224 120 1276 136
rect 1408 120 1450 136
rect 1584 120 1618 176
rect 1790 202 1928 210
rect 1224 86 1240 120
rect 1274 86 1412 120
rect 1446 86 1584 120
rect 1224 70 1618 86
rect 1654 152 1720 168
rect 1654 118 1670 152
rect 1704 118 1720 152
rect 1654 17 1720 118
rect 1756 120 1790 176
rect 1962 176 1978 210
rect 1756 70 1790 86
rect 1826 152 1892 168
rect 1826 118 1842 152
rect 1876 118 1892 152
rect 1826 17 1892 118
rect 1928 120 1978 176
rect 1962 86 1978 120
rect 1928 70 1978 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a2111oi_4
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 2699382
string GDS_START 2683270
<< end >>
