magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 1 49 821 167
rect 0 0 864 49
<< scnmos >>
rect 84 57 114 141
rect 162 57 192 141
rect 361 57 391 141
rect 439 57 469 141
rect 517 57 547 141
rect 636 57 666 141
rect 708 57 738 141
<< scpmoshvt >>
rect 87 408 137 608
rect 305 409 355 609
rect 411 409 461 609
rect 517 409 567 609
rect 644 409 694 609
<< ndiff >>
rect 27 116 84 141
rect 27 82 39 116
rect 73 82 84 116
rect 27 57 84 82
rect 114 57 162 141
rect 192 116 249 141
rect 192 82 203 116
rect 237 82 249 116
rect 192 57 249 82
rect 304 116 361 141
rect 304 82 316 116
rect 350 82 361 116
rect 304 57 361 82
rect 391 57 439 141
rect 469 57 517 141
rect 547 107 636 141
rect 547 73 558 107
rect 592 73 636 107
rect 547 57 636 73
rect 666 57 708 141
rect 738 116 795 141
rect 738 82 749 116
rect 783 82 795 116
rect 738 57 795 82
<< pdiff >>
rect 30 596 87 608
rect 30 562 42 596
rect 76 562 87 596
rect 30 525 87 562
rect 30 491 42 525
rect 76 491 87 525
rect 30 454 87 491
rect 30 420 42 454
rect 76 420 87 454
rect 30 408 87 420
rect 137 596 194 608
rect 137 562 148 596
rect 182 562 194 596
rect 137 525 194 562
rect 137 491 148 525
rect 182 491 194 525
rect 137 454 194 491
rect 137 420 148 454
rect 182 420 194 454
rect 137 408 194 420
rect 248 597 305 609
rect 248 563 260 597
rect 294 563 305 597
rect 248 526 305 563
rect 248 492 260 526
rect 294 492 305 526
rect 248 455 305 492
rect 248 421 260 455
rect 294 421 305 455
rect 248 409 305 421
rect 355 597 411 609
rect 355 563 366 597
rect 400 563 411 597
rect 355 524 411 563
rect 355 490 366 524
rect 400 490 411 524
rect 355 409 411 490
rect 461 597 517 609
rect 461 563 472 597
rect 506 563 517 597
rect 461 526 517 563
rect 461 492 472 526
rect 506 492 517 526
rect 461 455 517 492
rect 461 421 472 455
rect 506 421 517 455
rect 461 409 517 421
rect 567 597 644 609
rect 567 563 578 597
rect 612 563 644 597
rect 567 524 644 563
rect 567 490 578 524
rect 612 490 644 524
rect 567 409 644 490
rect 694 597 751 609
rect 694 563 705 597
rect 739 563 751 597
rect 694 526 751 563
rect 694 492 705 526
rect 739 492 751 526
rect 694 455 751 492
rect 694 421 705 455
rect 739 421 751 455
rect 694 409 751 421
<< ndiffc >>
rect 39 82 73 116
rect 203 82 237 116
rect 316 82 350 116
rect 558 73 592 107
rect 749 82 783 116
<< pdiffc >>
rect 42 562 76 596
rect 42 491 76 525
rect 42 420 76 454
rect 148 562 182 596
rect 148 491 182 525
rect 148 420 182 454
rect 260 563 294 597
rect 260 492 294 526
rect 260 421 294 455
rect 366 563 400 597
rect 366 490 400 524
rect 472 563 506 597
rect 472 492 506 526
rect 472 421 506 455
rect 578 563 612 597
rect 578 490 612 524
rect 705 563 739 597
rect 705 492 739 526
rect 705 421 739 455
<< poly >>
rect 87 608 137 634
rect 305 609 355 635
rect 411 609 461 635
rect 517 609 567 635
rect 644 609 694 635
rect 87 315 137 408
rect 305 368 355 409
rect 411 368 461 409
rect 517 368 567 409
rect 25 299 137 315
rect 25 265 41 299
rect 75 285 137 299
rect 211 352 355 368
rect 211 318 227 352
rect 261 318 355 352
rect 75 265 117 285
rect 25 231 117 265
rect 211 284 355 318
rect 211 250 227 284
rect 261 250 355 284
rect 211 234 355 250
rect 403 352 469 368
rect 403 318 419 352
rect 453 318 469 352
rect 403 284 469 318
rect 403 250 419 284
rect 453 250 469 284
rect 403 234 469 250
rect 25 197 41 231
rect 75 197 117 231
rect 25 186 117 197
rect 325 186 355 234
rect 25 156 192 186
rect 325 156 391 186
rect 84 141 114 156
rect 162 141 192 156
rect 361 141 391 156
rect 439 141 469 234
rect 517 352 583 368
rect 517 318 533 352
rect 567 318 583 352
rect 517 284 583 318
rect 644 298 694 409
rect 517 250 533 284
rect 567 250 583 284
rect 517 234 583 250
rect 631 282 738 298
rect 631 248 647 282
rect 681 248 738 282
rect 517 141 547 234
rect 631 214 738 248
rect 631 180 647 214
rect 681 180 738 214
rect 631 164 738 180
rect 636 141 666 164
rect 708 141 738 164
rect 84 31 114 57
rect 162 31 192 57
rect 361 31 391 57
rect 439 31 469 57
rect 517 31 547 57
rect 636 31 666 57
rect 708 31 738 57
<< polycont >>
rect 41 265 75 299
rect 227 318 261 352
rect 227 250 261 284
rect 419 318 453 352
rect 419 250 453 284
rect 41 197 75 231
rect 533 318 567 352
rect 533 250 567 284
rect 647 248 681 282
rect 647 180 681 214
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 26 596 92 649
rect 26 562 42 596
rect 76 562 92 596
rect 26 525 92 562
rect 26 491 42 525
rect 76 491 92 525
rect 26 454 92 491
rect 26 420 42 454
rect 76 420 92 454
rect 26 404 92 420
rect 132 596 198 612
rect 132 562 148 596
rect 182 562 198 596
rect 132 525 198 562
rect 132 491 148 525
rect 182 491 198 525
rect 132 454 198 491
rect 132 420 148 454
rect 182 420 198 454
rect 132 404 198 420
rect 244 597 310 613
rect 244 563 260 597
rect 294 563 310 597
rect 244 526 310 563
rect 244 492 260 526
rect 294 492 310 526
rect 244 455 310 492
rect 350 597 416 649
rect 350 563 366 597
rect 400 563 416 597
rect 350 524 416 563
rect 350 490 366 524
rect 400 490 416 524
rect 350 474 416 490
rect 456 597 522 613
rect 456 563 472 597
rect 506 563 522 597
rect 456 526 522 563
rect 456 492 472 526
rect 506 492 522 526
rect 244 421 260 455
rect 294 438 310 455
rect 456 455 522 492
rect 562 597 628 649
rect 562 563 578 597
rect 612 563 628 597
rect 562 524 628 563
rect 562 490 578 524
rect 612 490 628 524
rect 562 474 628 490
rect 689 597 839 613
rect 689 563 705 597
rect 739 563 839 597
rect 689 526 839 563
rect 689 492 705 526
rect 739 492 839 526
rect 456 438 472 455
rect 294 421 472 438
rect 506 438 522 455
rect 689 455 839 492
rect 506 421 653 438
rect 244 404 653 421
rect 689 421 705 455
rect 739 421 839 455
rect 689 405 839 421
rect 164 368 198 404
rect 25 299 91 356
rect 25 265 41 299
rect 75 265 91 299
rect 25 231 91 265
rect 25 197 41 231
rect 75 197 91 231
rect 25 181 91 197
rect 164 352 277 368
rect 164 318 227 352
rect 261 318 277 352
rect 164 284 277 318
rect 164 250 227 284
rect 261 250 277 284
rect 164 234 277 250
rect 313 352 469 368
rect 313 318 419 352
rect 453 318 469 352
rect 313 284 469 318
rect 313 250 419 284
rect 453 250 469 284
rect 313 234 469 250
rect 505 352 583 368
rect 505 318 533 352
rect 567 318 583 352
rect 505 284 583 318
rect 505 250 533 284
rect 567 250 583 284
rect 505 234 583 250
rect 619 298 653 404
rect 619 282 697 298
rect 619 248 647 282
rect 681 248 697 282
rect 23 116 89 145
rect 23 82 39 116
rect 73 82 89 116
rect 23 17 89 82
rect 164 116 253 234
rect 619 214 697 248
rect 619 198 647 214
rect 164 82 203 116
rect 237 82 253 116
rect 164 53 253 82
rect 300 180 647 198
rect 681 180 697 214
rect 300 164 697 180
rect 733 236 839 405
rect 300 116 366 164
rect 300 82 316 116
rect 350 82 366 116
rect 300 53 366 82
rect 542 107 608 128
rect 542 73 558 107
rect 592 73 608 107
rect 542 17 608 73
rect 733 116 799 236
rect 733 82 749 116
rect 783 82 799 116
rect 733 53 799 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and3b_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6373036
string GDS_START 6364868
<< end >>
