magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 1 157 275 208
rect 1 49 663 157
rect 0 0 672 49
<< scnmos >>
rect 80 98 110 182
rect 166 98 196 182
rect 367 47 397 131
rect 469 47 499 131
rect 547 47 577 131
<< scpmoshvt >>
rect 80 529 110 613
rect 166 529 196 613
rect 389 439 419 523
rect 475 439 505 523
rect 561 439 591 523
<< ndiff >>
rect 27 144 80 182
rect 27 110 35 144
rect 69 110 80 144
rect 27 98 80 110
rect 110 144 166 182
rect 110 110 121 144
rect 155 110 166 144
rect 110 98 166 110
rect 196 153 249 182
rect 196 119 207 153
rect 241 119 249 153
rect 196 98 249 119
rect 314 93 367 131
rect 314 59 322 93
rect 356 59 367 93
rect 314 47 367 59
rect 397 95 469 131
rect 397 61 424 95
rect 458 61 469 95
rect 397 47 469 61
rect 499 47 547 131
rect 577 93 637 131
rect 577 59 595 93
rect 629 59 637 93
rect 577 47 637 59
<< pdiff >>
rect 27 587 80 613
rect 27 553 35 587
rect 69 553 80 587
rect 27 529 80 553
rect 110 601 166 613
rect 110 567 121 601
rect 155 567 166 601
rect 110 529 166 567
rect 196 589 249 613
rect 196 555 207 589
rect 241 555 249 589
rect 196 529 249 555
rect 336 485 389 523
rect 336 451 344 485
rect 378 451 389 485
rect 336 439 389 451
rect 419 485 475 523
rect 419 451 430 485
rect 464 451 475 485
rect 419 439 475 451
rect 505 515 561 523
rect 505 481 516 515
rect 550 481 561 515
rect 505 439 561 481
rect 591 485 644 523
rect 591 451 602 485
rect 636 451 644 485
rect 591 439 644 451
<< ndiffc >>
rect 35 110 69 144
rect 121 110 155 144
rect 207 119 241 153
rect 322 59 356 93
rect 424 61 458 95
rect 595 59 629 93
<< pdiffc >>
rect 35 553 69 587
rect 121 567 155 601
rect 207 555 241 589
rect 344 451 378 485
rect 430 451 464 485
rect 516 481 550 515
rect 602 451 636 485
<< poly >>
rect 80 613 110 639
rect 166 613 196 639
rect 281 605 347 621
rect 281 571 297 605
rect 331 571 347 605
rect 281 555 347 571
rect 80 429 110 529
rect 166 507 196 529
rect 166 477 237 507
rect 80 413 151 429
rect 80 379 101 413
rect 135 379 151 413
rect 80 345 151 379
rect 80 311 101 345
rect 135 311 151 345
rect 80 295 151 311
rect 207 339 237 477
rect 291 417 321 555
rect 389 523 419 549
rect 475 523 505 549
rect 561 523 591 549
rect 389 417 419 439
rect 291 387 419 417
rect 207 323 273 339
rect 80 182 110 295
rect 207 289 223 323
rect 257 289 273 323
rect 207 255 273 289
rect 207 235 223 255
rect 166 221 223 235
rect 257 221 273 255
rect 166 205 273 221
rect 325 287 355 387
rect 475 287 505 439
rect 325 271 397 287
rect 325 237 341 271
rect 375 237 397 271
rect 166 182 196 205
rect 325 203 397 237
rect 325 169 341 203
rect 375 169 397 203
rect 325 153 397 169
rect 439 271 505 287
rect 439 237 455 271
rect 489 237 505 271
rect 439 203 505 237
rect 439 169 455 203
rect 489 169 505 203
rect 561 302 591 439
rect 561 286 645 302
rect 561 252 595 286
rect 629 252 645 286
rect 561 218 645 252
rect 561 198 595 218
rect 439 153 505 169
rect 547 184 595 198
rect 629 184 645 218
rect 547 168 645 184
rect 367 131 397 153
rect 469 131 499 153
rect 547 131 577 168
rect 80 72 110 98
rect 166 72 196 98
rect 367 21 397 47
rect 469 21 499 47
rect 547 21 577 47
<< polycont >>
rect 297 571 331 605
rect 101 379 135 413
rect 101 311 135 345
rect 223 289 257 323
rect 223 221 257 255
rect 341 237 375 271
rect 341 169 375 203
rect 455 237 489 271
rect 455 169 489 203
rect 595 252 629 286
rect 595 184 629 218
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 31 587 73 603
rect 31 553 35 587
rect 69 553 73 587
rect 31 537 73 553
rect 117 601 159 649
rect 117 567 121 601
rect 155 567 159 601
rect 117 551 159 567
rect 203 589 297 605
rect 203 555 207 589
rect 241 571 297 589
rect 331 571 347 605
rect 241 555 347 571
rect 203 539 347 555
rect 31 160 65 537
rect 512 515 554 649
rect 101 485 382 501
rect 101 467 344 485
rect 101 413 135 467
rect 340 451 344 467
rect 378 451 382 485
rect 101 345 135 379
rect 101 295 135 311
rect 223 323 257 424
rect 340 359 382 451
rect 426 485 468 501
rect 426 451 430 485
rect 464 451 468 485
rect 512 481 516 515
rect 550 481 554 515
rect 512 465 554 481
rect 598 485 640 501
rect 426 429 468 451
rect 598 451 602 485
rect 636 451 640 485
rect 598 429 640 451
rect 426 395 640 429
rect 340 325 559 359
rect 223 255 257 289
rect 223 205 257 221
rect 341 271 375 287
rect 341 203 375 237
rect 31 144 73 160
rect 31 110 35 144
rect 69 110 73 144
rect 31 94 73 110
rect 117 144 159 160
rect 117 110 121 144
rect 155 110 159 144
rect 117 17 159 110
rect 203 153 375 169
rect 415 271 489 287
rect 415 237 455 271
rect 415 203 489 237
rect 415 169 455 203
rect 415 153 489 169
rect 203 119 207 153
rect 241 135 375 153
rect 241 119 245 135
rect 203 103 245 119
rect 525 99 559 325
rect 595 286 641 350
rect 629 252 641 286
rect 595 218 641 252
rect 629 184 641 218
rect 595 168 641 184
rect 306 93 372 97
rect 306 59 322 93
rect 356 59 372 93
rect 306 17 372 59
rect 408 95 559 99
rect 408 61 424 95
rect 458 61 559 95
rect 408 57 559 61
rect 595 93 633 109
rect 629 59 633 93
rect 595 17 633 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21bo_m
flabel comment s 337 306 337 306 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3752326
string GDS_START 3744600
<< end >>
