magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 178 420 229
rect 1 49 765 178
rect 0 0 768 49
<< scnmos >>
rect 84 119 114 203
rect 156 119 186 203
rect 242 119 272 203
rect 314 119 344 203
rect 416 68 446 152
rect 494 68 524 152
rect 580 68 610 152
rect 652 68 682 152
<< scpmoshvt >>
rect 109 419 159 619
rect 215 419 265 619
rect 321 419 371 619
rect 540 412 590 612
rect 632 412 682 612
<< ndiff >>
rect 27 178 84 203
rect 27 144 39 178
rect 73 144 84 178
rect 27 119 84 144
rect 114 119 156 203
rect 186 178 242 203
rect 186 144 197 178
rect 231 144 242 178
rect 186 119 242 144
rect 272 119 314 203
rect 344 152 394 203
rect 344 127 416 152
rect 344 119 371 127
rect 359 93 371 119
rect 405 93 416 127
rect 359 68 416 93
rect 446 68 494 152
rect 524 127 580 152
rect 524 93 535 127
rect 569 93 580 127
rect 524 68 580 93
rect 610 68 652 152
rect 682 114 739 152
rect 682 80 693 114
rect 727 80 739 114
rect 682 68 739 80
<< pdiff >>
rect 49 597 109 619
rect 49 563 61 597
rect 95 563 109 597
rect 49 465 109 563
rect 49 431 61 465
rect 95 431 109 465
rect 49 419 109 431
rect 159 597 215 619
rect 159 563 170 597
rect 204 563 215 597
rect 159 528 215 563
rect 159 494 170 528
rect 204 494 215 528
rect 159 419 215 494
rect 265 602 321 619
rect 265 568 276 602
rect 310 568 321 602
rect 265 419 321 568
rect 371 597 428 619
rect 371 563 382 597
rect 416 563 428 597
rect 371 528 428 563
rect 371 494 382 528
rect 416 494 428 528
rect 371 419 428 494
rect 483 597 540 612
rect 483 563 495 597
rect 529 563 540 597
rect 483 527 540 563
rect 483 493 495 527
rect 529 493 540 527
rect 483 458 540 493
rect 483 424 495 458
rect 529 424 540 458
rect 483 412 540 424
rect 590 412 632 612
rect 682 600 739 612
rect 682 566 693 600
rect 727 566 739 600
rect 682 528 739 566
rect 682 494 693 528
rect 727 494 739 528
rect 682 412 739 494
<< ndiffc >>
rect 39 144 73 178
rect 197 144 231 178
rect 371 93 405 127
rect 535 93 569 127
rect 693 80 727 114
<< pdiffc >>
rect 61 563 95 597
rect 61 431 95 465
rect 170 563 204 597
rect 170 494 204 528
rect 276 568 310 602
rect 382 563 416 597
rect 382 494 416 528
rect 495 563 529 597
rect 495 493 529 527
rect 495 424 529 458
rect 693 566 727 600
rect 693 494 727 528
<< poly >>
rect 109 619 159 645
rect 215 619 265 645
rect 321 619 371 645
rect 540 612 590 638
rect 632 612 682 638
rect 109 379 159 419
rect 215 391 265 419
rect 84 363 173 379
rect 84 329 123 363
rect 157 343 173 363
rect 157 329 186 343
rect 84 313 186 329
rect 84 203 114 313
rect 156 203 186 313
rect 235 325 265 391
rect 321 397 371 419
rect 540 397 590 412
rect 321 367 590 397
rect 235 309 380 325
rect 235 295 330 309
rect 314 275 330 295
rect 364 275 380 309
rect 314 259 380 275
rect 458 302 488 367
rect 632 302 682 412
rect 458 286 524 302
rect 242 203 272 229
rect 314 203 344 259
rect 458 252 474 286
rect 508 252 524 286
rect 458 197 524 252
rect 416 167 524 197
rect 416 152 446 167
rect 494 152 524 167
rect 580 286 682 302
rect 580 252 603 286
rect 637 252 682 286
rect 580 236 682 252
rect 580 152 610 236
rect 652 152 682 236
rect 84 93 114 119
rect 156 93 186 119
rect 242 51 272 119
rect 314 93 344 119
rect 416 51 446 68
rect 242 21 446 51
rect 494 42 524 68
rect 580 42 610 68
rect 652 42 682 68
<< polycont >>
rect 123 329 157 363
rect 330 275 364 309
rect 474 252 508 286
rect 603 252 637 286
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 25 597 111 613
rect 25 563 61 597
rect 95 563 111 597
rect 25 465 111 563
rect 154 597 220 613
rect 154 563 170 597
rect 204 563 220 597
rect 154 528 220 563
rect 260 602 326 649
rect 260 568 276 602
rect 310 568 326 602
rect 260 548 326 568
rect 366 597 432 613
rect 366 563 382 597
rect 416 563 432 597
rect 154 494 170 528
rect 204 512 220 528
rect 366 528 432 563
rect 366 512 382 528
rect 204 494 382 512
rect 416 494 432 528
rect 154 478 432 494
rect 479 597 545 613
rect 479 563 495 597
rect 529 563 545 597
rect 479 527 545 563
rect 479 493 495 527
rect 529 493 545 527
rect 25 431 61 465
rect 95 431 111 465
rect 479 458 545 493
rect 677 600 743 649
rect 677 566 693 600
rect 727 566 743 600
rect 677 528 743 566
rect 677 494 693 528
rect 727 494 743 528
rect 677 478 743 494
rect 479 442 495 458
rect 25 415 111 431
rect 147 424 495 442
rect 529 442 545 458
rect 529 424 723 442
rect 25 277 71 415
rect 147 408 723 424
rect 147 379 181 408
rect 107 363 181 379
rect 107 329 123 363
rect 157 329 181 363
rect 107 313 181 329
rect 217 338 653 372
rect 217 309 380 338
rect 25 243 181 277
rect 217 275 330 309
rect 364 275 380 309
rect 217 259 380 275
rect 458 286 551 302
rect 147 207 181 243
rect 458 252 474 286
rect 508 252 551 286
rect 458 236 551 252
rect 587 286 653 338
rect 587 252 603 286
rect 637 252 653 286
rect 587 236 653 252
rect 23 178 89 207
rect 23 144 39 178
rect 73 144 89 178
rect 23 17 89 144
rect 147 178 247 207
rect 689 200 723 408
rect 147 144 197 178
rect 231 144 247 178
rect 519 166 723 200
rect 147 115 247 144
rect 355 127 421 156
rect 355 93 371 127
rect 405 93 421 127
rect 355 17 421 93
rect 519 127 585 166
rect 519 93 535 127
rect 569 93 585 127
rect 519 64 585 93
rect 677 114 743 130
rect 677 80 693 114
rect 727 80 743 114
rect 677 17 743 80
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xor2_lp
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2087068
string GDS_START 2080844
<< end >>
