magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 47 49 837 250
rect 0 0 864 49
<< scnmos >>
rect 126 56 156 224
rect 212 56 242 224
rect 298 56 328 224
rect 384 56 414 224
rect 470 56 500 224
rect 556 56 586 224
rect 642 56 672 224
rect 728 56 758 224
<< scpmoshvt >>
rect 126 367 156 619
rect 212 367 242 619
rect 298 367 328 619
rect 384 367 414 619
rect 470 367 500 619
rect 556 367 586 619
rect 642 367 672 619
rect 728 367 758 619
<< ndiff >>
rect 73 208 126 224
rect 73 174 81 208
rect 115 174 126 208
rect 73 102 126 174
rect 73 68 81 102
rect 115 68 126 102
rect 73 56 126 68
rect 156 192 212 224
rect 156 158 167 192
rect 201 158 212 192
rect 156 103 212 158
rect 156 69 167 103
rect 201 69 212 103
rect 156 56 212 69
rect 242 138 298 224
rect 242 104 253 138
rect 287 104 298 138
rect 242 56 298 104
rect 328 212 384 224
rect 328 178 339 212
rect 373 178 384 212
rect 328 103 384 178
rect 328 69 339 103
rect 373 69 384 103
rect 328 56 384 69
rect 414 215 470 224
rect 414 181 425 215
rect 459 181 470 215
rect 414 102 470 181
rect 414 68 425 102
rect 459 68 470 102
rect 414 56 470 68
rect 500 212 556 224
rect 500 178 511 212
rect 545 178 556 212
rect 500 103 556 178
rect 500 69 511 103
rect 545 69 556 103
rect 500 56 556 69
rect 586 183 642 224
rect 586 149 597 183
rect 631 149 642 183
rect 586 102 642 149
rect 586 68 597 102
rect 631 68 642 102
rect 586 56 642 68
rect 672 212 728 224
rect 672 178 683 212
rect 717 178 728 212
rect 672 103 728 178
rect 672 69 683 103
rect 717 69 728 103
rect 672 56 728 69
rect 758 212 811 224
rect 758 178 769 212
rect 803 178 811 212
rect 758 102 811 178
rect 758 68 769 102
rect 803 68 811 102
rect 758 56 811 68
<< pdiff >>
rect 73 599 126 619
rect 73 565 81 599
rect 115 565 126 599
rect 73 509 126 565
rect 73 475 81 509
rect 115 475 126 509
rect 73 413 126 475
rect 73 379 81 413
rect 115 379 126 413
rect 73 367 126 379
rect 156 607 212 619
rect 156 573 167 607
rect 201 573 212 607
rect 156 528 212 573
rect 156 494 167 528
rect 201 494 212 528
rect 156 453 212 494
rect 156 419 167 453
rect 201 419 212 453
rect 156 367 212 419
rect 242 599 298 619
rect 242 565 253 599
rect 287 565 298 599
rect 242 509 298 565
rect 242 475 253 509
rect 287 475 298 509
rect 242 413 298 475
rect 242 379 253 413
rect 287 379 298 413
rect 242 367 298 379
rect 328 607 384 619
rect 328 573 339 607
rect 373 573 384 607
rect 328 524 384 573
rect 328 490 339 524
rect 373 490 384 524
rect 328 453 384 490
rect 328 419 339 453
rect 373 419 384 453
rect 328 367 384 419
rect 414 599 470 619
rect 414 565 425 599
rect 459 565 470 599
rect 414 512 470 565
rect 414 478 425 512
rect 459 478 470 512
rect 414 413 470 478
rect 414 379 425 413
rect 459 379 470 413
rect 414 367 470 379
rect 500 531 556 619
rect 500 497 511 531
rect 545 497 556 531
rect 500 440 556 497
rect 500 406 511 440
rect 545 406 556 440
rect 500 367 556 406
rect 586 599 642 619
rect 586 565 597 599
rect 631 565 642 599
rect 586 510 642 565
rect 586 476 597 510
rect 631 476 642 510
rect 586 367 642 476
rect 672 531 728 619
rect 672 497 683 531
rect 717 497 728 531
rect 672 440 728 497
rect 672 406 683 440
rect 717 406 728 440
rect 672 367 728 406
rect 758 599 811 619
rect 758 565 769 599
rect 803 565 811 599
rect 758 516 811 565
rect 758 482 769 516
rect 803 482 811 516
rect 758 436 811 482
rect 758 402 769 436
rect 803 402 811 436
rect 758 367 811 402
<< ndiffc >>
rect 81 174 115 208
rect 81 68 115 102
rect 167 158 201 192
rect 167 69 201 103
rect 253 104 287 138
rect 339 178 373 212
rect 339 69 373 103
rect 425 181 459 215
rect 425 68 459 102
rect 511 178 545 212
rect 511 69 545 103
rect 597 149 631 183
rect 597 68 631 102
rect 683 178 717 212
rect 683 69 717 103
rect 769 178 803 212
rect 769 68 803 102
<< pdiffc >>
rect 81 565 115 599
rect 81 475 115 509
rect 81 379 115 413
rect 167 573 201 607
rect 167 494 201 528
rect 167 419 201 453
rect 253 565 287 599
rect 253 475 287 509
rect 253 379 287 413
rect 339 573 373 607
rect 339 490 373 524
rect 339 419 373 453
rect 425 565 459 599
rect 425 478 459 512
rect 425 379 459 413
rect 511 497 545 531
rect 511 406 545 440
rect 597 565 631 599
rect 597 476 631 510
rect 683 497 717 531
rect 683 406 717 440
rect 769 565 803 599
rect 769 482 803 516
rect 769 402 803 436
<< poly >>
rect 126 619 156 645
rect 212 619 242 645
rect 298 619 328 645
rect 384 619 414 645
rect 470 619 500 645
rect 556 619 586 645
rect 642 619 672 645
rect 728 619 758 645
rect 126 312 156 367
rect 212 312 242 367
rect 298 312 328 367
rect 384 312 414 367
rect 119 296 414 312
rect 119 262 135 296
rect 169 262 203 296
rect 237 262 271 296
rect 305 262 414 296
rect 119 246 414 262
rect 126 224 156 246
rect 212 224 242 246
rect 298 224 328 246
rect 384 224 414 246
rect 470 335 500 367
rect 556 335 586 367
rect 642 335 672 367
rect 728 335 758 367
rect 470 319 795 335
rect 470 285 597 319
rect 631 285 665 319
rect 699 285 733 319
rect 767 285 795 319
rect 470 269 795 285
rect 470 246 586 269
rect 470 224 500 246
rect 556 224 586 246
rect 642 224 672 269
rect 728 224 758 269
rect 126 30 156 56
rect 212 30 242 56
rect 298 30 328 56
rect 384 30 414 56
rect 470 30 500 56
rect 556 30 586 56
rect 642 30 672 56
rect 728 30 758 56
<< polycont >>
rect 135 262 169 296
rect 203 262 237 296
rect 271 262 305 296
rect 597 285 631 319
rect 665 285 699 319
rect 733 285 767 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 65 599 117 615
rect 65 565 81 599
rect 115 565 117 599
rect 65 509 117 565
rect 65 475 81 509
rect 115 475 117 509
rect 65 413 117 475
rect 151 607 217 649
rect 151 573 167 607
rect 201 573 217 607
rect 151 528 217 573
rect 151 494 167 528
rect 201 494 217 528
rect 151 453 217 494
rect 151 419 167 453
rect 201 419 217 453
rect 251 599 289 615
rect 251 565 253 599
rect 287 565 289 599
rect 251 509 289 565
rect 251 475 253 509
rect 287 475 289 509
rect 65 379 81 413
rect 115 385 117 413
rect 251 413 289 475
rect 323 607 389 649
rect 323 573 339 607
rect 373 573 389 607
rect 323 524 389 573
rect 323 490 339 524
rect 373 490 389 524
rect 323 453 389 490
rect 323 419 339 453
rect 373 419 389 453
rect 423 599 819 615
rect 423 565 425 599
rect 459 581 597 599
rect 459 565 467 581
rect 423 512 467 565
rect 590 565 597 581
rect 631 581 769 599
rect 631 565 641 581
rect 423 478 425 512
rect 459 478 467 512
rect 251 385 253 413
rect 115 379 253 385
rect 287 385 289 413
rect 423 413 467 478
rect 423 385 425 413
rect 287 379 425 385
rect 459 379 467 413
rect 65 346 467 379
rect 501 531 556 547
rect 501 497 511 531
rect 545 497 556 531
rect 501 440 556 497
rect 590 510 641 565
rect 761 565 769 581
rect 803 565 819 599
rect 590 476 597 510
rect 631 476 641 510
rect 590 458 641 476
rect 675 531 727 547
rect 675 497 683 531
rect 717 497 727 531
rect 501 406 511 440
rect 545 424 556 440
rect 675 440 727 497
rect 675 424 683 440
rect 545 406 683 424
rect 717 406 727 440
rect 501 390 727 406
rect 761 516 819 565
rect 761 482 769 516
rect 803 482 819 516
rect 761 436 819 482
rect 761 402 769 436
rect 803 402 819 436
rect 501 312 547 390
rect 761 386 819 402
rect 20 296 305 312
rect 20 262 135 296
rect 169 262 203 296
rect 237 262 271 296
rect 20 242 305 262
rect 339 265 547 312
rect 581 319 833 352
rect 581 285 597 319
rect 631 285 665 319
rect 699 285 733 319
rect 767 285 833 319
rect 339 212 382 265
rect 502 251 547 265
rect 65 174 81 208
rect 115 174 131 208
rect 65 102 131 174
rect 65 68 81 102
rect 115 68 131 102
rect 65 17 131 68
rect 165 192 339 208
rect 165 158 167 192
rect 201 178 339 192
rect 373 178 382 212
rect 201 174 382 178
rect 201 158 203 174
rect 165 103 203 158
rect 165 69 167 103
rect 201 69 203 103
rect 165 53 203 69
rect 237 138 303 140
rect 237 104 253 138
rect 287 104 303 138
rect 237 17 303 104
rect 337 103 382 174
rect 337 69 339 103
rect 373 69 382 103
rect 337 53 382 69
rect 416 215 468 231
rect 416 181 425 215
rect 459 181 468 215
rect 416 102 468 181
rect 416 68 425 102
rect 459 68 468 102
rect 416 17 468 68
rect 502 217 725 251
rect 502 212 547 217
rect 502 178 511 212
rect 545 178 547 212
rect 681 212 725 217
rect 502 103 547 178
rect 502 69 511 103
rect 545 69 547 103
rect 502 53 547 69
rect 581 149 597 183
rect 631 149 647 183
rect 581 102 647 149
rect 581 68 597 102
rect 631 68 647 102
rect 581 17 647 68
rect 681 178 683 212
rect 717 178 725 212
rect 681 103 725 178
rect 681 69 683 103
rect 717 69 725 103
rect 681 53 725 69
rect 759 212 819 228
rect 759 178 769 212
rect 803 178 819 212
rect 759 102 819 178
rect 759 68 769 102
rect 803 68 819 102
rect 759 17 819 68
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor2_4
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5321850
string GDS_START 5313444
<< end >>
