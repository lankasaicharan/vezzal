magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4466 1975
<< nwell >>
rect -38 331 3206 704
rect 726 316 2370 331
rect 726 311 2011 316
<< pwell >>
rect 1101 235 1445 265
rect 1833 258 2117 265
rect 1833 235 2133 258
rect 28 176 678 235
rect 1101 176 2133 235
rect 28 167 2133 176
rect 2484 167 2903 237
rect 28 49 3167 167
rect 0 0 3168 49
<< scnmos >>
rect 111 125 141 209
rect 189 125 219 209
rect 307 125 337 209
rect 385 125 415 209
rect 493 125 523 209
rect 565 125 595 209
rect 1248 155 1278 239
rect 1336 155 1366 239
rect 759 66 789 150
rect 831 66 861 150
rect 917 66 947 150
rect 989 66 1019 150
rect 1532 125 1562 209
rect 1644 125 1674 209
rect 1716 125 1746 209
rect 1912 155 1942 239
rect 2011 155 2041 239
rect 2215 57 2245 141
rect 2301 57 2331 141
rect 2373 57 2403 141
rect 2563 127 2593 211
rect 2635 127 2665 211
rect 2721 127 2751 211
rect 2793 127 2823 211
rect 2985 57 3015 141
rect 3057 57 3087 141
<< scpmoshvt >>
rect 81 409 131 609
rect 293 417 343 617
rect 399 417 449 617
rect 493 417 543 617
rect 599 417 649 617
rect 819 347 869 547
rect 925 347 975 547
rect 1326 347 1376 547
rect 1432 347 1482 547
rect 1530 347 1580 547
rect 1704 347 1754 547
rect 1852 347 1902 547
rect 1990 352 2040 552
rect 2089 352 2139 552
rect 2227 361 2277 561
rect 2558 401 2608 601
rect 2664 401 2714 601
rect 2898 409 2948 609
<< ndiff >>
rect 54 184 111 209
rect 54 150 66 184
rect 100 150 111 184
rect 54 125 111 150
rect 141 125 189 209
rect 219 176 307 209
rect 219 142 246 176
rect 280 142 307 176
rect 219 125 307 142
rect 337 125 385 209
rect 415 181 493 209
rect 415 147 448 181
rect 482 147 493 181
rect 415 125 493 147
rect 523 125 565 209
rect 595 184 652 209
rect 595 150 606 184
rect 640 150 652 184
rect 1127 205 1248 239
rect 1127 171 1135 205
rect 1169 171 1248 205
rect 1127 155 1248 171
rect 1278 227 1336 239
rect 1278 193 1291 227
rect 1325 193 1336 227
rect 1278 155 1336 193
rect 1366 214 1419 239
rect 1366 180 1377 214
rect 1411 180 1419 214
rect 1366 155 1419 180
rect 595 125 652 150
rect 706 125 759 150
rect 706 91 714 125
rect 748 91 759 125
rect 706 66 759 91
rect 789 66 831 150
rect 861 113 917 150
rect 861 79 872 113
rect 906 79 917 113
rect 861 66 917 79
rect 947 66 989 150
rect 1019 113 1073 150
rect 1019 79 1030 113
rect 1064 79 1073 113
rect 1019 66 1073 79
rect 1479 175 1532 209
rect 1479 141 1487 175
rect 1521 141 1532 175
rect 1479 125 1532 141
rect 1562 127 1644 209
rect 1562 125 1586 127
rect 1577 93 1586 125
rect 1620 125 1644 127
rect 1674 125 1716 209
rect 1746 184 1799 209
rect 1746 150 1757 184
rect 1791 150 1799 184
rect 1746 125 1799 150
rect 1620 93 1629 125
rect 1577 81 1629 93
rect 1859 214 1912 239
rect 1859 180 1867 214
rect 1901 180 1912 214
rect 1859 155 1912 180
rect 1942 227 2011 239
rect 1942 193 1966 227
rect 2000 193 2011 227
rect 1942 155 2011 193
rect 2041 232 2091 239
rect 2041 155 2107 232
rect 2056 87 2107 155
rect 2510 186 2563 211
rect 2510 152 2518 186
rect 2552 152 2563 186
rect 2056 53 2065 87
rect 2099 53 2107 87
rect 2161 116 2215 141
rect 2161 82 2170 116
rect 2204 82 2215 116
rect 2161 57 2215 82
rect 2245 103 2301 141
rect 2245 69 2256 103
rect 2290 69 2301 103
rect 2245 57 2301 69
rect 2331 57 2373 141
rect 2403 116 2456 141
rect 2510 127 2563 152
rect 2593 127 2635 211
rect 2665 186 2721 211
rect 2665 152 2676 186
rect 2710 152 2721 186
rect 2665 127 2721 152
rect 2751 127 2793 211
rect 2823 186 2877 211
rect 2823 152 2834 186
rect 2868 152 2877 186
rect 2823 127 2877 152
rect 2403 82 2414 116
rect 2448 82 2456 116
rect 2931 116 2985 141
rect 2403 57 2456 82
rect 2931 82 2940 116
rect 2974 82 2985 116
rect 2931 57 2985 82
rect 3015 57 3057 141
rect 3087 116 3141 141
rect 3087 82 3098 116
rect 3132 82 3141 116
rect 3087 57 3141 82
rect 2056 41 2107 53
<< pdiff >>
rect 27 597 81 609
rect 27 563 36 597
rect 70 563 81 597
rect 27 526 81 563
rect 27 492 36 526
rect 70 492 81 526
rect 27 455 81 492
rect 27 421 36 455
rect 70 421 81 455
rect 27 409 81 421
rect 131 597 185 609
rect 131 563 142 597
rect 176 563 185 597
rect 131 526 185 563
rect 131 492 142 526
rect 176 492 185 526
rect 131 455 185 492
rect 131 421 142 455
rect 176 421 185 455
rect 131 409 185 421
rect 239 597 293 617
rect 239 563 248 597
rect 282 563 293 597
rect 239 463 293 563
rect 239 429 248 463
rect 282 429 293 463
rect 239 417 293 429
rect 343 464 399 617
rect 343 430 354 464
rect 388 430 399 464
rect 343 417 399 430
rect 449 417 493 617
rect 543 605 599 617
rect 543 571 554 605
rect 588 571 599 605
rect 543 417 599 571
rect 649 574 706 617
rect 649 540 660 574
rect 694 540 706 574
rect 649 417 706 540
rect 762 394 819 547
rect 762 360 774 394
rect 808 360 819 394
rect 762 347 819 360
rect 869 535 925 547
rect 869 501 880 535
rect 914 501 925 535
rect 869 347 925 501
rect 975 394 1032 547
rect 2501 589 2558 601
rect 2154 552 2227 561
rect 1917 547 1990 552
rect 975 360 986 394
rect 1020 360 1032 394
rect 975 347 1032 360
rect 1269 535 1326 547
rect 1269 501 1281 535
rect 1315 501 1326 535
rect 1269 467 1326 501
rect 1269 433 1281 467
rect 1315 433 1326 467
rect 1269 399 1326 433
rect 1269 365 1281 399
rect 1315 365 1326 399
rect 1269 347 1326 365
rect 1376 535 1432 547
rect 1376 501 1387 535
rect 1421 501 1432 535
rect 1376 464 1432 501
rect 1376 430 1387 464
rect 1421 430 1432 464
rect 1376 393 1432 430
rect 1376 359 1387 393
rect 1421 359 1432 393
rect 1376 347 1432 359
rect 1482 347 1530 547
rect 1580 535 1704 547
rect 1580 501 1591 535
rect 1625 501 1704 535
rect 1580 453 1704 501
rect 1580 419 1591 453
rect 1625 419 1704 453
rect 1580 347 1704 419
rect 1754 535 1852 547
rect 1754 501 1765 535
rect 1799 501 1852 535
rect 1754 464 1852 501
rect 1754 430 1765 464
rect 1799 430 1852 464
rect 1754 393 1852 430
rect 1754 359 1765 393
rect 1799 359 1852 393
rect 1754 347 1852 359
rect 1902 540 1990 547
rect 1902 506 1929 540
rect 1963 506 1990 540
rect 1902 466 1990 506
rect 1902 432 1929 466
rect 1963 432 1990 466
rect 1902 393 1990 432
rect 1902 359 1929 393
rect 1963 359 1990 393
rect 1902 352 1990 359
rect 2040 352 2089 552
rect 2139 549 2227 552
rect 2139 515 2166 549
rect 2200 515 2227 549
rect 2139 476 2227 515
rect 2139 442 2166 476
rect 2200 442 2227 476
rect 2139 361 2227 442
rect 2277 549 2334 561
rect 2277 515 2288 549
rect 2322 515 2334 549
rect 2277 476 2334 515
rect 2277 442 2288 476
rect 2322 442 2334 476
rect 2277 361 2334 442
rect 2501 555 2513 589
rect 2547 555 2558 589
rect 2501 518 2558 555
rect 2501 484 2513 518
rect 2547 484 2558 518
rect 2501 447 2558 484
rect 2501 413 2513 447
rect 2547 413 2558 447
rect 2501 401 2558 413
rect 2608 589 2664 601
rect 2608 555 2619 589
rect 2653 555 2664 589
rect 2608 518 2664 555
rect 2608 484 2619 518
rect 2653 484 2664 518
rect 2608 447 2664 484
rect 2608 413 2619 447
rect 2653 413 2664 447
rect 2608 401 2664 413
rect 2714 589 2771 601
rect 2714 555 2725 589
rect 2759 555 2771 589
rect 2714 518 2771 555
rect 2714 484 2725 518
rect 2759 484 2771 518
rect 2714 447 2771 484
rect 2714 413 2725 447
rect 2759 413 2771 447
rect 2714 401 2771 413
rect 2841 597 2898 609
rect 2841 563 2853 597
rect 2887 563 2898 597
rect 2841 517 2898 563
rect 2841 483 2853 517
rect 2887 483 2898 517
rect 2841 409 2898 483
rect 2948 597 3005 609
rect 2948 563 2959 597
rect 2993 563 3005 597
rect 2948 526 3005 563
rect 2948 492 2959 526
rect 2993 492 3005 526
rect 2948 455 3005 492
rect 2948 421 2959 455
rect 2993 421 3005 455
rect 2948 409 3005 421
rect 2139 352 2212 361
rect 1902 347 1975 352
<< ndiffc >>
rect 66 150 100 184
rect 246 142 280 176
rect 448 147 482 181
rect 606 150 640 184
rect 1135 171 1169 205
rect 1291 193 1325 227
rect 1377 180 1411 214
rect 714 91 748 125
rect 872 79 906 113
rect 1030 79 1064 113
rect 1487 141 1521 175
rect 1586 93 1620 127
rect 1757 150 1791 184
rect 1867 180 1901 214
rect 1966 193 2000 227
rect 2518 152 2552 186
rect 2065 53 2099 87
rect 2170 82 2204 116
rect 2256 69 2290 103
rect 2676 152 2710 186
rect 2834 152 2868 186
rect 2414 82 2448 116
rect 2940 82 2974 116
rect 3098 82 3132 116
<< pdiffc >>
rect 36 563 70 597
rect 36 492 70 526
rect 36 421 70 455
rect 142 563 176 597
rect 142 492 176 526
rect 142 421 176 455
rect 248 563 282 597
rect 248 429 282 463
rect 354 430 388 464
rect 554 571 588 605
rect 660 540 694 574
rect 774 360 808 394
rect 880 501 914 535
rect 986 360 1020 394
rect 1281 501 1315 535
rect 1281 433 1315 467
rect 1281 365 1315 399
rect 1387 501 1421 535
rect 1387 430 1421 464
rect 1387 359 1421 393
rect 1591 501 1625 535
rect 1591 419 1625 453
rect 1765 501 1799 535
rect 1765 430 1799 464
rect 1765 359 1799 393
rect 1929 506 1963 540
rect 1929 432 1963 466
rect 1929 359 1963 393
rect 2166 515 2200 549
rect 2166 442 2200 476
rect 2288 515 2322 549
rect 2288 442 2322 476
rect 2513 555 2547 589
rect 2513 484 2547 518
rect 2513 413 2547 447
rect 2619 555 2653 589
rect 2619 484 2653 518
rect 2619 413 2653 447
rect 2725 555 2759 589
rect 2725 484 2759 518
rect 2725 413 2759 447
rect 2853 563 2887 597
rect 2853 483 2887 517
rect 2959 563 2993 597
rect 2959 492 2993 526
rect 2959 421 2993 455
<< poly >>
rect 81 609 131 635
rect 293 617 343 643
rect 399 617 449 643
rect 493 617 543 643
rect 599 617 649 643
rect 1103 615 2040 645
rect 819 547 869 573
rect 925 547 975 573
rect 81 369 131 409
rect 81 353 172 369
rect 293 367 343 417
rect 399 377 449 417
rect 81 319 122 353
rect 156 333 172 353
rect 271 351 337 367
rect 156 319 219 333
rect 81 303 219 319
rect 111 209 141 303
rect 189 209 219 303
rect 271 317 287 351
rect 321 317 337 351
rect 271 283 337 317
rect 271 249 287 283
rect 321 249 337 283
rect 271 233 337 249
rect 307 209 337 233
rect 385 361 451 377
rect 385 327 401 361
rect 435 327 451 361
rect 385 293 451 327
rect 385 259 401 293
rect 435 259 451 293
rect 385 243 451 259
rect 493 327 543 417
rect 599 383 649 417
rect 591 367 657 383
rect 591 333 607 367
rect 641 333 657 367
rect 1103 395 1133 615
rect 1326 547 1376 615
rect 1432 547 1482 573
rect 1530 547 1580 573
rect 1704 547 1754 573
rect 1852 547 1902 573
rect 1990 552 2040 615
rect 2558 601 2608 627
rect 2664 601 2714 627
rect 2898 609 2948 635
rect 2089 552 2139 578
rect 2227 561 2277 587
rect 1067 379 1133 395
rect 385 209 415 243
rect 493 209 523 327
rect 591 299 657 333
rect 819 302 869 347
rect 925 306 975 347
rect 1067 345 1083 379
rect 1117 345 1133 379
rect 2558 361 2608 401
rect 2664 361 2714 401
rect 1067 311 1133 345
rect 1326 321 1376 347
rect 591 279 607 299
rect 565 265 607 279
rect 641 265 657 299
rect 565 249 657 265
rect 759 286 869 302
rect 759 252 775 286
rect 809 252 869 286
rect 565 209 595 249
rect 759 236 869 252
rect 917 290 1019 306
rect 917 256 933 290
rect 967 256 1019 290
rect 1067 277 1083 311
rect 1117 291 1133 311
rect 1117 277 1278 291
rect 1067 261 1278 277
rect 759 150 789 236
rect 831 150 861 236
rect 917 222 1019 256
rect 1248 239 1278 261
rect 1336 239 1366 265
rect 1432 254 1482 347
rect 1530 297 1580 347
rect 1704 315 1754 347
rect 1644 299 1754 315
rect 1530 281 1596 297
rect 917 188 933 222
rect 967 188 1019 222
rect 917 172 1019 188
rect 917 150 947 172
rect 989 150 1019 172
rect 111 99 141 125
rect 189 51 219 125
rect 307 99 337 125
rect 385 99 415 125
rect 493 51 523 125
rect 565 99 595 125
rect 1248 129 1278 155
rect 189 21 523 51
rect 759 40 789 66
rect 831 40 861 66
rect 917 40 947 66
rect 989 51 1019 66
rect 1336 51 1366 155
rect 1434 51 1464 254
rect 1530 247 1546 281
rect 1580 247 1596 281
rect 1530 231 1596 247
rect 1644 265 1660 299
rect 1694 265 1754 299
rect 1852 284 1902 347
rect 1990 310 2040 352
rect 2089 320 2139 352
rect 2227 329 2277 361
rect 2495 345 2833 361
rect 1644 249 1754 265
rect 1814 254 1942 284
rect 1990 280 2041 310
rect 1532 209 1562 231
rect 1644 209 1674 249
rect 1716 209 1746 249
rect 1532 99 1562 125
rect 1644 99 1674 125
rect 1716 99 1746 125
rect 1814 51 1844 254
rect 1912 239 1942 254
rect 2011 239 2041 280
rect 2089 304 2179 320
rect 2089 270 2129 304
rect 2163 270 2179 304
rect 2089 254 2179 270
rect 2227 313 2331 329
rect 2227 279 2260 313
rect 2294 279 2331 313
rect 2495 311 2511 345
rect 2545 311 2579 345
rect 2613 311 2647 345
rect 2681 311 2715 345
rect 2749 311 2783 345
rect 2817 311 2833 345
rect 2495 295 2833 311
rect 2898 315 2948 409
rect 2898 299 3015 315
rect 2227 263 2331 279
rect 2149 215 2179 254
rect 2149 185 2245 215
rect 1912 129 1942 155
rect 2011 129 2041 155
rect 989 21 1844 51
rect 2215 141 2245 185
rect 2301 186 2331 263
rect 2563 211 2593 295
rect 2635 211 2665 295
rect 2721 211 2751 295
rect 2793 211 2823 295
rect 2898 265 2915 299
rect 2949 265 3015 299
rect 2898 231 3015 265
rect 2301 156 2403 186
rect 2301 141 2331 156
rect 2373 141 2403 156
rect 2898 197 2915 231
rect 2949 211 3015 231
rect 2949 197 3087 211
rect 2898 181 3087 197
rect 2985 141 3015 181
rect 3057 141 3087 181
rect 2563 101 2593 127
rect 2635 101 2665 127
rect 2721 101 2751 127
rect 2793 101 2823 127
rect 2215 31 2245 57
rect 2301 31 2331 57
rect 2373 31 2403 57
rect 2985 31 3015 57
rect 3057 31 3087 57
<< polycont >>
rect 122 319 156 353
rect 287 317 321 351
rect 287 249 321 283
rect 401 327 435 361
rect 401 259 435 293
rect 607 333 641 367
rect 1083 345 1117 379
rect 607 265 641 299
rect 775 252 809 286
rect 933 256 967 290
rect 1083 277 1117 311
rect 933 188 967 222
rect 1546 247 1580 281
rect 1660 265 1694 299
rect 2129 270 2163 304
rect 2260 279 2294 313
rect 2511 311 2545 345
rect 2579 311 2613 345
rect 2647 311 2681 345
rect 2715 311 2749 345
rect 2783 311 2817 345
rect 2915 265 2949 299
rect 2915 197 2949 231
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 20 597 70 613
rect 20 563 36 597
rect 20 526 70 563
rect 20 492 36 526
rect 20 455 70 492
rect 20 421 36 455
rect 20 267 70 421
rect 126 597 192 649
rect 126 563 142 597
rect 176 563 192 597
rect 126 526 192 563
rect 126 492 142 526
rect 176 492 192 526
rect 126 455 192 492
rect 126 421 142 455
rect 176 421 192 455
rect 126 405 192 421
rect 232 597 298 613
rect 232 563 248 597
rect 282 563 298 597
rect 538 605 604 649
rect 538 571 554 605
rect 588 571 604 605
rect 644 574 710 613
rect 232 535 298 563
rect 644 540 660 574
rect 694 540 710 574
rect 644 535 710 540
rect 232 501 710 535
rect 864 535 930 649
rect 864 501 880 535
rect 914 501 930 535
rect 1205 535 1331 551
rect 1205 501 1281 535
rect 1315 501 1331 535
rect 232 463 298 501
rect 1205 467 1331 501
rect 1205 465 1281 467
rect 232 429 248 463
rect 282 429 298 463
rect 232 413 298 429
rect 338 464 1281 465
rect 338 430 354 464
rect 388 433 1281 464
rect 1315 433 1331 467
rect 388 431 1331 433
rect 388 430 525 431
rect 338 413 525 430
rect 106 353 172 369
rect 106 319 122 353
rect 156 319 172 353
rect 106 303 172 319
rect 271 351 337 367
rect 271 317 287 351
rect 321 317 337 351
rect 271 283 337 317
rect 271 267 287 283
rect 20 249 287 267
rect 321 249 337 283
rect 20 233 337 249
rect 385 361 455 377
rect 385 327 401 361
rect 435 327 455 361
rect 385 293 455 327
rect 385 259 401 293
rect 435 259 455 293
rect 385 243 455 259
rect 20 184 116 233
rect 491 207 525 413
rect 1205 399 1331 431
rect 758 394 909 395
rect 591 367 657 383
rect 591 333 607 367
rect 641 333 657 367
rect 758 360 774 394
rect 808 360 909 394
rect 758 343 909 360
rect 970 394 1132 395
rect 970 360 986 394
rect 1020 379 1132 394
rect 1020 360 1083 379
rect 970 345 1083 360
rect 1117 345 1132 379
rect 970 343 1132 345
rect 591 299 657 333
rect 875 306 909 343
rect 1046 311 1132 343
rect 591 265 607 299
rect 641 265 657 299
rect 591 249 657 265
rect 697 286 839 302
rect 697 252 775 286
rect 809 252 839 286
rect 697 236 839 252
rect 875 290 982 306
rect 875 256 933 290
rect 967 256 982 290
rect 875 222 982 256
rect 20 150 66 184
rect 100 150 116 184
rect 20 121 116 150
rect 230 176 296 197
rect 230 142 246 176
rect 280 142 296 176
rect 230 17 296 142
rect 432 181 525 207
rect 432 147 448 181
rect 482 147 525 181
rect 432 121 525 147
rect 590 184 656 213
rect 875 200 933 222
rect 590 150 606 184
rect 640 150 656 184
rect 590 17 656 150
rect 698 188 933 200
rect 967 188 982 222
rect 698 166 982 188
rect 1046 277 1083 311
rect 1117 277 1132 311
rect 1046 261 1132 277
rect 1205 365 1281 399
rect 1315 365 1331 399
rect 1205 349 1331 365
rect 1371 535 1437 551
rect 1371 501 1387 535
rect 1421 501 1437 535
rect 1371 464 1437 501
rect 1371 430 1387 464
rect 1421 430 1437 464
rect 1371 393 1437 430
rect 1575 535 1641 649
rect 1575 501 1591 535
rect 1625 501 1641 535
rect 1575 453 1641 501
rect 1575 419 1591 453
rect 1625 419 1641 453
rect 1575 403 1641 419
rect 1749 535 1815 551
rect 1749 501 1765 535
rect 1799 501 1815 535
rect 1749 464 1815 501
rect 1749 430 1765 464
rect 1799 430 1815 464
rect 1371 359 1387 393
rect 1421 367 1437 393
rect 1749 393 1815 430
rect 1421 359 1710 367
rect 698 125 764 166
rect 1046 130 1080 261
rect 698 91 714 125
rect 748 91 764 125
rect 698 62 764 91
rect 856 113 922 130
rect 856 79 872 113
rect 906 79 922 113
rect 856 17 922 79
rect 1014 113 1080 130
rect 1014 79 1030 113
rect 1064 79 1080 113
rect 1014 62 1080 79
rect 1119 205 1169 225
rect 1119 171 1135 205
rect 1119 87 1169 171
rect 1205 157 1239 349
rect 1371 333 1710 359
rect 1371 313 1437 333
rect 1275 279 1437 313
rect 1644 299 1710 333
rect 1530 281 1596 297
rect 1275 227 1341 279
rect 1530 247 1546 281
rect 1580 247 1596 281
rect 1644 265 1660 299
rect 1694 265 1710 299
rect 1644 249 1710 265
rect 1749 359 1765 393
rect 1799 359 1815 393
rect 1275 193 1291 227
rect 1325 193 1341 227
rect 1377 214 1427 243
rect 1530 231 1596 247
rect 1411 180 1427 214
rect 1562 213 1596 231
rect 1749 213 1815 359
rect 1913 540 1979 556
rect 1913 506 1929 540
rect 1963 506 1979 540
rect 1913 466 1979 506
rect 1913 432 1929 466
rect 1963 432 1979 466
rect 1913 393 1979 432
rect 2150 549 2216 649
rect 2425 589 2567 605
rect 2150 515 2166 549
rect 2200 515 2216 549
rect 2150 476 2216 515
rect 2150 442 2166 476
rect 2200 442 2216 476
rect 2150 426 2216 442
rect 2272 549 2338 565
rect 2272 515 2288 549
rect 2322 515 2338 549
rect 2272 476 2338 515
rect 2272 442 2288 476
rect 2322 460 2338 476
rect 2425 555 2513 589
rect 2547 555 2567 589
rect 2425 518 2567 555
rect 2425 484 2513 518
rect 2547 484 2567 518
rect 2322 442 2380 460
rect 2272 426 2380 442
rect 1913 359 1929 393
rect 1963 390 1979 393
rect 1963 359 2310 390
rect 1913 356 2310 359
rect 1913 343 2016 356
rect 1377 157 1427 180
rect 1205 123 1427 157
rect 1471 175 1521 195
rect 1562 184 1815 213
rect 1562 179 1757 184
rect 1471 141 1487 175
rect 1741 150 1757 179
rect 1791 150 1815 184
rect 1471 87 1521 141
rect 1119 53 1521 87
rect 1570 127 1636 143
rect 1570 93 1586 127
rect 1620 93 1636 127
rect 1570 17 1636 93
rect 1741 87 1815 150
rect 1851 214 1901 243
rect 1851 180 1867 214
rect 1950 227 2016 343
rect 1950 193 1966 227
rect 2000 193 2016 227
rect 2113 304 2179 320
rect 2113 270 2129 304
rect 2163 270 2179 304
rect 2113 227 2179 270
rect 2244 313 2310 356
rect 2244 279 2260 313
rect 2294 279 2310 313
rect 2244 263 2310 279
rect 2346 227 2380 426
rect 2113 193 2380 227
rect 2425 447 2567 484
rect 2425 413 2513 447
rect 2547 413 2567 447
rect 2425 397 2567 413
rect 2603 589 2669 649
rect 2603 555 2619 589
rect 2653 555 2669 589
rect 2603 518 2669 555
rect 2603 484 2619 518
rect 2653 484 2669 518
rect 2603 447 2669 484
rect 2603 413 2619 447
rect 2653 413 2669 447
rect 2603 397 2669 413
rect 2709 589 2775 605
rect 2709 555 2725 589
rect 2759 555 2775 589
rect 2709 518 2775 555
rect 2709 484 2725 518
rect 2759 484 2775 518
rect 2709 447 2775 484
rect 2837 597 2903 649
rect 2837 563 2853 597
rect 2887 563 2903 597
rect 2837 517 2903 563
rect 2837 483 2853 517
rect 2887 483 2903 517
rect 2837 467 2903 483
rect 2943 597 3148 613
rect 2943 563 2959 597
rect 2993 563 3148 597
rect 2943 526 3148 563
rect 2943 492 2959 526
rect 2993 492 3148 526
rect 2709 413 2725 447
rect 2759 431 2775 447
rect 2943 455 3148 492
rect 2759 413 2903 431
rect 2709 397 2903 413
rect 2425 259 2459 397
rect 2495 345 2833 361
rect 2495 311 2511 345
rect 2545 311 2579 345
rect 2613 311 2647 345
rect 2681 311 2715 345
rect 2749 311 2783 345
rect 2817 311 2833 345
rect 2495 295 2833 311
rect 2869 315 2903 397
rect 2943 421 2959 455
rect 2993 421 3148 455
rect 2943 384 3148 421
rect 2869 299 2965 315
rect 2425 225 2552 259
rect 1851 157 1901 180
rect 2346 189 2380 193
rect 1851 123 2220 157
rect 2346 155 2464 189
rect 2154 116 2220 123
rect 1741 53 2065 87
rect 2099 53 2115 87
rect 2154 82 2170 116
rect 2204 82 2220 116
rect 2154 53 2220 82
rect 2256 103 2306 119
rect 2290 69 2306 103
rect 2256 17 2306 69
rect 2398 116 2464 155
rect 2502 186 2552 225
rect 2502 152 2518 186
rect 2502 123 2552 152
rect 2398 82 2414 116
rect 2448 87 2464 116
rect 2588 87 2622 295
rect 2869 265 2915 299
rect 2949 265 2965 299
rect 2869 231 2965 265
rect 2869 215 2915 231
rect 2448 82 2622 87
rect 2398 53 2622 82
rect 2660 186 2726 215
rect 2660 152 2676 186
rect 2710 152 2726 186
rect 2660 17 2726 152
rect 2818 197 2915 215
rect 2949 197 2965 231
rect 2818 186 2965 197
rect 2818 152 2834 186
rect 2868 181 2965 186
rect 2868 152 2884 181
rect 2818 123 2884 152
rect 2924 116 2990 145
rect 2924 82 2940 116
rect 2974 82 2990 116
rect 2924 17 2990 82
rect 3082 116 3148 384
rect 3082 82 3098 116
rect 3132 82 3148 116
rect 3082 53 3148 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
<< metal1 >>
rect 0 683 3168 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 0 617 3168 649
rect 0 17 3168 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
rect 0 -49 3168 -17
<< labels >>
flabel pwell s 0 0 3168 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 3168 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfxbp_lp
flabel metal1 s 0 617 3168 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 3168 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2431 464 2465 498 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2431 538 2465 572 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2527 464 2561 498 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2527 538 2561 572 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 3007 390 3041 424 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 3007 464 3041 498 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 3007 538 3041 572 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 3103 390 3137 424 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 3103 464 3137 498 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 3103 538 3137 572 0 FreeSans 340 0 0 0 Q_N
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3168 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6323682
string GDS_START 6303548
<< end >>
