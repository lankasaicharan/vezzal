magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 14 49 629 241
rect 0 0 672 49
<< scnmos >>
rect 93 131 123 215
rect 262 47 292 215
rect 348 47 378 215
rect 434 47 464 215
rect 520 47 550 215
<< scpmoshvt >>
rect 148 367 178 451
rect 253 367 283 619
rect 339 367 369 619
rect 425 367 455 619
rect 511 367 541 619
<< ndiff >>
rect 40 190 93 215
rect 40 156 48 190
rect 82 156 93 190
rect 40 131 93 156
rect 123 187 262 215
rect 123 153 134 187
rect 168 161 262 187
rect 168 153 217 161
rect 123 131 217 153
rect 141 127 217 131
rect 251 127 262 161
rect 141 93 262 127
rect 141 59 149 93
rect 183 59 217 93
rect 251 59 262 93
rect 141 47 262 59
rect 292 181 348 215
rect 292 147 303 181
rect 337 147 348 181
rect 292 101 348 147
rect 292 67 303 101
rect 337 67 348 101
rect 292 47 348 67
rect 378 105 434 215
rect 378 71 389 105
rect 423 71 434 105
rect 378 47 434 71
rect 464 181 520 215
rect 464 147 475 181
rect 509 147 520 181
rect 464 101 520 147
rect 464 67 475 101
rect 509 67 520 101
rect 464 47 520 67
rect 550 105 603 215
rect 550 71 561 105
rect 595 71 603 105
rect 550 47 603 71
<< pdiff >>
rect 200 607 253 619
rect 200 573 208 607
rect 242 573 253 607
rect 200 526 253 573
rect 200 492 208 526
rect 242 492 253 526
rect 200 451 253 492
rect 95 426 148 451
rect 95 392 103 426
rect 137 392 148 426
rect 95 367 148 392
rect 178 439 253 451
rect 178 405 189 439
rect 223 405 253 439
rect 178 367 253 405
rect 283 599 339 619
rect 283 565 294 599
rect 328 565 339 599
rect 283 529 339 565
rect 283 495 294 529
rect 328 495 339 529
rect 283 455 339 495
rect 283 421 294 455
rect 328 421 339 455
rect 283 367 339 421
rect 369 539 425 619
rect 369 505 380 539
rect 414 505 425 539
rect 369 439 425 505
rect 369 405 380 439
rect 414 405 425 439
rect 369 367 425 405
rect 455 599 511 619
rect 455 565 466 599
rect 500 565 511 599
rect 455 523 511 565
rect 455 489 466 523
rect 500 489 511 523
rect 455 367 511 489
rect 541 607 594 619
rect 541 573 552 607
rect 586 573 594 607
rect 541 511 594 573
rect 541 477 552 511
rect 586 477 594 511
rect 541 367 594 477
<< ndiffc >>
rect 48 156 82 190
rect 134 153 168 187
rect 217 127 251 161
rect 149 59 183 93
rect 217 59 251 93
rect 303 147 337 181
rect 303 67 337 101
rect 389 71 423 105
rect 475 147 509 181
rect 475 67 509 101
rect 561 71 595 105
<< pdiffc >>
rect 208 573 242 607
rect 208 492 242 526
rect 103 392 137 426
rect 189 405 223 439
rect 294 565 328 599
rect 294 495 328 529
rect 294 421 328 455
rect 380 505 414 539
rect 380 405 414 439
rect 466 565 500 599
rect 466 489 500 523
rect 552 573 586 607
rect 552 477 586 511
<< poly >>
rect 253 619 283 645
rect 339 619 369 645
rect 425 619 455 645
rect 511 619 541 645
rect 148 451 178 477
rect 148 303 178 367
rect 253 303 283 367
rect 339 335 369 367
rect 425 335 455 367
rect 339 319 455 335
rect 93 287 178 303
rect 93 253 127 287
rect 161 253 178 287
rect 93 237 178 253
rect 220 287 297 303
rect 220 253 236 287
rect 270 253 297 287
rect 339 285 405 319
rect 439 299 455 319
rect 511 303 541 367
rect 439 285 464 299
rect 339 269 464 285
rect 339 267 378 269
rect 220 237 297 253
rect 93 215 123 237
rect 262 215 292 237
rect 348 215 378 267
rect 434 215 464 269
rect 511 287 577 303
rect 511 253 527 287
rect 561 253 577 287
rect 511 237 577 253
rect 520 215 550 237
rect 93 105 123 131
rect 262 21 292 47
rect 348 21 378 47
rect 434 21 464 47
rect 520 21 550 47
<< polycont >>
rect 127 253 161 287
rect 236 253 270 287
rect 405 285 439 319
rect 527 253 561 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 173 607 250 649
rect 173 573 208 607
rect 242 573 250 607
rect 173 526 250 573
rect 173 492 208 526
rect 242 492 250 526
rect 32 426 139 442
rect 32 392 103 426
rect 137 392 139 426
rect 173 439 250 492
rect 173 405 189 439
rect 223 405 250 439
rect 284 599 502 615
rect 284 565 294 599
rect 328 579 466 599
rect 328 565 330 579
rect 284 529 330 565
rect 464 565 466 579
rect 500 565 502 599
rect 284 495 294 529
rect 328 495 330 529
rect 284 455 330 495
rect 284 421 294 455
rect 328 421 330 455
rect 284 405 330 421
rect 364 539 430 543
rect 364 505 380 539
rect 414 505 430 539
rect 364 439 430 505
rect 464 523 502 565
rect 464 489 466 523
rect 500 489 502 523
rect 464 473 502 489
rect 536 607 602 649
rect 536 573 552 607
rect 586 573 602 607
rect 536 511 602 573
rect 536 477 552 511
rect 586 477 602 511
rect 536 473 602 477
rect 364 405 380 439
rect 414 405 655 439
rect 32 371 139 392
rect 32 337 455 371
rect 32 190 86 337
rect 389 319 455 337
rect 120 287 177 303
rect 120 253 127 287
rect 161 253 177 287
rect 120 237 177 253
rect 211 253 236 287
rect 270 253 355 287
rect 389 285 405 319
rect 439 285 455 319
rect 389 283 455 285
rect 511 287 563 303
rect 211 249 355 253
rect 511 253 527 287
rect 561 253 563 287
rect 511 249 563 253
rect 211 215 563 249
rect 32 156 48 190
rect 82 156 86 190
rect 32 140 86 156
rect 124 187 179 203
rect 124 153 134 187
rect 168 177 179 187
rect 597 181 655 405
rect 168 161 253 177
rect 168 153 217 161
rect 124 127 217 153
rect 251 127 253 161
rect 124 93 253 127
rect 124 59 149 93
rect 183 59 217 93
rect 251 59 253 93
rect 124 17 253 59
rect 287 147 303 181
rect 337 147 475 181
rect 509 147 655 181
rect 287 101 339 147
rect 287 67 303 101
rect 337 67 339 101
rect 287 51 339 67
rect 373 105 439 113
rect 373 71 389 105
rect 423 71 439 105
rect 373 17 439 71
rect 473 101 511 147
rect 473 67 475 101
rect 509 67 511 101
rect 473 51 511 67
rect 545 105 611 113
rect 545 71 561 105
rect 595 71 611 105
rect 545 17 611 71
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 isobufsrc_2
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 SLEEP
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 SLEEP
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y
string GDS_END 1259016
string GDS_START 1252668
<< end >>
