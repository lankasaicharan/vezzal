magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1778 1975
<< nwell >>
rect -38 331 518 704
<< pwell >>
rect 6 49 438 161
rect 0 0 480 49
<< scnmos >>
rect 89 51 119 135
rect 161 51 191 135
rect 247 51 277 135
rect 325 51 355 135
<< scpmoshvt >>
rect 113 419 163 619
rect 219 419 269 619
rect 325 419 375 619
<< ndiff >>
rect 32 113 89 135
rect 32 79 44 113
rect 78 79 89 113
rect 32 51 89 79
rect 119 51 161 135
rect 191 110 247 135
rect 191 76 202 110
rect 236 76 247 110
rect 191 51 247 76
rect 277 51 325 135
rect 355 113 412 135
rect 355 79 366 113
rect 400 79 412 113
rect 355 51 412 79
<< pdiff >>
rect 56 597 113 619
rect 56 563 68 597
rect 102 563 113 597
rect 56 465 113 563
rect 56 431 68 465
rect 102 431 113 465
rect 56 419 113 431
rect 163 607 219 619
rect 163 573 174 607
rect 208 573 219 607
rect 163 536 219 573
rect 163 502 174 536
rect 208 502 219 536
rect 163 465 219 502
rect 163 431 174 465
rect 208 431 219 465
rect 163 419 219 431
rect 269 597 325 619
rect 269 563 280 597
rect 314 563 325 597
rect 269 465 325 563
rect 269 431 280 465
rect 314 431 325 465
rect 269 419 325 431
rect 375 607 445 619
rect 375 573 399 607
rect 433 573 445 607
rect 375 516 445 573
rect 375 482 399 516
rect 433 482 445 516
rect 375 419 445 482
<< ndiffc >>
rect 44 79 78 113
rect 202 76 236 110
rect 366 79 400 113
<< pdiffc >>
rect 68 563 102 597
rect 68 431 102 465
rect 174 573 208 607
rect 174 502 208 536
rect 174 431 208 465
rect 280 563 314 597
rect 280 431 314 465
rect 399 573 433 607
rect 399 482 433 516
<< poly >>
rect 113 619 163 645
rect 219 619 269 645
rect 325 619 375 645
rect 113 379 163 419
rect 219 379 269 419
rect 89 363 163 379
rect 89 329 113 363
rect 147 329 163 363
rect 89 295 163 329
rect 89 261 113 295
rect 147 261 163 295
rect 89 245 163 261
rect 211 363 277 379
rect 211 329 227 363
rect 261 329 277 363
rect 211 295 277 329
rect 211 261 227 295
rect 261 261 277 295
rect 211 245 277 261
rect 89 180 119 245
rect 89 150 191 180
rect 89 135 119 150
rect 161 135 191 150
rect 247 135 277 245
rect 325 309 375 419
rect 325 293 391 309
rect 325 259 341 293
rect 375 259 391 293
rect 325 225 391 259
rect 325 191 341 225
rect 375 191 391 225
rect 325 175 391 191
rect 325 135 355 175
rect 89 25 119 51
rect 161 25 191 51
rect 247 25 277 51
rect 325 25 355 51
<< polycont >>
rect 113 329 147 363
rect 113 261 147 295
rect 227 329 261 363
rect 227 261 261 295
rect 341 259 375 293
rect 341 191 375 225
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 27 597 118 613
rect 27 563 68 597
rect 102 563 118 597
rect 27 465 118 563
rect 27 431 68 465
rect 102 431 118 465
rect 27 415 118 431
rect 158 607 224 649
rect 158 573 174 607
rect 208 573 224 607
rect 158 536 224 573
rect 158 502 174 536
rect 208 502 224 536
rect 158 465 224 502
rect 158 431 174 465
rect 208 431 224 465
rect 158 415 224 431
rect 264 597 347 613
rect 264 563 280 597
rect 314 563 347 597
rect 264 465 347 563
rect 383 607 449 649
rect 383 573 399 607
rect 433 573 449 607
rect 383 516 449 573
rect 383 482 399 516
rect 433 482 449 516
rect 383 466 449 482
rect 264 431 280 465
rect 314 431 347 465
rect 264 430 347 431
rect 264 415 461 430
rect 27 209 61 415
rect 313 384 461 415
rect 97 363 167 379
rect 97 329 113 363
rect 147 329 167 363
rect 97 295 167 329
rect 97 261 113 295
rect 147 261 167 295
rect 97 245 167 261
rect 211 363 277 379
rect 211 329 227 363
rect 261 329 277 363
rect 211 295 277 329
rect 211 261 227 295
rect 261 261 277 295
rect 211 245 277 261
rect 325 293 391 309
rect 325 259 341 293
rect 375 259 391 293
rect 325 225 391 259
rect 325 209 341 225
rect 27 191 341 209
rect 375 191 391 225
rect 27 175 391 191
rect 27 113 94 175
rect 427 139 461 384
rect 27 79 44 113
rect 78 79 94 113
rect 27 53 94 79
rect 186 110 252 139
rect 186 76 202 110
rect 236 76 252 110
rect 186 17 252 76
rect 350 113 461 139
rect 350 79 366 113
rect 400 79 461 113
rect 350 53 461 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2b_lp
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4445084
string GDS_START 4440370
<< end >>
