magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3122 1975
<< nwell >>
rect -38 331 1862 704
<< pwell >>
rect 3 49 1765 241
rect 0 0 1824 49
<< scnmos >>
rect 82 47 112 215
rect 178 47 208 215
rect 264 47 294 215
rect 360 47 390 215
rect 446 47 476 215
rect 602 47 632 215
rect 688 47 718 215
rect 774 47 804 215
rect 860 47 890 215
rect 1046 47 1076 215
rect 1132 47 1162 215
rect 1218 47 1248 215
rect 1304 47 1334 215
rect 1392 47 1422 215
rect 1484 47 1514 215
rect 1570 47 1600 215
rect 1656 47 1686 215
<< scpmoshvt >>
rect 80 367 110 619
rect 270 367 300 619
rect 356 367 386 619
rect 442 367 472 619
rect 528 367 558 619
rect 614 367 644 619
rect 700 367 730 619
rect 786 367 816 619
rect 872 367 902 619
rect 1062 367 1092 619
rect 1148 367 1178 619
rect 1234 367 1264 619
rect 1320 367 1350 619
rect 1406 367 1436 619
rect 1492 367 1522 619
rect 1578 367 1608 619
rect 1664 367 1694 619
<< ndiff >>
rect 29 203 82 215
rect 29 169 37 203
rect 71 169 82 203
rect 29 101 82 169
rect 29 67 37 101
rect 71 67 82 101
rect 29 47 82 67
rect 112 163 178 215
rect 112 129 123 163
rect 157 129 178 163
rect 112 89 178 129
rect 112 55 123 89
rect 157 55 178 89
rect 112 47 178 55
rect 208 203 264 215
rect 208 169 219 203
rect 253 169 264 203
rect 208 101 264 169
rect 208 67 219 101
rect 253 67 264 101
rect 208 47 264 67
rect 294 159 360 215
rect 294 125 309 159
rect 343 125 360 159
rect 294 89 360 125
rect 294 55 309 89
rect 343 55 360 89
rect 294 47 360 55
rect 390 203 446 215
rect 390 169 401 203
rect 435 169 446 203
rect 390 101 446 169
rect 390 67 401 101
rect 435 67 446 101
rect 390 47 446 67
rect 476 157 602 215
rect 476 123 487 157
rect 521 123 557 157
rect 591 123 602 157
rect 476 89 602 123
rect 476 55 487 89
rect 521 55 557 89
rect 591 55 602 89
rect 476 47 602 55
rect 632 203 688 215
rect 632 169 643 203
rect 677 169 688 203
rect 632 101 688 169
rect 632 67 643 101
rect 677 67 688 101
rect 632 47 688 67
rect 718 127 774 215
rect 718 93 729 127
rect 763 93 774 127
rect 718 47 774 93
rect 804 186 860 215
rect 804 152 815 186
rect 849 152 860 186
rect 804 101 860 152
rect 804 67 815 101
rect 849 67 860 101
rect 804 47 860 67
rect 890 123 1046 215
rect 890 89 901 123
rect 935 89 1001 123
rect 1035 89 1046 123
rect 890 47 1046 89
rect 1076 198 1132 215
rect 1076 164 1087 198
rect 1121 164 1132 198
rect 1076 101 1132 164
rect 1076 67 1087 101
rect 1121 67 1132 101
rect 1076 47 1132 67
rect 1162 167 1218 215
rect 1162 133 1173 167
rect 1207 133 1218 167
rect 1162 93 1218 133
rect 1162 59 1173 93
rect 1207 59 1218 93
rect 1162 47 1218 59
rect 1248 203 1304 215
rect 1248 169 1259 203
rect 1293 169 1304 203
rect 1248 101 1304 169
rect 1248 67 1259 101
rect 1293 67 1304 101
rect 1248 47 1304 67
rect 1334 167 1392 215
rect 1334 133 1345 167
rect 1379 133 1392 167
rect 1334 93 1392 133
rect 1334 59 1345 93
rect 1379 59 1392 93
rect 1334 47 1392 59
rect 1422 203 1484 215
rect 1422 169 1435 203
rect 1469 169 1484 203
rect 1422 101 1484 169
rect 1422 67 1435 101
rect 1469 67 1484 101
rect 1422 47 1484 67
rect 1514 124 1570 215
rect 1514 90 1525 124
rect 1559 90 1570 124
rect 1514 47 1570 90
rect 1600 192 1656 215
rect 1600 158 1611 192
rect 1645 158 1656 192
rect 1600 101 1656 158
rect 1600 67 1611 101
rect 1645 67 1656 101
rect 1600 47 1656 67
rect 1686 203 1739 215
rect 1686 169 1697 203
rect 1731 169 1739 203
rect 1686 93 1739 169
rect 1686 59 1697 93
rect 1731 59 1739 93
rect 1686 47 1739 59
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 521 80 565
rect 27 487 35 521
rect 69 487 80 521
rect 27 436 80 487
rect 27 402 35 436
rect 69 402 80 436
rect 27 367 80 402
rect 110 607 163 619
rect 110 573 121 607
rect 155 573 163 607
rect 110 497 163 573
rect 110 463 121 497
rect 155 463 163 497
rect 110 367 163 463
rect 217 599 270 619
rect 217 565 225 599
rect 259 565 270 599
rect 217 510 270 565
rect 217 476 225 510
rect 259 476 270 510
rect 217 413 270 476
rect 217 379 225 413
rect 259 379 270 413
rect 217 367 270 379
rect 300 547 356 619
rect 300 513 311 547
rect 345 513 356 547
rect 300 477 356 513
rect 300 443 311 477
rect 345 443 356 477
rect 300 409 356 443
rect 300 375 311 409
rect 345 375 356 409
rect 300 367 356 375
rect 386 599 442 619
rect 386 565 397 599
rect 431 565 442 599
rect 386 521 442 565
rect 386 487 397 521
rect 431 487 442 521
rect 386 451 442 487
rect 386 417 397 451
rect 431 417 442 451
rect 386 367 442 417
rect 472 547 528 619
rect 472 513 483 547
rect 517 513 528 547
rect 472 477 528 513
rect 472 443 483 477
rect 517 443 528 477
rect 472 409 528 443
rect 472 375 483 409
rect 517 375 528 409
rect 472 367 528 375
rect 558 599 614 619
rect 558 565 569 599
rect 603 565 614 599
rect 558 521 614 565
rect 558 487 569 521
rect 603 487 614 521
rect 558 451 614 487
rect 558 417 569 451
rect 603 417 614 451
rect 558 367 614 417
rect 644 543 700 619
rect 644 509 655 543
rect 689 509 700 543
rect 644 439 700 509
rect 644 405 655 439
rect 689 405 700 439
rect 644 367 700 405
rect 730 599 786 619
rect 730 565 741 599
rect 775 565 786 599
rect 730 521 786 565
rect 730 487 741 521
rect 775 487 786 521
rect 730 367 786 487
rect 816 531 872 619
rect 816 497 827 531
rect 861 497 872 531
rect 816 437 872 497
rect 816 403 827 437
rect 861 403 872 437
rect 816 367 872 403
rect 902 599 955 619
rect 902 565 913 599
rect 947 565 955 599
rect 902 509 955 565
rect 902 475 913 509
rect 947 475 955 509
rect 902 367 955 475
rect 1009 607 1062 619
rect 1009 573 1017 607
rect 1051 573 1062 607
rect 1009 511 1062 573
rect 1009 477 1017 511
rect 1051 477 1062 511
rect 1009 367 1062 477
rect 1092 531 1148 619
rect 1092 497 1103 531
rect 1137 497 1148 531
rect 1092 437 1148 497
rect 1092 403 1103 437
rect 1137 403 1148 437
rect 1092 367 1148 403
rect 1178 599 1234 619
rect 1178 565 1189 599
rect 1223 565 1234 599
rect 1178 521 1234 565
rect 1178 487 1189 521
rect 1223 487 1234 521
rect 1178 367 1234 487
rect 1264 543 1320 619
rect 1264 509 1275 543
rect 1309 509 1320 543
rect 1264 437 1320 509
rect 1264 403 1275 437
rect 1309 403 1320 437
rect 1264 367 1320 403
rect 1350 599 1406 619
rect 1350 565 1361 599
rect 1395 565 1406 599
rect 1350 506 1406 565
rect 1350 472 1361 506
rect 1395 472 1406 506
rect 1350 413 1406 472
rect 1350 379 1361 413
rect 1395 379 1406 413
rect 1350 367 1406 379
rect 1436 607 1492 619
rect 1436 573 1447 607
rect 1481 573 1492 607
rect 1436 530 1492 573
rect 1436 496 1447 530
rect 1481 496 1492 530
rect 1436 455 1492 496
rect 1436 421 1447 455
rect 1481 421 1492 455
rect 1436 367 1492 421
rect 1522 599 1578 619
rect 1522 565 1533 599
rect 1567 565 1578 599
rect 1522 506 1578 565
rect 1522 472 1533 506
rect 1567 472 1578 506
rect 1522 413 1578 472
rect 1522 379 1533 413
rect 1567 379 1578 413
rect 1522 367 1578 379
rect 1608 607 1664 619
rect 1608 573 1619 607
rect 1653 573 1664 607
rect 1608 530 1664 573
rect 1608 496 1619 530
rect 1653 496 1664 530
rect 1608 455 1664 496
rect 1608 421 1619 455
rect 1653 421 1664 455
rect 1608 367 1664 421
rect 1694 599 1747 619
rect 1694 565 1705 599
rect 1739 565 1747 599
rect 1694 506 1747 565
rect 1694 472 1705 506
rect 1739 472 1747 506
rect 1694 413 1747 472
rect 1694 379 1705 413
rect 1739 379 1747 413
rect 1694 367 1747 379
<< ndiffc >>
rect 37 169 71 203
rect 37 67 71 101
rect 123 129 157 163
rect 123 55 157 89
rect 219 169 253 203
rect 219 67 253 101
rect 309 125 343 159
rect 309 55 343 89
rect 401 169 435 203
rect 401 67 435 101
rect 487 123 521 157
rect 557 123 591 157
rect 487 55 521 89
rect 557 55 591 89
rect 643 169 677 203
rect 643 67 677 101
rect 729 93 763 127
rect 815 152 849 186
rect 815 67 849 101
rect 901 89 935 123
rect 1001 89 1035 123
rect 1087 164 1121 198
rect 1087 67 1121 101
rect 1173 133 1207 167
rect 1173 59 1207 93
rect 1259 169 1293 203
rect 1259 67 1293 101
rect 1345 133 1379 167
rect 1345 59 1379 93
rect 1435 169 1469 203
rect 1435 67 1469 101
rect 1525 90 1559 124
rect 1611 158 1645 192
rect 1611 67 1645 101
rect 1697 169 1731 203
rect 1697 59 1731 93
<< pdiffc >>
rect 35 565 69 599
rect 35 487 69 521
rect 35 402 69 436
rect 121 573 155 607
rect 121 463 155 497
rect 225 565 259 599
rect 225 476 259 510
rect 225 379 259 413
rect 311 513 345 547
rect 311 443 345 477
rect 311 375 345 409
rect 397 565 431 599
rect 397 487 431 521
rect 397 417 431 451
rect 483 513 517 547
rect 483 443 517 477
rect 483 375 517 409
rect 569 565 603 599
rect 569 487 603 521
rect 569 417 603 451
rect 655 509 689 543
rect 655 405 689 439
rect 741 565 775 599
rect 741 487 775 521
rect 827 497 861 531
rect 827 403 861 437
rect 913 565 947 599
rect 913 475 947 509
rect 1017 573 1051 607
rect 1017 477 1051 511
rect 1103 497 1137 531
rect 1103 403 1137 437
rect 1189 565 1223 599
rect 1189 487 1223 521
rect 1275 509 1309 543
rect 1275 403 1309 437
rect 1361 565 1395 599
rect 1361 472 1395 506
rect 1361 379 1395 413
rect 1447 573 1481 607
rect 1447 496 1481 530
rect 1447 421 1481 455
rect 1533 565 1567 599
rect 1533 472 1567 506
rect 1533 379 1567 413
rect 1619 573 1653 607
rect 1619 496 1653 530
rect 1619 421 1653 455
rect 1705 565 1739 599
rect 1705 472 1739 506
rect 1705 379 1739 413
<< poly >>
rect 80 619 110 645
rect 270 619 300 645
rect 356 619 386 645
rect 442 619 472 645
rect 528 619 558 645
rect 614 619 644 645
rect 700 619 730 645
rect 786 619 816 645
rect 872 619 902 645
rect 1062 619 1092 645
rect 1148 619 1178 645
rect 1234 619 1264 645
rect 1320 619 1350 645
rect 1406 619 1436 645
rect 1492 619 1522 645
rect 1578 619 1608 645
rect 1664 619 1694 645
rect 80 325 110 367
rect 44 309 112 325
rect 270 313 300 367
rect 356 313 386 367
rect 442 313 472 367
rect 528 313 558 367
rect 614 313 644 367
rect 700 313 730 367
rect 786 313 816 367
rect 872 313 902 367
rect 1062 335 1092 367
rect 1148 335 1178 367
rect 1234 335 1264 367
rect 1320 335 1350 367
rect 1046 319 1350 335
rect 1406 321 1436 367
rect 1492 321 1522 367
rect 1578 321 1608 367
rect 1664 321 1694 367
rect 44 275 60 309
rect 94 275 112 309
rect 44 259 112 275
rect 82 215 112 259
rect 154 297 560 313
rect 154 263 170 297
rect 204 263 238 297
rect 272 263 306 297
rect 340 263 374 297
rect 408 263 442 297
rect 476 263 510 297
rect 544 263 560 297
rect 154 247 560 263
rect 602 297 940 313
rect 602 263 618 297
rect 652 263 686 297
rect 720 263 754 297
rect 788 263 822 297
rect 856 263 890 297
rect 924 263 940 297
rect 602 247 940 263
rect 1046 285 1062 319
rect 1096 285 1130 319
rect 1164 285 1198 319
rect 1232 285 1266 319
rect 1300 285 1350 319
rect 1046 269 1350 285
rect 1392 305 1798 321
rect 1392 271 1408 305
rect 1442 271 1476 305
rect 1510 271 1544 305
rect 1578 271 1612 305
rect 1646 271 1680 305
rect 1714 271 1748 305
rect 1782 271 1798 305
rect 178 215 208 247
rect 264 215 294 247
rect 360 215 390 247
rect 446 215 476 247
rect 602 215 632 247
rect 688 215 718 247
rect 774 215 804 247
rect 860 215 890 247
rect 1046 215 1076 269
rect 1132 215 1162 269
rect 1218 215 1248 269
rect 1304 215 1334 269
rect 1392 255 1798 271
rect 1392 215 1422 255
rect 1484 215 1514 255
rect 1570 215 1600 255
rect 1656 215 1686 255
rect 82 21 112 47
rect 178 21 208 47
rect 264 21 294 47
rect 360 21 390 47
rect 446 21 476 47
rect 602 21 632 47
rect 688 21 718 47
rect 774 21 804 47
rect 860 21 890 47
rect 1046 21 1076 47
rect 1132 21 1162 47
rect 1218 21 1248 47
rect 1304 21 1334 47
rect 1392 21 1422 47
rect 1484 21 1514 47
rect 1570 21 1600 47
rect 1656 21 1686 47
<< polycont >>
rect 60 275 94 309
rect 170 263 204 297
rect 238 263 272 297
rect 306 263 340 297
rect 374 263 408 297
rect 442 263 476 297
rect 510 263 544 297
rect 618 263 652 297
rect 686 263 720 297
rect 754 263 788 297
rect 822 263 856 297
rect 890 263 924 297
rect 1062 285 1096 319
rect 1130 285 1164 319
rect 1198 285 1232 319
rect 1266 285 1300 319
rect 1408 271 1442 305
rect 1476 271 1510 305
rect 1544 271 1578 305
rect 1612 271 1646 305
rect 1680 271 1714 305
rect 1748 271 1782 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 19 599 71 615
rect 19 565 35 599
rect 69 565 71 599
rect 19 521 71 565
rect 19 487 35 521
rect 69 487 71 521
rect 19 436 71 487
rect 105 607 171 649
rect 105 573 121 607
rect 155 573 171 607
rect 105 497 171 573
rect 105 463 121 497
rect 155 463 171 497
rect 105 454 171 463
rect 219 599 963 615
rect 219 565 225 599
rect 259 581 397 599
rect 259 565 261 581
rect 219 510 261 565
rect 395 565 397 581
rect 431 581 569 599
rect 431 565 433 581
rect 219 476 225 510
rect 259 476 261 510
rect 19 402 35 436
rect 69 420 71 436
rect 69 402 185 420
rect 19 386 185 402
rect 17 309 110 352
rect 17 275 60 309
rect 94 275 110 309
rect 17 265 110 275
rect 144 297 185 386
rect 219 413 261 476
rect 219 379 225 413
rect 259 379 261 413
rect 219 363 261 379
rect 295 513 311 547
rect 345 513 361 547
rect 295 477 361 513
rect 295 443 311 477
rect 345 443 361 477
rect 295 409 361 443
rect 295 375 311 409
rect 345 375 361 409
rect 395 521 433 565
rect 567 565 569 581
rect 603 581 741 599
rect 603 565 605 581
rect 395 487 397 521
rect 431 487 433 521
rect 395 451 433 487
rect 395 417 397 451
rect 431 417 433 451
rect 395 401 433 417
rect 467 513 483 547
rect 517 513 533 547
rect 467 477 533 513
rect 467 443 483 477
rect 517 443 533 477
rect 467 409 533 443
rect 295 367 361 375
rect 467 375 483 409
rect 517 375 533 409
rect 567 521 605 565
rect 739 565 741 581
rect 775 581 913 599
rect 775 565 779 581
rect 567 487 569 521
rect 603 487 605 521
rect 567 451 605 487
rect 567 417 569 451
rect 603 417 605 451
rect 567 401 605 417
rect 639 543 705 547
rect 639 509 655 543
rect 689 509 705 543
rect 639 439 705 509
rect 739 521 779 565
rect 897 565 913 581
rect 947 565 963 599
rect 739 487 741 521
rect 775 487 779 521
rect 739 471 779 487
rect 823 531 863 547
rect 823 497 827 531
rect 861 497 863 531
rect 639 405 655 439
rect 689 437 705 439
rect 823 437 863 497
rect 897 509 963 565
rect 897 475 913 509
rect 947 475 963 509
rect 897 471 963 475
rect 1001 607 1397 615
rect 1001 573 1017 607
rect 1051 599 1397 607
rect 1051 581 1189 599
rect 1051 573 1067 581
rect 1001 511 1067 573
rect 1180 565 1189 581
rect 1223 581 1361 599
rect 1223 565 1225 581
rect 1001 477 1017 511
rect 1051 477 1067 511
rect 1001 471 1067 477
rect 1101 531 1146 547
rect 1101 497 1103 531
rect 1137 497 1146 531
rect 1101 437 1146 497
rect 1180 521 1225 565
rect 1359 565 1361 581
rect 1395 565 1397 599
rect 1180 487 1189 521
rect 1223 487 1225 521
rect 1180 471 1225 487
rect 1259 543 1325 547
rect 1259 509 1275 543
rect 1309 509 1325 543
rect 1259 437 1325 509
rect 689 405 827 437
rect 639 403 827 405
rect 861 403 1103 437
rect 1137 403 1275 437
rect 1309 403 1325 437
rect 639 401 1325 403
rect 1359 506 1397 565
rect 1359 472 1361 506
rect 1395 472 1397 506
rect 1359 413 1397 472
rect 1431 607 1497 649
rect 1431 573 1447 607
rect 1481 573 1497 607
rect 1431 530 1497 573
rect 1431 496 1447 530
rect 1481 496 1497 530
rect 1431 455 1497 496
rect 1431 421 1447 455
rect 1481 421 1497 455
rect 1531 599 1569 615
rect 1531 565 1533 599
rect 1567 565 1569 599
rect 1531 506 1569 565
rect 1531 472 1533 506
rect 1567 472 1569 506
rect 467 367 533 375
rect 1359 379 1361 413
rect 1395 385 1397 413
rect 1531 413 1569 472
rect 1603 607 1669 649
rect 1603 573 1619 607
rect 1653 573 1669 607
rect 1603 530 1669 573
rect 1603 496 1619 530
rect 1653 496 1669 530
rect 1603 455 1669 496
rect 1603 421 1619 455
rect 1653 421 1669 455
rect 1703 599 1755 615
rect 1703 565 1705 599
rect 1739 565 1755 599
rect 1703 506 1755 565
rect 1703 472 1705 506
rect 1739 472 1755 506
rect 1531 385 1533 413
rect 1395 379 1533 385
rect 1567 385 1569 413
rect 1703 413 1755 472
rect 1703 385 1705 413
rect 1567 379 1705 385
rect 1739 379 1755 413
rect 295 333 1012 367
rect 144 263 170 297
rect 204 263 238 297
rect 272 263 306 297
rect 340 263 374 297
rect 408 263 442 297
rect 476 263 510 297
rect 544 263 560 297
rect 602 263 618 297
rect 652 263 686 297
rect 720 263 754 297
rect 788 263 822 297
rect 856 263 890 297
rect 924 263 940 297
rect 144 231 185 263
rect 777 242 940 263
rect 21 203 185 231
rect 974 237 1012 333
rect 1046 319 1325 367
rect 1359 339 1755 379
rect 1046 285 1062 319
rect 1096 285 1130 319
rect 1164 285 1198 319
rect 1232 285 1266 319
rect 1300 285 1325 319
rect 1046 271 1325 285
rect 1392 271 1408 305
rect 1442 271 1476 305
rect 1510 271 1544 305
rect 1578 271 1612 305
rect 1646 271 1680 305
rect 1714 271 1748 305
rect 1782 271 1806 305
rect 1547 242 1806 271
rect 21 169 37 203
rect 71 197 185 203
rect 219 208 681 229
rect 974 208 1485 237
rect 219 203 1647 208
rect 71 169 73 197
rect 21 101 73 169
rect 253 193 401 203
rect 253 169 259 193
rect 21 67 37 101
rect 71 67 73 101
rect 21 51 73 67
rect 107 129 123 163
rect 157 129 173 163
rect 107 89 173 129
rect 107 55 123 89
rect 157 55 173 89
rect 107 17 173 55
rect 219 101 259 169
rect 393 169 401 193
rect 435 193 643 203
rect 435 169 437 193
rect 253 67 259 101
rect 219 51 259 67
rect 293 125 309 159
rect 343 125 359 159
rect 293 89 359 125
rect 293 55 309 89
rect 343 55 359 89
rect 293 17 359 55
rect 393 101 437 169
rect 641 169 643 193
rect 677 201 1259 203
rect 677 198 1123 201
rect 677 186 1087 198
rect 677 169 815 186
rect 641 168 815 169
rect 393 67 401 101
rect 435 67 437 101
rect 393 51 437 67
rect 471 123 487 157
rect 521 123 557 157
rect 591 123 607 157
rect 471 89 607 123
rect 471 55 487 89
rect 521 55 557 89
rect 591 55 607 89
rect 471 17 607 55
rect 641 101 679 168
rect 813 152 815 168
rect 849 168 1087 186
rect 849 152 851 168
rect 641 67 643 101
rect 677 67 679 101
rect 641 51 679 67
rect 713 127 779 134
rect 713 93 729 127
rect 763 93 779 127
rect 713 17 779 93
rect 813 101 851 152
rect 1085 164 1087 168
rect 1121 164 1123 198
rect 1257 169 1259 201
rect 1293 201 1435 203
rect 1293 169 1295 201
rect 813 67 815 101
rect 849 67 851 101
rect 813 51 851 67
rect 885 123 1051 134
rect 885 89 901 123
rect 935 89 1001 123
rect 1035 89 1051 123
rect 885 17 1051 89
rect 1085 101 1123 164
rect 1085 67 1087 101
rect 1121 67 1123 101
rect 1085 51 1123 67
rect 1157 133 1173 167
rect 1207 133 1223 167
rect 1157 93 1223 133
rect 1157 59 1173 93
rect 1207 59 1223 93
rect 1157 17 1223 59
rect 1257 101 1295 169
rect 1429 169 1435 201
rect 1469 192 1647 203
rect 1469 174 1611 192
rect 1469 169 1475 174
rect 1257 67 1259 101
rect 1293 67 1295 101
rect 1257 51 1295 67
rect 1329 133 1345 167
rect 1379 133 1395 167
rect 1329 93 1395 133
rect 1329 59 1345 93
rect 1379 59 1395 93
rect 1329 17 1395 59
rect 1429 101 1475 169
rect 1609 158 1611 174
rect 1645 158 1647 192
rect 1429 67 1435 101
rect 1469 67 1475 101
rect 1429 51 1475 67
rect 1509 124 1575 140
rect 1509 90 1525 124
rect 1559 90 1575 124
rect 1509 17 1575 90
rect 1609 101 1647 158
rect 1609 67 1611 101
rect 1645 67 1647 101
rect 1609 51 1647 67
rect 1681 203 1747 208
rect 1681 169 1697 203
rect 1731 169 1747 203
rect 1681 93 1747 169
rect 1681 59 1697 93
rect 1731 59 1747 93
rect 1681 17 1747 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4b_4
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 991 168 1025 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1809128
string GDS_START 1793346
<< end >>
