magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
<< pwell >>
rect 549 243 1219 259
rect 11 49 1219 243
rect 0 0 1248 49
<< scnmos >>
rect 94 49 124 217
rect 180 49 210 217
rect 266 49 296 217
rect 352 49 382 217
rect 438 49 468 217
rect 644 65 674 233
rect 730 65 760 233
rect 832 65 862 233
rect 934 65 964 233
rect 1020 65 1050 233
rect 1106 65 1136 233
<< scpmoshvt >>
rect 102 367 132 619
rect 188 367 218 619
rect 274 367 304 619
rect 361 367 391 619
rect 447 367 477 619
rect 608 367 638 619
rect 694 367 724 619
rect 848 367 878 619
rect 934 367 964 619
rect 1020 367 1050 619
rect 1106 367 1136 619
<< ndiff >>
rect 37 190 94 217
rect 37 156 45 190
rect 79 156 94 190
rect 37 101 94 156
rect 37 67 45 101
rect 79 67 94 101
rect 37 49 94 67
rect 124 190 180 217
rect 124 156 135 190
rect 169 156 180 190
rect 124 95 180 156
rect 124 61 135 95
rect 169 61 180 95
rect 124 49 180 61
rect 210 205 266 217
rect 210 171 221 205
rect 255 171 266 205
rect 210 101 266 171
rect 210 67 221 101
rect 255 67 266 101
rect 210 49 266 67
rect 296 181 352 217
rect 296 147 307 181
rect 341 147 352 181
rect 296 95 352 147
rect 296 61 307 95
rect 341 61 352 95
rect 296 49 352 61
rect 382 205 438 217
rect 382 171 393 205
rect 427 171 438 205
rect 382 101 438 171
rect 382 67 393 101
rect 427 67 438 101
rect 382 49 438 67
rect 468 181 521 217
rect 468 147 479 181
rect 513 147 521 181
rect 468 95 521 147
rect 468 61 479 95
rect 513 61 521 95
rect 575 179 644 233
rect 575 145 585 179
rect 619 145 644 179
rect 575 111 644 145
rect 575 77 585 111
rect 619 77 644 111
rect 575 65 644 77
rect 674 225 730 233
rect 674 191 685 225
rect 719 191 730 225
rect 674 155 730 191
rect 674 121 685 155
rect 719 121 730 155
rect 674 65 730 121
rect 760 179 832 233
rect 760 145 787 179
rect 821 145 832 179
rect 760 107 832 145
rect 760 73 787 107
rect 821 73 832 107
rect 760 65 832 73
rect 862 107 934 233
rect 862 73 887 107
rect 921 73 934 107
rect 862 65 934 73
rect 964 221 1020 233
rect 964 187 975 221
rect 1009 187 1020 221
rect 964 109 1020 187
rect 964 75 975 109
rect 1009 75 1020 109
rect 964 65 1020 75
rect 1050 181 1106 233
rect 1050 147 1061 181
rect 1095 147 1106 181
rect 1050 107 1106 147
rect 1050 73 1061 107
rect 1095 73 1106 107
rect 1050 65 1106 73
rect 1136 221 1193 233
rect 1136 187 1151 221
rect 1185 187 1193 221
rect 1136 111 1193 187
rect 1136 77 1151 111
rect 1185 77 1193 111
rect 1136 65 1193 77
rect 468 49 521 61
<< pdiff >>
rect 49 599 102 619
rect 49 565 57 599
rect 91 565 102 599
rect 49 518 102 565
rect 49 484 57 518
rect 91 484 102 518
rect 49 434 102 484
rect 49 400 57 434
rect 91 400 102 434
rect 49 367 102 400
rect 132 596 188 619
rect 132 562 143 596
rect 177 562 188 596
rect 132 367 188 562
rect 218 436 274 619
rect 218 402 229 436
rect 263 402 274 436
rect 218 367 274 402
rect 304 596 361 619
rect 304 562 315 596
rect 349 562 361 596
rect 304 367 361 562
rect 391 436 447 619
rect 391 402 402 436
rect 436 402 447 436
rect 391 367 447 402
rect 477 611 608 619
rect 477 606 563 611
rect 477 572 488 606
rect 522 577 563 606
rect 597 577 608 611
rect 522 572 608 577
rect 477 543 608 572
rect 477 509 563 543
rect 597 509 608 543
rect 477 473 608 509
rect 477 439 563 473
rect 597 439 608 473
rect 477 367 608 439
rect 638 599 694 619
rect 638 565 649 599
rect 683 565 694 599
rect 638 509 694 565
rect 638 475 649 509
rect 683 475 694 509
rect 638 413 694 475
rect 638 379 649 413
rect 683 379 694 413
rect 638 367 694 379
rect 724 607 848 619
rect 724 573 735 607
rect 769 573 803 607
rect 837 573 848 607
rect 724 506 848 573
rect 724 472 735 506
rect 769 472 848 506
rect 724 413 848 472
rect 724 379 735 413
rect 769 379 848 413
rect 724 367 848 379
rect 878 584 934 619
rect 878 550 889 584
rect 923 550 934 584
rect 878 367 934 550
rect 964 424 1020 619
rect 964 390 975 424
rect 1009 390 1020 424
rect 964 367 1020 390
rect 1050 584 1106 619
rect 1050 550 1061 584
rect 1095 550 1106 584
rect 1050 367 1106 550
rect 1136 607 1199 619
rect 1136 573 1155 607
rect 1189 573 1199 607
rect 1136 509 1199 573
rect 1136 475 1155 509
rect 1189 475 1199 509
rect 1136 413 1199 475
rect 1136 379 1155 413
rect 1189 379 1199 413
rect 1136 367 1199 379
<< ndiffc >>
rect 45 156 79 190
rect 45 67 79 101
rect 135 156 169 190
rect 135 61 169 95
rect 221 171 255 205
rect 221 67 255 101
rect 307 147 341 181
rect 307 61 341 95
rect 393 171 427 205
rect 393 67 427 101
rect 479 147 513 181
rect 479 61 513 95
rect 585 145 619 179
rect 585 77 619 111
rect 685 191 719 225
rect 685 121 719 155
rect 787 145 821 179
rect 787 73 821 107
rect 887 73 921 107
rect 975 187 1009 221
rect 975 75 1009 109
rect 1061 147 1095 181
rect 1061 73 1095 107
rect 1151 187 1185 221
rect 1151 77 1185 111
<< pdiffc >>
rect 57 565 91 599
rect 57 484 91 518
rect 57 400 91 434
rect 143 562 177 596
rect 229 402 263 436
rect 315 562 349 596
rect 402 402 436 436
rect 488 572 522 606
rect 563 577 597 611
rect 563 509 597 543
rect 563 439 597 473
rect 649 565 683 599
rect 649 475 683 509
rect 649 379 683 413
rect 735 573 769 607
rect 803 573 837 607
rect 735 472 769 506
rect 735 379 769 413
rect 889 550 923 584
rect 975 390 1009 424
rect 1061 550 1095 584
rect 1155 573 1189 607
rect 1155 475 1189 509
rect 1155 379 1189 413
<< poly >>
rect 102 619 132 645
rect 188 619 218 645
rect 274 619 304 645
rect 361 619 391 645
rect 447 619 477 645
rect 608 619 638 645
rect 694 619 724 645
rect 848 619 878 645
rect 934 619 964 645
rect 1020 619 1050 645
rect 1106 619 1136 645
rect 102 308 132 367
rect 188 335 218 367
rect 274 335 304 367
rect 361 335 391 367
rect 447 335 477 367
rect 608 335 638 367
rect 694 335 724 367
rect 848 335 878 367
rect 188 319 477 335
rect 72 292 138 308
rect 188 299 291 319
rect 72 258 88 292
rect 122 258 138 292
rect 72 242 138 258
rect 180 285 291 299
rect 325 285 359 319
rect 393 285 427 319
rect 461 285 477 319
rect 180 269 477 285
rect 536 319 760 335
rect 536 285 552 319
rect 586 305 760 319
rect 586 285 602 305
rect 536 269 602 285
rect 94 217 124 242
rect 180 217 210 269
rect 266 217 296 269
rect 352 217 382 269
rect 438 217 468 269
rect 644 233 674 305
rect 730 233 760 305
rect 803 319 878 335
rect 803 285 819 319
rect 853 285 878 319
rect 803 269 878 285
rect 934 335 964 367
rect 1020 335 1050 367
rect 934 319 1050 335
rect 934 285 1000 319
rect 1034 285 1050 319
rect 934 269 1050 285
rect 832 233 862 269
rect 934 233 964 269
rect 1020 233 1050 269
rect 1106 335 1136 367
rect 1106 319 1172 335
rect 1106 285 1122 319
rect 1156 285 1172 319
rect 1106 269 1172 285
rect 1106 233 1136 269
rect 94 23 124 49
rect 180 23 210 49
rect 266 23 296 49
rect 352 23 382 49
rect 438 23 468 49
rect 644 39 674 65
rect 730 39 760 65
rect 832 39 862 65
rect 934 39 964 65
rect 1020 39 1050 65
rect 1106 39 1136 65
<< polycont >>
rect 88 258 122 292
rect 291 285 325 319
rect 359 285 393 319
rect 427 285 461 319
rect 552 285 586 319
rect 819 285 853 319
rect 1000 285 1034 319
rect 1122 285 1156 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 17 599 93 615
rect 17 565 57 599
rect 91 565 93 599
rect 17 522 93 565
rect 127 596 193 649
rect 127 562 143 596
rect 177 562 193 596
rect 127 556 193 562
rect 299 596 365 649
rect 299 562 315 596
rect 349 562 365 596
rect 299 556 365 562
rect 472 611 607 649
rect 472 606 563 611
rect 472 572 488 606
rect 522 577 563 606
rect 597 577 607 611
rect 522 572 607 577
rect 472 556 607 572
rect 553 543 607 556
rect 17 518 519 522
rect 17 484 57 518
rect 91 486 519 518
rect 17 434 91 484
rect 17 400 57 434
rect 17 384 91 400
rect 125 436 451 452
rect 125 402 229 436
rect 263 402 402 436
rect 436 402 451 436
rect 125 386 451 402
rect 485 389 519 486
rect 553 509 563 543
rect 597 509 607 543
rect 553 473 607 509
rect 553 439 563 473
rect 597 439 607 473
rect 553 423 607 439
rect 641 599 685 615
rect 641 565 649 599
rect 683 565 685 599
rect 641 509 685 565
rect 641 475 649 509
rect 683 475 685 509
rect 641 413 685 475
rect 125 384 241 386
rect 17 206 52 384
rect 86 292 173 350
rect 86 258 88 292
rect 122 258 173 292
rect 86 240 173 258
rect 207 249 241 384
rect 485 355 602 389
rect 275 319 497 321
rect 275 285 291 319
rect 325 285 359 319
rect 393 285 427 319
rect 461 285 497 319
rect 275 283 497 285
rect 536 319 602 355
rect 536 285 552 319
rect 586 285 602 319
rect 536 283 602 285
rect 641 379 649 413
rect 683 379 685 413
rect 463 249 497 283
rect 641 249 685 379
rect 719 607 853 649
rect 719 573 735 607
rect 769 573 803 607
rect 837 573 853 607
rect 1155 607 1205 649
rect 719 557 853 573
rect 887 584 1099 600
rect 719 506 781 557
rect 887 550 889 584
rect 923 550 1061 584
rect 1095 550 1099 584
rect 887 534 1099 550
rect 1189 573 1205 607
rect 719 472 735 506
rect 769 472 781 506
rect 1155 509 1205 573
rect 719 413 781 472
rect 719 379 735 413
rect 769 379 781 413
rect 719 363 781 379
rect 815 462 1121 500
rect 815 335 869 462
rect 803 319 869 335
rect 803 285 819 319
rect 853 285 869 319
rect 803 283 869 285
rect 905 424 1025 428
rect 905 390 975 424
rect 1009 390 1025 424
rect 905 386 1025 390
rect 905 249 939 386
rect 984 319 1050 352
rect 984 285 1000 319
rect 1034 285 1050 319
rect 984 283 1050 285
rect 1087 329 1121 462
rect 1189 475 1205 509
rect 1155 413 1205 475
rect 1189 379 1205 413
rect 1155 363 1205 379
rect 1087 319 1172 329
rect 1087 285 1122 319
rect 1156 285 1172 319
rect 1087 283 1172 285
rect 207 215 429 249
rect 463 225 939 249
rect 463 215 685 225
rect 17 190 85 206
rect 17 156 45 190
rect 79 156 85 190
rect 17 101 85 156
rect 17 67 45 101
rect 79 67 85 101
rect 17 51 85 67
rect 119 190 173 206
rect 119 156 135 190
rect 169 156 173 190
rect 119 95 173 156
rect 119 61 135 95
rect 169 61 173 95
rect 119 17 173 61
rect 207 205 257 215
rect 207 171 221 205
rect 255 171 257 205
rect 391 205 429 215
rect 207 101 257 171
rect 207 67 221 101
rect 255 67 257 101
rect 207 51 257 67
rect 291 147 307 181
rect 341 147 357 181
rect 291 95 357 147
rect 291 61 307 95
rect 341 61 357 95
rect 291 17 357 61
rect 391 171 393 205
rect 427 171 429 205
rect 669 191 685 215
rect 719 215 939 225
rect 973 221 1201 249
rect 719 191 735 215
rect 391 101 429 171
rect 391 67 393 101
rect 427 67 429 101
rect 391 51 429 67
rect 463 147 479 181
rect 513 147 529 181
rect 463 95 529 147
rect 463 61 479 95
rect 513 61 529 95
rect 463 17 529 61
rect 567 179 635 181
rect 567 145 585 179
rect 619 145 635 179
rect 567 111 635 145
rect 669 155 735 191
rect 973 187 975 221
rect 1009 215 1151 221
rect 1009 187 1011 215
rect 973 179 1011 187
rect 1147 187 1151 215
rect 1185 187 1201 221
rect 669 121 685 155
rect 719 121 735 155
rect 771 145 787 179
rect 821 145 1011 179
rect 567 77 585 111
rect 619 87 635 111
rect 771 107 837 145
rect 771 87 787 107
rect 619 77 787 87
rect 567 73 787 77
rect 821 73 837 107
rect 567 53 837 73
rect 871 107 939 111
rect 871 73 887 107
rect 921 73 939 107
rect 871 17 939 73
rect 973 109 1011 145
rect 973 75 975 109
rect 1009 75 1011 109
rect 973 59 1011 75
rect 1045 147 1061 181
rect 1095 147 1111 181
rect 1045 107 1111 147
rect 1045 73 1061 107
rect 1095 73 1111 107
rect 1045 17 1111 73
rect 1147 111 1201 187
rect 1147 77 1151 111
rect 1185 77 1201 111
rect 1147 61 1201 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21ba_4
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 895 464 929 498 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 464 1025 498 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 464 1121 498 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6510724
string GDS_START 6500230
<< end >>
