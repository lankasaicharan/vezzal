magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3794 1975
<< nwell >>
rect -38 331 2534 704
<< pwell >>
rect 1 241 447 243
rect 1 49 2495 241
rect 0 0 2496 49
<< scnmos >>
rect 80 49 110 217
rect 166 49 196 217
rect 252 49 282 217
rect 338 49 368 217
rect 580 47 610 215
rect 666 47 696 215
rect 752 47 782 215
rect 838 47 868 215
rect 924 47 954 215
rect 1010 47 1040 215
rect 1096 47 1126 215
rect 1182 47 1212 215
rect 1268 47 1298 215
rect 1354 47 1384 215
rect 1440 47 1470 215
rect 1526 47 1556 215
rect 1612 47 1642 215
rect 1698 47 1728 215
rect 1784 47 1814 215
rect 1870 47 1900 215
rect 1956 47 1986 215
rect 2042 47 2072 215
rect 2128 47 2158 215
rect 2214 47 2244 215
rect 2300 47 2330 215
rect 2386 47 2416 215
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 252 367 282 619
rect 338 367 368 619
rect 580 367 610 619
rect 666 367 696 619
rect 752 367 782 619
rect 838 367 868 619
rect 924 367 954 619
rect 1010 367 1040 619
rect 1096 367 1126 619
rect 1182 367 1212 619
rect 1268 367 1298 619
rect 1354 367 1384 619
rect 1440 367 1470 619
rect 1526 367 1556 619
rect 1612 367 1642 619
rect 1698 367 1728 619
rect 1784 367 1814 619
rect 1870 367 1900 619
rect 1956 367 1986 619
rect 2042 367 2072 619
rect 2128 367 2158 619
rect 2214 367 2244 619
rect 2300 367 2330 619
rect 2386 367 2416 619
<< ndiff >>
rect 27 185 80 217
rect 27 151 35 185
rect 69 151 80 185
rect 27 101 80 151
rect 27 67 35 101
rect 69 67 80 101
rect 27 49 80 67
rect 110 163 166 217
rect 110 129 121 163
rect 155 129 166 163
rect 110 95 166 129
rect 110 61 121 95
rect 155 61 166 95
rect 110 49 166 61
rect 196 184 252 217
rect 196 150 207 184
rect 241 150 252 184
rect 196 101 252 150
rect 196 67 207 101
rect 241 67 252 101
rect 196 49 252 67
rect 282 170 338 217
rect 282 136 293 170
rect 327 136 338 170
rect 282 102 338 136
rect 282 68 293 102
rect 327 68 338 102
rect 282 49 338 68
rect 368 184 421 217
rect 368 150 379 184
rect 413 150 421 184
rect 368 101 421 150
rect 368 67 379 101
rect 413 67 421 101
rect 368 49 421 67
rect 527 163 580 215
rect 527 129 535 163
rect 569 129 580 163
rect 527 95 580 129
rect 527 61 535 95
rect 569 61 580 95
rect 527 47 580 61
rect 610 189 666 215
rect 610 155 621 189
rect 655 155 666 189
rect 610 107 666 155
rect 610 73 621 107
rect 655 73 666 107
rect 610 47 666 73
rect 696 159 752 215
rect 696 125 707 159
rect 741 125 752 159
rect 696 91 752 125
rect 696 57 707 91
rect 741 57 752 91
rect 696 47 752 57
rect 782 189 838 215
rect 782 155 793 189
rect 827 155 838 189
rect 782 107 838 155
rect 782 73 793 107
rect 827 73 838 107
rect 782 47 838 73
rect 868 159 924 215
rect 868 125 879 159
rect 913 125 924 159
rect 868 91 924 125
rect 868 57 879 91
rect 913 57 924 91
rect 868 47 924 57
rect 954 189 1010 215
rect 954 155 965 189
rect 999 155 1010 189
rect 954 107 1010 155
rect 954 73 965 107
rect 999 73 1010 107
rect 954 47 1010 73
rect 1040 159 1096 215
rect 1040 125 1051 159
rect 1085 125 1096 159
rect 1040 91 1096 125
rect 1040 57 1051 91
rect 1085 57 1096 91
rect 1040 47 1096 57
rect 1126 189 1182 215
rect 1126 155 1137 189
rect 1171 155 1182 189
rect 1126 107 1182 155
rect 1126 73 1137 107
rect 1171 73 1182 107
rect 1126 47 1182 73
rect 1212 189 1268 215
rect 1212 155 1223 189
rect 1257 155 1268 189
rect 1212 107 1268 155
rect 1212 73 1223 107
rect 1257 73 1268 107
rect 1212 47 1268 73
rect 1298 189 1354 215
rect 1298 155 1309 189
rect 1343 155 1354 189
rect 1298 107 1354 155
rect 1298 73 1309 107
rect 1343 73 1354 107
rect 1298 47 1354 73
rect 1384 189 1440 215
rect 1384 155 1395 189
rect 1429 155 1440 189
rect 1384 107 1440 155
rect 1384 73 1395 107
rect 1429 73 1440 107
rect 1384 47 1440 73
rect 1470 189 1526 215
rect 1470 155 1481 189
rect 1515 155 1526 189
rect 1470 107 1526 155
rect 1470 73 1481 107
rect 1515 73 1526 107
rect 1470 47 1526 73
rect 1556 189 1612 215
rect 1556 155 1567 189
rect 1601 155 1612 189
rect 1556 107 1612 155
rect 1556 73 1567 107
rect 1601 73 1612 107
rect 1556 47 1612 73
rect 1642 189 1698 215
rect 1642 155 1653 189
rect 1687 155 1698 189
rect 1642 107 1698 155
rect 1642 73 1653 107
rect 1687 73 1698 107
rect 1642 47 1698 73
rect 1728 189 1784 215
rect 1728 155 1739 189
rect 1773 155 1784 189
rect 1728 107 1784 155
rect 1728 73 1739 107
rect 1773 73 1784 107
rect 1728 47 1784 73
rect 1814 189 1870 215
rect 1814 155 1825 189
rect 1859 155 1870 189
rect 1814 107 1870 155
rect 1814 73 1825 107
rect 1859 73 1870 107
rect 1814 47 1870 73
rect 1900 189 1956 215
rect 1900 155 1911 189
rect 1945 155 1956 189
rect 1900 107 1956 155
rect 1900 73 1911 107
rect 1945 73 1956 107
rect 1900 47 1956 73
rect 1986 189 2042 215
rect 1986 155 1997 189
rect 2031 155 2042 189
rect 1986 107 2042 155
rect 1986 73 1997 107
rect 2031 73 2042 107
rect 1986 47 2042 73
rect 2072 189 2128 215
rect 2072 155 2083 189
rect 2117 155 2128 189
rect 2072 107 2128 155
rect 2072 73 2083 107
rect 2117 73 2128 107
rect 2072 47 2128 73
rect 2158 189 2214 215
rect 2158 155 2169 189
rect 2203 155 2214 189
rect 2158 107 2214 155
rect 2158 73 2169 107
rect 2203 73 2214 107
rect 2158 47 2214 73
rect 2244 189 2300 215
rect 2244 155 2255 189
rect 2289 155 2300 189
rect 2244 107 2300 155
rect 2244 73 2255 107
rect 2289 73 2300 107
rect 2244 47 2300 73
rect 2330 189 2386 215
rect 2330 155 2341 189
rect 2375 155 2386 189
rect 2330 107 2386 155
rect 2330 73 2341 107
rect 2375 73 2386 107
rect 2330 47 2386 73
rect 2416 189 2469 215
rect 2416 155 2427 189
rect 2461 155 2469 189
rect 2416 107 2469 155
rect 2416 73 2427 107
rect 2461 73 2469 107
rect 2416 47 2469 73
<< pdiff >>
rect 27 590 80 619
rect 27 556 35 590
rect 69 556 80 590
rect 27 511 80 556
rect 27 477 35 511
rect 69 477 80 511
rect 27 434 80 477
rect 27 400 35 434
rect 69 400 80 434
rect 27 367 80 400
rect 110 570 166 619
rect 110 536 121 570
rect 155 536 166 570
rect 110 502 166 536
rect 110 468 121 502
rect 155 468 166 502
rect 110 367 166 468
rect 196 590 252 619
rect 196 556 207 590
rect 241 556 252 590
rect 196 506 252 556
rect 196 472 207 506
rect 241 472 252 506
rect 196 422 252 472
rect 196 388 207 422
rect 241 388 252 422
rect 196 367 252 388
rect 282 603 338 619
rect 282 569 293 603
rect 327 569 338 603
rect 282 535 338 569
rect 282 501 293 535
rect 327 501 338 535
rect 282 467 338 501
rect 282 433 293 467
rect 327 433 338 467
rect 282 367 338 433
rect 368 590 421 619
rect 368 556 379 590
rect 413 556 421 590
rect 368 506 421 556
rect 368 472 379 506
rect 413 472 421 506
rect 368 422 421 472
rect 368 388 379 422
rect 413 388 421 422
rect 368 367 421 388
rect 527 598 580 619
rect 527 564 535 598
rect 569 564 580 598
rect 527 530 580 564
rect 527 496 535 530
rect 569 496 580 530
rect 527 462 580 496
rect 527 428 535 462
rect 569 428 580 462
rect 527 367 580 428
rect 610 594 666 619
rect 610 560 621 594
rect 655 560 666 594
rect 610 510 666 560
rect 610 476 621 510
rect 655 476 666 510
rect 610 426 666 476
rect 610 392 621 426
rect 655 392 666 426
rect 610 367 666 392
rect 696 605 752 619
rect 696 571 707 605
rect 741 571 752 605
rect 696 537 752 571
rect 696 503 707 537
rect 741 503 752 537
rect 696 469 752 503
rect 696 435 707 469
rect 741 435 752 469
rect 696 367 752 435
rect 782 594 838 619
rect 782 560 793 594
rect 827 560 838 594
rect 782 510 838 560
rect 782 476 793 510
rect 827 476 838 510
rect 782 426 838 476
rect 782 392 793 426
rect 827 392 838 426
rect 782 367 838 392
rect 868 605 924 619
rect 868 571 879 605
rect 913 571 924 605
rect 868 537 924 571
rect 868 503 879 537
rect 913 503 924 537
rect 868 469 924 503
rect 868 435 879 469
rect 913 435 924 469
rect 868 367 924 435
rect 954 594 1010 619
rect 954 560 965 594
rect 999 560 1010 594
rect 954 510 1010 560
rect 954 476 965 510
rect 999 476 1010 510
rect 954 426 1010 476
rect 954 392 965 426
rect 999 392 1010 426
rect 954 367 1010 392
rect 1040 605 1096 619
rect 1040 571 1051 605
rect 1085 571 1096 605
rect 1040 537 1096 571
rect 1040 503 1051 537
rect 1085 503 1096 537
rect 1040 469 1096 503
rect 1040 435 1051 469
rect 1085 435 1096 469
rect 1040 367 1096 435
rect 1126 594 1182 619
rect 1126 560 1137 594
rect 1171 560 1182 594
rect 1126 510 1182 560
rect 1126 476 1137 510
rect 1171 476 1182 510
rect 1126 426 1182 476
rect 1126 392 1137 426
rect 1171 392 1182 426
rect 1126 367 1182 392
rect 1212 598 1268 619
rect 1212 564 1223 598
rect 1257 564 1268 598
rect 1212 516 1268 564
rect 1212 482 1223 516
rect 1257 482 1268 516
rect 1212 435 1268 482
rect 1212 401 1223 435
rect 1257 401 1268 435
rect 1212 367 1268 401
rect 1298 594 1354 619
rect 1298 560 1309 594
rect 1343 560 1354 594
rect 1298 510 1354 560
rect 1298 476 1309 510
rect 1343 476 1354 510
rect 1298 426 1354 476
rect 1298 392 1309 426
rect 1343 392 1354 426
rect 1298 367 1354 392
rect 1384 598 1440 619
rect 1384 564 1395 598
rect 1429 564 1440 598
rect 1384 516 1440 564
rect 1384 482 1395 516
rect 1429 482 1440 516
rect 1384 435 1440 482
rect 1384 401 1395 435
rect 1429 401 1440 435
rect 1384 367 1440 401
rect 1470 594 1526 619
rect 1470 560 1481 594
rect 1515 560 1526 594
rect 1470 510 1526 560
rect 1470 476 1481 510
rect 1515 476 1526 510
rect 1470 426 1526 476
rect 1470 392 1481 426
rect 1515 392 1526 426
rect 1470 367 1526 392
rect 1556 598 1612 619
rect 1556 564 1567 598
rect 1601 564 1612 598
rect 1556 516 1612 564
rect 1556 482 1567 516
rect 1601 482 1612 516
rect 1556 435 1612 482
rect 1556 401 1567 435
rect 1601 401 1612 435
rect 1556 367 1612 401
rect 1642 594 1698 619
rect 1642 560 1653 594
rect 1687 560 1698 594
rect 1642 510 1698 560
rect 1642 476 1653 510
rect 1687 476 1698 510
rect 1642 426 1698 476
rect 1642 392 1653 426
rect 1687 392 1698 426
rect 1642 367 1698 392
rect 1728 598 1784 619
rect 1728 564 1739 598
rect 1773 564 1784 598
rect 1728 516 1784 564
rect 1728 482 1739 516
rect 1773 482 1784 516
rect 1728 435 1784 482
rect 1728 401 1739 435
rect 1773 401 1784 435
rect 1728 367 1784 401
rect 1814 594 1870 619
rect 1814 560 1825 594
rect 1859 560 1870 594
rect 1814 510 1870 560
rect 1814 476 1825 510
rect 1859 476 1870 510
rect 1814 426 1870 476
rect 1814 392 1825 426
rect 1859 392 1870 426
rect 1814 367 1870 392
rect 1900 598 1956 619
rect 1900 564 1911 598
rect 1945 564 1956 598
rect 1900 516 1956 564
rect 1900 482 1911 516
rect 1945 482 1956 516
rect 1900 435 1956 482
rect 1900 401 1911 435
rect 1945 401 1956 435
rect 1900 367 1956 401
rect 1986 594 2042 619
rect 1986 560 1997 594
rect 2031 560 2042 594
rect 1986 510 2042 560
rect 1986 476 1997 510
rect 2031 476 2042 510
rect 1986 426 2042 476
rect 1986 392 1997 426
rect 2031 392 2042 426
rect 1986 367 2042 392
rect 2072 598 2128 619
rect 2072 564 2083 598
rect 2117 564 2128 598
rect 2072 516 2128 564
rect 2072 482 2083 516
rect 2117 482 2128 516
rect 2072 435 2128 482
rect 2072 401 2083 435
rect 2117 401 2128 435
rect 2072 367 2128 401
rect 2158 594 2214 619
rect 2158 560 2169 594
rect 2203 560 2214 594
rect 2158 510 2214 560
rect 2158 476 2169 510
rect 2203 476 2214 510
rect 2158 426 2214 476
rect 2158 392 2169 426
rect 2203 392 2214 426
rect 2158 367 2214 392
rect 2244 598 2300 619
rect 2244 564 2255 598
rect 2289 564 2300 598
rect 2244 516 2300 564
rect 2244 482 2255 516
rect 2289 482 2300 516
rect 2244 435 2300 482
rect 2244 401 2255 435
rect 2289 401 2300 435
rect 2244 367 2300 401
rect 2330 594 2386 619
rect 2330 560 2341 594
rect 2375 560 2386 594
rect 2330 510 2386 560
rect 2330 476 2341 510
rect 2375 476 2386 510
rect 2330 426 2386 476
rect 2330 392 2341 426
rect 2375 392 2386 426
rect 2330 367 2386 392
rect 2416 598 2469 619
rect 2416 564 2427 598
rect 2461 564 2469 598
rect 2416 516 2469 564
rect 2416 482 2427 516
rect 2461 482 2469 516
rect 2416 435 2469 482
rect 2416 401 2427 435
rect 2461 401 2469 435
rect 2416 367 2469 401
<< ndiffc >>
rect 35 151 69 185
rect 35 67 69 101
rect 121 129 155 163
rect 121 61 155 95
rect 207 150 241 184
rect 207 67 241 101
rect 293 136 327 170
rect 293 68 327 102
rect 379 150 413 184
rect 379 67 413 101
rect 535 129 569 163
rect 535 61 569 95
rect 621 155 655 189
rect 621 73 655 107
rect 707 125 741 159
rect 707 57 741 91
rect 793 155 827 189
rect 793 73 827 107
rect 879 125 913 159
rect 879 57 913 91
rect 965 155 999 189
rect 965 73 999 107
rect 1051 125 1085 159
rect 1051 57 1085 91
rect 1137 155 1171 189
rect 1137 73 1171 107
rect 1223 155 1257 189
rect 1223 73 1257 107
rect 1309 155 1343 189
rect 1309 73 1343 107
rect 1395 155 1429 189
rect 1395 73 1429 107
rect 1481 155 1515 189
rect 1481 73 1515 107
rect 1567 155 1601 189
rect 1567 73 1601 107
rect 1653 155 1687 189
rect 1653 73 1687 107
rect 1739 155 1773 189
rect 1739 73 1773 107
rect 1825 155 1859 189
rect 1825 73 1859 107
rect 1911 155 1945 189
rect 1911 73 1945 107
rect 1997 155 2031 189
rect 1997 73 2031 107
rect 2083 155 2117 189
rect 2083 73 2117 107
rect 2169 155 2203 189
rect 2169 73 2203 107
rect 2255 155 2289 189
rect 2255 73 2289 107
rect 2341 155 2375 189
rect 2341 73 2375 107
rect 2427 155 2461 189
rect 2427 73 2461 107
<< pdiffc >>
rect 35 556 69 590
rect 35 477 69 511
rect 35 400 69 434
rect 121 536 155 570
rect 121 468 155 502
rect 207 556 241 590
rect 207 472 241 506
rect 207 388 241 422
rect 293 569 327 603
rect 293 501 327 535
rect 293 433 327 467
rect 379 556 413 590
rect 379 472 413 506
rect 379 388 413 422
rect 535 564 569 598
rect 535 496 569 530
rect 535 428 569 462
rect 621 560 655 594
rect 621 476 655 510
rect 621 392 655 426
rect 707 571 741 605
rect 707 503 741 537
rect 707 435 741 469
rect 793 560 827 594
rect 793 476 827 510
rect 793 392 827 426
rect 879 571 913 605
rect 879 503 913 537
rect 879 435 913 469
rect 965 560 999 594
rect 965 476 999 510
rect 965 392 999 426
rect 1051 571 1085 605
rect 1051 503 1085 537
rect 1051 435 1085 469
rect 1137 560 1171 594
rect 1137 476 1171 510
rect 1137 392 1171 426
rect 1223 564 1257 598
rect 1223 482 1257 516
rect 1223 401 1257 435
rect 1309 560 1343 594
rect 1309 476 1343 510
rect 1309 392 1343 426
rect 1395 564 1429 598
rect 1395 482 1429 516
rect 1395 401 1429 435
rect 1481 560 1515 594
rect 1481 476 1515 510
rect 1481 392 1515 426
rect 1567 564 1601 598
rect 1567 482 1601 516
rect 1567 401 1601 435
rect 1653 560 1687 594
rect 1653 476 1687 510
rect 1653 392 1687 426
rect 1739 564 1773 598
rect 1739 482 1773 516
rect 1739 401 1773 435
rect 1825 560 1859 594
rect 1825 476 1859 510
rect 1825 392 1859 426
rect 1911 564 1945 598
rect 1911 482 1945 516
rect 1911 401 1945 435
rect 1997 560 2031 594
rect 1997 476 2031 510
rect 1997 392 2031 426
rect 2083 564 2117 598
rect 2083 482 2117 516
rect 2083 401 2117 435
rect 2169 560 2203 594
rect 2169 476 2203 510
rect 2169 392 2203 426
rect 2255 564 2289 598
rect 2255 482 2289 516
rect 2255 401 2289 435
rect 2341 560 2375 594
rect 2341 476 2375 510
rect 2341 392 2375 426
rect 2427 564 2461 598
rect 2427 482 2461 516
rect 2427 401 2461 435
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 252 619 282 645
rect 338 619 368 645
rect 580 619 610 645
rect 666 619 696 645
rect 752 619 782 645
rect 838 619 868 645
rect 924 619 954 645
rect 1010 619 1040 645
rect 1096 619 1126 645
rect 1182 619 1212 645
rect 1268 619 1298 645
rect 1354 619 1384 645
rect 1440 619 1470 645
rect 1526 619 1556 645
rect 1612 619 1642 645
rect 1698 619 1728 645
rect 1784 619 1814 645
rect 1870 619 1900 645
rect 1956 619 1986 645
rect 2042 619 2072 645
rect 2128 619 2158 645
rect 2214 619 2244 645
rect 2300 619 2330 645
rect 2386 619 2416 645
rect 80 325 110 367
rect 31 309 110 325
rect 31 275 47 309
rect 81 275 110 309
rect 31 259 110 275
rect 80 217 110 259
rect 166 331 196 367
rect 252 331 282 367
rect 338 331 368 367
rect 166 315 436 331
rect 580 329 610 367
rect 666 329 696 367
rect 752 329 782 367
rect 838 329 868 367
rect 924 329 954 367
rect 1010 329 1040 367
rect 166 281 182 315
rect 216 281 250 315
rect 284 281 318 315
rect 352 281 386 315
rect 420 281 436 315
rect 166 265 436 281
rect 553 313 1040 329
rect 553 279 569 313
rect 603 279 637 313
rect 671 279 705 313
rect 739 279 773 313
rect 807 279 841 313
rect 875 279 909 313
rect 943 279 977 313
rect 1011 279 1040 313
rect 166 217 196 265
rect 252 217 282 265
rect 338 217 368 265
rect 553 263 1040 279
rect 580 215 610 263
rect 666 215 696 263
rect 752 215 782 263
rect 838 215 868 263
rect 924 215 954 263
rect 1010 215 1040 263
rect 1096 329 1126 367
rect 1182 329 1212 367
rect 1268 329 1298 367
rect 1354 329 1384 367
rect 1440 329 1470 367
rect 1526 329 1556 367
rect 1612 329 1642 367
rect 1698 329 1728 367
rect 1784 329 1814 367
rect 1870 329 1900 367
rect 1956 329 1986 367
rect 2042 329 2072 367
rect 2128 329 2158 367
rect 2214 329 2244 367
rect 2300 329 2330 367
rect 2386 329 2416 367
rect 1096 313 2416 329
rect 1096 279 1223 313
rect 1257 279 1395 313
rect 1429 279 1567 313
rect 1601 279 1739 313
rect 1773 279 1911 313
rect 1945 279 2083 313
rect 2117 279 2255 313
rect 2289 279 2416 313
rect 1096 263 2416 279
rect 1096 215 1126 263
rect 1182 215 1212 263
rect 1268 215 1298 263
rect 1354 215 1384 263
rect 1440 215 1470 263
rect 1526 215 1556 263
rect 1612 215 1642 263
rect 1698 215 1728 263
rect 1784 215 1814 263
rect 1870 215 1900 263
rect 1956 215 1986 263
rect 2042 215 2072 263
rect 2128 215 2158 263
rect 2214 215 2244 263
rect 2300 215 2330 263
rect 2386 215 2416 263
rect 80 23 110 49
rect 166 23 196 49
rect 252 23 282 49
rect 338 23 368 49
rect 580 21 610 47
rect 666 21 696 47
rect 752 21 782 47
rect 838 21 868 47
rect 924 21 954 47
rect 1010 21 1040 47
rect 1096 21 1126 47
rect 1182 21 1212 47
rect 1268 21 1298 47
rect 1354 21 1384 47
rect 1440 21 1470 47
rect 1526 21 1556 47
rect 1612 21 1642 47
rect 1698 21 1728 47
rect 1784 21 1814 47
rect 1870 21 1900 47
rect 1956 21 1986 47
rect 2042 21 2072 47
rect 2128 21 2158 47
rect 2214 21 2244 47
rect 2300 21 2330 47
rect 2386 21 2416 47
<< polycont >>
rect 47 275 81 309
rect 182 281 216 315
rect 250 281 284 315
rect 318 281 352 315
rect 386 281 420 315
rect 569 279 603 313
rect 637 279 671 313
rect 705 279 739 313
rect 773 279 807 313
rect 841 279 875 313
rect 909 279 943 313
rect 977 279 1011 313
rect 1223 279 1257 313
rect 1395 279 1429 313
rect 1567 279 1601 313
rect 1739 279 1773 313
rect 1911 279 1945 313
rect 2083 279 2117 313
rect 2255 279 2289 313
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 19 590 78 615
rect 19 556 35 590
rect 69 556 78 590
rect 19 511 78 556
rect 19 477 35 511
rect 69 477 78 511
rect 19 434 78 477
rect 112 570 164 649
rect 112 536 121 570
rect 155 536 164 570
rect 112 502 164 536
rect 112 468 121 502
rect 155 468 164 502
rect 112 452 164 468
rect 201 590 243 615
rect 201 556 207 590
rect 241 556 243 590
rect 201 506 243 556
rect 201 472 207 506
rect 241 472 243 506
rect 19 400 35 434
rect 69 418 78 434
rect 201 422 243 472
rect 277 603 343 649
rect 277 569 293 603
rect 327 569 343 603
rect 277 535 343 569
rect 277 501 293 535
rect 327 501 343 535
rect 277 467 343 501
rect 277 433 293 467
rect 327 433 343 467
rect 277 423 343 433
rect 377 590 429 615
rect 377 556 379 590
rect 413 556 429 590
rect 377 506 429 556
rect 377 472 379 506
rect 413 472 429 506
rect 69 400 167 418
rect 19 384 167 400
rect 31 309 97 350
rect 31 275 47 309
rect 81 275 97 309
rect 31 271 97 275
rect 133 318 167 384
rect 201 388 207 422
rect 241 389 243 422
rect 377 422 429 472
rect 377 389 379 422
rect 241 388 379 389
rect 413 388 429 422
rect 519 598 585 649
rect 519 564 535 598
rect 569 564 585 598
rect 519 530 585 564
rect 519 496 535 530
rect 569 496 585 530
rect 519 462 585 496
rect 519 428 535 462
rect 569 428 585 462
rect 519 420 585 428
rect 619 594 664 615
rect 619 560 621 594
rect 655 560 664 594
rect 619 510 664 560
rect 619 476 621 510
rect 655 476 664 510
rect 619 426 664 476
rect 201 386 429 388
rect 619 392 621 426
rect 655 392 664 426
rect 698 605 750 649
rect 698 571 707 605
rect 741 571 750 605
rect 698 537 750 571
rect 698 503 707 537
rect 741 503 750 537
rect 698 469 750 503
rect 698 435 707 469
rect 741 435 750 469
rect 698 419 750 435
rect 784 594 836 615
rect 784 560 793 594
rect 827 560 836 594
rect 784 510 836 560
rect 784 476 793 510
rect 827 476 836 510
rect 784 426 836 476
rect 201 352 504 386
rect 133 315 436 318
rect 133 281 182 315
rect 216 281 250 315
rect 284 281 318 315
rect 352 281 386 315
rect 420 281 436 315
rect 470 315 504 352
rect 619 385 664 392
rect 784 392 793 426
rect 827 392 836 426
rect 870 605 922 649
rect 870 571 879 605
rect 913 571 922 605
rect 870 537 922 571
rect 870 503 879 537
rect 913 503 922 537
rect 870 469 922 503
rect 870 435 879 469
rect 913 435 922 469
rect 870 419 922 435
rect 956 594 1008 615
rect 956 560 965 594
rect 999 560 1008 594
rect 956 510 1008 560
rect 956 476 965 510
rect 999 476 1008 510
rect 956 426 1008 476
rect 784 385 836 392
rect 956 392 965 426
rect 999 392 1008 426
rect 1042 605 1094 649
rect 1042 571 1051 605
rect 1085 571 1094 605
rect 1042 537 1094 571
rect 1042 503 1051 537
rect 1085 503 1094 537
rect 1042 469 1094 503
rect 1042 435 1051 469
rect 1085 435 1094 469
rect 1042 419 1094 435
rect 1133 594 1180 615
rect 1133 560 1137 594
rect 1171 560 1180 594
rect 1133 510 1180 560
rect 1133 476 1137 510
rect 1171 476 1180 510
rect 1133 426 1180 476
rect 956 385 1008 392
rect 1133 390 1137 426
rect 1171 390 1180 426
rect 619 350 1099 385
rect 619 349 1063 350
rect 1061 316 1063 349
rect 1097 316 1099 350
rect 470 313 1027 315
rect 133 237 167 281
rect 470 279 569 313
rect 603 279 637 313
rect 671 279 705 313
rect 739 279 773 313
rect 807 279 841 313
rect 875 279 909 313
rect 943 279 977 313
rect 1011 279 1027 313
rect 470 277 1027 279
rect 470 247 571 277
rect 19 203 167 237
rect 205 213 571 247
rect 1061 243 1099 316
rect 19 185 71 203
rect 19 151 35 185
rect 69 151 71 185
rect 205 184 243 213
rect 19 101 71 151
rect 19 67 35 101
rect 69 67 71 101
rect 19 51 71 67
rect 105 163 171 169
rect 105 129 121 163
rect 155 129 171 163
rect 105 95 171 129
rect 105 61 121 95
rect 155 61 171 95
rect 105 17 171 61
rect 205 150 207 184
rect 241 150 243 184
rect 377 184 429 213
rect 205 101 243 150
rect 205 67 207 101
rect 241 67 243 101
rect 205 51 243 67
rect 277 170 343 179
rect 277 136 293 170
rect 327 136 343 170
rect 277 102 343 136
rect 277 68 293 102
rect 327 68 343 102
rect 277 17 343 68
rect 377 150 379 184
rect 413 150 429 184
rect 611 209 1099 243
rect 611 189 657 209
rect 377 101 429 150
rect 377 67 379 101
rect 413 67 429 101
rect 377 51 429 67
rect 519 163 577 179
rect 519 129 535 163
rect 569 129 577 163
rect 519 95 577 129
rect 519 61 535 95
rect 569 61 577 95
rect 519 17 577 61
rect 611 155 621 189
rect 655 155 657 189
rect 784 189 836 209
rect 611 107 657 155
rect 611 73 621 107
rect 655 73 657 107
rect 611 51 657 73
rect 691 159 750 175
rect 691 125 707 159
rect 741 125 750 159
rect 691 91 750 125
rect 691 57 707 91
rect 741 57 750 91
rect 691 17 750 57
rect 784 155 793 189
rect 827 155 836 189
rect 956 189 1008 209
rect 784 107 836 155
rect 784 73 793 107
rect 827 73 836 107
rect 784 51 836 73
rect 870 159 922 175
rect 870 125 879 159
rect 913 125 922 159
rect 870 91 922 125
rect 870 57 879 91
rect 913 57 922 91
rect 870 17 922 57
rect 956 155 965 189
rect 999 155 1008 189
rect 1133 189 1180 390
rect 1214 598 1266 649
rect 1214 564 1223 598
rect 1257 564 1266 598
rect 1214 516 1266 564
rect 1214 482 1223 516
rect 1257 482 1266 516
rect 1214 435 1266 482
rect 1214 401 1223 435
rect 1257 401 1266 435
rect 1214 385 1266 401
rect 1300 594 1352 615
rect 1300 560 1309 594
rect 1343 560 1352 594
rect 1300 510 1352 560
rect 1300 476 1309 510
rect 1343 476 1352 510
rect 1300 426 1352 476
rect 1300 390 1309 426
rect 1343 390 1352 426
rect 1214 350 1266 351
rect 1214 316 1223 350
rect 1257 316 1266 350
rect 1214 313 1266 316
rect 1214 279 1223 313
rect 1257 279 1266 313
rect 1214 263 1266 279
rect 956 107 1008 155
rect 956 73 965 107
rect 999 73 1008 107
rect 956 51 1008 73
rect 1042 159 1094 175
rect 1042 125 1051 159
rect 1085 125 1094 159
rect 1042 91 1094 125
rect 1042 57 1051 91
rect 1085 57 1094 91
rect 1042 17 1094 57
rect 1133 155 1137 189
rect 1171 155 1180 189
rect 1133 107 1180 155
rect 1133 73 1137 107
rect 1171 73 1180 107
rect 1133 51 1180 73
rect 1214 189 1266 215
rect 1214 155 1223 189
rect 1257 155 1266 189
rect 1214 107 1266 155
rect 1214 73 1223 107
rect 1257 73 1266 107
rect 1214 17 1266 73
rect 1300 189 1352 390
rect 1386 598 1438 649
rect 1386 564 1395 598
rect 1429 564 1438 598
rect 1386 516 1438 564
rect 1386 482 1395 516
rect 1429 482 1438 516
rect 1386 435 1438 482
rect 1386 401 1395 435
rect 1429 401 1438 435
rect 1386 385 1438 401
rect 1472 594 1524 615
rect 1472 560 1481 594
rect 1515 560 1524 594
rect 1472 510 1524 560
rect 1472 476 1481 510
rect 1515 476 1524 510
rect 1472 426 1524 476
rect 1472 390 1481 426
rect 1515 390 1524 426
rect 1386 350 1438 351
rect 1386 316 1395 350
rect 1429 316 1438 350
rect 1386 313 1438 316
rect 1386 279 1395 313
rect 1429 279 1438 313
rect 1386 263 1438 279
rect 1300 155 1309 189
rect 1343 155 1352 189
rect 1300 107 1352 155
rect 1300 73 1309 107
rect 1343 73 1352 107
rect 1300 51 1352 73
rect 1386 189 1438 215
rect 1386 155 1395 189
rect 1429 155 1438 189
rect 1386 107 1438 155
rect 1386 73 1395 107
rect 1429 73 1438 107
rect 1386 17 1438 73
rect 1472 189 1524 390
rect 1558 598 1610 649
rect 1558 564 1567 598
rect 1601 564 1610 598
rect 1558 516 1610 564
rect 1558 482 1567 516
rect 1601 482 1610 516
rect 1558 435 1610 482
rect 1558 401 1567 435
rect 1601 401 1610 435
rect 1558 385 1610 401
rect 1644 594 1696 615
rect 1644 560 1653 594
rect 1687 560 1696 594
rect 1644 510 1696 560
rect 1644 476 1653 510
rect 1687 476 1696 510
rect 1644 426 1696 476
rect 1644 390 1653 426
rect 1687 390 1696 426
rect 1558 350 1610 351
rect 1558 316 1567 350
rect 1601 316 1610 350
rect 1558 313 1610 316
rect 1558 279 1567 313
rect 1601 279 1610 313
rect 1558 263 1610 279
rect 1472 155 1481 189
rect 1515 155 1524 189
rect 1472 107 1524 155
rect 1472 73 1481 107
rect 1515 73 1524 107
rect 1472 51 1524 73
rect 1558 189 1610 215
rect 1558 155 1567 189
rect 1601 155 1610 189
rect 1558 107 1610 155
rect 1558 73 1567 107
rect 1601 73 1610 107
rect 1558 17 1610 73
rect 1644 189 1696 390
rect 1730 598 1782 649
rect 1730 564 1739 598
rect 1773 564 1782 598
rect 1730 516 1782 564
rect 1730 482 1739 516
rect 1773 482 1782 516
rect 1730 435 1782 482
rect 1730 401 1739 435
rect 1773 401 1782 435
rect 1730 385 1782 401
rect 1816 594 1868 615
rect 1816 560 1825 594
rect 1859 560 1868 594
rect 1816 510 1868 560
rect 1816 476 1825 510
rect 1859 476 1868 510
rect 1816 426 1868 476
rect 1816 390 1825 426
rect 1859 390 1868 426
rect 1730 350 1782 351
rect 1730 316 1739 350
rect 1773 316 1782 350
rect 1730 313 1782 316
rect 1730 279 1739 313
rect 1773 279 1782 313
rect 1730 263 1782 279
rect 1644 155 1653 189
rect 1687 155 1696 189
rect 1644 107 1696 155
rect 1644 73 1653 107
rect 1687 73 1696 107
rect 1644 51 1696 73
rect 1730 189 1782 215
rect 1730 155 1739 189
rect 1773 155 1782 189
rect 1730 107 1782 155
rect 1730 73 1739 107
rect 1773 73 1782 107
rect 1730 17 1782 73
rect 1816 189 1868 390
rect 1902 598 1954 649
rect 1902 564 1911 598
rect 1945 564 1954 598
rect 1902 516 1954 564
rect 1902 482 1911 516
rect 1945 482 1954 516
rect 1902 435 1954 482
rect 1902 401 1911 435
rect 1945 401 1954 435
rect 1902 385 1954 401
rect 1988 594 2040 615
rect 1988 560 1997 594
rect 2031 560 2040 594
rect 1988 510 2040 560
rect 1988 476 1997 510
rect 2031 476 2040 510
rect 1988 426 2040 476
rect 1988 390 1997 426
rect 2031 390 2040 426
rect 1902 350 1954 351
rect 1902 316 1911 350
rect 1945 316 1954 350
rect 1902 313 1954 316
rect 1902 279 1911 313
rect 1945 279 1954 313
rect 1902 263 1954 279
rect 1816 155 1825 189
rect 1859 155 1868 189
rect 1816 107 1868 155
rect 1816 73 1825 107
rect 1859 73 1868 107
rect 1816 51 1868 73
rect 1902 189 1954 215
rect 1902 155 1911 189
rect 1945 155 1954 189
rect 1902 107 1954 155
rect 1902 73 1911 107
rect 1945 73 1954 107
rect 1902 17 1954 73
rect 1988 189 2040 390
rect 2074 598 2126 649
rect 2074 564 2083 598
rect 2117 564 2126 598
rect 2074 516 2126 564
rect 2074 482 2083 516
rect 2117 482 2126 516
rect 2074 435 2126 482
rect 2074 401 2083 435
rect 2117 401 2126 435
rect 2074 385 2126 401
rect 2160 594 2212 615
rect 2160 560 2169 594
rect 2203 560 2212 594
rect 2160 510 2212 560
rect 2160 476 2169 510
rect 2203 476 2212 510
rect 2160 426 2212 476
rect 2160 390 2169 426
rect 2203 390 2212 426
rect 2074 350 2126 351
rect 2074 316 2083 350
rect 2117 316 2126 350
rect 2074 313 2126 316
rect 2074 279 2083 313
rect 2117 279 2126 313
rect 2074 263 2126 279
rect 1988 155 1997 189
rect 2031 155 2040 189
rect 1988 107 2040 155
rect 1988 73 1997 107
rect 2031 73 2040 107
rect 1988 51 2040 73
rect 2074 189 2126 215
rect 2074 155 2083 189
rect 2117 155 2126 189
rect 2074 107 2126 155
rect 2074 73 2083 107
rect 2117 73 2126 107
rect 2074 17 2126 73
rect 2160 189 2212 390
rect 2246 598 2298 649
rect 2246 564 2255 598
rect 2289 564 2298 598
rect 2246 516 2298 564
rect 2246 482 2255 516
rect 2289 482 2298 516
rect 2246 435 2298 482
rect 2246 401 2255 435
rect 2289 401 2298 435
rect 2246 385 2298 401
rect 2332 594 2384 615
rect 2332 560 2341 594
rect 2375 560 2384 594
rect 2332 510 2384 560
rect 2332 476 2341 510
rect 2375 476 2384 510
rect 2332 426 2384 476
rect 2332 390 2341 426
rect 2375 390 2384 426
rect 2246 350 2298 351
rect 2246 316 2255 350
rect 2289 316 2298 350
rect 2246 313 2298 316
rect 2246 279 2255 313
rect 2289 279 2298 313
rect 2246 263 2298 279
rect 2160 155 2169 189
rect 2203 155 2212 189
rect 2160 107 2212 155
rect 2160 73 2169 107
rect 2203 73 2212 107
rect 2160 51 2212 73
rect 2246 189 2298 215
rect 2246 155 2255 189
rect 2289 155 2298 189
rect 2246 107 2298 155
rect 2246 73 2255 107
rect 2289 73 2298 107
rect 2246 17 2298 73
rect 2332 189 2384 390
rect 2418 598 2477 649
rect 2418 564 2427 598
rect 2461 564 2477 598
rect 2418 516 2477 564
rect 2418 482 2427 516
rect 2461 482 2477 516
rect 2418 435 2477 482
rect 2418 401 2427 435
rect 2461 401 2477 435
rect 2418 385 2477 401
rect 2332 155 2341 189
rect 2375 155 2384 189
rect 2332 107 2384 155
rect 2332 73 2341 107
rect 2375 73 2384 107
rect 2332 51 2384 73
rect 2418 189 2477 215
rect 2418 155 2427 189
rect 2461 155 2477 189
rect 2418 107 2477 155
rect 2418 73 2427 107
rect 2461 73 2477 107
rect 2418 17 2477 73
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 1137 392 1171 424
rect 1137 390 1171 392
rect 1063 316 1097 350
rect 1309 392 1343 424
rect 1309 390 1343 392
rect 1223 316 1257 350
rect 1481 392 1515 424
rect 1481 390 1515 392
rect 1395 316 1429 350
rect 1653 392 1687 424
rect 1653 390 1687 392
rect 1567 316 1601 350
rect 1825 392 1859 424
rect 1825 390 1859 392
rect 1739 316 1773 350
rect 1997 392 2031 424
rect 1997 390 2031 392
rect 1911 316 1945 350
rect 2169 392 2203 424
rect 2169 390 2203 392
rect 2083 316 2117 350
rect 2341 392 2375 424
rect 2341 390 2375 392
rect 2255 316 2289 350
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 683 2496 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 0 617 2496 649
rect 1125 424 2387 430
rect 1125 390 1137 424
rect 1171 390 1309 424
rect 1343 390 1481 424
rect 1515 390 1653 424
rect 1687 390 1825 424
rect 1859 390 1997 424
rect 2031 390 2169 424
rect 2203 390 2341 424
rect 2375 390 2387 424
rect 1125 384 2387 390
rect 1051 350 2301 356
rect 1051 316 1063 350
rect 1097 316 1223 350
rect 1257 316 1395 350
rect 1429 316 1567 350
rect 1601 316 1739 350
rect 1773 316 1911 350
rect 1945 316 2083 350
rect 2117 316 2255 350
rect 2289 316 2301 350
rect 1051 310 2301 316
rect 0 17 2496 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
rect 0 -49 2496 -17
<< labels >>
flabel pwell s 0 0 2496 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 2496 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 bufbuf_16
flabel metal1 s 1125 384 2387 430 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel metal1 s 0 617 2496 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 2496 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2496 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6888368
string GDS_START 6867588
<< end >>
