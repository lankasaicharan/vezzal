magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 3 157 565 161
rect 3 49 863 157
rect 0 0 864 49
<< scnmos >>
rect 86 51 116 135
rect 188 51 218 135
rect 296 51 326 135
rect 374 51 404 135
rect 452 51 482 135
rect 678 47 708 131
rect 750 47 780 131
<< scpmoshvt >>
rect 84 419 134 619
rect 182 419 232 619
rect 296 419 346 619
rect 466 419 516 619
rect 576 419 626 619
rect 682 419 732 619
<< ndiff >>
rect 29 113 86 135
rect 29 79 41 113
rect 75 79 86 113
rect 29 51 86 79
rect 116 110 188 135
rect 116 76 127 110
rect 161 76 188 110
rect 116 51 188 76
rect 218 113 296 135
rect 218 79 229 113
rect 263 79 296 113
rect 218 51 296 79
rect 326 51 374 135
rect 404 51 452 135
rect 482 99 539 135
rect 482 65 493 99
rect 527 65 539 99
rect 482 51 539 65
rect 621 97 678 131
rect 621 63 633 97
rect 667 63 678 97
rect 621 47 678 63
rect 708 47 750 131
rect 780 111 837 131
rect 780 77 791 111
rect 825 77 837 111
rect 780 47 837 77
<< pdiff >>
rect 27 607 84 619
rect 27 573 39 607
rect 73 573 84 607
rect 27 536 84 573
rect 27 502 39 536
rect 73 502 84 536
rect 27 465 84 502
rect 27 431 39 465
rect 73 431 84 465
rect 27 419 84 431
rect 134 419 182 619
rect 232 597 296 619
rect 232 563 251 597
rect 285 563 296 597
rect 232 465 296 563
rect 232 431 251 465
rect 285 431 296 465
rect 232 419 296 431
rect 346 596 466 619
rect 346 562 357 596
rect 391 562 466 596
rect 346 419 466 562
rect 516 597 576 619
rect 516 563 531 597
rect 565 563 576 597
rect 516 465 576 563
rect 516 431 531 465
rect 565 431 576 465
rect 516 419 576 431
rect 626 607 682 619
rect 626 573 637 607
rect 671 573 682 607
rect 626 536 682 573
rect 626 502 637 536
rect 671 502 682 536
rect 626 465 682 502
rect 626 431 637 465
rect 671 431 682 465
rect 626 419 682 431
rect 732 597 789 619
rect 732 563 743 597
rect 777 563 789 597
rect 732 465 789 563
rect 732 431 743 465
rect 777 431 789 465
rect 732 419 789 431
<< ndiffc >>
rect 41 79 75 113
rect 127 76 161 110
rect 229 79 263 113
rect 493 65 527 99
rect 633 63 667 97
rect 791 77 825 111
<< pdiffc >>
rect 39 573 73 607
rect 39 502 73 536
rect 39 431 73 465
rect 251 563 285 597
rect 251 431 285 465
rect 357 562 391 596
rect 531 563 565 597
rect 531 431 565 465
rect 637 573 671 607
rect 637 502 671 536
rect 637 431 671 465
rect 743 563 777 597
rect 743 431 777 465
<< poly >>
rect 84 619 134 645
rect 182 619 232 645
rect 296 619 346 645
rect 466 619 516 645
rect 576 619 626 645
rect 682 619 732 645
rect 84 379 134 419
rect 68 363 134 379
rect 68 329 84 363
rect 118 329 134 363
rect 68 295 134 329
rect 68 261 84 295
rect 118 261 134 295
rect 68 245 134 261
rect 182 379 232 419
rect 296 379 346 419
rect 466 387 516 419
rect 182 363 248 379
rect 182 329 198 363
rect 232 329 248 363
rect 182 295 248 329
rect 182 261 198 295
rect 232 261 248 295
rect 182 245 248 261
rect 296 363 365 379
rect 296 329 315 363
rect 349 329 365 363
rect 296 313 365 329
rect 413 371 516 387
rect 413 337 429 371
rect 463 337 516 371
rect 86 135 116 245
rect 188 135 218 245
rect 296 135 326 313
rect 413 265 516 337
rect 374 235 516 265
rect 374 135 404 235
rect 576 219 626 419
rect 682 377 732 419
rect 678 361 749 377
rect 678 327 699 361
rect 733 327 749 361
rect 678 293 749 327
rect 678 259 699 293
rect 733 273 749 293
rect 733 259 780 273
rect 678 243 780 259
rect 564 203 630 219
rect 564 183 580 203
rect 452 169 580 183
rect 614 169 630 203
rect 452 153 630 169
rect 452 135 482 153
rect 678 131 708 243
rect 750 131 780 243
rect 86 25 116 51
rect 188 25 218 51
rect 296 25 326 51
rect 374 25 404 51
rect 452 25 482 51
rect 678 21 708 47
rect 750 21 780 47
<< polycont >>
rect 84 329 118 363
rect 84 261 118 295
rect 198 329 232 363
rect 198 261 232 295
rect 315 329 349 363
rect 429 337 463 371
rect 699 327 733 361
rect 699 259 733 293
rect 580 169 614 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 23 607 89 649
rect 23 573 39 607
rect 73 573 89 607
rect 23 536 89 573
rect 23 502 39 536
rect 73 502 89 536
rect 23 465 89 502
rect 23 431 39 465
rect 73 431 89 465
rect 23 415 89 431
rect 235 597 301 613
rect 235 563 251 597
rect 285 563 301 597
rect 235 500 301 563
rect 341 596 407 649
rect 341 562 357 596
rect 391 562 407 596
rect 341 536 407 562
rect 515 597 581 613
rect 515 563 531 597
rect 565 563 581 597
rect 515 500 581 563
rect 235 466 581 500
rect 235 465 301 466
rect 235 431 251 465
rect 285 431 301 465
rect 235 415 301 431
rect 515 465 581 466
rect 515 431 531 465
rect 565 431 581 465
rect 25 363 134 379
rect 25 329 84 363
rect 118 329 134 363
rect 25 295 134 329
rect 25 261 84 295
rect 118 261 134 295
rect 25 245 134 261
rect 182 363 263 379
rect 182 329 198 363
rect 232 329 263 363
rect 182 295 263 329
rect 182 261 198 295
rect 232 261 263 295
rect 182 245 263 261
rect 299 363 365 379
rect 299 329 315 363
rect 349 329 365 363
rect 25 175 263 209
rect 25 113 75 175
rect 25 79 41 113
rect 25 53 75 79
rect 111 110 177 139
rect 111 76 127 110
rect 161 76 177 110
rect 111 17 177 76
rect 213 113 263 175
rect 213 79 229 113
rect 299 88 365 329
rect 409 371 479 430
rect 409 337 429 371
rect 463 337 479 371
rect 409 323 479 337
rect 515 377 581 431
rect 621 607 687 649
rect 621 573 637 607
rect 671 573 687 607
rect 621 536 687 573
rect 621 502 637 536
rect 671 502 687 536
rect 621 465 687 502
rect 621 431 637 465
rect 671 431 687 465
rect 621 415 687 431
rect 727 597 841 613
rect 727 563 743 597
rect 777 563 841 597
rect 727 465 841 563
rect 727 431 743 465
rect 777 431 841 465
rect 727 415 841 431
rect 515 361 749 377
rect 515 343 699 361
rect 515 287 549 343
rect 435 253 549 287
rect 683 327 699 343
rect 733 327 749 361
rect 683 293 749 327
rect 683 259 699 293
rect 733 259 749 293
rect 435 117 469 253
rect 683 243 749 259
rect 505 203 647 217
rect 505 169 580 203
rect 614 169 647 203
rect 505 153 647 169
rect 793 135 841 415
rect 435 99 543 117
rect 213 53 263 79
rect 435 65 493 99
rect 527 65 543 99
rect 435 63 543 65
rect 617 97 683 117
rect 617 63 633 97
rect 667 63 683 97
rect 617 17 683 63
rect 775 111 841 135
rect 775 77 791 111
rect 825 77 841 111
rect 775 53 841 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2111a_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4240668
string GDS_START 4232268
<< end >>
