magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4466 1975
<< nwell >>
rect -38 331 3206 704
rect 2545 311 2815 331
<< pwell >>
rect 1158 218 2105 235
rect 724 176 2105 218
rect 724 167 2363 176
rect 724 157 3167 167
rect 31 49 3167 157
rect 0 0 3168 49
<< scnmos >>
rect 114 47 144 131
rect 186 47 216 131
rect 338 47 368 131
rect 416 47 446 131
rect 502 47 532 131
rect 580 47 610 131
rect 807 108 837 192
rect 885 108 915 192
rect 971 108 1001 192
rect 1043 108 1073 192
rect 1241 125 1271 209
rect 1353 125 1383 209
rect 1425 125 1455 209
rect 1706 125 1736 209
rect 1784 125 1814 209
rect 1898 125 1928 209
rect 1976 125 2006 209
rect 2094 66 2124 150
rect 2172 66 2202 150
rect 2250 66 2280 150
rect 2554 57 2584 141
rect 2626 57 2656 141
rect 2824 57 2854 141
rect 2896 57 2926 141
rect 2982 57 3012 141
rect 3054 57 3084 141
<< scpmoshvt >>
rect 84 409 134 609
rect 302 406 352 606
rect 408 406 458 606
rect 506 406 556 606
rect 612 406 662 606
rect 830 409 880 609
rect 936 409 986 609
rect 1149 419 1199 619
rect 1321 419 1371 619
rect 1427 419 1477 619
rect 1607 419 1657 619
rect 1713 419 1763 619
rect 1878 419 1928 619
rect 1976 419 2026 619
rect 2156 419 2206 619
rect 2264 419 2314 619
rect 2420 419 2470 619
rect 2638 347 2688 547
rect 2890 374 2940 574
rect 2996 374 3046 574
<< ndiff >>
rect 750 176 807 192
rect 750 142 762 176
rect 796 142 807 176
rect 57 111 114 131
rect 57 77 69 111
rect 103 77 114 111
rect 57 47 114 77
rect 144 47 186 131
rect 216 106 338 131
rect 216 72 227 106
rect 261 72 338 106
rect 216 47 338 72
rect 368 47 416 131
rect 446 106 502 131
rect 446 72 457 106
rect 491 72 502 106
rect 446 47 502 72
rect 532 47 580 131
rect 610 96 667 131
rect 750 108 807 142
rect 837 108 885 192
rect 915 167 971 192
rect 915 133 926 167
rect 960 133 971 167
rect 915 108 971 133
rect 1001 108 1043 192
rect 1073 176 1130 192
rect 1073 142 1084 176
rect 1118 142 1130 176
rect 1073 108 1130 142
rect 1184 184 1241 209
rect 1184 150 1196 184
rect 1230 150 1241 184
rect 1184 125 1241 150
rect 1271 184 1353 209
rect 1271 150 1295 184
rect 1329 150 1353 184
rect 1271 125 1353 150
rect 1383 125 1425 209
rect 1455 125 1525 209
rect 1649 185 1706 209
rect 1649 151 1661 185
rect 1695 151 1706 185
rect 1649 125 1706 151
rect 1736 125 1784 209
rect 1814 184 1898 209
rect 1814 150 1833 184
rect 1867 150 1898 184
rect 1814 125 1898 150
rect 1928 125 1976 209
rect 2006 197 2079 209
rect 2006 163 2033 197
rect 2067 163 2079 197
rect 2006 150 2079 163
rect 2006 125 2094 150
rect 610 62 621 96
rect 655 62 667 96
rect 610 47 667 62
rect 1470 121 1525 125
rect 1470 87 1479 121
rect 1513 87 1525 121
rect 2021 112 2094 125
rect 1470 75 1525 87
rect 2021 78 2033 112
rect 2067 78 2094 112
rect 2021 66 2094 78
rect 2124 66 2172 150
rect 2202 66 2250 150
rect 2280 121 2337 150
rect 2280 87 2291 121
rect 2325 87 2337 121
rect 2280 66 2337 87
rect 2497 116 2554 141
rect 2497 82 2509 116
rect 2543 82 2554 116
rect 2497 57 2554 82
rect 2584 57 2626 141
rect 2656 116 2713 141
rect 2656 82 2667 116
rect 2701 82 2713 116
rect 2656 57 2713 82
rect 2767 116 2824 141
rect 2767 82 2779 116
rect 2813 82 2824 116
rect 2767 57 2824 82
rect 2854 57 2896 141
rect 2926 116 2982 141
rect 2926 82 2937 116
rect 2971 82 2982 116
rect 2926 57 2982 82
rect 3012 57 3054 141
rect 3084 116 3141 141
rect 3084 82 3095 116
rect 3129 82 3141 116
rect 3084 57 3141 82
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 526 84 563
rect 27 492 39 526
rect 73 492 84 526
rect 27 455 84 492
rect 27 421 39 455
rect 73 421 84 455
rect 27 409 84 421
rect 134 597 191 609
rect 1492 621 1550 633
rect 1492 619 1504 621
rect 134 563 145 597
rect 179 563 191 597
rect 134 526 191 563
rect 134 492 145 526
rect 179 492 191 526
rect 134 455 191 492
rect 134 421 145 455
rect 179 421 191 455
rect 134 409 191 421
rect 245 594 302 606
rect 245 560 257 594
rect 291 560 302 594
rect 245 523 302 560
rect 245 489 257 523
rect 291 489 302 523
rect 245 452 302 489
rect 245 418 257 452
rect 291 418 302 452
rect 245 406 302 418
rect 352 527 408 606
rect 352 493 363 527
rect 397 493 408 527
rect 352 452 408 493
rect 352 418 363 452
rect 397 418 408 452
rect 352 406 408 418
rect 458 406 506 606
rect 556 589 612 606
rect 556 555 567 589
rect 601 555 612 589
rect 556 406 612 555
rect 662 594 719 606
rect 662 560 673 594
rect 707 560 719 594
rect 662 523 719 560
rect 662 489 673 523
rect 707 489 719 523
rect 662 452 719 489
rect 662 418 673 452
rect 707 418 719 452
rect 662 406 719 418
rect 773 597 830 609
rect 773 563 785 597
rect 819 563 830 597
rect 773 526 830 563
rect 773 492 785 526
rect 819 492 830 526
rect 773 455 830 492
rect 773 421 785 455
rect 819 421 830 455
rect 773 409 830 421
rect 880 597 936 609
rect 880 563 891 597
rect 925 563 936 597
rect 880 524 936 563
rect 880 490 891 524
rect 925 490 936 524
rect 880 409 936 490
rect 986 597 1040 609
rect 986 563 997 597
rect 1031 563 1040 597
rect 986 524 1040 563
rect 986 490 997 524
rect 1031 490 1040 524
rect 986 409 1040 490
rect 1094 496 1149 619
rect 1094 462 1104 496
rect 1138 462 1149 496
rect 1094 419 1149 462
rect 1199 496 1321 619
rect 1199 462 1276 496
rect 1310 462 1321 496
rect 1199 419 1321 462
rect 1371 419 1427 619
rect 1477 587 1504 619
rect 1538 619 1550 621
rect 1538 587 1607 619
rect 1477 419 1607 587
rect 1657 465 1713 619
rect 1657 431 1668 465
rect 1702 431 1713 465
rect 1657 419 1713 431
rect 1763 606 1878 619
rect 1763 572 1774 606
rect 1808 572 1878 606
rect 1763 419 1878 572
rect 1928 419 1976 619
rect 2026 597 2156 619
rect 2026 563 2064 597
rect 2098 563 2156 597
rect 2026 465 2156 563
rect 2026 431 2064 465
rect 2098 431 2156 465
rect 2026 419 2156 431
rect 2206 419 2264 619
rect 2314 596 2420 619
rect 2314 562 2325 596
rect 2359 562 2420 596
rect 2314 419 2420 562
rect 2470 597 2527 619
rect 2470 563 2481 597
rect 2515 563 2527 597
rect 2470 516 2527 563
rect 2833 562 2890 574
rect 2470 482 2481 516
rect 2515 482 2527 516
rect 2470 419 2527 482
rect 2581 527 2638 547
rect 2581 493 2593 527
rect 2627 493 2638 527
rect 2581 393 2638 493
rect 2581 359 2593 393
rect 2627 359 2638 393
rect 2581 347 2638 359
rect 2688 535 2779 547
rect 2688 501 2733 535
rect 2767 501 2779 535
rect 2688 401 2779 501
rect 2688 367 2733 401
rect 2767 367 2779 401
rect 2833 528 2845 562
rect 2879 528 2890 562
rect 2833 491 2890 528
rect 2833 457 2845 491
rect 2879 457 2890 491
rect 2833 420 2890 457
rect 2833 386 2845 420
rect 2879 386 2890 420
rect 2833 374 2890 386
rect 2940 562 2996 574
rect 2940 528 2951 562
rect 2985 528 2996 562
rect 2940 491 2996 528
rect 2940 457 2951 491
rect 2985 457 2996 491
rect 2940 420 2996 457
rect 2940 386 2951 420
rect 2985 386 2996 420
rect 2940 374 2996 386
rect 3046 562 3103 574
rect 3046 528 3057 562
rect 3091 528 3103 562
rect 3046 491 3103 528
rect 3046 457 3057 491
rect 3091 457 3103 491
rect 3046 420 3103 457
rect 3046 386 3057 420
rect 3091 386 3103 420
rect 3046 374 3103 386
rect 2688 347 2779 367
<< ndiffc >>
rect 762 142 796 176
rect 69 77 103 111
rect 227 72 261 106
rect 457 72 491 106
rect 926 133 960 167
rect 1084 142 1118 176
rect 1196 150 1230 184
rect 1295 150 1329 184
rect 1661 151 1695 185
rect 1833 150 1867 184
rect 2033 163 2067 197
rect 621 62 655 96
rect 1479 87 1513 121
rect 2033 78 2067 112
rect 2291 87 2325 121
rect 2509 82 2543 116
rect 2667 82 2701 116
rect 2779 82 2813 116
rect 2937 82 2971 116
rect 3095 82 3129 116
<< pdiffc >>
rect 39 563 73 597
rect 39 492 73 526
rect 39 421 73 455
rect 145 563 179 597
rect 145 492 179 526
rect 145 421 179 455
rect 257 560 291 594
rect 257 489 291 523
rect 257 418 291 452
rect 363 493 397 527
rect 363 418 397 452
rect 567 555 601 589
rect 673 560 707 594
rect 673 489 707 523
rect 673 418 707 452
rect 785 563 819 597
rect 785 492 819 526
rect 785 421 819 455
rect 891 563 925 597
rect 891 490 925 524
rect 997 563 1031 597
rect 997 490 1031 524
rect 1104 462 1138 496
rect 1276 462 1310 496
rect 1504 587 1538 621
rect 1668 431 1702 465
rect 1774 572 1808 606
rect 2064 563 2098 597
rect 2064 431 2098 465
rect 2325 562 2359 596
rect 2481 563 2515 597
rect 2481 482 2515 516
rect 2593 493 2627 527
rect 2593 359 2627 393
rect 2733 501 2767 535
rect 2733 367 2767 401
rect 2845 528 2879 562
rect 2845 457 2879 491
rect 2845 386 2879 420
rect 2951 528 2985 562
rect 2951 457 2985 491
rect 2951 386 2985 420
rect 3057 528 3091 562
rect 3057 457 3091 491
rect 3057 386 3091 420
<< poly >>
rect 84 609 134 635
rect 302 606 352 632
rect 408 606 458 632
rect 506 606 556 632
rect 612 606 662 632
rect 830 609 880 635
rect 936 609 986 635
rect 1149 619 1199 645
rect 1321 619 1371 645
rect 1427 619 1477 645
rect 84 237 134 409
rect 1607 619 1657 645
rect 1713 619 1763 645
rect 1878 619 1928 645
rect 1976 619 2026 645
rect 2156 619 2206 645
rect 2264 619 2314 645
rect 2420 619 2470 645
rect 2890 574 2940 600
rect 2996 574 3046 600
rect 2638 547 2688 573
rect 302 358 352 406
rect 408 358 458 406
rect 506 358 556 406
rect 612 366 662 406
rect 830 368 880 409
rect 936 377 986 409
rect 211 342 352 358
rect 211 308 227 342
rect 261 308 352 342
rect 211 292 352 308
rect 394 342 460 358
rect 394 308 410 342
rect 444 308 460 342
rect 394 292 460 308
rect 502 342 568 358
rect 502 308 518 342
rect 552 308 568 342
rect 84 221 216 237
rect 84 187 166 221
rect 200 187 216 221
rect 84 171 216 187
rect 114 131 144 171
rect 186 131 216 171
rect 322 176 352 292
rect 322 146 368 176
rect 338 131 368 146
rect 416 131 446 292
rect 502 274 568 308
rect 502 240 518 274
rect 552 240 568 274
rect 502 224 568 240
rect 612 350 738 366
rect 612 316 688 350
rect 722 316 738 350
rect 612 282 738 316
rect 612 248 688 282
rect 722 248 738 282
rect 612 232 738 248
rect 807 352 894 368
rect 807 318 844 352
rect 878 318 894 352
rect 807 263 894 318
rect 936 361 1025 377
rect 1149 368 1199 419
rect 1321 404 1371 419
rect 936 327 975 361
rect 1009 327 1025 361
rect 936 311 1025 327
rect 1133 352 1199 368
rect 1133 318 1149 352
rect 1183 318 1199 352
rect 807 233 915 263
rect 502 131 532 224
rect 612 176 642 232
rect 807 192 837 233
rect 885 192 915 233
rect 971 254 1001 311
rect 1133 302 1199 318
rect 1241 374 1371 404
rect 1427 377 1477 419
rect 1607 379 1657 419
rect 1713 387 1763 419
rect 1241 254 1271 374
rect 1427 361 1551 377
rect 1427 327 1501 361
rect 1535 327 1551 361
rect 1313 310 1379 326
rect 1313 276 1329 310
rect 1363 290 1379 310
rect 1427 293 1551 327
rect 1599 363 1665 379
rect 1599 329 1615 363
rect 1649 329 1665 363
rect 1599 313 1665 329
rect 1713 371 1820 387
rect 1878 383 1928 419
rect 1713 337 1770 371
rect 1804 337 1820 371
rect 1713 321 1820 337
rect 1862 367 1928 383
rect 1976 404 2026 419
rect 1976 374 2108 404
rect 2156 387 2206 419
rect 1862 333 1878 367
rect 1912 333 1928 367
rect 1363 276 1383 290
rect 1313 260 1383 276
rect 1427 273 1501 293
rect 971 224 1271 254
rect 971 192 1001 224
rect 1043 192 1073 224
rect 1241 209 1271 224
rect 1353 209 1383 260
rect 1425 259 1501 273
rect 1535 259 1551 293
rect 1425 243 1551 259
rect 1635 273 1665 313
rect 1635 243 1736 273
rect 1425 209 1455 243
rect 1706 209 1736 243
rect 1784 209 1814 321
rect 1862 299 1928 333
rect 1862 265 1878 299
rect 1912 265 1928 299
rect 1862 249 1928 265
rect 1970 310 2036 326
rect 1970 276 1986 310
rect 2020 276 2036 310
rect 1970 260 2036 276
rect 1898 209 1928 249
rect 1976 209 2006 260
rect 2078 254 2108 374
rect 2150 371 2216 387
rect 2150 337 2166 371
rect 2200 337 2216 371
rect 2150 321 2216 337
rect 2264 377 2314 419
rect 2420 387 2470 419
rect 2264 361 2378 377
rect 2264 327 2328 361
rect 2362 327 2378 361
rect 2264 293 2378 327
rect 2264 273 2328 293
rect 2172 259 2328 273
rect 2362 259 2378 293
rect 2078 224 2124 254
rect 580 146 642 176
rect 580 131 610 146
rect 2094 150 2124 224
rect 2172 243 2378 259
rect 2420 371 2486 387
rect 2420 337 2436 371
rect 2470 337 2486 371
rect 2420 303 2486 337
rect 2420 269 2436 303
rect 2470 269 2486 303
rect 2172 150 2202 243
rect 2420 195 2486 269
rect 2638 315 2688 347
rect 2890 315 2940 374
rect 2996 332 3046 374
rect 2638 299 2940 315
rect 2638 265 2679 299
rect 2713 285 2940 299
rect 2982 316 3048 332
rect 2713 265 2729 285
rect 2638 231 2729 265
rect 2638 197 2679 231
rect 2713 197 2729 231
rect 2638 195 2729 197
rect 2250 165 2486 195
rect 2554 165 2729 195
rect 2250 150 2280 165
rect 807 82 837 108
rect 885 82 915 108
rect 971 82 1001 108
rect 1043 82 1073 108
rect 1241 51 1271 125
rect 1353 99 1383 125
rect 1425 99 1455 125
rect 1706 99 1736 125
rect 1784 99 1814 125
rect 1898 99 1928 125
rect 1976 99 2006 125
rect 2554 141 2584 165
rect 2626 141 2656 165
rect 2824 141 2854 285
rect 2896 141 2926 285
rect 2982 282 2998 316
rect 3032 282 3048 316
rect 2982 248 3048 282
rect 2982 214 2998 248
rect 3032 228 3048 248
rect 3032 214 3084 228
rect 2982 198 3084 214
rect 2982 141 3012 198
rect 3054 141 3084 198
rect 2094 51 2124 66
rect 114 21 144 47
rect 186 21 216 47
rect 338 21 368 47
rect 416 21 446 47
rect 502 21 532 47
rect 580 21 610 47
rect 1241 21 2124 51
rect 2172 40 2202 66
rect 2250 40 2280 66
rect 2554 31 2584 57
rect 2626 31 2656 57
rect 2824 31 2854 57
rect 2896 31 2926 57
rect 2982 31 3012 57
rect 3054 31 3084 57
<< polycont >>
rect 227 308 261 342
rect 410 308 444 342
rect 518 308 552 342
rect 166 187 200 221
rect 518 240 552 274
rect 688 316 722 350
rect 688 248 722 282
rect 844 318 878 352
rect 975 327 1009 361
rect 1149 318 1183 352
rect 1501 327 1535 361
rect 1329 276 1363 310
rect 1615 329 1649 363
rect 1770 337 1804 371
rect 1878 333 1912 367
rect 1501 259 1535 293
rect 1878 265 1912 299
rect 1986 276 2020 310
rect 2166 337 2200 371
rect 2328 327 2362 361
rect 2328 259 2362 293
rect 2436 337 2470 371
rect 2436 269 2470 303
rect 2679 265 2713 299
rect 2679 197 2713 231
rect 2998 282 3032 316
rect 2998 214 3032 248
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 526 89 563
rect 23 492 39 526
rect 73 492 89 526
rect 23 455 89 492
rect 23 421 39 455
rect 73 421 89 455
rect 23 358 89 421
rect 129 597 195 649
rect 129 563 145 597
rect 179 563 195 597
rect 129 526 195 563
rect 129 492 145 526
rect 179 492 195 526
rect 129 455 195 492
rect 129 421 145 455
rect 179 421 195 455
rect 129 405 195 421
rect 241 594 483 613
rect 241 560 257 594
rect 291 579 483 594
rect 291 560 307 579
rect 241 523 307 560
rect 241 489 257 523
rect 291 489 307 523
rect 241 452 307 489
rect 241 418 257 452
rect 291 418 307 452
rect 241 402 307 418
rect 347 527 413 543
rect 347 493 363 527
rect 397 493 413 527
rect 347 452 413 493
rect 449 498 483 579
rect 551 589 617 649
rect 551 555 567 589
rect 601 555 617 589
rect 551 534 617 555
rect 673 594 723 610
rect 707 560 723 594
rect 673 523 723 560
rect 449 489 673 498
rect 707 489 723 523
rect 449 464 723 489
rect 347 418 363 452
rect 397 428 413 452
rect 673 452 723 464
rect 397 418 637 428
rect 347 394 637 418
rect 707 418 723 452
rect 673 402 723 418
rect 769 597 835 613
rect 769 563 785 597
rect 819 563 835 597
rect 769 526 835 563
rect 769 492 785 526
rect 819 492 835 526
rect 769 455 835 492
rect 875 597 941 649
rect 1488 621 1554 649
rect 875 563 891 597
rect 925 563 941 597
rect 875 524 941 563
rect 875 490 891 524
rect 925 490 941 524
rect 875 474 941 490
rect 981 597 1396 613
rect 981 563 997 597
rect 1031 579 1396 597
rect 1031 563 1047 579
rect 981 524 1047 563
rect 981 490 997 524
rect 1031 490 1047 524
rect 981 474 1047 490
rect 1088 496 1154 543
rect 769 421 785 455
rect 819 438 835 455
rect 1088 462 1104 496
rect 1138 462 1154 496
rect 1088 438 1154 462
rect 819 421 1020 438
rect 769 404 1020 421
rect 23 342 277 358
rect 23 308 227 342
rect 261 308 277 342
rect 23 292 277 308
rect 313 342 460 358
rect 313 308 410 342
rect 444 308 460 342
rect 313 292 460 308
rect 502 342 567 358
rect 502 308 518 342
rect 552 308 567 342
rect 23 135 89 292
rect 502 274 567 308
rect 502 256 518 274
rect 313 240 518 256
rect 552 240 567 274
rect 313 237 567 240
rect 150 222 567 237
rect 150 221 455 222
rect 150 187 166 221
rect 200 187 455 221
rect 150 171 455 187
rect 603 186 637 394
rect 673 350 737 366
rect 673 316 688 350
rect 722 316 737 350
rect 673 282 737 316
rect 673 248 688 282
rect 722 248 737 282
rect 673 232 737 248
rect 773 196 807 404
rect 843 352 929 368
rect 843 318 844 352
rect 878 318 929 352
rect 843 302 929 318
rect 965 361 1020 404
rect 965 327 975 361
rect 1009 327 1020 361
rect 965 311 1020 327
rect 1056 404 1154 438
rect 1056 266 1090 404
rect 1190 368 1224 579
rect 1260 496 1326 543
rect 1362 535 1396 579
rect 1488 587 1504 621
rect 1538 587 1554 621
rect 1488 571 1554 587
rect 1758 606 1824 649
rect 1758 572 1774 606
rect 1808 572 1824 606
rect 1758 571 1824 572
rect 2048 597 2114 613
rect 2048 563 2064 597
rect 2098 563 2114 597
rect 1362 501 2004 535
rect 1260 462 1276 496
rect 1310 462 1326 496
rect 1260 449 1326 462
rect 1260 415 1449 449
rect 848 232 1090 266
rect 1126 352 1224 368
rect 1126 318 1149 352
rect 1183 326 1224 352
rect 1183 318 1379 326
rect 1126 310 1379 318
rect 1126 276 1329 310
rect 1363 276 1379 310
rect 1126 260 1379 276
rect 313 162 455 171
rect 491 152 725 186
rect 23 111 119 135
rect 23 77 69 111
rect 103 77 119 111
rect 23 53 119 77
rect 211 106 277 135
rect 491 126 525 152
rect 211 72 227 106
rect 261 72 277 106
rect 211 17 277 72
rect 441 106 525 126
rect 441 72 457 106
rect 491 72 525 106
rect 441 53 525 72
rect 605 96 655 116
rect 605 62 621 96
rect 605 17 655 62
rect 691 87 725 152
rect 762 176 812 196
rect 796 142 812 176
rect 762 123 812 142
rect 848 87 882 232
rect 691 53 882 87
rect 926 167 960 196
rect 926 17 960 133
rect 998 87 1032 232
rect 1126 196 1160 260
rect 1415 213 1449 415
rect 1485 431 1668 465
rect 1702 431 1718 465
rect 1485 415 1718 431
rect 1759 424 1820 430
rect 1485 361 1551 415
rect 1793 390 1820 424
rect 1485 327 1501 361
rect 1535 327 1551 361
rect 1485 293 1551 327
rect 1599 363 1723 379
rect 1599 329 1615 363
rect 1649 329 1723 363
rect 1599 313 1723 329
rect 1759 371 1820 390
rect 1759 337 1770 371
rect 1804 337 1820 371
rect 1759 321 1820 337
rect 1862 367 1928 383
rect 1862 333 1878 367
rect 1912 333 1928 367
rect 1485 259 1501 293
rect 1535 277 1551 293
rect 1689 283 1723 313
rect 1862 299 1928 333
rect 1862 283 1878 299
rect 1535 259 1653 277
rect 1485 243 1653 259
rect 1689 265 1878 283
rect 1912 265 1928 299
rect 1689 249 1928 265
rect 1970 326 2004 501
rect 2048 500 2114 563
rect 2309 596 2375 649
rect 2309 562 2325 596
rect 2359 562 2375 596
rect 2309 536 2375 562
rect 2465 597 2697 613
rect 2465 563 2481 597
rect 2515 579 2697 597
rect 2515 563 2531 579
rect 2465 516 2531 563
rect 2465 500 2481 516
rect 2048 482 2481 500
rect 2515 482 2531 516
rect 2048 466 2531 482
rect 2577 527 2627 543
rect 2577 493 2593 527
rect 2048 465 2114 466
rect 2048 431 2064 465
rect 2098 431 2114 465
rect 2048 415 2114 431
rect 2150 371 2211 387
rect 2150 337 2166 371
rect 2200 337 2211 371
rect 2150 326 2211 337
rect 1970 310 2211 326
rect 1970 276 1986 310
rect 2020 292 2211 310
rect 2020 276 2036 292
rect 1970 260 2036 276
rect 1068 176 1160 196
rect 1068 142 1084 176
rect 1118 142 1160 176
rect 1068 123 1160 142
rect 1196 184 1230 213
rect 1196 87 1230 150
rect 1279 207 1449 213
rect 1619 213 1653 243
rect 1279 184 1583 207
rect 1279 150 1295 184
rect 1329 173 1583 184
rect 1329 150 1345 173
rect 1279 121 1345 150
rect 1463 121 1513 137
rect 998 53 1230 87
rect 1463 87 1479 121
rect 1463 17 1513 87
rect 1549 87 1583 173
rect 1619 185 1711 213
rect 1619 151 1661 185
rect 1695 151 1711 185
rect 1619 123 1711 151
rect 1747 87 1781 249
rect 2247 217 2281 466
rect 2420 424 2486 430
rect 2420 390 2431 424
rect 2465 390 2486 424
rect 1549 53 1781 87
rect 1817 184 1883 213
rect 1817 150 1833 184
rect 1867 150 1883 184
rect 1817 17 1883 150
rect 2017 197 2281 217
rect 2017 163 2033 197
rect 2067 183 2281 197
rect 2317 361 2378 377
rect 2317 327 2328 361
rect 2362 327 2378 361
rect 2317 293 2378 327
rect 2317 259 2328 293
rect 2362 259 2378 293
rect 2317 217 2378 259
rect 2420 371 2486 390
rect 2420 337 2436 371
rect 2470 337 2486 371
rect 2420 303 2486 337
rect 2420 269 2436 303
rect 2470 269 2486 303
rect 2420 253 2486 269
rect 2577 393 2627 493
rect 2577 359 2593 393
rect 2577 217 2627 359
rect 2317 183 2627 217
rect 2663 315 2697 579
rect 2733 535 2783 649
rect 2767 501 2783 535
rect 2733 401 2783 501
rect 2767 367 2783 401
rect 2733 351 2783 367
rect 2819 562 2895 578
rect 2819 528 2845 562
rect 2879 528 2895 562
rect 2819 491 2895 528
rect 2819 457 2845 491
rect 2879 457 2895 491
rect 2819 420 2895 457
rect 2819 386 2845 420
rect 2879 386 2895 420
rect 2663 299 2729 315
rect 2663 265 2679 299
rect 2713 265 2729 299
rect 2663 231 2729 265
rect 2663 197 2679 231
rect 2713 197 2729 231
rect 2067 163 2106 183
rect 2017 112 2106 163
rect 2017 78 2033 112
rect 2067 78 2106 112
rect 2017 62 2106 78
rect 2275 121 2341 147
rect 2275 87 2291 121
rect 2325 87 2341 121
rect 2275 17 2341 87
rect 2493 116 2559 183
rect 2663 181 2729 197
rect 2819 232 2895 386
rect 2935 562 3001 649
rect 2935 528 2951 562
rect 2985 528 3001 562
rect 2935 491 3001 528
rect 2935 457 2951 491
rect 2985 457 3001 491
rect 2935 420 3001 457
rect 2935 386 2951 420
rect 2985 386 3001 420
rect 2935 370 3001 386
rect 3041 562 3145 578
rect 3041 528 3057 562
rect 3091 528 3145 562
rect 3041 491 3145 528
rect 3041 457 3057 491
rect 3091 457 3145 491
rect 3041 420 3145 457
rect 3041 386 3057 420
rect 3091 386 3145 420
rect 3041 370 3145 386
rect 2982 316 3048 332
rect 2982 282 2998 316
rect 3032 282 3048 316
rect 2982 248 3048 282
rect 2982 232 2998 248
rect 2819 214 2998 232
rect 3032 214 3048 248
rect 2819 198 3048 214
rect 2819 145 2853 198
rect 3097 145 3145 370
rect 2493 82 2509 116
rect 2543 82 2559 116
rect 2493 53 2559 82
rect 2651 116 2717 145
rect 2651 82 2667 116
rect 2701 82 2717 116
rect 2651 17 2717 82
rect 2763 116 2853 145
rect 2763 82 2779 116
rect 2813 82 2853 116
rect 2763 53 2853 82
rect 2921 116 2987 145
rect 2921 82 2937 116
rect 2971 82 2987 116
rect 2921 17 2987 82
rect 3079 116 3145 145
rect 3079 82 3095 116
rect 3129 82 3145 116
rect 3079 53 3145 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 1759 390 1793 424
rect 2431 390 2465 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
<< metal1 >>
rect 0 683 3168 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 0 617 3168 649
rect 1747 424 1805 430
rect 1747 390 1759 424
rect 1793 421 1805 424
rect 2419 424 2477 430
rect 2419 421 2431 424
rect 1793 393 2431 421
rect 1793 390 1805 393
rect 1747 384 1805 390
rect 2419 390 2431 393
rect 2465 390 2477 424
rect 2419 384 2477 390
rect 0 17 3168 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
rect 0 -49 3168 -17
<< labels >>
flabel pwell s 0 0 3168 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 3168 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfstp_lp
flabel metal1 s 2431 390 2465 424 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel metal1 s 0 617 3168 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 3168 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 3103 242 3137 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3103 316 3137 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3103 390 3137 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3103 464 3137 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3103 538 3137 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3168 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 173800
string GDS_START 152836
<< end >>
