magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
<< pwell >>
rect 292 241 1222 263
rect 16 49 1222 241
rect 0 0 1248 49
<< scnmos >>
rect 95 47 125 215
rect 181 47 211 215
rect 375 69 405 237
rect 461 69 491 237
rect 547 69 577 237
rect 633 69 663 237
rect 855 69 885 237
rect 941 69 971 237
rect 1027 69 1057 237
rect 1113 69 1143 237
<< scpmoshvt >>
rect 156 367 186 619
rect 242 367 272 619
rect 328 367 358 619
rect 447 367 477 619
rect 533 367 563 619
rect 735 367 765 619
rect 821 367 851 619
rect 941 367 971 619
rect 1027 367 1057 619
rect 1113 367 1143 619
<< ndiff >>
rect 42 203 95 215
rect 42 169 50 203
rect 84 169 95 203
rect 42 93 95 169
rect 42 59 50 93
rect 84 59 95 93
rect 42 47 95 59
rect 125 185 181 215
rect 125 151 136 185
rect 170 151 181 185
rect 125 101 181 151
rect 125 67 136 101
rect 170 67 181 101
rect 125 47 181 67
rect 211 132 264 215
rect 211 98 222 132
rect 256 98 264 132
rect 211 47 264 98
rect 318 124 375 237
rect 318 90 326 124
rect 360 90 375 124
rect 318 69 375 90
rect 405 229 461 237
rect 405 195 416 229
rect 450 195 461 229
rect 405 153 461 195
rect 405 119 416 153
rect 450 119 461 153
rect 405 69 461 119
rect 491 225 547 237
rect 491 191 502 225
rect 536 191 547 225
rect 491 115 547 191
rect 491 81 502 115
rect 536 81 547 115
rect 491 69 547 81
rect 577 183 633 237
rect 577 149 588 183
rect 622 149 633 183
rect 577 111 633 149
rect 577 77 588 111
rect 622 77 633 111
rect 577 69 633 77
rect 663 225 730 237
rect 663 191 688 225
rect 722 191 730 225
rect 663 153 730 191
rect 663 119 688 153
rect 722 119 730 153
rect 663 69 730 119
rect 788 225 855 237
rect 788 191 796 225
rect 830 191 855 225
rect 788 153 855 191
rect 788 119 796 153
rect 830 119 855 153
rect 788 69 855 119
rect 885 132 941 237
rect 885 98 896 132
rect 930 98 941 132
rect 885 69 941 98
rect 971 225 1027 237
rect 971 191 982 225
rect 1016 191 1027 225
rect 971 115 1027 191
rect 971 81 982 115
rect 1016 81 1027 115
rect 971 69 1027 81
rect 1057 183 1113 237
rect 1057 149 1068 183
rect 1102 149 1113 183
rect 1057 111 1113 149
rect 1057 77 1068 111
rect 1102 77 1113 111
rect 1057 69 1113 77
rect 1143 225 1196 237
rect 1143 191 1154 225
rect 1188 191 1196 225
rect 1143 115 1196 191
rect 1143 81 1154 115
rect 1188 81 1196 115
rect 1143 69 1196 81
<< pdiff >>
rect 103 599 156 619
rect 103 565 111 599
rect 145 565 156 599
rect 103 518 156 565
rect 103 484 111 518
rect 145 484 156 518
rect 103 434 156 484
rect 103 400 111 434
rect 145 400 156 434
rect 103 367 156 400
rect 186 545 242 619
rect 186 511 197 545
rect 231 511 242 545
rect 186 477 242 511
rect 186 443 197 477
rect 231 443 242 477
rect 186 409 242 443
rect 186 375 197 409
rect 231 375 242 409
rect 186 367 242 375
rect 272 611 328 619
rect 272 577 283 611
rect 317 577 328 611
rect 272 542 328 577
rect 272 508 283 542
rect 317 508 328 542
rect 272 474 328 508
rect 272 440 283 474
rect 317 440 328 474
rect 272 367 328 440
rect 358 607 447 619
rect 358 573 385 607
rect 419 573 447 607
rect 358 531 447 573
rect 358 497 385 531
rect 419 497 447 531
rect 358 367 447 497
rect 477 605 533 619
rect 477 571 488 605
rect 522 571 533 605
rect 477 535 533 571
rect 477 501 488 535
rect 522 501 533 535
rect 477 458 533 501
rect 477 424 488 458
rect 522 424 533 458
rect 477 367 533 424
rect 563 607 735 619
rect 563 573 590 607
rect 624 573 690 607
rect 724 573 735 607
rect 563 539 735 573
rect 563 505 590 539
rect 624 505 690 539
rect 724 505 735 539
rect 563 367 735 505
rect 765 599 821 619
rect 765 565 776 599
rect 810 565 821 599
rect 765 506 821 565
rect 765 472 776 506
rect 810 472 821 506
rect 765 413 821 472
rect 765 379 776 413
rect 810 379 821 413
rect 765 367 821 379
rect 851 607 941 619
rect 851 573 879 607
rect 913 573 941 607
rect 851 527 941 573
rect 851 493 879 527
rect 913 493 941 527
rect 851 445 941 493
rect 851 411 879 445
rect 913 411 941 445
rect 851 367 941 411
rect 971 599 1027 619
rect 971 565 982 599
rect 1016 565 1027 599
rect 971 506 1027 565
rect 971 472 982 506
rect 1016 472 1027 506
rect 971 413 1027 472
rect 971 379 982 413
rect 1016 379 1027 413
rect 971 367 1027 379
rect 1057 607 1113 619
rect 1057 573 1068 607
rect 1102 573 1113 607
rect 1057 494 1113 573
rect 1057 460 1068 494
rect 1102 460 1113 494
rect 1057 367 1113 460
rect 1143 599 1196 619
rect 1143 565 1154 599
rect 1188 565 1196 599
rect 1143 518 1196 565
rect 1143 484 1154 518
rect 1188 484 1196 518
rect 1143 435 1196 484
rect 1143 401 1154 435
rect 1188 401 1196 435
rect 1143 367 1196 401
<< ndiffc >>
rect 50 169 84 203
rect 50 59 84 93
rect 136 151 170 185
rect 136 67 170 101
rect 222 98 256 132
rect 326 90 360 124
rect 416 195 450 229
rect 416 119 450 153
rect 502 191 536 225
rect 502 81 536 115
rect 588 149 622 183
rect 588 77 622 111
rect 688 191 722 225
rect 688 119 722 153
rect 796 191 830 225
rect 796 119 830 153
rect 896 98 930 132
rect 982 191 1016 225
rect 982 81 1016 115
rect 1068 149 1102 183
rect 1068 77 1102 111
rect 1154 191 1188 225
rect 1154 81 1188 115
<< pdiffc >>
rect 111 565 145 599
rect 111 484 145 518
rect 111 400 145 434
rect 197 511 231 545
rect 197 443 231 477
rect 197 375 231 409
rect 283 577 317 611
rect 283 508 317 542
rect 283 440 317 474
rect 385 573 419 607
rect 385 497 419 531
rect 488 571 522 605
rect 488 501 522 535
rect 488 424 522 458
rect 590 573 624 607
rect 690 573 724 607
rect 590 505 624 539
rect 690 505 724 539
rect 776 565 810 599
rect 776 472 810 506
rect 776 379 810 413
rect 879 573 913 607
rect 879 493 913 527
rect 879 411 913 445
rect 982 565 1016 599
rect 982 472 1016 506
rect 982 379 1016 413
rect 1068 573 1102 607
rect 1068 460 1102 494
rect 1154 565 1188 599
rect 1154 484 1188 518
rect 1154 401 1188 435
<< poly >>
rect 156 619 186 645
rect 242 619 272 645
rect 328 619 358 645
rect 447 619 477 645
rect 533 619 563 645
rect 735 619 765 645
rect 821 619 851 645
rect 941 619 971 645
rect 1027 619 1057 645
rect 1113 619 1143 645
rect 156 303 186 367
rect 242 303 272 367
rect 328 325 358 367
rect 447 325 477 367
rect 95 287 272 303
rect 95 253 111 287
rect 145 253 272 287
rect 314 309 477 325
rect 314 275 330 309
rect 364 289 477 309
rect 533 335 563 367
rect 735 335 765 367
rect 533 319 765 335
rect 364 275 491 289
rect 314 259 491 275
rect 533 285 619 319
rect 653 285 687 319
rect 721 285 765 319
rect 533 269 765 285
rect 821 325 851 367
rect 941 325 971 367
rect 821 309 971 325
rect 821 275 837 309
rect 871 275 907 309
rect 941 275 971 309
rect 95 237 272 253
rect 375 237 405 259
rect 461 237 491 259
rect 547 237 577 269
rect 633 237 663 269
rect 821 259 971 275
rect 855 237 885 259
rect 941 237 971 259
rect 1027 335 1057 367
rect 1113 335 1143 367
rect 1027 319 1143 335
rect 1027 285 1068 319
rect 1102 285 1143 319
rect 1027 269 1143 285
rect 1027 237 1057 269
rect 1113 237 1143 269
rect 95 215 125 237
rect 181 215 211 237
rect 95 21 125 47
rect 181 21 211 47
rect 375 43 405 69
rect 461 43 491 69
rect 547 43 577 69
rect 633 43 663 69
rect 855 43 885 69
rect 941 43 971 69
rect 1027 43 1057 69
rect 1113 43 1143 69
<< polycont >>
rect 111 253 145 287
rect 330 275 364 309
rect 619 285 653 319
rect 687 285 721 319
rect 837 275 871 309
rect 907 275 941 309
rect 1068 285 1102 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 95 611 333 615
rect 95 599 283 611
rect 95 565 111 599
rect 145 579 283 599
rect 145 565 147 579
rect 267 577 283 579
rect 317 577 333 611
rect 95 518 147 565
rect 95 484 111 518
rect 145 484 147 518
rect 95 434 147 484
rect 95 400 111 434
rect 145 400 147 434
rect 95 384 147 400
rect 181 511 197 545
rect 231 511 247 545
rect 181 477 247 511
rect 181 443 197 477
rect 231 443 247 477
rect 181 409 247 443
rect 281 542 333 577
rect 281 508 283 542
rect 317 508 333 542
rect 281 474 333 508
rect 369 607 435 649
rect 369 573 385 607
rect 419 573 435 607
rect 369 531 435 573
rect 369 497 385 531
rect 419 497 435 531
rect 369 492 435 497
rect 472 605 538 615
rect 472 571 488 605
rect 522 571 538 605
rect 472 535 538 571
rect 472 501 488 535
rect 522 501 538 535
rect 572 607 740 649
rect 572 573 590 607
rect 624 573 690 607
rect 724 573 740 607
rect 572 539 740 573
rect 572 505 590 539
rect 624 505 690 539
rect 724 505 740 539
rect 572 501 740 505
rect 774 599 826 615
rect 774 565 776 599
rect 810 565 826 599
rect 774 506 826 565
rect 281 440 283 474
rect 317 458 333 474
rect 472 465 538 501
rect 774 472 776 506
rect 810 472 826 506
rect 774 465 826 472
rect 472 458 826 465
rect 317 440 488 458
rect 281 424 488 440
rect 522 424 826 458
rect 181 378 197 409
rect 195 375 197 378
rect 231 390 247 409
rect 771 413 826 424
rect 231 375 560 390
rect 195 356 560 375
rect 771 379 776 413
rect 810 379 826 413
rect 863 607 929 649
rect 863 573 879 607
rect 913 573 929 607
rect 863 527 929 573
rect 863 493 879 527
rect 913 493 929 527
rect 863 445 929 493
rect 863 411 879 445
rect 913 411 929 445
rect 966 599 1018 615
rect 966 565 982 599
rect 1016 565 1018 599
rect 966 506 1018 565
rect 966 472 982 506
rect 1016 472 1018 506
rect 966 419 1018 472
rect 1052 607 1118 649
rect 1052 573 1068 607
rect 1102 573 1118 607
rect 1052 494 1118 573
rect 1052 460 1068 494
rect 1102 460 1118 494
rect 1052 453 1118 460
rect 1152 599 1204 615
rect 1152 565 1154 599
rect 1188 565 1204 599
rect 1152 518 1204 565
rect 1152 484 1154 518
rect 1188 484 1204 518
rect 1152 435 1204 484
rect 1152 419 1154 435
rect 966 413 1154 419
rect 771 377 826 379
rect 966 379 982 413
rect 1016 401 1154 413
rect 1188 401 1204 435
rect 1016 385 1204 401
rect 966 377 1016 379
rect 17 287 161 350
rect 17 253 111 287
rect 145 253 161 287
rect 17 242 161 253
rect 223 309 380 322
rect 223 275 330 309
rect 364 275 380 309
rect 223 242 380 275
rect 414 285 560 356
rect 594 319 737 366
rect 771 343 1016 377
rect 594 285 619 319
rect 653 285 687 319
rect 721 285 737 319
rect 1050 319 1231 350
rect 414 229 466 285
rect 821 275 837 309
rect 871 275 907 309
rect 941 275 957 309
rect 1050 285 1068 319
rect 1102 285 1231 319
rect 414 208 416 229
rect 34 203 100 208
rect 34 169 50 203
rect 84 169 100 203
rect 34 93 100 169
rect 34 59 50 93
rect 84 59 100 93
rect 34 17 100 59
rect 134 195 416 208
rect 450 195 466 229
rect 134 185 466 195
rect 134 151 136 185
rect 170 174 466 185
rect 170 151 172 174
rect 134 101 172 151
rect 400 153 466 174
rect 134 67 136 101
rect 170 67 172 101
rect 134 51 172 67
rect 206 132 272 140
rect 206 98 222 132
rect 256 98 272 132
rect 206 17 272 98
rect 310 124 366 140
rect 310 90 326 124
rect 360 90 366 124
rect 400 119 416 153
rect 450 119 466 153
rect 500 225 738 251
rect 880 242 946 275
rect 500 191 502 225
rect 536 217 688 225
rect 536 191 538 217
rect 310 85 366 90
rect 500 115 538 191
rect 672 191 688 217
rect 722 191 738 225
rect 500 85 502 115
rect 310 81 502 85
rect 536 81 538 115
rect 310 51 538 81
rect 572 149 588 183
rect 622 149 638 183
rect 572 111 638 149
rect 672 153 738 191
rect 672 119 688 153
rect 722 119 738 153
rect 780 225 846 241
rect 780 191 796 225
rect 830 208 846 225
rect 982 225 1204 251
rect 830 191 982 208
rect 1016 217 1154 225
rect 1016 191 1018 217
rect 780 174 1018 191
rect 1152 191 1154 217
rect 1188 191 1204 225
rect 780 153 846 174
rect 780 119 796 153
rect 830 119 846 153
rect 880 132 946 140
rect 572 77 588 111
rect 622 85 638 111
rect 880 98 896 132
rect 930 98 946 132
rect 880 85 946 98
rect 622 77 946 85
rect 572 51 946 77
rect 980 115 1018 174
rect 980 81 982 115
rect 1016 81 1018 115
rect 980 65 1018 81
rect 1052 149 1068 183
rect 1102 149 1118 183
rect 1052 111 1118 149
rect 1052 77 1068 111
rect 1102 77 1118 111
rect 1052 17 1118 77
rect 1152 115 1204 191
rect 1152 81 1154 115
rect 1188 81 1204 115
rect 1152 65 1204 81
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a41oi_2
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1384452
string GDS_START 1373328
<< end >>
