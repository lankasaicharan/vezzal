magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3506 1975
<< nwell >>
rect -38 331 2246 704
<< pwell >>
rect 599 229 829 235
rect 1725 233 2207 251
rect 599 223 1056 229
rect 31 199 1056 223
rect 1402 199 2207 233
rect 31 49 2207 199
rect 0 0 2208 49
<< scnmos >>
rect 114 113 144 197
rect 186 113 216 197
rect 400 113 430 197
rect 478 113 508 197
rect 580 113 610 197
rect 723 125 753 209
rect 825 66 855 150
rect 943 119 973 203
rect 1215 89 1245 173
rect 1287 89 1317 173
rect 1495 123 1525 207
rect 1587 123 1617 207
rect 1830 141 1860 225
rect 1902 141 1932 225
rect 2016 141 2046 225
rect 2094 141 2124 225
<< scpmoshvt >>
rect 126 419 176 619
rect 338 419 388 619
rect 444 419 494 619
rect 657 419 707 619
rect 831 419 881 619
rect 939 419 989 619
rect 1175 396 1225 596
rect 1409 406 1459 606
rect 1515 406 1565 606
rect 1808 413 1858 613
rect 1980 413 2030 613
<< ndiff >>
rect 625 197 723 209
rect 57 172 114 197
rect 57 138 69 172
rect 103 138 114 172
rect 57 113 114 138
rect 144 113 186 197
rect 216 163 400 197
rect 216 129 227 163
rect 261 129 400 163
rect 216 113 400 129
rect 430 113 478 197
rect 508 172 580 197
rect 508 138 519 172
rect 553 138 580 172
rect 508 113 580 138
rect 610 185 723 197
rect 610 151 637 185
rect 671 151 723 185
rect 610 125 723 151
rect 753 150 803 209
rect 870 191 943 203
rect 870 157 882 191
rect 916 157 943 191
rect 870 150 943 157
rect 753 125 825 150
rect 610 113 683 125
rect 768 116 825 125
rect 768 82 780 116
rect 814 82 825 116
rect 768 66 825 82
rect 855 119 943 150
rect 973 178 1030 203
rect 973 144 984 178
rect 1018 144 1030 178
rect 1428 182 1495 207
rect 973 119 1030 144
rect 1158 148 1215 173
rect 855 112 928 119
rect 855 78 882 112
rect 916 78 928 112
rect 855 66 928 78
rect 1158 114 1170 148
rect 1204 114 1215 148
rect 1158 89 1215 114
rect 1245 89 1287 173
rect 1317 148 1374 173
rect 1317 114 1328 148
rect 1362 114 1374 148
rect 1428 148 1440 182
rect 1474 148 1495 182
rect 1428 123 1495 148
rect 1525 182 1587 207
rect 1525 148 1542 182
rect 1576 148 1587 182
rect 1525 123 1587 148
rect 1617 184 1690 207
rect 1617 150 1644 184
rect 1678 150 1690 184
rect 1617 123 1690 150
rect 1751 200 1830 225
rect 1751 166 1763 200
rect 1797 166 1830 200
rect 1751 141 1830 166
rect 1860 141 1902 225
rect 1932 194 2016 225
rect 1932 160 1971 194
rect 2005 160 2016 194
rect 1932 141 2016 160
rect 2046 141 2094 225
rect 2124 200 2181 225
rect 2124 166 2135 200
rect 2169 166 2181 200
rect 2124 141 2181 166
rect 1317 89 1374 114
<< pdiff >>
rect 69 597 126 619
rect 69 563 81 597
rect 115 563 126 597
rect 69 465 126 563
rect 69 431 81 465
rect 115 431 126 465
rect 69 419 126 431
rect 176 596 338 619
rect 176 562 187 596
rect 221 562 338 596
rect 176 419 338 562
rect 388 496 444 619
rect 388 462 399 496
rect 433 462 444 496
rect 388 419 444 462
rect 494 496 657 619
rect 494 462 505 496
rect 539 462 657 496
rect 494 419 657 462
rect 707 566 831 619
rect 707 532 718 566
rect 752 532 831 566
rect 707 419 831 532
rect 881 519 939 619
rect 881 485 894 519
rect 928 485 939 519
rect 881 419 939 485
rect 989 496 1046 619
rect 989 462 1000 496
rect 1034 462 1046 496
rect 989 419 1046 462
rect 1100 527 1175 596
rect 1100 493 1112 527
rect 1146 493 1175 527
rect 1100 442 1175 493
rect 1100 408 1112 442
rect 1146 408 1175 442
rect 1100 396 1175 408
rect 1225 584 1298 596
rect 1225 550 1252 584
rect 1286 550 1298 584
rect 1225 513 1298 550
rect 1225 479 1252 513
rect 1286 479 1298 513
rect 1225 442 1298 479
rect 1225 408 1252 442
rect 1286 408 1298 442
rect 1225 396 1298 408
rect 1352 594 1409 606
rect 1352 560 1364 594
rect 1398 560 1409 594
rect 1352 523 1409 560
rect 1352 489 1364 523
rect 1398 489 1409 523
rect 1352 452 1409 489
rect 1352 418 1364 452
rect 1398 418 1409 452
rect 1352 406 1409 418
rect 1459 594 1515 606
rect 1459 560 1470 594
rect 1504 560 1515 594
rect 1459 523 1515 560
rect 1459 489 1470 523
rect 1504 489 1515 523
rect 1459 452 1515 489
rect 1459 418 1470 452
rect 1504 418 1515 452
rect 1459 406 1515 418
rect 1565 527 1622 606
rect 1565 493 1576 527
rect 1610 493 1622 527
rect 1565 452 1622 493
rect 1565 418 1576 452
rect 1610 418 1622 452
rect 1565 406 1622 418
rect 1751 527 1808 613
rect 1751 493 1763 527
rect 1797 493 1808 527
rect 1751 459 1808 493
rect 1751 425 1763 459
rect 1797 425 1808 459
rect 1751 413 1808 425
rect 1858 601 1980 613
rect 1858 567 1935 601
rect 1969 567 1980 601
rect 1858 469 1980 567
rect 1858 435 1935 469
rect 1969 435 1980 469
rect 1858 413 1980 435
rect 2030 597 2087 613
rect 2030 563 2041 597
rect 2075 563 2087 597
rect 2030 469 2087 563
rect 2030 435 2041 469
rect 2075 435 2087 469
rect 2030 413 2087 435
<< ndiffc >>
rect 69 138 103 172
rect 227 129 261 163
rect 519 138 553 172
rect 637 151 671 185
rect 882 157 916 191
rect 780 82 814 116
rect 984 144 1018 178
rect 882 78 916 112
rect 1170 114 1204 148
rect 1328 114 1362 148
rect 1440 148 1474 182
rect 1542 148 1576 182
rect 1644 150 1678 184
rect 1763 166 1797 200
rect 1971 160 2005 194
rect 2135 166 2169 200
<< pdiffc >>
rect 81 563 115 597
rect 81 431 115 465
rect 187 562 221 596
rect 399 462 433 496
rect 505 462 539 496
rect 718 532 752 566
rect 894 485 928 519
rect 1000 462 1034 496
rect 1112 493 1146 527
rect 1112 408 1146 442
rect 1252 550 1286 584
rect 1252 479 1286 513
rect 1252 408 1286 442
rect 1364 560 1398 594
rect 1364 489 1398 523
rect 1364 418 1398 452
rect 1470 560 1504 594
rect 1470 489 1504 523
rect 1470 418 1504 452
rect 1576 493 1610 527
rect 1576 418 1610 452
rect 1763 493 1797 527
rect 1763 425 1797 459
rect 1935 567 1969 601
rect 1935 435 1969 469
rect 2041 563 2075 597
rect 2041 435 2075 469
<< poly >>
rect 126 619 176 645
rect 338 619 388 645
rect 444 619 494 645
rect 657 619 707 645
rect 831 619 881 645
rect 939 619 989 645
rect 1175 596 1225 622
rect 1409 606 1459 632
rect 1515 606 1565 632
rect 1808 613 1858 639
rect 1980 613 2030 639
rect 126 387 176 419
rect 114 371 233 387
rect 114 337 183 371
rect 217 337 233 371
rect 114 321 233 337
rect 114 197 144 321
rect 186 197 216 321
rect 338 285 388 419
rect 444 379 494 419
rect 444 363 609 379
rect 657 375 707 419
rect 444 329 559 363
rect 593 329 609 363
rect 444 313 609 329
rect 651 345 707 375
rect 831 379 881 419
rect 939 391 989 419
rect 831 363 897 379
rect 281 269 388 285
rect 281 235 297 269
rect 331 249 388 269
rect 651 254 681 345
rect 831 329 847 363
rect 881 329 897 363
rect 831 313 897 329
rect 959 356 989 391
rect 959 340 1127 356
rect 959 326 1077 340
rect 331 235 508 249
rect 281 219 508 235
rect 400 197 430 219
rect 478 197 508 219
rect 580 224 681 254
rect 723 281 789 297
rect 723 247 739 281
rect 773 247 789 281
rect 723 231 789 247
rect 867 248 897 313
rect 1061 306 1077 326
rect 1111 306 1127 340
rect 1061 290 1127 306
rect 1175 248 1225 396
rect 1409 366 1459 406
rect 1515 391 1565 406
rect 1808 391 1858 413
rect 1393 350 1459 366
rect 1393 316 1409 350
rect 1443 316 1459 350
rect 1393 300 1459 316
rect 1501 361 1896 391
rect 1501 252 1531 361
rect 1866 313 1896 361
rect 1980 381 2030 413
rect 1980 365 2093 381
rect 1980 331 2043 365
rect 2077 331 2093 365
rect 580 197 610 224
rect 723 209 753 231
rect 867 218 1317 248
rect 943 203 973 218
rect 825 150 855 176
rect 114 87 144 113
rect 186 87 216 113
rect 400 87 430 113
rect 478 87 508 113
rect 580 51 610 113
rect 723 99 753 125
rect 1215 173 1245 218
rect 1287 173 1317 218
rect 1495 222 1531 252
rect 1573 297 1639 313
rect 1573 263 1589 297
rect 1623 277 1639 297
rect 1706 297 1788 313
rect 1706 277 1738 297
rect 1623 263 1738 277
rect 1772 263 1788 297
rect 1866 297 1932 313
rect 1866 277 1882 297
rect 1573 247 1788 263
rect 1830 263 1882 277
rect 1916 263 1932 297
rect 1830 247 1932 263
rect 1980 297 2093 331
rect 1980 263 2043 297
rect 2077 277 2093 297
rect 2077 263 2124 277
rect 1980 247 2124 263
rect 1495 207 1525 222
rect 1587 207 1617 247
rect 1830 225 1860 247
rect 1902 225 1932 247
rect 2016 225 2046 247
rect 2094 225 2124 247
rect 943 93 973 119
rect 1070 103 1136 119
rect 1070 69 1086 103
rect 1120 69 1136 103
rect 1495 97 1525 123
rect 1587 97 1617 123
rect 1830 115 1860 141
rect 1902 115 1932 141
rect 2016 119 2046 141
rect 1974 103 2046 119
rect 2094 115 2124 141
rect 825 51 855 66
rect 1070 51 1136 69
rect 1215 63 1245 89
rect 1287 63 1317 89
rect 1974 69 1990 103
rect 2024 69 2046 103
rect 1974 53 2046 69
rect 580 21 1136 51
<< polycont >>
rect 183 337 217 371
rect 559 329 593 363
rect 297 235 331 269
rect 847 329 881 363
rect 739 247 773 281
rect 1077 306 1111 340
rect 1409 316 1443 350
rect 2043 331 2077 365
rect 1589 263 1623 297
rect 1738 263 1772 297
rect 1882 263 1916 297
rect 2043 263 2077 297
rect 1086 69 1120 103
rect 1990 69 2024 103
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 53 597 131 613
rect 53 563 81 597
rect 115 563 131 597
rect 53 500 131 563
rect 171 596 237 649
rect 171 562 187 596
rect 221 562 237 596
rect 171 536 237 562
rect 273 579 768 613
rect 273 500 307 579
rect 702 566 768 579
rect 53 466 307 500
rect 383 496 449 543
rect 53 465 131 466
rect 53 431 81 465
rect 115 431 131 465
rect 53 285 131 431
rect 383 462 399 496
rect 433 462 449 496
rect 167 371 263 430
rect 167 337 183 371
rect 217 337 263 371
rect 167 321 263 337
rect 53 269 347 285
rect 53 235 297 269
rect 331 235 347 269
rect 53 219 347 235
rect 53 172 119 219
rect 53 138 69 172
rect 103 138 119 172
rect 53 109 119 138
rect 211 163 277 183
rect 211 129 227 163
rect 261 129 277 163
rect 211 17 277 129
rect 313 87 347 219
rect 383 202 449 462
rect 485 496 555 543
rect 485 462 505 496
rect 539 462 555 496
rect 702 532 718 566
rect 752 532 768 566
rect 702 485 768 532
rect 804 579 1216 613
rect 485 449 555 462
rect 804 449 838 579
rect 878 519 955 543
rect 878 485 894 519
rect 928 498 955 519
rect 878 464 895 485
rect 929 464 955 498
rect 878 462 955 464
rect 485 415 838 449
rect 485 271 519 415
rect 555 363 885 379
rect 555 329 559 363
rect 593 329 847 363
rect 881 329 885 363
rect 555 313 885 329
rect 555 310 647 313
rect 723 281 789 313
rect 485 237 687 271
rect 383 168 415 202
rect 449 172 569 201
rect 449 168 519 172
rect 383 162 519 168
rect 503 138 519 162
rect 553 138 569 172
rect 503 125 569 138
rect 621 185 687 237
rect 723 247 739 281
rect 773 247 789 281
rect 921 277 955 462
rect 723 231 789 247
rect 866 243 955 277
rect 991 496 1050 543
rect 991 462 1000 496
rect 1034 462 1050 496
rect 991 392 1050 462
rect 1096 527 1146 543
rect 1096 493 1112 527
rect 1096 442 1146 493
rect 1096 408 1112 442
rect 621 151 637 185
rect 671 151 687 185
rect 621 123 687 151
rect 866 207 900 243
rect 991 208 1025 392
rect 1096 356 1146 408
rect 1061 340 1146 356
rect 1061 306 1077 340
rect 1111 306 1146 340
rect 1061 290 1146 306
rect 991 207 1034 208
rect 866 191 932 207
rect 866 157 882 191
rect 916 157 932 191
rect 764 116 830 137
rect 764 87 780 116
rect 313 82 780 87
rect 814 82 830 116
rect 313 53 830 82
rect 866 112 932 157
rect 968 202 1034 207
rect 968 178 991 202
rect 968 144 984 178
rect 1025 168 1034 202
rect 1018 144 1034 168
rect 968 115 1034 144
rect 1112 177 1146 290
rect 1182 264 1216 579
rect 1252 584 1286 649
rect 1252 513 1286 550
rect 1252 442 1286 479
rect 1252 392 1286 408
rect 1323 594 1414 610
rect 1323 560 1364 594
rect 1398 560 1414 594
rect 1323 523 1414 560
rect 1323 489 1364 523
rect 1398 489 1414 523
rect 1323 452 1414 489
rect 1323 418 1364 452
rect 1398 418 1414 452
rect 1323 402 1414 418
rect 1454 594 1883 613
rect 1454 560 1470 594
rect 1504 579 1883 594
rect 1504 560 1520 579
rect 1454 523 1520 560
rect 1454 489 1470 523
rect 1504 489 1520 523
rect 1454 452 1520 489
rect 1454 418 1470 452
rect 1504 418 1520 452
rect 1454 402 1520 418
rect 1560 527 1697 543
rect 1560 498 1576 527
rect 1560 464 1567 498
rect 1610 493 1697 527
rect 1601 464 1697 493
rect 1560 452 1697 464
rect 1560 418 1576 452
rect 1610 418 1697 452
rect 1560 402 1697 418
rect 1323 264 1357 402
rect 1393 350 1528 366
rect 1393 316 1409 350
rect 1443 316 1528 350
rect 1393 313 1528 316
rect 1393 300 1627 313
rect 1494 297 1627 300
rect 1182 230 1458 264
rect 1494 263 1589 297
rect 1623 263 1627 297
rect 1494 247 1627 263
rect 1424 211 1458 230
rect 1663 211 1697 402
rect 1424 182 1490 211
rect 1112 148 1220 177
rect 1112 119 1170 148
rect 866 78 882 112
rect 916 78 932 112
rect 866 62 932 78
rect 1070 114 1170 119
rect 1204 114 1220 148
rect 1070 103 1220 114
rect 1070 69 1086 103
rect 1120 85 1220 103
rect 1312 148 1378 177
rect 1312 114 1328 148
rect 1362 114 1378 148
rect 1424 148 1440 182
rect 1474 148 1490 182
rect 1424 119 1490 148
rect 1526 182 1592 211
rect 1526 148 1542 182
rect 1576 148 1592 182
rect 1120 69 1146 85
rect 1070 53 1146 69
rect 1312 17 1378 114
rect 1526 87 1592 148
rect 1628 184 1697 211
rect 1628 150 1644 184
rect 1678 150 1697 184
rect 1628 123 1697 150
rect 1733 527 1813 543
rect 1733 493 1763 527
rect 1797 493 1813 527
rect 1733 459 1813 493
rect 1733 425 1763 459
rect 1797 425 1813 459
rect 1733 297 1813 425
rect 1849 383 1883 579
rect 1919 601 1985 649
rect 1919 567 1935 601
rect 1969 567 1985 601
rect 1919 469 1985 567
rect 1919 435 1935 469
rect 1969 435 1985 469
rect 1919 419 1985 435
rect 2025 597 2091 613
rect 2025 563 2041 597
rect 2075 563 2091 597
rect 2025 469 2091 563
rect 2025 435 2041 469
rect 2075 453 2091 469
rect 2135 453 2185 578
rect 2075 435 2185 453
rect 2025 419 2185 435
rect 1849 365 2093 383
rect 1849 349 2043 365
rect 2027 331 2043 349
rect 2077 331 2093 365
rect 1733 263 1738 297
rect 1772 263 1813 297
rect 1733 200 1813 263
rect 1849 297 1991 313
rect 1849 263 1882 297
rect 1916 263 1991 297
rect 1849 236 1991 263
rect 2027 297 2093 331
rect 2027 263 2043 297
rect 2077 263 2093 297
rect 2027 247 2093 263
rect 2135 200 2185 419
rect 1733 166 1763 200
rect 1797 166 1813 200
rect 1733 137 1813 166
rect 1955 194 2099 200
rect 1955 160 1971 194
rect 2005 160 2099 194
rect 1955 155 2099 160
rect 1974 103 2029 119
rect 1974 87 1990 103
rect 1526 69 1990 87
rect 2024 69 2029 103
rect 1526 53 2029 69
rect 2065 17 2099 155
rect 2169 166 2185 200
rect 2135 137 2185 166
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 895 485 928 498
rect 928 485 929 498
rect 895 464 929 485
rect 415 168 449 202
rect 991 178 1025 202
rect 991 168 1018 178
rect 1018 168 1025 178
rect 1567 493 1576 498
rect 1576 493 1601 498
rect 1567 464 1601 493
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 883 498 941 504
rect 883 464 895 498
rect 929 495 941 498
rect 1555 498 1613 504
rect 1555 495 1567 498
rect 929 467 1567 495
rect 929 464 941 467
rect 883 458 941 464
rect 1555 464 1567 467
rect 1601 464 1613 498
rect 1555 458 1613 464
rect 403 202 461 208
rect 403 168 415 202
rect 449 199 461 202
rect 979 202 1037 208
rect 979 199 991 202
rect 449 171 991 199
rect 449 168 461 171
rect 403 162 461 168
rect 979 168 991 171
rect 1025 168 1037 202
rect 979 162 1037 168
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xor3_lp
flabel comment s 2046 261 2046 261 0 FreeSans 200 180 0 0 no_jumper_check
flabel comment s 1664 261 1664 261 0 FreeSans 200 180 0 0 no_jumper_check
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 2143 242 2177 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 2143 316 2177 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 2143 390 2177 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 2143 464 2177 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 2143 538 2177 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4647838
string GDS_START 4633234
<< end >>
