magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 60 49 644 167
rect 0 0 672 49
<< scnmos >>
rect 143 57 173 141
rect 215 57 245 141
rect 301 57 331 141
rect 373 57 403 141
rect 459 57 489 141
rect 531 57 561 141
<< scpmoshvt >>
rect 247 409 297 609
rect 345 409 395 609
rect 459 409 509 609
<< ndiff >>
rect 86 116 143 141
rect 86 82 98 116
rect 132 82 143 116
rect 86 57 143 82
rect 173 57 215 141
rect 245 108 301 141
rect 245 74 256 108
rect 290 74 301 108
rect 245 57 301 74
rect 331 57 373 141
rect 403 116 459 141
rect 403 82 414 116
rect 448 82 459 116
rect 403 57 459 82
rect 489 57 531 141
rect 561 116 618 141
rect 561 82 572 116
rect 606 82 618 116
rect 561 57 618 82
<< pdiff >>
rect 190 597 247 609
rect 190 563 202 597
rect 236 563 247 597
rect 190 526 247 563
rect 190 492 202 526
rect 236 492 247 526
rect 190 455 247 492
rect 190 421 202 455
rect 236 421 247 455
rect 190 409 247 421
rect 297 409 345 609
rect 395 409 459 609
rect 509 597 566 609
rect 509 563 520 597
rect 554 563 566 597
rect 509 526 566 563
rect 509 492 520 526
rect 554 492 566 526
rect 509 455 566 492
rect 509 421 520 455
rect 554 421 566 455
rect 509 409 566 421
<< ndiffc >>
rect 98 82 132 116
rect 256 74 290 108
rect 414 82 448 116
rect 572 82 606 116
<< pdiffc >>
rect 202 563 236 597
rect 202 492 236 526
rect 202 421 236 455
rect 520 563 554 597
rect 520 492 554 526
rect 520 421 554 455
<< poly >>
rect 247 609 297 635
rect 345 609 395 635
rect 459 609 509 635
rect 247 369 297 409
rect 345 370 395 409
rect 459 383 509 409
rect 211 353 277 369
rect 211 319 227 353
rect 261 319 277 353
rect 211 285 277 319
rect 211 265 227 285
rect 143 251 227 265
rect 261 251 277 285
rect 143 235 277 251
rect 345 354 411 370
rect 345 320 361 354
rect 395 320 411 354
rect 345 286 411 320
rect 345 252 361 286
rect 395 252 411 286
rect 345 236 411 252
rect 459 335 489 383
rect 459 319 571 335
rect 459 285 521 319
rect 555 285 571 319
rect 459 251 571 285
rect 143 141 173 235
rect 215 141 245 235
rect 345 186 375 236
rect 459 217 521 251
rect 555 217 571 251
rect 459 201 571 217
rect 301 156 403 186
rect 301 141 331 156
rect 373 141 403 156
rect 459 141 489 201
rect 531 141 561 201
rect 143 31 173 57
rect 215 31 245 57
rect 301 31 331 57
rect 373 31 403 57
rect 459 31 489 57
rect 531 31 561 57
<< polycont >>
rect 227 319 261 353
rect 227 251 261 285
rect 361 320 395 354
rect 361 252 395 286
rect 521 285 555 319
rect 521 217 555 251
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 186 597 252 613
rect 186 578 202 597
rect 25 563 202 578
rect 236 563 252 597
rect 504 597 570 649
rect 25 526 252 563
rect 25 492 202 526
rect 236 492 252 526
rect 25 455 252 492
rect 25 421 202 455
rect 236 421 252 455
rect 25 405 252 421
rect 25 236 167 405
rect 82 199 167 236
rect 211 353 277 369
rect 211 319 227 353
rect 261 319 277 353
rect 211 285 277 319
rect 211 251 227 285
rect 261 251 277 285
rect 211 235 277 251
rect 313 354 455 578
rect 504 563 520 597
rect 554 563 570 597
rect 504 526 570 563
rect 504 492 520 526
rect 554 492 570 526
rect 504 455 570 492
rect 504 421 520 455
rect 554 421 570 455
rect 504 405 570 421
rect 313 320 361 354
rect 395 320 455 354
rect 313 286 455 320
rect 313 252 361 286
rect 395 252 455 286
rect 313 236 455 252
rect 505 319 647 356
rect 505 285 521 319
rect 555 285 647 319
rect 505 251 647 285
rect 505 217 521 251
rect 555 217 647 251
rect 505 201 647 217
rect 82 165 432 199
rect 82 116 148 165
rect 398 145 432 165
rect 82 82 98 116
rect 132 82 148 116
rect 82 53 148 82
rect 240 108 306 129
rect 240 74 256 108
rect 290 74 306 108
rect 240 17 306 74
rect 398 116 464 145
rect 398 82 414 116
rect 448 82 464 116
rect 398 53 464 82
rect 556 116 622 145
rect 556 82 572 116
rect 606 82 622 116
rect 556 17 622 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor3_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2507026
string GDS_START 2499272
<< end >>
