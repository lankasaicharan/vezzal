magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 760 241
rect 0 0 768 49
<< scnmos >>
rect 80 47 110 215
rect 233 47 263 215
rect 326 47 356 215
rect 423 47 453 215
rect 579 47 609 215
rect 651 47 681 215
<< scpmoshvt >>
rect 118 367 148 619
rect 219 367 249 619
rect 305 367 335 619
rect 471 367 501 619
rect 557 367 587 619
rect 651 367 681 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 101 80 169
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 137 233 215
rect 110 103 188 137
rect 222 103 233 137
rect 110 93 233 103
rect 110 59 121 93
rect 155 59 233 93
rect 110 47 233 59
rect 263 47 326 215
rect 356 47 423 215
rect 453 203 579 215
rect 453 169 464 203
rect 498 169 534 203
rect 568 169 579 203
rect 453 93 579 169
rect 453 59 464 93
rect 498 59 534 93
rect 568 59 579 93
rect 453 47 579 59
rect 609 47 651 215
rect 681 203 734 215
rect 681 169 692 203
rect 726 169 734 203
rect 681 93 734 169
rect 681 59 692 93
rect 726 59 734 93
rect 681 47 734 59
<< pdiff >>
rect 65 599 118 619
rect 65 565 73 599
rect 107 565 118 599
rect 65 520 118 565
rect 65 486 73 520
rect 107 486 118 520
rect 65 420 118 486
rect 65 386 73 420
rect 107 386 118 420
rect 65 367 118 386
rect 148 607 219 619
rect 148 573 160 607
rect 194 573 219 607
rect 148 532 219 573
rect 148 498 160 532
rect 194 498 219 532
rect 148 455 219 498
rect 148 421 160 455
rect 194 421 219 455
rect 148 367 219 421
rect 249 597 305 619
rect 249 563 260 597
rect 294 563 305 597
rect 249 522 305 563
rect 249 488 260 522
rect 294 488 305 522
rect 249 443 305 488
rect 249 409 260 443
rect 294 409 305 443
rect 249 367 305 409
rect 335 607 471 619
rect 335 573 346 607
rect 380 573 426 607
rect 460 573 471 607
rect 335 517 471 573
rect 335 483 346 517
rect 380 483 426 517
rect 460 483 471 517
rect 335 367 471 483
rect 501 599 557 619
rect 501 565 512 599
rect 546 565 557 599
rect 501 529 557 565
rect 501 495 512 529
rect 546 495 557 529
rect 501 461 557 495
rect 501 427 512 461
rect 546 427 557 461
rect 501 367 557 427
rect 587 543 651 619
rect 587 509 600 543
rect 634 509 651 543
rect 587 413 651 509
rect 587 379 600 413
rect 634 379 651 413
rect 587 367 651 379
rect 681 599 734 619
rect 681 565 692 599
rect 726 565 734 599
rect 681 517 734 565
rect 681 483 692 517
rect 726 483 734 517
rect 681 436 734 483
rect 681 402 692 436
rect 726 402 734 436
rect 681 367 734 402
<< ndiffc >>
rect 35 169 69 203
rect 35 67 69 101
rect 188 103 222 137
rect 121 59 155 93
rect 464 169 498 203
rect 534 169 568 203
rect 464 59 498 93
rect 534 59 568 93
rect 692 169 726 203
rect 692 59 726 93
<< pdiffc >>
rect 73 565 107 599
rect 73 486 107 520
rect 73 386 107 420
rect 160 573 194 607
rect 160 498 194 532
rect 160 421 194 455
rect 260 563 294 597
rect 260 488 294 522
rect 260 409 294 443
rect 346 573 380 607
rect 426 573 460 607
rect 346 483 380 517
rect 426 483 460 517
rect 512 565 546 599
rect 512 495 546 529
rect 512 427 546 461
rect 600 509 634 543
rect 600 379 634 413
rect 692 565 726 599
rect 692 483 726 517
rect 692 402 726 436
<< poly >>
rect 118 619 148 645
rect 219 619 249 645
rect 305 619 335 645
rect 471 619 501 645
rect 557 619 587 645
rect 651 619 681 645
rect 118 303 148 367
rect 219 305 249 367
rect 80 287 153 303
rect 80 253 103 287
rect 137 253 153 287
rect 80 237 153 253
rect 195 289 263 305
rect 195 255 213 289
rect 247 255 263 289
rect 195 239 263 255
rect 80 215 110 237
rect 233 215 263 239
rect 305 303 335 367
rect 471 305 501 367
rect 305 287 375 303
rect 305 253 322 287
rect 356 253 375 287
rect 305 237 375 253
rect 423 289 501 305
rect 557 303 587 367
rect 651 308 681 367
rect 423 255 439 289
rect 473 255 501 289
rect 423 239 501 255
rect 543 287 609 303
rect 543 253 559 287
rect 593 253 609 287
rect 326 215 356 237
rect 423 215 453 239
rect 543 237 609 253
rect 579 215 609 237
rect 651 292 744 308
rect 651 258 694 292
rect 728 258 744 292
rect 651 242 744 258
rect 651 215 681 242
rect 80 21 110 47
rect 233 21 263 47
rect 326 21 356 47
rect 423 21 453 47
rect 579 21 609 47
rect 651 21 681 47
<< polycont >>
rect 103 253 137 287
rect 213 255 247 289
rect 322 253 356 287
rect 439 255 473 289
rect 559 253 593 287
rect 694 258 728 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 19 599 109 615
rect 19 565 73 599
rect 107 565 109 599
rect 19 520 109 565
rect 19 486 73 520
rect 107 486 109 520
rect 19 420 109 486
rect 144 607 210 649
rect 144 573 160 607
rect 194 573 210 607
rect 144 532 210 573
rect 144 498 160 532
rect 194 498 210 532
rect 144 455 210 498
rect 144 421 160 455
rect 194 421 210 455
rect 244 597 296 613
rect 244 563 260 597
rect 294 563 296 597
rect 244 522 296 563
rect 244 488 260 522
rect 294 488 296 522
rect 244 443 296 488
rect 330 607 476 649
rect 330 573 346 607
rect 380 573 426 607
rect 460 573 476 607
rect 330 517 476 573
rect 330 483 346 517
rect 380 483 426 517
rect 460 483 476 517
rect 330 477 476 483
rect 510 599 742 615
rect 510 565 512 599
rect 546 581 692 599
rect 546 565 550 581
rect 510 529 550 565
rect 684 565 692 581
rect 726 565 742 599
rect 510 495 512 529
rect 546 495 550 529
rect 510 461 550 495
rect 510 443 512 461
rect 19 386 73 420
rect 107 386 109 420
rect 244 409 260 443
rect 294 427 512 443
rect 546 427 550 461
rect 294 409 550 427
rect 584 543 650 547
rect 584 509 600 543
rect 634 509 650 543
rect 584 413 650 509
rect 19 370 109 386
rect 584 379 600 413
rect 634 379 650 413
rect 684 517 742 565
rect 684 483 692 517
rect 726 483 742 517
rect 684 436 742 483
rect 684 402 692 436
rect 726 402 742 436
rect 684 386 742 402
rect 584 375 650 379
rect 19 203 69 370
rect 143 341 650 375
rect 143 303 177 341
rect 19 169 35 203
rect 103 287 177 303
rect 137 253 177 287
rect 103 205 177 253
rect 211 289 270 305
rect 211 255 213 289
rect 247 255 270 289
rect 211 239 270 255
rect 305 287 375 305
rect 305 253 322 287
rect 356 253 375 287
rect 305 239 375 253
rect 415 289 473 305
rect 415 255 439 289
rect 415 239 473 255
rect 511 287 650 303
rect 511 253 559 287
rect 593 253 650 287
rect 511 239 650 253
rect 684 292 751 350
rect 684 258 694 292
rect 728 258 751 292
rect 684 242 751 258
rect 103 203 584 205
rect 103 171 464 203
rect 19 101 69 169
rect 448 169 464 171
rect 498 169 534 203
rect 568 169 584 203
rect 19 67 35 101
rect 19 51 69 67
rect 109 103 188 137
rect 222 103 239 137
rect 109 93 239 103
rect 109 59 121 93
rect 155 59 239 93
rect 109 17 239 59
rect 448 93 584 169
rect 448 59 464 93
rect 498 59 534 93
rect 568 59 584 93
rect 448 51 584 59
rect 676 203 742 208
rect 676 169 692 203
rect 726 169 742 203
rect 676 93 742 169
rect 676 59 692 93
rect 726 59 742 93
rect 676 17 742 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a32o_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2161124
string GDS_START 2153076
<< end >>
