magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 1 49 767 248
rect 0 0 768 49
<< scpmos >>
rect 112 368 142 592
rect 294 368 324 592
rect 378 368 408 592
rect 492 368 522 592
rect 606 368 636 592
<< nmoslvt >>
rect 84 74 114 222
rect 296 74 326 222
rect 396 74 426 222
rect 496 74 526 222
rect 654 74 684 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 138 185 222
rect 114 104 125 138
rect 159 104 185 138
rect 114 74 185 104
rect 239 210 296 222
rect 239 176 251 210
rect 285 176 296 210
rect 239 74 296 176
rect 326 143 396 222
rect 326 109 351 143
rect 385 109 396 143
rect 326 74 396 109
rect 426 210 496 222
rect 426 176 451 210
rect 485 176 496 210
rect 426 120 496 176
rect 426 86 451 120
rect 485 86 496 120
rect 426 74 496 86
rect 526 142 654 222
rect 526 108 537 142
rect 571 108 609 142
rect 643 108 654 142
rect 526 74 654 108
rect 684 210 741 222
rect 684 176 695 210
rect 729 176 741 210
rect 684 120 741 176
rect 684 86 695 120
rect 729 86 741 120
rect 684 74 741 86
<< pdiff >>
rect 53 580 112 592
rect 53 546 65 580
rect 99 546 112 580
rect 53 510 112 546
rect 53 476 65 510
rect 99 476 112 510
rect 53 440 112 476
rect 53 406 65 440
rect 99 406 112 440
rect 53 368 112 406
rect 142 580 294 592
rect 142 546 155 580
rect 189 546 247 580
rect 281 546 294 580
rect 142 508 294 546
rect 142 474 155 508
rect 189 492 294 508
rect 189 474 247 492
rect 142 458 247 474
rect 281 458 294 492
rect 142 368 294 458
rect 324 368 378 592
rect 408 580 492 592
rect 408 546 421 580
rect 455 546 492 580
rect 408 510 492 546
rect 408 476 421 510
rect 455 476 492 510
rect 408 440 492 476
rect 408 406 421 440
rect 455 406 492 440
rect 408 368 492 406
rect 522 368 606 592
rect 636 580 695 592
rect 636 546 649 580
rect 683 546 695 580
rect 636 510 695 546
rect 636 476 649 510
rect 683 476 695 510
rect 636 440 695 476
rect 636 406 649 440
rect 683 406 695 440
rect 636 368 695 406
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 104 159 138
rect 251 176 285 210
rect 351 109 385 143
rect 451 176 485 210
rect 451 86 485 120
rect 537 108 571 142
rect 609 108 643 142
rect 695 176 729 210
rect 695 86 729 120
<< pdiffc >>
rect 65 546 99 580
rect 65 476 99 510
rect 65 406 99 440
rect 155 546 189 580
rect 247 546 281 580
rect 155 474 189 508
rect 247 458 281 492
rect 421 546 455 580
rect 421 476 455 510
rect 421 406 455 440
rect 649 546 683 580
rect 649 476 683 510
rect 649 406 683 440
<< poly >>
rect 112 592 142 618
rect 294 592 324 618
rect 378 592 408 618
rect 492 592 522 618
rect 606 592 636 618
rect 112 353 142 368
rect 294 353 324 368
rect 378 353 408 368
rect 492 353 522 368
rect 606 353 636 368
rect 109 326 145 353
rect 291 336 327 353
rect 21 310 145 326
rect 21 276 37 310
rect 71 296 145 310
rect 193 320 327 336
rect 71 276 114 296
rect 21 260 114 276
rect 193 286 209 320
rect 243 286 277 320
rect 311 286 327 320
rect 193 270 327 286
rect 375 336 411 353
rect 489 336 525 353
rect 375 320 441 336
rect 375 286 391 320
rect 425 286 441 320
rect 375 270 441 286
rect 489 320 555 336
rect 489 286 505 320
rect 539 286 555 320
rect 489 270 555 286
rect 603 326 639 353
rect 603 310 737 326
rect 603 276 619 310
rect 653 276 687 310
rect 721 276 737 310
rect 84 222 114 260
rect 296 222 326 270
rect 396 222 426 270
rect 496 222 526 270
rect 603 260 737 276
rect 654 222 684 260
rect 84 48 114 74
rect 296 48 326 74
rect 396 48 426 74
rect 496 48 526 74
rect 654 48 684 74
<< polycont >>
rect 37 276 71 310
rect 209 286 243 320
rect 277 286 311 320
rect 391 286 425 320
rect 505 286 539 320
rect 619 276 653 310
rect 687 276 721 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 65 580 115 596
rect 99 546 115 580
rect 65 510 115 546
rect 99 476 115 510
rect 65 440 115 476
rect 149 580 312 649
rect 149 546 155 580
rect 189 546 247 580
rect 281 546 312 580
rect 149 508 312 546
rect 149 474 155 508
rect 189 492 312 508
rect 189 474 247 492
rect 149 458 247 474
rect 281 458 312 492
rect 405 580 471 596
rect 405 546 421 580
rect 455 546 471 580
rect 633 580 699 649
rect 405 510 471 546
rect 405 476 421 510
rect 455 476 471 510
rect 99 424 115 440
rect 405 440 471 476
rect 405 424 421 440
rect 99 406 421 424
rect 455 406 471 440
rect 65 390 471 406
rect 21 310 87 356
rect 21 276 37 310
rect 71 276 87 310
rect 21 260 87 276
rect 121 226 155 390
rect 193 320 327 356
rect 193 286 209 320
rect 243 286 277 320
rect 311 286 327 320
rect 193 270 327 286
rect 375 320 455 356
rect 505 336 555 578
rect 633 546 649 580
rect 683 546 699 580
rect 633 510 699 546
rect 633 476 649 510
rect 683 476 699 510
rect 633 440 699 476
rect 633 406 649 440
rect 683 406 699 440
rect 633 390 699 406
rect 375 286 391 320
rect 425 286 455 320
rect 375 270 455 286
rect 489 320 555 336
rect 489 286 505 320
rect 539 286 555 320
rect 489 270 555 286
rect 601 310 743 356
rect 601 276 619 310
rect 653 276 687 310
rect 721 276 743 310
rect 601 260 743 276
rect 23 210 155 226
rect 23 176 39 210
rect 73 192 155 210
rect 235 226 501 236
rect 235 210 745 226
rect 73 176 89 192
rect 23 120 89 176
rect 235 176 251 210
rect 285 202 451 210
rect 285 176 301 202
rect 235 160 301 176
rect 435 176 451 202
rect 485 192 695 210
rect 485 176 501 192
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 138 189 154
rect 123 104 125 138
rect 159 104 189 138
rect 335 143 401 159
rect 335 109 351 143
rect 385 109 401 143
rect 335 104 401 109
rect 123 70 401 104
rect 435 120 501 176
rect 679 176 695 192
rect 729 176 745 210
rect 435 86 451 120
rect 485 86 501 120
rect 435 70 501 86
rect 535 142 645 158
rect 535 108 537 142
rect 571 108 609 142
rect 643 108 645 142
rect 535 17 645 108
rect 679 120 745 176
rect 679 86 695 120
rect 729 86 745 120
rect 679 70 745 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o221ai_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 3836220
string GDS_START 3828756
<< end >>
