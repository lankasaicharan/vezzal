magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 1244 241 1518 243
rect 4 49 1518 241
rect 0 0 1536 49
<< scnmos >>
rect 83 47 113 215
rect 169 47 199 215
rect 255 47 285 215
rect 341 47 371 215
rect 427 47 457 215
rect 513 47 543 215
rect 703 47 733 215
rect 789 47 819 215
rect 875 47 905 215
rect 961 47 991 215
rect 1047 47 1077 215
rect 1133 47 1163 215
rect 1323 49 1353 217
rect 1409 49 1439 217
<< scpmoshvt >>
rect 83 367 113 619
rect 169 367 199 619
rect 255 367 285 619
rect 341 367 371 619
rect 427 367 457 619
rect 513 367 543 619
rect 599 367 629 619
rect 685 367 715 619
rect 875 367 905 619
rect 961 367 991 619
rect 1047 367 1077 619
rect 1133 367 1163 619
rect 1219 367 1249 619
rect 1305 367 1335 619
<< ndiff >>
rect 30 178 83 215
rect 30 144 38 178
rect 72 144 83 178
rect 30 93 83 144
rect 30 59 38 93
rect 72 59 83 93
rect 30 47 83 59
rect 113 203 169 215
rect 113 169 124 203
rect 158 169 169 203
rect 113 101 169 169
rect 113 67 124 101
rect 158 67 169 101
rect 113 47 169 67
rect 199 175 255 215
rect 199 141 210 175
rect 244 141 255 175
rect 199 89 255 141
rect 199 55 210 89
rect 244 55 255 89
rect 199 47 255 55
rect 285 203 341 215
rect 285 169 296 203
rect 330 169 341 203
rect 285 101 341 169
rect 285 67 296 101
rect 330 67 341 101
rect 285 47 341 67
rect 371 199 427 215
rect 371 165 382 199
rect 416 165 427 199
rect 371 93 427 165
rect 371 59 382 93
rect 416 59 427 93
rect 371 47 427 59
rect 457 187 513 215
rect 457 153 468 187
rect 502 153 513 187
rect 457 101 513 153
rect 457 67 468 101
rect 502 67 513 101
rect 457 47 513 67
rect 543 119 596 215
rect 543 85 554 119
rect 588 85 596 119
rect 543 47 596 85
rect 650 119 703 215
rect 650 85 658 119
rect 692 85 703 119
rect 650 47 703 85
rect 733 169 789 215
rect 733 135 744 169
rect 778 135 789 169
rect 733 47 789 135
rect 819 189 875 215
rect 819 155 830 189
rect 864 155 875 189
rect 819 101 875 155
rect 819 67 830 101
rect 864 67 875 101
rect 819 47 875 67
rect 905 121 961 215
rect 905 87 916 121
rect 950 87 961 121
rect 905 47 961 87
rect 991 189 1047 215
rect 991 155 1002 189
rect 1036 155 1047 189
rect 991 101 1047 155
rect 991 67 1002 101
rect 1036 67 1047 101
rect 991 47 1047 67
rect 1077 187 1133 215
rect 1077 153 1088 187
rect 1122 153 1133 187
rect 1077 47 1133 153
rect 1163 97 1216 215
rect 1163 63 1174 97
rect 1208 63 1216 97
rect 1163 47 1216 63
rect 1270 205 1323 217
rect 1270 171 1278 205
rect 1312 171 1323 205
rect 1270 101 1323 171
rect 1270 67 1278 101
rect 1312 67 1323 101
rect 1270 49 1323 67
rect 1353 179 1409 217
rect 1353 145 1364 179
rect 1398 145 1409 179
rect 1353 95 1409 145
rect 1353 61 1364 95
rect 1398 61 1409 95
rect 1353 49 1409 61
rect 1439 205 1492 217
rect 1439 171 1450 205
rect 1484 171 1492 205
rect 1439 101 1492 171
rect 1439 67 1450 101
rect 1484 67 1492 101
rect 1439 49 1492 67
<< pdiff >>
rect 30 607 83 619
rect 30 573 38 607
rect 72 573 83 607
rect 30 532 83 573
rect 30 498 38 532
rect 72 498 83 532
rect 30 453 83 498
rect 30 419 38 453
rect 72 419 83 453
rect 30 367 83 419
rect 113 599 169 619
rect 113 565 124 599
rect 158 565 169 599
rect 113 514 169 565
rect 113 480 124 514
rect 158 480 169 514
rect 113 413 169 480
rect 113 379 124 413
rect 158 379 169 413
rect 113 367 169 379
rect 199 607 255 619
rect 199 573 210 607
rect 244 573 255 607
rect 199 530 255 573
rect 199 496 210 530
rect 244 496 255 530
rect 199 453 255 496
rect 199 419 210 453
rect 244 419 255 453
rect 199 367 255 419
rect 285 599 341 619
rect 285 565 296 599
rect 330 565 341 599
rect 285 514 341 565
rect 285 480 296 514
rect 330 480 341 514
rect 285 413 341 480
rect 285 379 296 413
rect 330 379 341 413
rect 285 367 341 379
rect 371 607 427 619
rect 371 573 382 607
rect 416 573 427 607
rect 371 524 427 573
rect 371 490 382 524
rect 416 490 427 524
rect 371 443 427 490
rect 371 409 382 443
rect 416 409 427 443
rect 371 367 427 409
rect 457 599 513 619
rect 457 565 468 599
rect 502 565 513 599
rect 457 529 513 565
rect 457 495 468 529
rect 502 495 513 529
rect 457 459 513 495
rect 457 425 468 459
rect 502 425 513 459
rect 457 367 513 425
rect 543 607 599 619
rect 543 573 554 607
rect 588 573 599 607
rect 543 513 599 573
rect 543 479 554 513
rect 588 479 599 513
rect 543 367 599 479
rect 629 597 685 619
rect 629 563 640 597
rect 674 563 685 597
rect 629 529 685 563
rect 629 495 640 529
rect 674 495 685 529
rect 629 459 685 495
rect 629 425 640 459
rect 674 425 685 459
rect 629 367 685 425
rect 715 607 768 619
rect 715 573 726 607
rect 760 573 768 607
rect 715 511 768 573
rect 715 477 726 511
rect 760 477 768 511
rect 715 367 768 477
rect 822 597 875 619
rect 822 563 830 597
rect 864 563 875 597
rect 822 367 875 563
rect 905 445 961 619
rect 905 411 916 445
rect 950 411 961 445
rect 905 367 961 411
rect 991 597 1047 619
rect 991 563 1002 597
rect 1036 563 1047 597
rect 991 367 1047 563
rect 1077 507 1133 619
rect 1077 473 1088 507
rect 1122 473 1133 507
rect 1077 413 1133 473
rect 1077 379 1088 413
rect 1122 379 1133 413
rect 1077 367 1133 379
rect 1163 597 1219 619
rect 1163 563 1174 597
rect 1208 563 1219 597
rect 1163 524 1219 563
rect 1163 490 1174 524
rect 1208 490 1219 524
rect 1163 446 1219 490
rect 1163 412 1174 446
rect 1208 412 1219 446
rect 1163 367 1219 412
rect 1249 529 1305 619
rect 1249 495 1260 529
rect 1294 495 1305 529
rect 1249 413 1305 495
rect 1249 379 1260 413
rect 1294 379 1305 413
rect 1249 367 1305 379
rect 1335 597 1388 619
rect 1335 563 1346 597
rect 1380 563 1388 597
rect 1335 506 1388 563
rect 1335 472 1346 506
rect 1380 472 1388 506
rect 1335 418 1388 472
rect 1335 384 1346 418
rect 1380 384 1388 418
rect 1335 367 1388 384
<< ndiffc >>
rect 38 144 72 178
rect 38 59 72 93
rect 124 169 158 203
rect 124 67 158 101
rect 210 141 244 175
rect 210 55 244 89
rect 296 169 330 203
rect 296 67 330 101
rect 382 165 416 199
rect 382 59 416 93
rect 468 153 502 187
rect 468 67 502 101
rect 554 85 588 119
rect 658 85 692 119
rect 744 135 778 169
rect 830 155 864 189
rect 830 67 864 101
rect 916 87 950 121
rect 1002 155 1036 189
rect 1002 67 1036 101
rect 1088 153 1122 187
rect 1174 63 1208 97
rect 1278 171 1312 205
rect 1278 67 1312 101
rect 1364 145 1398 179
rect 1364 61 1398 95
rect 1450 171 1484 205
rect 1450 67 1484 101
<< pdiffc >>
rect 38 573 72 607
rect 38 498 72 532
rect 38 419 72 453
rect 124 565 158 599
rect 124 480 158 514
rect 124 379 158 413
rect 210 573 244 607
rect 210 496 244 530
rect 210 419 244 453
rect 296 565 330 599
rect 296 480 330 514
rect 296 379 330 413
rect 382 573 416 607
rect 382 490 416 524
rect 382 409 416 443
rect 468 565 502 599
rect 468 495 502 529
rect 468 425 502 459
rect 554 573 588 607
rect 554 479 588 513
rect 640 563 674 597
rect 640 495 674 529
rect 640 425 674 459
rect 726 573 760 607
rect 726 477 760 511
rect 830 563 864 597
rect 916 411 950 445
rect 1002 563 1036 597
rect 1088 473 1122 507
rect 1088 379 1122 413
rect 1174 563 1208 597
rect 1174 490 1208 524
rect 1174 412 1208 446
rect 1260 495 1294 529
rect 1260 379 1294 413
rect 1346 563 1380 597
rect 1346 472 1380 506
rect 1346 384 1380 418
<< poly >>
rect 83 619 113 645
rect 169 619 199 645
rect 255 619 285 645
rect 341 619 371 645
rect 427 619 457 645
rect 513 619 543 645
rect 599 619 629 645
rect 685 619 715 645
rect 875 619 905 645
rect 961 619 991 645
rect 1047 619 1077 645
rect 1133 619 1163 645
rect 1219 619 1249 645
rect 1305 619 1335 645
rect 83 331 113 367
rect 169 331 199 367
rect 255 331 285 367
rect 341 331 371 367
rect 83 315 371 331
rect 83 281 117 315
rect 151 281 185 315
rect 219 281 253 315
rect 287 281 321 315
rect 355 281 371 315
rect 427 303 457 367
rect 513 304 543 367
rect 513 303 557 304
rect 83 265 371 281
rect 83 215 113 265
rect 169 215 199 265
rect 255 215 285 265
rect 341 215 371 265
rect 422 287 557 303
rect 422 253 439 287
rect 473 253 507 287
rect 541 253 557 287
rect 422 237 557 253
rect 599 303 629 367
rect 685 303 715 367
rect 875 305 905 367
rect 961 305 991 367
rect 1047 305 1077 367
rect 1133 305 1163 367
rect 1219 335 1249 367
rect 1305 335 1335 367
rect 1219 315 1460 335
rect 599 287 819 303
rect 599 253 682 287
rect 716 253 750 287
rect 784 253 819 287
rect 599 237 819 253
rect 427 215 457 237
rect 513 215 543 237
rect 703 215 733 237
rect 789 215 819 237
rect 875 289 991 305
rect 875 255 927 289
rect 961 255 991 289
rect 875 239 991 255
rect 1043 289 1177 305
rect 1043 255 1059 289
rect 1093 255 1127 289
rect 1161 255 1177 289
rect 1219 281 1342 315
rect 1376 281 1410 315
rect 1444 281 1460 315
rect 1219 269 1460 281
rect 1043 239 1177 255
rect 1323 265 1460 269
rect 875 215 905 239
rect 961 215 991 239
rect 1047 215 1077 239
rect 1133 215 1163 239
rect 1323 217 1353 265
rect 1409 217 1439 265
rect 83 21 113 47
rect 169 21 199 47
rect 255 21 285 47
rect 341 21 371 47
rect 427 21 457 47
rect 513 21 543 47
rect 703 21 733 47
rect 789 21 819 47
rect 875 21 905 47
rect 961 21 991 47
rect 1047 21 1077 47
rect 1133 21 1163 47
rect 1323 23 1353 49
rect 1409 23 1439 49
<< polycont >>
rect 117 281 151 315
rect 185 281 219 315
rect 253 281 287 315
rect 321 281 355 315
rect 439 253 473 287
rect 507 253 541 287
rect 682 253 716 287
rect 750 253 784 287
rect 927 255 961 289
rect 1059 255 1093 289
rect 1127 255 1161 289
rect 1342 281 1376 315
rect 1410 281 1444 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 22 607 88 649
rect 22 573 38 607
rect 72 573 88 607
rect 22 532 88 573
rect 22 498 38 532
rect 72 498 88 532
rect 22 453 88 498
rect 22 419 38 453
rect 72 419 88 453
rect 122 599 158 615
rect 122 565 124 599
rect 122 514 158 565
rect 122 480 124 514
rect 122 413 158 480
rect 194 607 260 649
rect 194 573 210 607
rect 244 573 260 607
rect 194 530 260 573
rect 194 496 210 530
rect 244 496 260 530
rect 194 453 260 496
rect 194 419 210 453
rect 244 419 260 453
rect 294 599 332 615
rect 294 565 296 599
rect 330 565 332 599
rect 294 514 332 565
rect 294 480 296 514
rect 330 480 332 514
rect 122 385 124 413
rect 22 379 124 385
rect 294 413 332 480
rect 294 385 296 413
rect 158 379 296 385
rect 330 379 332 413
rect 366 607 432 649
rect 366 573 382 607
rect 416 573 432 607
rect 366 524 432 573
rect 366 490 382 524
rect 416 490 432 524
rect 366 443 432 490
rect 366 409 382 443
rect 416 409 432 443
rect 466 599 504 615
rect 466 565 468 599
rect 502 565 504 599
rect 466 529 504 565
rect 466 495 468 529
rect 502 495 504 529
rect 466 459 504 495
rect 538 607 604 649
rect 538 573 554 607
rect 588 573 604 607
rect 538 513 604 573
rect 538 479 554 513
rect 588 479 604 513
rect 638 597 676 613
rect 638 563 640 597
rect 674 563 676 597
rect 638 529 676 563
rect 638 495 640 529
rect 674 495 676 529
rect 466 425 468 459
rect 502 445 504 459
rect 638 459 676 495
rect 710 607 776 649
rect 710 573 726 607
rect 760 573 776 607
rect 710 511 776 573
rect 814 597 1396 613
rect 814 563 830 597
rect 864 563 1002 597
rect 1036 563 1174 597
rect 1208 579 1346 597
rect 1208 563 1224 579
rect 814 557 1224 563
rect 1158 524 1224 557
rect 1330 563 1346 579
rect 1380 563 1396 597
rect 710 477 726 511
rect 760 477 776 511
rect 814 507 1124 523
rect 814 489 1088 507
rect 638 445 640 459
rect 502 425 640 445
rect 674 443 676 459
rect 814 443 863 489
rect 1072 473 1088 489
rect 1122 473 1124 507
rect 674 425 863 443
rect 466 409 863 425
rect 900 445 966 455
rect 900 411 916 445
rect 950 411 966 445
rect 22 351 332 379
rect 900 375 966 411
rect 22 246 67 351
rect 370 341 966 375
rect 1072 413 1124 473
rect 1072 379 1088 413
rect 1122 379 1124 413
rect 1158 490 1174 524
rect 1208 490 1224 524
rect 1158 446 1224 490
rect 1158 412 1174 446
rect 1208 412 1224 446
rect 1158 411 1224 412
rect 1258 529 1294 545
rect 1258 495 1260 529
rect 1258 413 1294 495
rect 1072 375 1124 379
rect 1258 379 1260 413
rect 1330 506 1396 563
rect 1330 472 1346 506
rect 1380 472 1396 506
rect 1330 418 1396 472
rect 1330 384 1346 418
rect 1380 384 1396 418
rect 1258 375 1294 379
rect 1072 341 1294 375
rect 370 338 859 341
rect 370 317 404 338
rect 101 315 404 317
rect 101 281 117 315
rect 151 281 185 315
rect 219 281 253 315
rect 287 281 321 315
rect 355 281 404 315
rect 101 280 404 281
rect 438 287 641 303
rect 438 253 439 287
rect 473 253 507 287
rect 541 253 641 287
rect 22 212 332 246
rect 438 237 641 253
rect 675 287 791 303
rect 675 253 682 287
rect 716 253 750 287
rect 784 253 791 287
rect 675 237 791 253
rect 122 209 332 212
rect 122 203 160 209
rect 22 144 38 178
rect 72 144 88 178
rect 22 93 88 144
rect 22 59 38 93
rect 72 59 88 93
rect 22 17 88 59
rect 122 169 124 203
rect 158 169 160 203
rect 294 203 332 209
rect 825 205 859 338
rect 1328 324 1505 350
rect 1326 315 1505 324
rect 893 289 1025 305
rect 893 255 927 289
rect 961 255 1025 289
rect 893 239 1025 255
rect 1059 289 1227 305
rect 1093 255 1127 289
rect 1161 255 1227 289
rect 1326 281 1342 315
rect 1376 281 1410 315
rect 1444 281 1505 315
rect 1059 239 1227 255
rect 1274 213 1500 247
rect 1274 205 1314 213
rect 122 101 160 169
rect 122 67 124 101
rect 158 67 160 101
rect 122 51 160 67
rect 194 141 210 175
rect 244 141 260 175
rect 194 89 260 141
rect 194 55 210 89
rect 244 55 260 89
rect 194 17 260 55
rect 294 169 296 203
rect 330 169 332 203
rect 294 101 332 169
rect 294 67 296 101
rect 330 67 332 101
rect 294 51 332 67
rect 366 199 432 203
rect 366 165 382 199
rect 416 165 432 199
rect 366 93 432 165
rect 366 59 382 93
rect 416 59 432 93
rect 366 17 432 59
rect 466 187 791 203
rect 466 153 468 187
rect 502 169 791 187
rect 502 153 504 169
rect 466 101 504 153
rect 740 135 744 169
rect 778 135 791 169
rect 466 67 468 101
rect 502 67 504 101
rect 466 51 504 67
rect 538 119 604 135
rect 538 85 554 119
rect 588 85 604 119
rect 538 17 604 85
rect 642 119 706 135
rect 740 119 791 135
rect 825 189 1047 205
rect 1274 203 1278 205
rect 825 155 830 189
rect 864 171 1002 189
rect 864 155 873 171
rect 642 85 658 119
rect 692 85 706 119
rect 825 101 873 155
rect 993 155 1002 171
rect 1036 155 1047 189
rect 825 85 830 101
rect 642 67 830 85
rect 864 67 873 101
rect 642 51 873 67
rect 907 121 959 137
rect 907 87 916 121
rect 950 87 959 121
rect 907 17 959 87
rect 993 103 1047 155
rect 1081 187 1278 203
rect 1081 153 1088 187
rect 1122 171 1278 187
rect 1312 171 1314 205
rect 1448 205 1500 213
rect 1122 153 1314 171
rect 1081 137 1314 153
rect 993 101 1224 103
rect 993 67 1002 101
rect 1036 97 1224 101
rect 1036 67 1174 97
rect 993 63 1174 67
rect 1208 63 1224 97
rect 993 51 1224 63
rect 1262 101 1314 137
rect 1262 67 1278 101
rect 1312 67 1314 101
rect 1262 51 1314 67
rect 1348 145 1364 179
rect 1398 145 1414 179
rect 1348 95 1414 145
rect 1348 61 1364 95
rect 1398 61 1414 95
rect 1348 17 1414 61
rect 1448 171 1450 205
rect 1484 171 1500 205
rect 1448 101 1500 171
rect 1448 67 1450 101
rect 1484 67 1500 101
rect 1448 51 1500 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a221o_4
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6134220
string GDS_START 6121252
<< end >>
