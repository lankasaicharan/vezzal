magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3890 1975
<< nwell >>
rect -38 331 2630 704
rect 1042 279 1582 331
<< pwell >>
rect 191 201 556 284
rect 1664 241 2030 284
rect 2394 241 2588 251
rect 1664 237 2588 241
rect 1151 207 2588 237
rect 984 201 2588 207
rect 191 179 2588 201
rect 1 49 2588 179
rect 0 0 2592 49
<< scnmos >>
rect 80 69 110 153
rect 270 130 300 258
rect 342 130 372 258
rect 447 174 477 258
rect 637 47 667 175
rect 709 47 739 175
rect 814 47 844 131
rect 886 47 916 131
rect 958 47 988 131
rect 1232 127 1262 211
rect 1339 127 1369 211
rect 1425 127 1455 211
rect 1527 127 1557 211
rect 1768 174 1798 258
rect 1846 174 1876 258
rect 1918 174 1948 258
rect 2114 131 2144 215
rect 2186 131 2216 215
rect 2272 131 2302 215
rect 2476 57 2506 225
<< scpmoshvt >>
rect 82 400 112 528
rect 189 400 219 568
rect 404 405 434 533
rect 598 451 628 619
rect 670 451 700 619
rect 780 419 830 619
rect 878 419 928 619
rect 1196 341 1246 541
rect 1294 341 1344 541
rect 1439 341 1489 541
rect 1765 466 1795 594
rect 1874 368 1904 496
rect 2006 368 2056 568
rect 2323 367 2353 495
rect 2476 367 2506 619
<< ndiff >>
rect 217 246 270 258
rect 217 212 225 246
rect 259 212 270 246
rect 217 176 270 212
rect 27 128 80 153
rect 27 94 35 128
rect 69 94 80 128
rect 27 69 80 94
rect 110 128 163 153
rect 217 142 225 176
rect 259 142 270 176
rect 217 130 270 142
rect 300 130 342 258
rect 372 212 447 258
rect 372 178 383 212
rect 417 178 447 212
rect 372 174 447 178
rect 477 227 530 258
rect 477 193 488 227
rect 522 193 530 227
rect 477 174 530 193
rect 372 130 425 174
rect 584 158 637 175
rect 110 94 121 128
rect 155 94 163 128
rect 584 124 592 158
rect 626 124 637 158
rect 110 69 163 94
rect 584 47 637 124
rect 667 47 709 175
rect 739 158 792 175
rect 739 124 750 158
rect 784 131 792 158
rect 1690 233 1768 258
rect 1010 169 1065 181
rect 1010 135 1019 169
rect 1053 135 1065 169
rect 1010 131 1065 135
rect 784 124 814 131
rect 739 47 814 124
rect 844 47 886 131
rect 916 47 958 131
rect 988 47 1065 131
rect 1177 173 1232 211
rect 1177 139 1187 173
rect 1221 139 1232 173
rect 1177 127 1232 139
rect 1262 186 1339 211
rect 1262 152 1294 186
rect 1328 152 1339 186
rect 1262 127 1339 152
rect 1369 180 1425 211
rect 1369 146 1380 180
rect 1414 146 1425 180
rect 1369 127 1425 146
rect 1455 127 1527 211
rect 1557 148 1636 211
rect 1690 199 1701 233
rect 1735 199 1768 233
rect 1690 174 1768 199
rect 1798 174 1846 258
rect 1876 174 1918 258
rect 1948 233 2004 258
rect 1948 199 1959 233
rect 1993 199 2004 233
rect 1948 174 2004 199
rect 2058 190 2114 215
rect 2058 156 2069 190
rect 2103 156 2114 190
rect 1557 127 1591 148
rect 1579 114 1591 127
rect 1625 114 1636 148
rect 2058 131 2114 156
rect 2144 131 2186 215
rect 2216 190 2272 215
rect 2216 156 2227 190
rect 2261 156 2272 190
rect 2216 131 2272 156
rect 2302 190 2358 215
rect 2302 156 2313 190
rect 2347 156 2358 190
rect 2302 131 2358 156
rect 2420 213 2476 225
rect 2420 179 2431 213
rect 2465 179 2476 213
rect 1579 72 1636 114
rect 2420 103 2476 179
rect 2420 69 2431 103
rect 2465 69 2476 103
rect 2420 57 2476 69
rect 2506 213 2562 225
rect 2506 179 2517 213
rect 2551 179 2562 213
rect 2506 103 2562 179
rect 2506 69 2517 103
rect 2551 69 2562 103
rect 2506 57 2562 69
<< pdiff >>
rect 328 619 382 631
rect 328 585 338 619
rect 372 585 382 619
rect 134 535 189 568
rect 134 528 144 535
rect 27 516 82 528
rect 27 482 37 516
rect 71 482 82 516
rect 27 446 82 482
rect 27 412 37 446
rect 71 412 82 446
rect 27 400 82 412
rect 112 501 144 528
rect 178 501 189 535
rect 112 400 189 501
rect 219 556 274 568
rect 219 522 230 556
rect 264 522 274 556
rect 219 446 274 522
rect 219 412 230 446
rect 264 412 274 446
rect 219 400 274 412
rect 328 533 382 585
rect 543 599 598 619
rect 543 565 553 599
rect 587 565 598 599
rect 328 405 404 533
rect 434 451 489 533
rect 543 503 598 565
rect 543 469 553 503
rect 587 469 598 503
rect 543 451 598 469
rect 628 451 670 619
rect 700 498 780 619
rect 700 464 734 498
rect 768 464 780 498
rect 700 451 780 464
rect 434 417 445 451
rect 479 417 489 451
rect 434 405 489 417
rect 722 419 780 451
rect 830 419 878 619
rect 928 590 984 619
rect 928 556 939 590
rect 973 556 984 590
rect 928 419 984 556
rect 1366 581 1424 593
rect 1366 547 1378 581
rect 1412 547 1424 581
rect 1366 541 1424 547
rect 2405 607 2476 619
rect 1708 582 1765 594
rect 1708 548 1720 582
rect 1754 548 1765 582
rect 1116 361 1196 541
rect 1116 327 1128 361
rect 1162 341 1196 361
rect 1246 341 1294 541
rect 1344 341 1439 541
rect 1489 400 1546 541
rect 1708 466 1765 548
rect 1795 496 1845 594
rect 1926 582 1984 594
rect 1926 548 1938 582
rect 1972 568 1984 582
rect 2405 573 2417 607
rect 2451 573 2476 607
rect 1972 548 2006 568
rect 1926 496 2006 548
rect 1795 466 1874 496
rect 1489 366 1500 400
rect 1534 366 1546 400
rect 1489 341 1546 366
rect 1162 327 1174 341
rect 1116 315 1174 327
rect 1817 414 1874 466
rect 1817 380 1829 414
rect 1863 380 1874 414
rect 1817 368 1874 380
rect 1904 368 2006 496
rect 2056 556 2113 568
rect 2056 522 2067 556
rect 2101 522 2113 556
rect 2056 485 2113 522
rect 2405 510 2476 573
rect 2405 495 2417 510
rect 2056 451 2067 485
rect 2101 451 2113 485
rect 2056 414 2113 451
rect 2266 483 2323 495
rect 2266 449 2278 483
rect 2312 449 2323 483
rect 2056 380 2067 414
rect 2101 380 2113 414
rect 2056 368 2113 380
rect 2266 413 2323 449
rect 2266 379 2278 413
rect 2312 379 2323 413
rect 2266 367 2323 379
rect 2353 476 2417 495
rect 2451 476 2476 510
rect 2353 413 2476 476
rect 2353 379 2417 413
rect 2451 379 2476 413
rect 2353 367 2476 379
rect 2506 599 2563 619
rect 2506 565 2517 599
rect 2551 565 2563 599
rect 2506 506 2563 565
rect 2506 472 2517 506
rect 2551 472 2563 506
rect 2506 413 2563 472
rect 2506 379 2517 413
rect 2551 379 2563 413
rect 2506 367 2563 379
<< ndiffc >>
rect 225 212 259 246
rect 35 94 69 128
rect 225 142 259 176
rect 383 178 417 212
rect 488 193 522 227
rect 121 94 155 128
rect 592 124 626 158
rect 750 124 784 158
rect 1019 135 1053 169
rect 1187 139 1221 173
rect 1294 152 1328 186
rect 1380 146 1414 180
rect 1701 199 1735 233
rect 1959 199 1993 233
rect 2069 156 2103 190
rect 1591 114 1625 148
rect 2227 156 2261 190
rect 2313 156 2347 190
rect 2431 179 2465 213
rect 2431 69 2465 103
rect 2517 179 2551 213
rect 2517 69 2551 103
<< pdiffc >>
rect 338 585 372 619
rect 37 482 71 516
rect 37 412 71 446
rect 144 501 178 535
rect 230 522 264 556
rect 230 412 264 446
rect 553 565 587 599
rect 553 469 587 503
rect 734 464 768 498
rect 445 417 479 451
rect 939 556 973 590
rect 1378 547 1412 581
rect 1720 548 1754 582
rect 1128 327 1162 361
rect 1938 548 1972 582
rect 2417 573 2451 607
rect 1500 366 1534 400
rect 1829 380 1863 414
rect 2067 522 2101 556
rect 2067 451 2101 485
rect 2278 449 2312 483
rect 2067 380 2101 414
rect 2278 379 2312 413
rect 2417 476 2451 510
rect 2417 379 2451 413
rect 2517 565 2551 599
rect 2517 472 2551 506
rect 2517 379 2551 413
<< poly >>
rect 598 619 628 645
rect 670 619 700 645
rect 780 619 830 645
rect 878 619 928 645
rect 189 568 219 594
rect 82 528 112 554
rect 404 533 434 559
rect 598 419 628 451
rect 670 419 700 451
rect 1294 615 1676 645
rect 1196 541 1246 567
rect 1294 541 1344 615
rect 1610 599 1676 615
rect 1439 541 1489 567
rect 1610 565 1626 599
rect 1660 565 1676 599
rect 1765 594 1795 620
rect 2476 619 2506 645
rect 1610 549 1676 565
rect 82 325 112 400
rect 189 362 219 400
rect 404 383 434 405
rect 598 403 700 419
rect 598 383 621 403
rect 404 369 621 383
rect 655 389 700 403
rect 655 369 671 389
rect 780 369 830 419
rect 25 309 112 325
rect 25 275 41 309
rect 75 275 112 309
rect 160 346 226 362
rect 404 353 671 369
rect 160 312 176 346
rect 210 326 226 346
rect 210 312 300 326
rect 160 296 300 312
rect 25 241 112 275
rect 270 258 300 296
rect 342 258 372 284
rect 447 258 477 353
rect 742 339 830 369
rect 878 387 928 419
rect 878 371 994 387
rect 878 357 944 371
rect 719 309 772 339
rect 928 337 944 357
rect 978 337 994 371
rect 928 321 994 337
rect 2006 568 2056 594
rect 1874 496 1904 522
rect 1657 414 1723 430
rect 1657 380 1673 414
rect 1707 380 1723 414
rect 1657 346 1723 380
rect 719 263 749 309
rect 25 207 41 241
rect 75 207 112 241
rect 25 191 112 207
rect 80 153 110 191
rect 566 247 749 263
rect 566 213 582 247
rect 616 233 749 247
rect 814 275 880 291
rect 814 241 830 275
rect 864 241 880 275
rect 616 213 667 233
rect 566 197 667 213
rect 637 175 667 197
rect 709 175 739 233
rect 814 225 880 241
rect 447 148 477 174
rect 270 104 300 130
rect 342 106 372 130
rect 342 90 462 106
rect 80 43 110 69
rect 342 56 412 90
rect 446 56 462 90
rect 342 40 462 56
rect 814 131 844 225
rect 958 183 988 321
rect 1196 263 1246 341
rect 1294 315 1344 341
rect 1314 299 1344 315
rect 1439 303 1489 341
rect 1314 269 1369 299
rect 1196 233 1262 263
rect 1232 211 1262 233
rect 1339 211 1369 269
rect 1417 287 1489 303
rect 1657 312 1673 346
rect 1707 326 1723 346
rect 1765 326 1795 466
rect 2323 495 2353 521
rect 2144 414 2211 430
rect 2144 380 2161 414
rect 2195 380 2211 414
rect 1874 326 1904 368
rect 2006 326 2056 368
rect 2144 346 2211 380
rect 2144 326 2161 346
rect 1707 312 1798 326
rect 1657 296 1798 312
rect 1417 253 1433 287
rect 1467 267 1489 287
rect 1467 253 1557 267
rect 1768 258 1798 296
rect 1846 312 2161 326
rect 2195 326 2211 346
rect 2195 312 2216 326
rect 1846 296 2216 312
rect 1846 258 1876 296
rect 1918 258 1948 296
rect 1417 237 1557 253
rect 1425 211 1455 237
rect 1527 211 1557 237
rect 886 153 988 183
rect 886 131 916 153
rect 958 131 988 153
rect 2114 215 2144 296
rect 2186 215 2216 296
rect 2323 267 2353 367
rect 2476 329 2506 367
rect 2272 237 2353 267
rect 2401 313 2506 329
rect 2401 279 2417 313
rect 2451 279 2506 313
rect 2401 263 2506 279
rect 2272 215 2302 237
rect 2476 225 2506 263
rect 1768 148 1798 174
rect 1846 148 1876 174
rect 1918 148 1948 174
rect 1087 96 1153 112
rect 1087 62 1103 96
rect 1137 76 1153 96
rect 1232 76 1262 127
rect 1339 101 1369 127
rect 1137 62 1262 76
rect 637 21 667 47
rect 709 21 739 47
rect 814 21 844 47
rect 886 21 916 47
rect 958 21 988 47
rect 1087 46 1262 62
rect 1425 57 1455 127
rect 1527 101 1557 127
rect 2114 105 2144 131
rect 2186 105 2216 131
rect 2272 57 2302 131
rect 1425 27 2302 57
rect 2476 31 2506 57
<< polycont >>
rect 1626 565 1660 599
rect 621 369 655 403
rect 41 275 75 309
rect 176 312 210 346
rect 944 337 978 371
rect 1673 380 1707 414
rect 41 207 75 241
rect 582 213 616 247
rect 830 241 864 275
rect 412 56 446 90
rect 1673 312 1707 346
rect 2161 380 2195 414
rect 1433 253 1467 287
rect 2161 312 2195 346
rect 2417 279 2451 313
rect 1103 62 1137 96
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 128 535 194 649
rect 322 619 388 649
rect 322 585 338 619
rect 372 585 388 619
rect 21 516 87 532
rect 21 482 37 516
rect 71 482 87 516
rect 21 446 87 482
rect 128 501 144 535
rect 178 501 194 535
rect 128 464 194 501
rect 230 556 280 572
rect 322 569 388 585
rect 537 599 603 615
rect 264 535 280 556
rect 537 565 553 599
rect 587 565 603 599
rect 537 535 603 565
rect 264 522 603 535
rect 230 503 603 522
rect 230 501 553 503
rect 21 412 37 446
rect 71 430 87 446
rect 230 446 294 501
rect 537 469 553 501
rect 587 469 603 503
rect 71 412 171 430
rect 21 396 171 412
rect 264 412 294 446
rect 230 396 294 412
rect 137 362 171 396
rect 25 309 91 356
rect 25 275 41 309
rect 75 275 91 309
rect 25 241 91 275
rect 25 207 41 241
rect 75 207 91 241
rect 25 191 91 207
rect 137 346 226 362
rect 137 312 176 346
rect 210 312 226 346
rect 137 296 226 312
rect 137 157 171 296
rect 260 262 294 396
rect 429 451 503 467
rect 429 417 445 451
rect 479 417 503 451
rect 429 296 503 417
rect 19 128 69 157
rect 19 94 35 128
rect 19 17 69 94
rect 105 128 171 157
rect 105 94 121 128
rect 155 94 171 128
rect 209 246 294 262
rect 209 212 225 246
rect 259 212 294 246
rect 209 176 294 212
rect 209 142 225 176
rect 259 142 294 176
rect 367 212 433 262
rect 367 178 383 212
rect 417 178 433 212
rect 367 163 433 178
rect 469 251 503 296
rect 537 453 603 469
rect 637 581 880 615
rect 537 319 571 453
rect 637 419 671 581
rect 605 403 671 419
rect 718 498 784 547
rect 718 464 734 498
rect 768 464 784 498
rect 718 415 784 464
rect 846 497 880 581
rect 923 590 1031 615
rect 1610 599 1686 615
rect 923 556 939 590
rect 973 581 1031 590
rect 973 556 991 581
rect 923 547 991 556
rect 1025 547 1031 581
rect 923 531 1031 547
rect 1362 581 1428 597
rect 1362 547 1375 581
rect 1412 547 1428 581
rect 1610 565 1626 599
rect 1660 565 1686 599
rect 2401 607 2467 649
rect 1610 549 1686 565
rect 1362 531 1428 547
rect 1652 498 1686 549
rect 1720 582 1799 598
rect 1754 581 1799 582
rect 1754 548 1759 581
rect 1720 547 1759 548
rect 1793 547 1799 581
rect 1720 532 1799 547
rect 1849 582 1988 598
rect 1849 581 1938 582
rect 1849 547 1855 581
rect 1889 548 1938 581
rect 1972 548 1988 582
rect 2401 573 2417 607
rect 2451 573 2467 607
rect 1889 547 1988 548
rect 1849 532 1988 547
rect 2051 556 2101 572
rect 2051 522 2067 556
rect 2051 498 2101 522
rect 2401 510 2467 573
rect 846 463 1618 497
rect 1652 485 2101 498
rect 1652 464 2067 485
rect 605 369 621 403
rect 655 369 671 403
rect 605 353 671 369
rect 537 285 700 319
rect 469 247 632 251
rect 469 227 582 247
rect 469 193 488 227
rect 522 213 582 227
rect 616 213 632 247
rect 522 197 632 213
rect 522 193 538 197
rect 469 170 538 193
rect 666 163 700 285
rect 209 126 294 142
rect 328 129 433 163
rect 576 158 700 163
rect 105 65 171 94
rect 328 17 362 129
rect 576 124 592 158
rect 626 124 700 158
rect 576 119 700 124
rect 734 179 768 415
rect 846 291 880 463
rect 928 400 1550 429
rect 928 395 1500 400
rect 928 371 994 395
rect 928 337 944 371
rect 978 337 994 371
rect 1484 366 1500 395
rect 1534 366 1550 400
rect 928 325 994 337
rect 1112 327 1128 361
rect 1162 327 1178 361
rect 1484 337 1550 366
rect 1112 325 1178 327
rect 1028 303 1450 325
rect 1028 291 1482 303
rect 814 275 880 291
rect 814 241 830 275
rect 864 241 880 275
rect 814 225 880 241
rect 914 257 1062 291
rect 1416 287 1482 291
rect 914 179 948 257
rect 1096 223 1328 257
rect 1416 253 1433 287
rect 1467 253 1482 287
rect 1416 237 1482 253
rect 1096 202 1130 223
rect 734 158 948 179
rect 734 124 750 158
rect 784 124 948 158
rect 734 119 948 124
rect 1003 169 1130 202
rect 1003 135 1019 169
rect 1053 168 1130 169
rect 1187 173 1237 189
rect 1003 119 1053 135
rect 1221 139 1237 173
rect 1087 112 1127 134
rect 1087 96 1153 112
rect 396 90 462 95
rect 396 56 412 90
rect 446 85 462 90
rect 1087 85 1103 96
rect 446 62 1103 85
rect 1137 62 1153 96
rect 446 56 1153 62
rect 396 51 1153 56
rect 1187 17 1237 139
rect 1278 186 1328 223
rect 1278 152 1294 186
rect 1278 123 1328 152
rect 1364 180 1430 203
rect 1364 146 1380 180
rect 1414 146 1430 180
rect 1516 194 1550 337
rect 1584 262 1618 463
rect 2051 451 2067 464
rect 1657 414 1723 430
rect 1657 380 1673 414
rect 1707 380 1723 414
rect 1657 346 1723 380
rect 1657 312 1673 346
rect 1707 312 1723 346
rect 1657 296 1723 312
rect 1813 414 1879 430
rect 1813 380 1829 414
rect 1863 380 1879 414
rect 1813 262 1879 380
rect 2051 414 2101 451
rect 2262 483 2328 499
rect 2262 449 2278 483
rect 2312 449 2328 483
rect 2051 380 2067 414
rect 1584 233 1879 262
rect 1584 228 1701 233
rect 1685 199 1701 228
rect 1735 228 1879 233
rect 1943 233 2009 262
rect 1735 199 1751 228
rect 1516 160 1641 194
rect 1685 170 1751 199
rect 1943 199 1959 233
rect 1993 199 2009 233
rect 1364 17 1430 146
rect 1575 148 1641 160
rect 1575 114 1591 148
rect 1625 114 1641 148
rect 1575 68 1641 114
rect 1943 17 2009 199
rect 2051 219 2101 380
rect 2137 414 2211 430
rect 2137 380 2161 414
rect 2195 380 2211 414
rect 2137 346 2211 380
rect 2137 312 2161 346
rect 2195 312 2211 346
rect 2137 296 2211 312
rect 2262 413 2328 449
rect 2262 379 2278 413
rect 2312 379 2328 413
rect 2262 329 2328 379
rect 2401 476 2417 510
rect 2451 476 2467 510
rect 2401 413 2467 476
rect 2401 379 2417 413
rect 2451 379 2467 413
rect 2401 363 2467 379
rect 2501 599 2567 615
rect 2501 565 2517 599
rect 2551 565 2567 599
rect 2501 506 2567 565
rect 2501 472 2517 506
rect 2551 472 2567 506
rect 2501 413 2567 472
rect 2501 379 2517 413
rect 2551 379 2567 413
rect 2262 313 2467 329
rect 2262 295 2417 313
rect 2297 279 2417 295
rect 2451 279 2467 313
rect 2297 263 2467 279
rect 2051 190 2119 219
rect 2051 156 2069 190
rect 2103 156 2119 190
rect 2051 127 2119 156
rect 2211 190 2261 219
rect 2211 156 2227 190
rect 2211 17 2261 156
rect 2297 190 2363 263
rect 2297 156 2313 190
rect 2347 156 2363 190
rect 2297 127 2363 156
rect 2415 213 2465 229
rect 2415 179 2431 213
rect 2415 103 2465 179
rect 2415 69 2431 103
rect 2415 17 2465 69
rect 2501 213 2567 379
rect 2501 179 2517 213
rect 2551 179 2567 213
rect 2501 103 2567 179
rect 2501 69 2517 103
rect 2551 69 2567 103
rect 2501 53 2567 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 991 547 1025 581
rect 1375 547 1378 581
rect 1378 547 1409 581
rect 1759 547 1793 581
rect 1855 547 1889 581
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
<< metal1 >>
rect 0 683 2592 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2592 683
rect 0 617 2592 649
rect 14 581 2578 589
rect 14 547 991 581
rect 1025 547 1375 581
rect 1409 547 1759 581
rect 1793 547 1855 581
rect 1889 547 2578 581
rect 14 535 2578 547
rect 0 17 2592 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2592 17
rect 0 -49 2592 -17
<< labels >>
flabel pwell s 0 0 2592 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2592 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 srdlstp_1
flabel metal1 s 14 535 2578 589 0 FreeSans 200 0 0 0 KAPWR
port 5 nsew power bidirectional
flabel metal1 s 0 617 2592 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2592 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1663 390 1697 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 2143 316 2177 350 0 FreeSans 340 0 0 0 SLEEP_B
port 4 nsew signal input
flabel locali s 2143 390 2177 424 0 FreeSans 340 0 0 0 SLEEP_B
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1087 94 1121 128 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 2527 94 2561 128 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2527 168 2561 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2527 242 2561 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2527 316 2561 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2527 390 2561 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2592 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3832836
string GDS_START 3815366
<< end >>
