magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 51 49 792 241
rect 0 0 864 49
<< scnmos >>
rect 130 47 160 215
rect 202 47 232 215
rect 310 47 340 215
rect 425 47 455 215
rect 511 47 541 215
rect 597 47 627 215
rect 683 47 713 215
<< scpmoshvt >>
rect 130 367 160 619
rect 232 367 262 619
rect 318 367 348 619
rect 425 367 455 619
rect 511 367 541 619
rect 597 367 627 619
rect 683 367 713 619
<< ndiff >>
rect 77 198 130 215
rect 77 164 85 198
rect 119 164 130 198
rect 77 93 130 164
rect 77 59 85 93
rect 119 59 130 93
rect 77 47 130 59
rect 160 47 202 215
rect 232 47 310 215
rect 340 129 425 215
rect 340 95 365 129
rect 399 95 425 129
rect 340 47 425 95
rect 455 203 511 215
rect 455 169 466 203
rect 500 169 511 203
rect 455 101 511 169
rect 455 67 466 101
rect 500 67 511 101
rect 455 47 511 67
rect 541 175 597 215
rect 541 141 552 175
rect 586 141 597 175
rect 541 93 597 141
rect 541 59 552 93
rect 586 59 597 93
rect 541 47 597 59
rect 627 203 683 215
rect 627 169 638 203
rect 672 169 683 203
rect 627 101 683 169
rect 627 67 638 101
rect 672 67 683 101
rect 627 47 683 67
rect 713 163 766 215
rect 713 129 724 163
rect 758 129 766 163
rect 713 93 766 129
rect 713 59 724 93
rect 758 59 766 93
rect 713 47 766 59
<< pdiff >>
rect 77 599 130 619
rect 77 565 85 599
rect 119 565 130 599
rect 77 512 130 565
rect 77 478 85 512
rect 119 478 130 512
rect 77 413 130 478
rect 77 379 85 413
rect 119 379 130 413
rect 77 367 130 379
rect 160 607 232 619
rect 160 573 179 607
rect 213 573 232 607
rect 160 527 232 573
rect 160 493 179 527
rect 213 493 232 527
rect 160 455 232 493
rect 160 421 179 455
rect 213 421 232 455
rect 160 367 232 421
rect 262 599 318 619
rect 262 565 273 599
rect 307 565 318 599
rect 262 512 318 565
rect 262 478 273 512
rect 307 478 318 512
rect 262 413 318 478
rect 262 379 273 413
rect 307 379 318 413
rect 262 367 318 379
rect 348 607 425 619
rect 348 573 369 607
rect 403 573 425 607
rect 348 527 425 573
rect 348 493 369 527
rect 403 493 425 527
rect 348 444 425 493
rect 348 410 369 444
rect 403 410 425 444
rect 348 367 425 410
rect 455 599 511 619
rect 455 565 466 599
rect 500 565 511 599
rect 455 512 511 565
rect 455 478 466 512
rect 500 478 511 512
rect 455 413 511 478
rect 455 379 466 413
rect 500 379 511 413
rect 455 367 511 379
rect 541 611 597 619
rect 541 577 552 611
rect 586 577 597 611
rect 541 532 597 577
rect 541 498 552 532
rect 586 498 597 532
rect 541 453 597 498
rect 541 419 552 453
rect 586 419 597 453
rect 541 367 597 419
rect 627 599 683 619
rect 627 565 638 599
rect 672 565 683 599
rect 627 512 683 565
rect 627 478 638 512
rect 672 478 683 512
rect 627 413 683 478
rect 627 379 638 413
rect 672 379 683 413
rect 627 367 683 379
rect 713 607 766 619
rect 713 573 724 607
rect 758 573 766 607
rect 713 532 766 573
rect 713 498 724 532
rect 758 498 766 532
rect 713 453 766 498
rect 713 419 724 453
rect 758 419 766 453
rect 713 367 766 419
<< ndiffc >>
rect 85 164 119 198
rect 85 59 119 93
rect 365 95 399 129
rect 466 169 500 203
rect 466 67 500 101
rect 552 141 586 175
rect 552 59 586 93
rect 638 169 672 203
rect 638 67 672 101
rect 724 129 758 163
rect 724 59 758 93
<< pdiffc >>
rect 85 565 119 599
rect 85 478 119 512
rect 85 379 119 413
rect 179 573 213 607
rect 179 493 213 527
rect 179 421 213 455
rect 273 565 307 599
rect 273 478 307 512
rect 273 379 307 413
rect 369 573 403 607
rect 369 493 403 527
rect 369 410 403 444
rect 466 565 500 599
rect 466 478 500 512
rect 466 379 500 413
rect 552 577 586 611
rect 552 498 586 532
rect 552 419 586 453
rect 638 565 672 599
rect 638 478 672 512
rect 638 379 672 413
rect 724 573 758 607
rect 724 498 758 532
rect 724 419 758 453
<< poly >>
rect 130 619 160 645
rect 232 619 262 645
rect 318 619 348 645
rect 425 619 455 645
rect 511 619 541 645
rect 597 619 627 645
rect 683 619 713 645
rect 130 303 160 367
rect 232 308 262 367
rect 318 308 348 367
rect 425 333 455 367
rect 511 333 541 367
rect 597 333 627 367
rect 683 333 713 367
rect 425 317 763 333
rect 94 287 160 303
rect 94 253 110 287
rect 144 253 160 287
rect 94 237 160 253
rect 130 215 160 237
rect 202 292 268 308
rect 202 258 218 292
rect 252 258 268 292
rect 202 242 268 258
rect 310 292 376 308
rect 310 258 326 292
rect 360 258 376 292
rect 310 242 376 258
rect 425 283 441 317
rect 475 283 509 317
rect 543 283 577 317
rect 611 283 645 317
rect 679 283 713 317
rect 747 283 763 317
rect 425 267 763 283
rect 202 215 232 242
rect 310 215 340 242
rect 425 215 455 267
rect 511 215 541 267
rect 597 215 627 267
rect 683 215 713 267
rect 130 21 160 47
rect 202 21 232 47
rect 310 21 340 47
rect 425 21 455 47
rect 511 21 541 47
rect 597 21 627 47
rect 683 21 713 47
<< polycont >>
rect 110 253 144 287
rect 218 258 252 292
rect 326 258 360 292
rect 441 283 475 317
rect 509 283 543 317
rect 577 283 611 317
rect 645 283 679 317
rect 713 283 747 317
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 69 599 123 615
rect 69 565 85 599
rect 119 565 123 599
rect 69 512 123 565
rect 69 478 85 512
rect 119 478 123 512
rect 69 413 123 478
rect 163 607 229 649
rect 163 573 179 607
rect 213 573 229 607
rect 163 527 229 573
rect 163 493 179 527
rect 213 493 229 527
rect 163 455 229 493
rect 163 421 179 455
rect 213 421 229 455
rect 270 599 319 615
rect 270 565 273 599
rect 307 565 319 599
rect 270 512 319 565
rect 270 478 273 512
rect 307 478 319 512
rect 69 379 85 413
rect 119 385 123 413
rect 270 413 319 478
rect 270 385 273 413
rect 119 379 273 385
rect 307 379 319 413
rect 353 607 419 649
rect 353 573 369 607
rect 403 573 419 607
rect 353 527 419 573
rect 353 493 369 527
rect 403 493 419 527
rect 353 444 419 493
rect 353 410 369 444
rect 403 410 419 444
rect 464 599 502 615
rect 464 565 466 599
rect 500 565 502 599
rect 464 512 502 565
rect 464 478 466 512
rect 500 478 502 512
rect 464 413 502 478
rect 536 611 602 649
rect 536 577 552 611
rect 586 577 602 611
rect 536 532 602 577
rect 536 498 552 532
rect 586 498 602 532
rect 536 453 602 498
rect 536 419 552 453
rect 586 419 602 453
rect 636 599 674 615
rect 636 565 638 599
rect 672 565 674 599
rect 636 512 674 565
rect 636 478 638 512
rect 672 478 674 512
rect 69 376 319 379
rect 464 379 466 413
rect 500 385 502 413
rect 636 413 674 478
rect 708 607 774 649
rect 708 573 724 607
rect 758 573 774 607
rect 708 532 774 573
rect 708 498 724 532
rect 758 498 774 532
rect 708 453 774 498
rect 708 419 724 453
rect 758 419 774 453
rect 636 385 638 413
rect 500 379 638 385
rect 672 385 674 413
rect 672 379 845 385
rect 69 342 430 376
rect 464 351 845 379
rect 396 317 430 342
rect 20 287 161 303
rect 20 253 110 287
rect 144 253 161 287
rect 20 242 161 253
rect 202 292 268 308
rect 202 258 218 292
rect 252 258 268 292
rect 202 242 268 258
rect 319 292 362 308
rect 319 258 326 292
rect 360 258 362 292
rect 319 242 362 258
rect 396 283 441 317
rect 475 283 509 317
rect 543 283 577 317
rect 611 283 645 317
rect 679 283 713 317
rect 747 283 763 317
rect 396 208 430 283
rect 799 247 845 351
rect 69 198 430 208
rect 69 164 85 198
rect 119 174 430 198
rect 464 213 845 247
rect 464 203 502 213
rect 119 164 135 174
rect 69 93 135 164
rect 464 169 466 203
rect 500 169 502 203
rect 636 203 674 213
rect 69 59 85 93
rect 119 59 135 93
rect 69 51 135 59
rect 349 129 415 140
rect 349 95 365 129
rect 399 95 415 129
rect 349 17 415 95
rect 464 101 502 169
rect 464 67 466 101
rect 500 67 502 101
rect 464 51 502 67
rect 536 175 602 179
rect 536 141 552 175
rect 586 141 602 175
rect 536 93 602 141
rect 536 59 552 93
rect 586 59 602 93
rect 536 17 602 59
rect 636 169 638 203
rect 672 169 674 203
rect 636 101 674 169
rect 636 67 638 101
rect 672 67 674 101
rect 636 51 674 67
rect 708 163 765 179
rect 708 129 724 163
rect 758 129 765 163
rect 708 93 765 129
rect 708 59 724 93
rect 758 59 765 93
rect 799 78 845 213
rect 708 17 765 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and3_4
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5182190
string GDS_START 5174338
<< end >>
