magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 718 251
rect 0 0 768 49
<< scnmos >>
rect 84 141 114 225
rect 156 141 186 225
rect 243 141 273 225
rect 329 141 359 225
rect 447 141 477 225
rect 533 141 563 225
rect 605 141 635 225
<< scpmoshvt >>
rect 87 419 137 619
rect 208 419 258 619
rect 306 419 356 619
rect 414 419 464 619
rect 522 419 572 619
rect 630 419 680 619
<< ndiff >>
rect 27 194 84 225
rect 27 160 39 194
rect 73 160 84 194
rect 27 141 84 160
rect 114 141 156 225
rect 186 194 243 225
rect 186 160 197 194
rect 231 160 243 194
rect 186 141 243 160
rect 273 200 329 225
rect 273 166 284 200
rect 318 166 329 200
rect 273 141 329 166
rect 359 187 447 225
rect 359 153 386 187
rect 420 153 447 187
rect 359 141 447 153
rect 477 200 533 225
rect 477 166 488 200
rect 522 166 533 200
rect 477 141 533 166
rect 563 141 605 225
rect 635 198 692 225
rect 635 164 646 198
rect 680 164 692 198
rect 635 141 692 164
<< pdiff >>
rect 30 597 87 619
rect 30 563 42 597
rect 76 563 87 597
rect 30 473 87 563
rect 30 439 42 473
rect 76 439 87 473
rect 30 419 87 439
rect 137 573 208 619
rect 137 539 148 573
rect 182 539 208 573
rect 137 419 208 539
rect 258 419 306 619
rect 356 419 414 619
rect 464 597 522 619
rect 464 563 475 597
rect 509 563 522 597
rect 464 470 522 563
rect 464 436 475 470
rect 509 436 522 470
rect 464 419 522 436
rect 572 573 630 619
rect 572 539 583 573
rect 617 539 630 573
rect 572 419 630 539
rect 680 597 737 619
rect 680 563 691 597
rect 725 563 737 597
rect 680 470 737 563
rect 680 436 691 470
rect 725 436 737 470
rect 680 419 737 436
<< ndiffc >>
rect 39 160 73 194
rect 197 160 231 194
rect 284 166 318 200
rect 386 153 420 187
rect 488 166 522 200
rect 646 164 680 198
<< pdiffc >>
rect 42 563 76 597
rect 42 439 76 473
rect 148 539 182 573
rect 475 563 509 597
rect 475 436 509 470
rect 583 539 617 573
rect 691 563 725 597
rect 691 436 725 470
<< poly >>
rect 87 619 137 645
rect 208 619 258 645
rect 306 619 356 645
rect 414 619 464 645
rect 522 619 572 645
rect 630 619 680 645
rect 87 387 137 419
rect 84 371 156 387
rect 208 384 258 419
rect 306 384 356 419
rect 84 337 106 371
rect 140 337 156 371
rect 84 303 156 337
rect 198 368 264 384
rect 198 334 214 368
rect 248 334 264 368
rect 198 318 264 334
rect 306 368 372 384
rect 306 334 322 368
rect 356 334 372 368
rect 306 318 372 334
rect 414 376 464 419
rect 522 384 572 419
rect 630 384 680 419
rect 414 360 480 376
rect 414 326 430 360
rect 464 326 480 360
rect 84 269 106 303
rect 140 270 156 303
rect 234 270 264 318
rect 140 269 186 270
rect 84 240 186 269
rect 234 240 273 270
rect 84 225 114 240
rect 156 225 186 240
rect 243 225 273 240
rect 329 225 359 318
rect 414 310 480 326
rect 522 368 588 384
rect 522 334 538 368
rect 572 334 588 368
rect 522 318 588 334
rect 630 368 696 384
rect 630 334 646 368
rect 680 334 696 368
rect 630 318 696 334
rect 447 225 477 310
rect 533 225 563 318
rect 630 270 660 318
rect 605 240 660 270
rect 605 225 635 240
rect 84 115 114 141
rect 156 115 186 141
rect 243 115 273 141
rect 329 115 359 141
rect 447 115 477 141
rect 533 115 563 141
rect 605 115 635 141
<< polycont >>
rect 106 337 140 371
rect 214 334 248 368
rect 322 334 356 368
rect 430 326 464 360
rect 106 269 140 303
rect 538 334 572 368
rect 646 334 680 368
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 20 597 92 613
rect 20 563 42 597
rect 76 563 92 597
rect 20 473 92 563
rect 132 573 198 649
rect 132 539 148 573
rect 182 539 198 573
rect 132 490 198 539
rect 459 597 525 613
rect 459 563 475 597
rect 509 563 525 597
rect 20 439 42 473
rect 76 439 92 473
rect 459 470 525 563
rect 567 573 633 649
rect 567 539 583 573
rect 617 539 633 573
rect 567 490 633 539
rect 691 597 750 613
rect 725 563 750 597
rect 459 454 475 470
rect 20 423 92 439
rect 128 436 475 454
rect 509 454 525 470
rect 691 470 750 563
rect 509 436 691 454
rect 725 436 750 470
rect 20 217 54 423
rect 128 420 750 436
rect 128 387 162 420
rect 90 371 162 387
rect 90 337 106 371
rect 140 337 162 371
rect 90 303 162 337
rect 198 368 264 384
rect 198 334 214 368
rect 248 334 264 368
rect 198 310 264 334
rect 306 368 372 384
rect 306 334 322 368
rect 356 334 372 368
rect 306 310 372 334
rect 409 360 472 376
rect 409 326 430 360
rect 464 326 472 360
rect 409 310 472 326
rect 506 368 572 384
rect 506 334 538 368
rect 506 310 572 334
rect 606 368 682 384
rect 606 334 646 368
rect 680 334 682 368
rect 606 310 682 334
rect 90 269 106 303
rect 140 269 162 303
rect 90 253 162 269
rect 300 240 538 274
rect 300 229 334 240
rect 20 194 89 217
rect 20 160 39 194
rect 73 160 89 194
rect 20 88 89 160
rect 181 194 231 217
rect 181 160 197 194
rect 181 17 231 160
rect 268 200 334 229
rect 268 166 284 200
rect 318 166 334 200
rect 268 137 334 166
rect 370 187 436 204
rect 370 153 386 187
rect 420 153 436 187
rect 370 17 436 153
rect 472 200 538 240
rect 716 214 750 420
rect 472 166 488 200
rect 522 166 538 200
rect 472 137 538 166
rect 630 198 750 214
rect 630 164 646 198
rect 680 164 750 198
rect 630 148 750 164
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o311a_lp
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4398902
string GDS_START 4392534
<< end >>
