magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 1 157 433 161
rect 1 49 1051 157
rect 0 0 1056 49
<< scnmos >>
rect 84 51 114 135
rect 156 51 186 135
rect 242 51 272 135
rect 320 51 350 135
rect 518 47 548 131
rect 596 47 626 131
rect 674 47 704 131
rect 752 47 782 131
rect 866 47 896 131
rect 938 47 968 131
<< scpmoshvt >>
rect 84 401 134 601
rect 348 409 398 609
rect 454 409 504 609
rect 560 409 610 609
rect 682 409 732 609
rect 788 409 838 609
rect 915 409 965 609
<< ndiff >>
rect 27 113 84 135
rect 27 79 39 113
rect 73 79 84 113
rect 27 51 84 79
rect 114 51 156 135
rect 186 101 242 135
rect 186 67 197 101
rect 231 67 242 101
rect 186 51 242 67
rect 272 51 320 135
rect 350 113 407 135
rect 350 79 361 113
rect 395 79 407 113
rect 350 51 407 79
rect 461 103 518 131
rect 461 69 473 103
rect 507 69 518 103
rect 461 47 518 69
rect 548 47 596 131
rect 626 47 674 131
rect 704 47 752 131
rect 782 97 866 131
rect 782 63 793 97
rect 827 63 866 97
rect 782 47 866 63
rect 896 47 938 131
rect 968 111 1025 131
rect 968 77 979 111
rect 1013 77 1025 111
rect 968 47 1025 77
<< pdiff >>
rect 27 589 84 601
rect 27 555 39 589
rect 73 555 84 589
rect 27 518 84 555
rect 27 484 39 518
rect 73 484 84 518
rect 27 447 84 484
rect 27 413 39 447
rect 73 413 84 447
rect 27 401 84 413
rect 134 589 191 601
rect 134 555 145 589
rect 179 555 191 589
rect 134 518 191 555
rect 134 484 145 518
rect 179 484 191 518
rect 134 447 191 484
rect 134 413 145 447
rect 179 413 191 447
rect 134 401 191 413
rect 291 597 348 609
rect 291 563 303 597
rect 337 563 348 597
rect 291 526 348 563
rect 291 492 303 526
rect 337 492 348 526
rect 291 455 348 492
rect 291 421 303 455
rect 337 421 348 455
rect 291 409 348 421
rect 398 597 454 609
rect 398 563 409 597
rect 443 563 454 597
rect 398 517 454 563
rect 398 483 409 517
rect 443 483 454 517
rect 398 409 454 483
rect 504 597 560 609
rect 504 563 515 597
rect 549 563 560 597
rect 504 517 560 563
rect 504 483 515 517
rect 549 483 560 517
rect 504 409 560 483
rect 610 592 682 609
rect 610 558 621 592
rect 655 558 682 592
rect 610 409 682 558
rect 732 597 788 609
rect 732 563 743 597
rect 777 563 788 597
rect 732 526 788 563
rect 732 492 743 526
rect 777 492 788 526
rect 732 455 788 492
rect 732 421 743 455
rect 777 421 788 455
rect 732 409 788 421
rect 838 597 915 609
rect 838 563 849 597
rect 883 563 915 597
rect 838 514 915 563
rect 838 480 849 514
rect 883 480 915 514
rect 838 409 915 480
rect 965 597 1022 609
rect 965 563 976 597
rect 1010 563 1022 597
rect 965 526 1022 563
rect 965 492 976 526
rect 1010 492 1022 526
rect 965 455 1022 492
rect 965 421 976 455
rect 1010 421 1022 455
rect 965 409 1022 421
<< ndiffc >>
rect 39 79 73 113
rect 197 67 231 101
rect 361 79 395 113
rect 473 69 507 103
rect 793 63 827 97
rect 979 77 1013 111
<< pdiffc >>
rect 39 555 73 589
rect 39 484 73 518
rect 39 413 73 447
rect 145 555 179 589
rect 145 484 179 518
rect 145 413 179 447
rect 303 563 337 597
rect 303 492 337 526
rect 303 421 337 455
rect 409 563 443 597
rect 409 483 443 517
rect 515 563 549 597
rect 515 483 549 517
rect 621 558 655 592
rect 743 563 777 597
rect 743 492 777 526
rect 743 421 777 455
rect 849 563 883 597
rect 849 480 883 514
rect 976 563 1010 597
rect 976 492 1010 526
rect 976 421 1010 455
<< poly >>
rect 84 601 134 627
rect 348 609 398 635
rect 454 609 504 635
rect 560 609 610 635
rect 682 609 732 635
rect 788 609 838 635
rect 915 609 965 635
rect 84 291 134 401
rect 348 291 398 409
rect 454 361 504 409
rect 560 377 610 409
rect 560 361 626 377
rect 84 275 191 291
rect 84 241 141 275
rect 175 241 191 275
rect 312 275 398 291
rect 312 255 328 275
rect 84 207 191 241
rect 84 173 141 207
rect 175 173 191 207
rect 84 157 191 173
rect 242 241 328 255
rect 362 261 398 275
rect 446 345 512 361
rect 446 311 462 345
rect 496 311 512 345
rect 446 277 512 311
rect 362 241 378 261
rect 242 225 378 241
rect 446 243 462 277
rect 496 243 512 277
rect 560 327 576 361
rect 610 327 626 361
rect 682 358 732 409
rect 788 358 838 409
rect 560 293 626 327
rect 560 259 576 293
rect 610 259 626 293
rect 560 243 626 259
rect 446 227 512 243
rect 84 135 114 157
rect 156 135 186 157
rect 242 135 272 225
rect 320 135 350 225
rect 482 195 512 227
rect 482 165 548 195
rect 518 131 548 165
rect 596 131 626 243
rect 674 342 740 358
rect 674 308 690 342
rect 724 308 740 342
rect 674 274 740 308
rect 674 240 690 274
rect 724 240 740 274
rect 674 224 740 240
rect 788 342 854 358
rect 788 308 804 342
rect 838 308 854 342
rect 915 322 965 409
rect 788 274 854 308
rect 788 240 804 274
rect 838 240 854 274
rect 788 224 854 240
rect 902 306 968 322
rect 902 272 918 306
rect 952 272 968 306
rect 902 238 968 272
rect 674 131 704 224
rect 788 176 818 224
rect 902 204 918 238
rect 952 204 968 238
rect 902 176 968 204
rect 752 146 818 176
rect 866 146 968 176
rect 752 131 782 146
rect 866 131 896 146
rect 938 131 968 146
rect 84 25 114 51
rect 156 25 186 51
rect 242 25 272 51
rect 320 25 350 51
rect 518 21 548 47
rect 596 21 626 47
rect 674 21 704 47
rect 752 21 782 47
rect 866 21 896 47
rect 938 21 968 47
<< polycont >>
rect 141 241 175 275
rect 141 173 175 207
rect 328 241 362 275
rect 462 311 496 345
rect 462 243 496 277
rect 576 327 610 361
rect 576 259 610 293
rect 690 308 724 342
rect 690 240 724 274
rect 804 308 838 342
rect 804 240 838 274
rect 918 272 952 306
rect 918 204 952 238
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 589 89 605
rect 23 555 39 589
rect 73 555 89 589
rect 23 518 89 555
rect 23 484 39 518
rect 73 484 89 518
rect 23 447 89 484
rect 23 413 39 447
rect 73 413 89 447
rect 23 361 89 413
rect 129 589 195 649
rect 129 555 145 589
rect 179 555 195 589
rect 129 518 195 555
rect 129 484 145 518
rect 179 484 195 518
rect 129 447 195 484
rect 129 413 145 447
rect 179 413 195 447
rect 129 397 195 413
rect 287 597 353 613
rect 287 563 303 597
rect 337 563 353 597
rect 287 526 353 563
rect 287 492 303 526
rect 337 492 353 526
rect 287 455 353 492
rect 393 597 459 649
rect 393 563 409 597
rect 443 563 459 597
rect 393 517 459 563
rect 393 483 409 517
rect 443 483 459 517
rect 393 467 459 483
rect 499 597 565 613
rect 499 563 515 597
rect 549 563 565 597
rect 499 517 565 563
rect 605 592 671 649
rect 605 558 621 592
rect 655 558 671 592
rect 605 537 671 558
rect 727 597 793 613
rect 727 563 743 597
rect 777 563 793 597
rect 499 483 515 517
rect 549 501 565 517
rect 727 526 793 563
rect 727 501 743 526
rect 549 492 743 501
rect 777 492 793 526
rect 549 483 793 492
rect 499 467 793 483
rect 287 421 303 455
rect 337 431 353 455
rect 727 455 793 467
rect 833 597 899 649
rect 833 563 849 597
rect 883 563 899 597
rect 833 514 899 563
rect 833 480 849 514
rect 883 480 899 514
rect 833 464 899 480
rect 960 597 1038 613
rect 960 563 976 597
rect 1010 563 1038 597
rect 960 526 1038 563
rect 960 492 976 526
rect 1010 492 1038 526
rect 337 421 594 431
rect 287 397 594 421
rect 560 377 594 397
rect 727 421 743 455
rect 777 428 793 455
rect 960 455 1038 492
rect 777 421 924 428
rect 727 394 924 421
rect 560 361 626 377
rect 23 345 512 361
rect 23 327 462 345
rect 23 113 89 327
rect 446 311 462 327
rect 496 311 512 345
rect 125 275 263 291
rect 125 241 141 275
rect 175 241 263 275
rect 125 207 263 241
rect 312 275 378 291
rect 312 241 328 275
rect 362 241 378 275
rect 312 225 378 241
rect 446 277 512 311
rect 446 243 462 277
rect 496 243 512 277
rect 446 227 512 243
rect 560 327 576 361
rect 610 327 626 361
rect 560 293 626 327
rect 560 259 576 293
rect 610 259 626 293
rect 560 243 626 259
rect 674 342 743 358
rect 674 308 690 342
rect 724 308 743 342
rect 674 274 743 308
rect 125 173 141 207
rect 175 173 263 207
rect 560 189 594 243
rect 674 240 690 274
rect 724 240 743 274
rect 674 224 743 240
rect 788 342 854 358
rect 788 308 804 342
rect 838 308 854 342
rect 788 274 854 308
rect 788 240 804 274
rect 838 240 854 274
rect 788 224 854 240
rect 890 322 924 394
rect 960 421 976 455
rect 1010 421 1038 455
rect 960 384 1038 421
rect 890 306 968 322
rect 890 272 918 306
rect 952 272 968 306
rect 890 238 968 272
rect 125 157 263 173
rect 345 155 594 189
rect 890 204 918 238
rect 952 204 968 238
rect 890 188 968 204
rect 23 79 39 113
rect 73 79 89 113
rect 23 53 89 79
rect 181 101 247 121
rect 181 67 197 101
rect 231 67 247 101
rect 181 17 247 67
rect 345 113 411 155
rect 662 154 924 188
rect 662 119 696 154
rect 1004 135 1038 384
rect 345 79 361 113
rect 395 79 411 113
rect 345 53 411 79
rect 457 103 696 119
rect 457 69 473 103
rect 507 69 696 103
rect 457 53 696 69
rect 777 97 843 118
rect 777 63 793 97
rect 827 63 843 97
rect 777 17 843 63
rect 963 111 1038 135
rect 963 77 979 111
rect 1013 77 1038 111
rect 963 53 1038 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4bb_lp
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 991 464 1025 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 991 538 1025 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5150578
string GDS_START 5141520
<< end >>
