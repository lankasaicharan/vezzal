magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 1 235 380 243
rect 1 49 959 235
rect 0 0 960 49
<< scnmos >>
rect 80 133 110 217
rect 185 49 215 217
rect 271 49 301 217
rect 486 125 516 209
rect 558 125 588 209
rect 666 125 696 209
rect 738 125 768 209
rect 846 125 876 209
<< scpmoshvt >>
rect 93 367 123 451
rect 198 367 228 619
rect 284 367 314 619
rect 486 415 516 499
rect 572 415 602 499
rect 666 415 696 499
rect 759 415 789 499
rect 846 415 876 499
<< ndiff >>
rect 27 192 80 217
rect 27 158 35 192
rect 69 158 80 192
rect 27 133 80 158
rect 110 181 185 217
rect 110 147 121 181
rect 155 147 185 181
rect 110 133 185 147
rect 132 95 185 133
rect 132 61 140 95
rect 174 61 185 95
rect 132 49 185 61
rect 215 205 271 217
rect 215 171 226 205
rect 260 171 271 205
rect 215 101 271 171
rect 215 67 226 101
rect 260 67 271 101
rect 215 49 271 67
rect 301 165 354 217
rect 301 131 312 165
rect 346 131 354 165
rect 301 95 354 131
rect 433 184 486 209
rect 433 150 441 184
rect 475 150 486 184
rect 433 125 486 150
rect 516 125 558 209
rect 588 125 666 209
rect 696 125 738 209
rect 768 198 846 209
rect 768 164 779 198
rect 813 164 846 198
rect 768 125 846 164
rect 876 201 933 209
rect 876 167 887 201
rect 921 167 933 201
rect 876 125 933 167
rect 301 61 312 95
rect 346 61 354 95
rect 301 49 354 61
<< pdiff >>
rect 145 583 198 619
rect 145 549 153 583
rect 187 549 198 583
rect 145 451 198 549
rect 40 434 93 451
rect 40 400 48 434
rect 82 400 93 434
rect 40 367 93 400
rect 123 367 198 451
rect 228 437 284 619
rect 228 403 239 437
rect 273 403 284 437
rect 228 367 284 403
rect 314 583 367 619
rect 314 549 325 583
rect 359 549 367 583
rect 314 499 367 549
rect 314 477 486 499
rect 314 443 401 477
rect 435 443 486 477
rect 314 415 486 443
rect 516 474 572 499
rect 516 440 527 474
rect 561 440 572 474
rect 516 415 572 440
rect 602 491 666 499
rect 602 457 613 491
rect 647 457 666 491
rect 602 415 666 457
rect 696 474 759 499
rect 696 440 707 474
rect 741 440 759 474
rect 696 415 759 440
rect 789 474 846 499
rect 789 440 800 474
rect 834 440 846 474
rect 789 415 846 440
rect 876 474 929 499
rect 876 440 887 474
rect 921 440 929 474
rect 876 415 929 440
rect 314 367 367 415
<< ndiffc >>
rect 35 158 69 192
rect 121 147 155 181
rect 140 61 174 95
rect 226 171 260 205
rect 226 67 260 101
rect 312 131 346 165
rect 441 150 475 184
rect 779 164 813 198
rect 887 167 921 201
rect 312 61 346 95
<< pdiffc >>
rect 153 549 187 583
rect 48 400 82 434
rect 239 403 273 437
rect 325 549 359 583
rect 401 443 435 477
rect 527 440 561 474
rect 613 457 647 491
rect 707 440 741 474
rect 800 440 834 474
rect 887 440 921 474
<< poly >>
rect 198 619 228 645
rect 284 619 314 645
rect 93 451 123 477
rect 651 588 717 604
rect 651 554 667 588
rect 701 554 717 588
rect 651 538 717 554
rect 486 499 516 525
rect 572 499 602 525
rect 666 499 696 538
rect 759 499 789 525
rect 846 499 876 525
rect 93 335 123 367
rect 44 319 123 335
rect 44 285 60 319
rect 94 305 123 319
rect 94 285 110 305
rect 198 287 228 367
rect 284 323 314 367
rect 486 335 516 415
rect 572 367 602 415
rect 284 307 350 323
rect 284 287 300 307
rect 44 269 110 285
rect 80 217 110 269
rect 185 273 300 287
rect 334 273 350 307
rect 185 257 350 273
rect 392 319 516 335
rect 392 285 408 319
rect 442 285 516 319
rect 392 269 516 285
rect 185 217 215 257
rect 271 217 301 257
rect 80 107 110 133
rect 486 209 516 269
rect 558 351 624 367
rect 558 317 574 351
rect 608 317 624 351
rect 558 283 624 317
rect 558 249 574 283
rect 608 249 624 283
rect 558 233 624 249
rect 558 209 588 233
rect 666 209 696 415
rect 759 297 789 415
rect 846 375 876 415
rect 846 345 882 375
rect 738 281 804 297
rect 738 247 754 281
rect 788 247 804 281
rect 852 261 882 345
rect 738 231 804 247
rect 846 231 882 261
rect 738 209 768 231
rect 846 209 876 231
rect 486 99 516 125
rect 558 99 588 125
rect 666 99 696 125
rect 738 99 768 125
rect 846 103 876 125
rect 828 87 894 103
rect 828 53 844 87
rect 878 53 894 87
rect 185 23 215 49
rect 271 23 301 49
rect 828 37 894 53
<< polycont >>
rect 667 554 701 588
rect 60 285 94 319
rect 300 273 334 307
rect 408 285 442 319
rect 574 317 608 351
rect 574 249 608 283
rect 754 247 788 281
rect 844 53 878 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 137 583 203 649
rect 137 549 153 583
rect 187 549 203 583
rect 137 545 203 549
rect 309 583 444 649
rect 309 549 325 583
rect 359 549 444 583
rect 309 545 444 549
rect 146 477 357 511
rect 32 434 180 477
rect 32 400 48 434
rect 82 400 180 434
rect 32 384 180 400
rect 17 319 110 350
rect 17 285 60 319
rect 94 285 110 319
rect 146 249 180 384
rect 19 215 180 249
rect 216 437 289 443
rect 216 403 239 437
rect 273 403 289 437
rect 216 387 289 403
rect 323 393 357 477
rect 391 477 444 545
rect 597 504 631 649
rect 667 588 747 604
rect 701 554 747 588
rect 667 538 747 554
rect 597 491 663 504
rect 391 443 401 477
rect 435 443 444 477
rect 391 427 444 443
rect 478 474 563 490
rect 478 440 527 474
rect 561 440 563 474
rect 597 457 613 491
rect 647 457 663 491
rect 597 455 663 457
rect 697 474 747 490
rect 478 421 563 440
rect 697 440 707 474
rect 741 440 747 474
rect 697 421 747 440
rect 781 474 837 649
rect 781 440 800 474
rect 834 440 837 474
rect 781 424 837 440
rect 871 474 937 490
rect 871 440 887 474
rect 921 440 937 474
rect 19 192 71 215
rect 19 158 35 192
rect 69 158 71 192
rect 216 205 262 387
rect 323 359 444 393
rect 19 142 71 158
rect 105 147 121 181
rect 155 147 182 181
rect 105 95 182 147
rect 105 61 140 95
rect 174 61 182 95
rect 105 17 182 61
rect 216 171 226 205
rect 260 171 262 205
rect 296 307 350 323
rect 296 273 300 307
rect 334 273 350 307
rect 296 235 350 273
rect 392 319 444 359
rect 392 285 408 319
rect 442 285 444 319
rect 392 269 444 285
rect 478 387 747 421
rect 478 235 512 387
rect 871 353 937 440
rect 558 351 937 353
rect 558 317 574 351
rect 608 317 937 351
rect 558 283 624 317
rect 558 249 574 283
rect 608 249 624 283
rect 682 281 837 283
rect 682 247 754 281
rect 788 247 837 281
rect 682 236 837 247
rect 296 199 512 235
rect 216 101 262 171
rect 425 184 512 199
rect 216 67 226 101
rect 260 67 262 101
rect 216 51 262 67
rect 296 131 312 165
rect 346 131 362 165
rect 425 150 441 184
rect 475 150 512 184
rect 425 134 512 150
rect 687 198 829 202
rect 687 164 779 198
rect 813 164 829 198
rect 871 201 937 317
rect 871 167 887 201
rect 921 167 937 201
rect 871 164 937 167
rect 296 95 362 131
rect 296 61 312 95
rect 346 61 362 95
rect 296 17 362 61
rect 687 17 755 164
rect 789 87 929 130
rect 789 53 844 87
rect 878 53 929 87
rect 789 51 929 53
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4bb_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 895 94 929 128 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5251790
string GDS_START 5243786
<< end >>
