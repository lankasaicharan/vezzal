magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 241 325 263
rect 1 49 707 241
rect 0 0 768 49
<< scnmos >>
rect 80 69 110 237
rect 212 153 242 237
rect 406 47 436 215
rect 526 47 556 215
rect 598 47 628 215
<< scpmoshvt >>
rect 102 367 132 619
rect 207 367 237 451
rect 406 367 436 619
rect 492 367 522 619
rect 598 367 628 619
<< ndiff >>
rect 27 225 80 237
rect 27 191 35 225
rect 69 191 80 225
rect 27 115 80 191
rect 27 81 35 115
rect 69 81 80 115
rect 27 69 80 81
rect 110 153 212 237
rect 242 229 299 237
rect 242 195 253 229
rect 287 195 299 229
rect 242 153 299 195
rect 110 93 190 153
rect 110 69 144 93
rect 132 59 144 69
rect 178 59 190 93
rect 132 43 190 59
rect 353 93 406 215
rect 353 59 361 93
rect 395 59 406 93
rect 353 47 406 59
rect 436 203 526 215
rect 436 169 465 203
rect 499 169 526 203
rect 436 93 526 169
rect 436 59 465 93
rect 499 59 526 93
rect 436 47 526 59
rect 556 47 598 215
rect 628 203 681 215
rect 628 169 639 203
rect 673 169 681 203
rect 628 93 681 169
rect 628 59 639 93
rect 673 59 681 93
rect 628 47 681 59
<< pdiff >>
rect 49 599 102 619
rect 49 565 57 599
rect 91 565 102 599
rect 49 509 102 565
rect 49 475 57 509
rect 91 475 102 509
rect 49 413 102 475
rect 49 379 57 413
rect 91 379 102 413
rect 49 367 102 379
rect 132 574 185 619
rect 132 540 143 574
rect 177 540 185 574
rect 132 451 185 540
rect 353 599 406 619
rect 353 565 361 599
rect 395 565 406 599
rect 353 508 406 565
rect 353 474 361 508
rect 395 474 406 508
rect 132 367 207 451
rect 237 424 290 451
rect 237 390 248 424
rect 282 390 290 424
rect 237 367 290 390
rect 353 419 406 474
rect 353 385 361 419
rect 395 385 406 419
rect 353 367 406 385
rect 436 599 492 619
rect 436 565 447 599
rect 481 565 492 599
rect 436 508 492 565
rect 436 474 447 508
rect 481 474 492 508
rect 436 413 492 474
rect 436 379 447 413
rect 481 379 492 413
rect 436 367 492 379
rect 522 607 598 619
rect 522 573 543 607
rect 577 573 598 607
rect 522 515 598 573
rect 522 481 543 515
rect 577 481 598 515
rect 522 428 598 481
rect 522 394 543 428
rect 577 394 598 428
rect 522 367 598 394
rect 628 599 681 619
rect 628 565 639 599
rect 673 565 681 599
rect 628 508 681 565
rect 628 474 639 508
rect 673 474 681 508
rect 628 413 681 474
rect 628 379 639 413
rect 673 379 681 413
rect 628 367 681 379
<< ndiffc >>
rect 35 191 69 225
rect 35 81 69 115
rect 253 195 287 229
rect 144 59 178 93
rect 361 59 395 93
rect 465 169 499 203
rect 465 59 499 93
rect 639 169 673 203
rect 639 59 673 93
<< pdiffc >>
rect 57 565 91 599
rect 57 475 91 509
rect 57 379 91 413
rect 143 540 177 574
rect 361 565 395 599
rect 361 474 395 508
rect 248 390 282 424
rect 361 385 395 419
rect 447 565 481 599
rect 447 474 481 508
rect 447 379 481 413
rect 543 573 577 607
rect 543 481 577 515
rect 543 394 577 428
rect 639 565 673 599
rect 639 474 673 508
rect 639 379 673 413
<< poly >>
rect 102 619 132 645
rect 406 619 436 645
rect 492 619 522 645
rect 598 619 628 645
rect 207 451 237 477
rect 102 325 132 367
rect 207 335 237 367
rect 406 335 436 367
rect 80 309 159 325
rect 80 275 109 309
rect 143 275 159 309
rect 80 259 159 275
rect 207 319 273 335
rect 207 285 223 319
rect 257 285 273 319
rect 207 269 273 285
rect 329 319 436 335
rect 329 285 345 319
rect 379 285 436 319
rect 492 303 522 367
rect 598 303 628 367
rect 329 269 436 285
rect 80 237 110 259
rect 212 237 242 269
rect 406 215 436 269
rect 490 287 556 303
rect 490 253 506 287
rect 540 253 556 287
rect 490 237 556 253
rect 526 215 556 237
rect 598 287 670 303
rect 598 253 620 287
rect 654 253 670 287
rect 598 237 670 253
rect 598 215 628 237
rect 212 127 242 153
rect 80 43 110 69
rect 406 21 436 47
rect 526 21 556 47
rect 598 21 628 47
<< polycont >>
rect 109 275 143 309
rect 223 285 257 319
rect 345 285 379 319
rect 506 253 540 287
rect 620 253 654 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 599 93 615
rect 17 565 57 599
rect 91 565 93 599
rect 17 509 93 565
rect 127 574 193 649
rect 127 540 143 574
rect 177 540 193 574
rect 127 532 193 540
rect 345 599 405 615
rect 345 565 361 599
rect 395 565 405 599
rect 17 475 57 509
rect 91 475 93 509
rect 345 508 405 565
rect 345 498 361 508
rect 17 413 93 475
rect 17 379 57 413
rect 91 379 93 413
rect 17 363 93 379
rect 131 474 361 498
rect 395 474 405 508
rect 131 464 405 474
rect 17 225 73 363
rect 131 325 165 464
rect 232 424 327 428
rect 232 390 248 424
rect 282 390 327 424
rect 232 386 327 390
rect 107 309 165 325
rect 107 275 109 309
rect 143 275 165 309
rect 107 259 165 275
rect 201 319 257 350
rect 201 285 223 319
rect 201 269 257 285
rect 293 335 327 386
rect 361 419 405 464
rect 395 385 405 419
rect 361 369 405 385
rect 439 599 491 615
rect 439 565 447 599
rect 481 565 491 599
rect 439 508 491 565
rect 439 474 447 508
rect 481 474 491 508
rect 439 413 491 474
rect 439 379 447 413
rect 481 379 491 413
rect 527 607 593 649
rect 527 573 543 607
rect 577 573 593 607
rect 527 515 593 573
rect 527 481 543 515
rect 577 481 593 515
rect 527 428 593 481
rect 527 394 543 428
rect 577 394 593 428
rect 635 599 683 615
rect 635 565 639 599
rect 673 565 683 599
rect 635 508 683 565
rect 635 474 639 508
rect 673 474 683 508
rect 635 413 683 474
rect 439 360 491 379
rect 635 379 639 413
rect 673 379 683 413
rect 635 360 683 379
rect 293 319 379 335
rect 439 326 683 360
rect 293 285 345 319
rect 293 269 379 285
rect 415 287 562 292
rect 17 191 35 225
rect 69 191 73 225
rect 17 115 73 191
rect 131 161 165 259
rect 293 235 327 269
rect 415 253 506 287
rect 540 253 562 287
rect 415 242 562 253
rect 604 287 751 292
rect 604 253 620 287
rect 654 253 751 287
rect 604 242 751 253
rect 237 229 327 235
rect 237 195 253 229
rect 287 195 327 229
rect 449 203 515 208
rect 449 169 465 203
rect 499 169 515 203
rect 449 161 515 169
rect 131 127 515 161
rect 17 81 35 115
rect 69 81 73 115
rect 449 93 515 127
rect 17 65 73 81
rect 128 59 144 93
rect 178 59 194 93
rect 128 17 194 59
rect 345 59 361 93
rect 395 59 411 93
rect 345 17 411 59
rect 449 59 465 93
rect 499 59 515 93
rect 449 51 515 59
rect 623 203 689 208
rect 623 169 639 203
rect 673 169 689 203
rect 623 93 689 169
rect 623 59 639 93
rect 673 59 689 93
rect 623 17 689 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21bo_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3770668
string GDS_START 3763218
<< end >>
