magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 502 243 1343 259
rect 22 49 1343 243
rect 0 0 1344 49
<< scnmos >>
rect 101 49 131 217
rect 187 49 217 217
rect 273 49 303 217
rect 359 49 389 217
rect 601 65 631 233
rect 687 65 717 233
rect 773 65 803 233
rect 859 65 889 233
rect 945 65 975 233
rect 1062 65 1092 233
rect 1148 65 1178 233
rect 1234 65 1264 233
<< scpmoshvt >>
rect 146 367 176 619
rect 232 367 262 619
rect 318 367 348 619
rect 404 367 434 619
rect 490 367 520 619
rect 576 367 606 619
rect 773 367 803 619
rect 859 367 889 619
rect 945 367 975 619
rect 1062 367 1092 619
rect 1148 367 1178 619
rect 1234 367 1264 619
<< ndiff >>
rect 48 177 101 217
rect 48 143 56 177
rect 90 143 101 177
rect 48 95 101 143
rect 48 61 56 95
rect 90 61 101 95
rect 48 49 101 61
rect 131 205 187 217
rect 131 171 142 205
rect 176 171 187 205
rect 131 101 187 171
rect 131 67 142 101
rect 176 67 187 101
rect 131 49 187 67
rect 217 177 273 217
rect 217 143 228 177
rect 262 143 273 177
rect 217 91 273 143
rect 217 57 228 91
rect 262 57 273 91
rect 217 49 273 57
rect 303 205 359 217
rect 303 171 314 205
rect 348 171 359 205
rect 303 101 359 171
rect 303 67 314 101
rect 348 67 359 101
rect 303 49 359 67
rect 389 205 442 217
rect 389 171 400 205
rect 434 171 442 205
rect 389 95 442 171
rect 389 61 400 95
rect 434 61 442 95
rect 528 181 601 233
rect 528 147 540 181
rect 574 147 601 181
rect 528 107 601 147
rect 528 73 540 107
rect 574 73 601 107
rect 528 65 601 73
rect 631 225 687 233
rect 631 191 642 225
rect 676 191 687 225
rect 631 155 687 191
rect 631 121 642 155
rect 676 121 687 155
rect 631 65 687 121
rect 717 221 773 233
rect 717 187 728 221
rect 762 187 773 221
rect 717 111 773 187
rect 717 77 728 111
rect 762 77 773 111
rect 717 65 773 77
rect 803 179 859 233
rect 803 145 814 179
rect 848 145 859 179
rect 803 107 859 145
rect 803 73 814 107
rect 848 73 859 107
rect 803 65 859 73
rect 889 221 945 233
rect 889 187 900 221
rect 934 187 945 221
rect 889 111 945 187
rect 889 77 900 111
rect 934 77 945 111
rect 889 65 945 77
rect 975 130 1062 233
rect 975 96 1001 130
rect 1035 96 1062 130
rect 975 65 1062 96
rect 1092 192 1148 233
rect 1092 158 1103 192
rect 1137 158 1148 192
rect 1092 111 1148 158
rect 1092 77 1103 111
rect 1137 77 1148 111
rect 1092 65 1148 77
rect 1178 111 1234 233
rect 1178 77 1189 111
rect 1223 77 1234 111
rect 1178 65 1234 77
rect 1264 192 1317 233
rect 1264 158 1275 192
rect 1309 158 1317 192
rect 1264 111 1317 158
rect 1264 77 1275 111
rect 1309 77 1317 111
rect 1264 65 1317 77
rect 389 49 442 61
<< pdiff >>
rect 93 607 146 619
rect 93 573 101 607
rect 135 573 146 607
rect 93 530 146 573
rect 93 496 101 530
rect 135 496 146 530
rect 93 453 146 496
rect 93 419 101 453
rect 135 419 146 453
rect 93 367 146 419
rect 176 599 232 619
rect 176 565 187 599
rect 221 565 232 599
rect 176 502 232 565
rect 176 468 187 502
rect 221 468 232 502
rect 176 413 232 468
rect 176 379 187 413
rect 221 379 232 413
rect 176 367 232 379
rect 262 607 318 619
rect 262 573 273 607
rect 307 573 318 607
rect 262 530 318 573
rect 262 496 273 530
rect 307 496 318 530
rect 262 453 318 496
rect 262 419 273 453
rect 307 419 318 453
rect 262 367 318 419
rect 348 599 404 619
rect 348 565 359 599
rect 393 565 404 599
rect 348 502 404 565
rect 348 468 359 502
rect 393 468 404 502
rect 348 413 404 468
rect 348 379 359 413
rect 393 379 404 413
rect 348 367 404 379
rect 434 607 490 619
rect 434 573 445 607
rect 479 573 490 607
rect 434 507 490 573
rect 434 473 445 507
rect 479 473 490 507
rect 434 413 490 473
rect 434 379 445 413
rect 479 379 490 413
rect 434 367 490 379
rect 520 599 576 619
rect 520 565 531 599
rect 565 565 576 599
rect 520 502 576 565
rect 520 468 531 502
rect 565 468 576 502
rect 520 413 576 468
rect 520 379 531 413
rect 565 379 576 413
rect 520 367 576 379
rect 606 567 659 619
rect 606 533 617 567
rect 651 533 659 567
rect 606 367 659 533
rect 720 420 773 619
rect 720 386 728 420
rect 762 386 773 420
rect 720 367 773 386
rect 803 599 859 619
rect 803 565 814 599
rect 848 565 859 599
rect 803 508 859 565
rect 803 474 814 508
rect 848 474 859 508
rect 803 367 859 474
rect 889 599 945 619
rect 889 565 900 599
rect 934 565 945 599
rect 889 504 945 565
rect 889 470 900 504
rect 934 470 945 504
rect 889 418 945 470
rect 889 384 900 418
rect 934 384 945 418
rect 889 367 945 384
rect 975 607 1062 619
rect 975 573 1001 607
rect 1035 573 1062 607
rect 975 526 1062 573
rect 975 492 1001 526
rect 1035 492 1062 526
rect 975 367 1062 492
rect 1092 529 1148 619
rect 1092 495 1103 529
rect 1137 495 1148 529
rect 1092 367 1148 495
rect 1178 607 1234 619
rect 1178 573 1189 607
rect 1223 573 1234 607
rect 1178 367 1234 573
rect 1264 449 1317 619
rect 1264 415 1275 449
rect 1309 415 1317 449
rect 1264 367 1317 415
<< ndiffc >>
rect 56 143 90 177
rect 56 61 90 95
rect 142 171 176 205
rect 142 67 176 101
rect 228 143 262 177
rect 228 57 262 91
rect 314 171 348 205
rect 314 67 348 101
rect 400 171 434 205
rect 400 61 434 95
rect 540 147 574 181
rect 540 73 574 107
rect 642 191 676 225
rect 642 121 676 155
rect 728 187 762 221
rect 728 77 762 111
rect 814 145 848 179
rect 814 73 848 107
rect 900 187 934 221
rect 900 77 934 111
rect 1001 96 1035 130
rect 1103 158 1137 192
rect 1103 77 1137 111
rect 1189 77 1223 111
rect 1275 158 1309 192
rect 1275 77 1309 111
<< pdiffc >>
rect 101 573 135 607
rect 101 496 135 530
rect 101 419 135 453
rect 187 565 221 599
rect 187 468 221 502
rect 187 379 221 413
rect 273 573 307 607
rect 273 496 307 530
rect 273 419 307 453
rect 359 565 393 599
rect 359 468 393 502
rect 359 379 393 413
rect 445 573 479 607
rect 445 473 479 507
rect 445 379 479 413
rect 531 565 565 599
rect 531 468 565 502
rect 531 379 565 413
rect 617 533 651 567
rect 728 386 762 420
rect 814 565 848 599
rect 814 474 848 508
rect 900 565 934 599
rect 900 470 934 504
rect 900 384 934 418
rect 1001 573 1035 607
rect 1001 492 1035 526
rect 1103 495 1137 529
rect 1189 573 1223 607
rect 1275 415 1309 449
<< poly >>
rect 146 619 176 645
rect 232 619 262 645
rect 318 619 348 645
rect 404 619 434 645
rect 490 619 520 645
rect 576 619 606 645
rect 773 619 803 645
rect 859 619 889 645
rect 945 619 975 645
rect 1062 619 1092 645
rect 1148 619 1178 645
rect 1234 619 1264 645
rect 146 331 176 367
rect 232 331 262 367
rect 318 331 348 367
rect 404 331 434 367
rect 101 315 439 331
rect 101 281 117 315
rect 151 281 185 315
rect 219 281 253 315
rect 287 281 321 315
rect 355 281 389 315
rect 423 281 439 315
rect 101 265 439 281
rect 490 299 520 367
rect 576 335 606 367
rect 773 335 803 367
rect 859 335 889 367
rect 576 319 667 335
rect 576 299 617 319
rect 490 285 617 299
rect 651 299 667 319
rect 773 319 889 335
rect 651 285 717 299
rect 490 269 717 285
rect 101 217 131 265
rect 187 217 217 265
rect 273 217 303 265
rect 359 217 389 265
rect 601 233 631 269
rect 687 233 717 269
rect 773 285 789 319
rect 823 285 889 319
rect 773 269 889 285
rect 773 233 803 269
rect 859 233 889 269
rect 945 335 975 367
rect 945 319 1020 335
rect 945 285 970 319
rect 1004 285 1020 319
rect 945 269 1020 285
rect 1062 321 1092 367
rect 1148 321 1178 367
rect 1062 305 1178 321
rect 1062 271 1128 305
rect 1162 271 1178 305
rect 945 233 975 269
rect 1062 255 1178 271
rect 1062 233 1092 255
rect 1148 233 1178 255
rect 1234 325 1264 367
rect 1234 309 1319 325
rect 1234 275 1269 309
rect 1303 275 1319 309
rect 1234 259 1319 275
rect 1234 233 1264 259
rect 101 23 131 49
rect 187 23 217 49
rect 273 23 303 49
rect 359 23 389 49
rect 601 39 631 65
rect 687 39 717 65
rect 773 39 803 65
rect 859 39 889 65
rect 945 39 975 65
rect 1062 39 1092 65
rect 1148 39 1178 65
rect 1234 39 1264 65
<< polycont >>
rect 117 281 151 315
rect 185 281 219 315
rect 253 281 287 315
rect 321 281 355 315
rect 389 281 423 315
rect 617 285 651 319
rect 789 285 823 319
rect 970 285 1004 319
rect 1128 271 1162 305
rect 1269 275 1303 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 85 607 151 649
rect 85 573 101 607
rect 135 573 151 607
rect 85 530 151 573
rect 85 496 101 530
rect 135 496 151 530
rect 85 453 151 496
rect 85 419 101 453
rect 135 419 151 453
rect 185 599 223 615
rect 185 565 187 599
rect 221 565 223 599
rect 185 502 223 565
rect 185 468 187 502
rect 221 468 223 502
rect 185 413 223 468
rect 257 607 323 649
rect 257 573 273 607
rect 307 573 323 607
rect 257 530 323 573
rect 257 496 273 530
rect 307 496 323 530
rect 257 453 323 496
rect 257 419 273 453
rect 307 419 323 453
rect 359 599 395 615
rect 393 565 395 599
rect 359 502 395 565
rect 393 468 395 502
rect 185 385 187 413
rect 17 379 187 385
rect 221 385 223 413
rect 359 413 395 468
rect 221 379 359 385
rect 393 379 395 413
rect 17 351 395 379
rect 429 607 495 649
rect 429 573 445 607
rect 479 573 495 607
rect 429 507 495 573
rect 429 473 445 507
rect 479 473 495 507
rect 429 413 495 473
rect 429 379 445 413
rect 479 379 495 413
rect 429 363 495 379
rect 529 599 565 615
rect 529 565 531 599
rect 529 502 565 565
rect 601 567 667 649
rect 601 533 617 567
rect 651 533 667 567
rect 601 526 667 533
rect 798 599 852 615
rect 798 565 814 599
rect 848 565 852 599
rect 529 468 531 502
rect 798 508 852 565
rect 798 492 814 508
rect 565 474 814 492
rect 848 474 852 508
rect 565 468 852 474
rect 529 458 852 468
rect 886 599 950 615
rect 886 565 900 599
rect 934 565 950 599
rect 886 504 950 565
rect 886 470 900 504
rect 934 470 950 504
rect 985 607 1239 615
rect 985 573 1001 607
rect 1035 573 1189 607
rect 1223 573 1239 607
rect 985 567 1239 573
rect 985 526 1051 567
rect 1273 533 1325 649
rect 985 492 1001 526
rect 1035 492 1051 526
rect 985 487 1051 492
rect 1085 529 1325 533
rect 1085 495 1103 529
rect 1137 495 1325 529
rect 1085 487 1325 495
rect 529 413 567 458
rect 886 453 950 470
rect 886 449 1325 453
rect 886 424 1275 449
rect 529 379 531 413
rect 565 379 567 413
rect 17 245 67 351
rect 529 315 567 379
rect 101 281 117 315
rect 151 281 185 315
rect 219 281 253 315
rect 287 281 321 315
rect 355 281 389 315
rect 423 281 567 315
rect 601 319 667 424
rect 712 420 1275 424
rect 712 386 728 420
rect 762 418 1275 420
rect 762 386 900 418
rect 712 384 900 386
rect 934 415 1275 418
rect 1309 415 1325 449
rect 934 409 1325 415
rect 934 384 950 409
rect 984 350 1319 375
rect 601 285 617 319
rect 651 285 667 319
rect 703 319 936 350
rect 703 285 789 319
rect 823 285 936 319
rect 970 341 1319 350
rect 970 319 1041 341
rect 1004 285 1041 319
rect 1253 309 1319 341
rect 527 249 567 281
rect 970 269 1041 285
rect 1075 305 1219 307
rect 1075 271 1128 305
rect 1162 271 1219 305
rect 17 211 350 245
rect 527 225 692 249
rect 140 205 178 211
rect 40 143 56 177
rect 90 143 106 177
rect 40 95 106 143
rect 40 61 56 95
rect 90 61 106 95
rect 40 17 106 61
rect 140 171 142 205
rect 176 171 178 205
rect 312 205 350 211
rect 140 101 178 171
rect 140 67 142 101
rect 176 67 178 101
rect 140 51 178 67
rect 212 143 228 177
rect 262 143 278 177
rect 212 91 278 143
rect 212 57 228 91
rect 262 57 278 91
rect 212 17 278 57
rect 312 171 314 205
rect 348 171 350 205
rect 312 101 350 171
rect 312 67 314 101
rect 348 67 350 101
rect 312 51 350 67
rect 384 205 450 221
rect 527 215 642 225
rect 384 171 400 205
rect 434 171 450 205
rect 626 191 642 215
rect 676 191 692 225
rect 384 95 450 171
rect 384 61 400 95
rect 434 61 450 95
rect 384 17 450 61
rect 524 147 540 181
rect 574 147 590 181
rect 524 107 590 147
rect 626 155 692 191
rect 626 121 642 155
rect 676 121 692 155
rect 726 221 942 249
rect 1075 242 1219 271
rect 1253 275 1269 309
rect 1303 275 1319 309
rect 1253 259 1319 275
rect 726 187 728 221
rect 762 215 900 221
rect 762 187 764 215
rect 524 73 540 107
rect 574 87 590 107
rect 726 111 764 187
rect 898 187 900 215
rect 934 208 942 221
rect 934 192 1325 208
rect 934 187 1103 192
rect 726 87 728 111
rect 574 77 728 87
rect 762 77 764 111
rect 574 73 764 77
rect 524 51 764 73
rect 798 145 814 179
rect 848 145 864 179
rect 798 107 864 145
rect 798 73 814 107
rect 848 73 864 107
rect 798 17 864 73
rect 898 174 1103 187
rect 898 111 950 174
rect 1087 158 1103 174
rect 1137 174 1275 192
rect 1137 158 1139 174
rect 898 77 900 111
rect 934 77 950 111
rect 898 61 950 77
rect 985 130 1051 140
rect 985 96 1001 130
rect 1035 96 1051 130
rect 985 17 1051 96
rect 1087 111 1139 158
rect 1273 158 1275 174
rect 1309 158 1325 192
rect 1087 77 1103 111
rect 1137 77 1139 111
rect 1087 61 1139 77
rect 1173 111 1239 140
rect 1173 77 1189 111
rect 1223 77 1239 111
rect 1173 17 1239 77
rect 1273 111 1325 158
rect 1273 77 1275 111
rect 1309 77 1325 111
rect 1273 61 1325 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o31a_4
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1192006
string GDS_START 1180654
<< end >>
