magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 2 49 830 241
rect 0 0 864 49
<< scnmos >>
rect 85 47 115 215
rect 171 47 201 215
rect 325 47 355 215
rect 397 47 427 215
rect 505 47 535 215
rect 613 47 643 215
rect 721 47 751 215
<< scpmoshvt >>
rect 100 367 130 619
rect 186 367 216 619
rect 311 367 341 619
rect 397 367 427 619
rect 541 367 571 619
rect 627 367 657 619
rect 721 367 751 619
<< ndiff >>
rect 28 203 85 215
rect 28 169 40 203
rect 74 169 85 203
rect 28 93 85 169
rect 28 59 40 93
rect 74 59 85 93
rect 28 47 85 59
rect 115 203 171 215
rect 115 169 126 203
rect 160 169 171 203
rect 115 101 171 169
rect 115 67 126 101
rect 160 67 171 101
rect 115 47 171 67
rect 201 127 325 215
rect 201 93 212 127
rect 246 93 280 127
rect 314 93 325 127
rect 201 47 325 93
rect 355 47 397 215
rect 427 47 505 215
rect 535 203 613 215
rect 535 169 557 203
rect 591 169 613 203
rect 535 93 613 169
rect 535 59 557 93
rect 591 59 613 93
rect 535 47 613 59
rect 643 127 721 215
rect 643 93 666 127
rect 700 93 721 127
rect 643 47 721 93
rect 751 203 804 215
rect 751 169 762 203
rect 796 169 804 203
rect 751 101 804 169
rect 751 67 762 101
rect 796 67 804 101
rect 751 47 804 67
<< pdiff >>
rect 47 607 100 619
rect 47 573 55 607
rect 89 573 100 607
rect 47 513 100 573
rect 47 479 55 513
rect 89 479 100 513
rect 47 413 100 479
rect 47 379 55 413
rect 89 379 100 413
rect 47 367 100 379
rect 130 599 186 619
rect 130 565 141 599
rect 175 565 186 599
rect 130 511 186 565
rect 130 477 141 511
rect 175 477 186 511
rect 130 420 186 477
rect 130 386 141 420
rect 175 386 186 420
rect 130 367 186 386
rect 216 607 311 619
rect 216 573 246 607
rect 280 573 311 607
rect 216 524 311 573
rect 216 490 246 524
rect 280 490 311 524
rect 216 443 311 490
rect 216 409 246 443
rect 280 409 311 443
rect 216 367 311 409
rect 341 607 397 619
rect 341 573 352 607
rect 386 573 397 607
rect 341 523 397 573
rect 341 489 352 523
rect 386 489 397 523
rect 341 443 397 489
rect 341 409 352 443
rect 386 409 397 443
rect 341 367 397 409
rect 427 607 541 619
rect 427 573 468 607
rect 502 573 541 607
rect 427 516 541 573
rect 427 482 468 516
rect 502 482 541 516
rect 427 367 541 482
rect 571 607 627 619
rect 571 573 582 607
rect 616 573 627 607
rect 571 523 627 573
rect 571 489 582 523
rect 616 489 627 523
rect 571 443 627 489
rect 571 409 582 443
rect 616 409 627 443
rect 571 367 627 409
rect 657 367 721 619
rect 751 607 804 619
rect 751 573 762 607
rect 796 573 804 607
rect 751 509 804 573
rect 751 475 762 509
rect 796 475 804 509
rect 751 413 804 475
rect 751 379 762 413
rect 796 379 804 413
rect 751 367 804 379
<< ndiffc >>
rect 40 169 74 203
rect 40 59 74 93
rect 126 169 160 203
rect 126 67 160 101
rect 212 93 246 127
rect 280 93 314 127
rect 557 169 591 203
rect 557 59 591 93
rect 666 93 700 127
rect 762 169 796 203
rect 762 67 796 101
<< pdiffc >>
rect 55 573 89 607
rect 55 479 89 513
rect 55 379 89 413
rect 141 565 175 599
rect 141 477 175 511
rect 141 386 175 420
rect 246 573 280 607
rect 246 490 280 524
rect 246 409 280 443
rect 352 573 386 607
rect 352 489 386 523
rect 352 409 386 443
rect 468 573 502 607
rect 468 482 502 516
rect 582 573 616 607
rect 582 489 616 523
rect 582 409 616 443
rect 762 573 796 607
rect 762 475 796 509
rect 762 379 796 413
<< poly >>
rect 100 619 130 645
rect 186 619 216 645
rect 311 619 341 645
rect 397 619 427 645
rect 541 619 571 645
rect 627 619 657 645
rect 721 619 751 645
rect 100 267 130 367
rect 186 303 216 367
rect 311 303 341 367
rect 397 305 427 367
rect 541 305 571 367
rect 172 287 247 303
rect 172 267 197 287
rect 85 253 197 267
rect 231 253 247 287
rect 85 237 247 253
rect 289 287 355 303
rect 289 253 305 287
rect 339 253 355 287
rect 289 237 355 253
rect 85 215 115 237
rect 171 215 201 237
rect 325 215 355 237
rect 397 289 463 305
rect 397 255 413 289
rect 447 255 463 289
rect 397 239 463 255
rect 505 289 571 305
rect 627 303 657 367
rect 721 305 751 367
rect 505 255 521 289
rect 555 255 571 289
rect 505 239 571 255
rect 613 287 679 303
rect 613 253 629 287
rect 663 253 679 287
rect 397 215 427 239
rect 505 215 535 239
rect 613 237 679 253
rect 721 289 823 305
rect 721 255 773 289
rect 807 255 823 289
rect 721 239 823 255
rect 613 215 643 237
rect 721 215 751 239
rect 85 21 115 47
rect 171 21 201 47
rect 325 21 355 47
rect 397 21 427 47
rect 505 21 535 47
rect 613 21 643 47
rect 721 21 751 47
<< polycont >>
rect 197 253 231 287
rect 305 253 339 287
rect 413 255 447 289
rect 521 255 555 289
rect 629 253 663 287
rect 773 255 807 289
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 39 607 93 649
rect 39 573 55 607
rect 89 573 93 607
rect 39 513 93 573
rect 39 479 55 513
rect 89 479 93 513
rect 39 413 93 479
rect 39 379 55 413
rect 89 379 93 413
rect 39 363 93 379
rect 127 599 181 615
rect 127 565 141 599
rect 175 565 181 599
rect 127 511 181 565
rect 127 477 141 511
rect 175 477 181 511
rect 127 420 181 477
rect 127 386 141 420
rect 175 386 181 420
rect 230 607 296 649
rect 230 573 246 607
rect 280 573 296 607
rect 230 524 296 573
rect 230 490 246 524
rect 280 490 296 524
rect 230 443 296 490
rect 230 409 246 443
rect 280 409 296 443
rect 336 607 402 613
rect 336 573 352 607
rect 386 573 402 607
rect 336 523 402 573
rect 336 489 352 523
rect 386 489 402 523
rect 336 443 402 489
rect 452 607 518 649
rect 452 573 468 607
rect 502 573 518 607
rect 452 516 518 573
rect 452 482 468 516
rect 502 482 518 516
rect 452 477 518 482
rect 566 607 632 613
rect 566 573 582 607
rect 616 573 632 607
rect 566 523 632 573
rect 566 489 582 523
rect 616 489 632 523
rect 566 443 632 489
rect 336 409 352 443
rect 386 409 582 443
rect 616 409 632 443
rect 746 607 812 615
rect 746 573 762 607
rect 796 573 812 607
rect 746 509 812 573
rect 746 475 762 509
rect 796 475 812 509
rect 746 413 812 475
rect 127 370 181 386
rect 746 379 762 413
rect 796 379 812 413
rect 746 375 812 379
rect 127 307 162 370
rect 24 203 82 219
rect 24 169 40 203
rect 74 169 82 203
rect 24 93 82 169
rect 24 59 40 93
rect 74 59 82 93
rect 24 17 82 59
rect 116 203 162 307
rect 215 339 812 375
rect 215 303 249 339
rect 116 169 126 203
rect 160 169 162 203
rect 197 287 249 303
rect 231 253 249 287
rect 197 203 249 253
rect 289 287 365 305
rect 289 253 305 287
rect 339 253 365 287
rect 289 237 365 253
rect 399 289 467 305
rect 399 255 413 289
rect 447 255 467 289
rect 399 237 467 255
rect 501 289 567 305
rect 501 255 521 289
rect 555 255 567 289
rect 501 237 567 255
rect 601 287 739 305
rect 601 253 629 287
rect 663 253 739 287
rect 601 237 739 253
rect 773 289 847 305
rect 807 255 847 289
rect 773 237 847 255
rect 197 169 557 203
rect 591 169 762 203
rect 796 169 812 203
rect 116 101 162 169
rect 116 67 126 101
rect 160 67 162 101
rect 116 51 162 67
rect 196 127 330 135
rect 196 93 212 127
rect 246 93 280 127
rect 314 93 330 127
rect 196 17 330 93
rect 541 93 607 169
rect 541 59 557 93
rect 591 59 607 93
rect 541 51 607 59
rect 650 127 716 135
rect 650 93 666 127
rect 700 93 716 127
rect 650 17 716 93
rect 750 101 812 169
rect 750 67 762 101
rect 796 67 812 101
rect 750 51 812 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a311o_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3891356
string GDS_START 3883128
<< end >>
