magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 135 49 1343 241
rect 0 0 1344 49
<< scnmos >>
rect 214 47 244 215
rect 300 47 330 215
rect 386 47 416 215
rect 475 47 505 215
rect 561 47 591 215
rect 650 47 680 215
rect 736 47 766 215
rect 822 47 852 215
rect 976 47 1006 215
rect 1062 47 1092 215
rect 1148 47 1178 215
rect 1234 47 1264 215
<< scpmoshvt >>
rect 103 367 133 619
rect 189 367 219 619
rect 275 367 305 619
rect 361 367 391 619
rect 580 367 610 619
rect 666 367 696 619
rect 752 367 782 619
rect 846 367 876 619
rect 954 367 984 619
rect 1062 367 1092 619
rect 1148 367 1178 619
rect 1234 367 1264 619
<< ndiff >>
rect 161 176 214 215
rect 161 142 169 176
rect 203 142 214 176
rect 161 93 214 142
rect 161 59 169 93
rect 203 59 214 93
rect 161 47 214 59
rect 244 203 300 215
rect 244 169 255 203
rect 289 169 300 203
rect 244 101 300 169
rect 244 67 255 101
rect 289 67 300 101
rect 244 47 300 67
rect 330 174 386 215
rect 330 140 341 174
rect 375 140 386 174
rect 330 89 386 140
rect 330 55 341 89
rect 375 55 386 89
rect 330 47 386 55
rect 416 203 475 215
rect 416 169 427 203
rect 461 169 475 203
rect 416 101 475 169
rect 416 67 427 101
rect 461 67 475 101
rect 416 47 475 67
rect 505 160 561 215
rect 505 126 516 160
rect 550 126 561 160
rect 505 89 561 126
rect 505 55 516 89
rect 550 55 561 89
rect 505 47 561 55
rect 591 203 650 215
rect 591 169 602 203
rect 636 169 650 203
rect 591 101 650 169
rect 591 67 602 101
rect 636 67 650 101
rect 591 47 650 67
rect 680 123 736 215
rect 680 89 691 123
rect 725 89 736 123
rect 680 47 736 89
rect 766 203 822 215
rect 766 169 777 203
rect 811 169 822 203
rect 766 101 822 169
rect 766 67 777 101
rect 811 67 822 101
rect 766 47 822 67
rect 852 161 976 215
rect 852 59 863 161
rect 965 59 976 161
rect 852 47 976 59
rect 1006 175 1062 215
rect 1006 141 1017 175
rect 1051 141 1062 175
rect 1006 93 1062 141
rect 1006 59 1017 93
rect 1051 59 1062 93
rect 1006 47 1062 59
rect 1092 169 1148 215
rect 1092 135 1103 169
rect 1137 135 1148 169
rect 1092 47 1148 135
rect 1178 203 1234 215
rect 1178 169 1189 203
rect 1223 169 1234 203
rect 1178 92 1234 169
rect 1178 58 1189 92
rect 1223 58 1234 92
rect 1178 47 1234 58
rect 1264 203 1317 215
rect 1264 169 1275 203
rect 1309 169 1317 203
rect 1264 93 1317 169
rect 1264 59 1275 93
rect 1309 59 1317 93
rect 1264 47 1317 59
<< pdiff >>
rect 50 607 103 619
rect 50 573 58 607
rect 92 573 103 607
rect 50 531 103 573
rect 50 497 58 531
rect 92 497 103 531
rect 50 453 103 497
rect 50 419 58 453
rect 92 419 103 453
rect 50 367 103 419
rect 133 599 189 619
rect 133 565 144 599
rect 178 565 189 599
rect 133 510 189 565
rect 133 476 144 510
rect 178 476 189 510
rect 133 413 189 476
rect 133 379 144 413
rect 178 379 189 413
rect 133 367 189 379
rect 219 607 275 619
rect 219 573 230 607
rect 264 573 275 607
rect 219 531 275 573
rect 219 497 230 531
rect 264 497 275 531
rect 219 455 275 497
rect 219 421 230 455
rect 264 421 275 455
rect 219 367 275 421
rect 305 599 361 619
rect 305 565 316 599
rect 350 565 361 599
rect 305 510 361 565
rect 305 476 316 510
rect 350 476 361 510
rect 305 413 361 476
rect 305 379 316 413
rect 350 379 361 413
rect 305 367 361 379
rect 391 607 444 619
rect 391 573 402 607
rect 436 573 444 607
rect 391 510 444 573
rect 391 476 402 510
rect 436 476 444 510
rect 391 413 444 476
rect 391 379 402 413
rect 436 379 444 413
rect 391 367 444 379
rect 527 599 580 619
rect 527 565 535 599
rect 569 565 580 599
rect 527 525 580 565
rect 527 491 535 525
rect 569 491 580 525
rect 527 367 580 491
rect 610 595 666 619
rect 610 561 621 595
rect 655 561 666 595
rect 610 367 666 561
rect 696 447 752 619
rect 696 413 707 447
rect 741 413 752 447
rect 696 367 752 413
rect 782 595 846 619
rect 782 561 793 595
rect 827 561 846 595
rect 782 367 846 561
rect 876 599 954 619
rect 876 565 896 599
rect 930 565 954 599
rect 876 519 954 565
rect 876 485 896 519
rect 930 485 954 519
rect 876 441 954 485
rect 876 407 896 441
rect 930 407 954 441
rect 876 367 954 407
rect 984 571 1062 619
rect 984 537 995 571
rect 1029 537 1062 571
rect 984 367 1062 537
rect 1092 599 1148 619
rect 1092 565 1103 599
rect 1137 565 1148 599
rect 1092 510 1148 565
rect 1092 476 1103 510
rect 1137 476 1148 510
rect 1092 367 1148 476
rect 1178 574 1234 619
rect 1178 540 1189 574
rect 1223 540 1234 574
rect 1178 367 1234 540
rect 1264 599 1317 619
rect 1264 565 1275 599
rect 1309 565 1317 599
rect 1264 502 1317 565
rect 1264 468 1275 502
rect 1309 468 1317 502
rect 1264 413 1317 468
rect 1264 379 1275 413
rect 1309 379 1317 413
rect 1264 367 1317 379
<< ndiffc >>
rect 169 142 203 176
rect 169 59 203 93
rect 255 169 289 203
rect 255 67 289 101
rect 341 140 375 174
rect 341 55 375 89
rect 427 169 461 203
rect 427 67 461 101
rect 516 126 550 160
rect 516 55 550 89
rect 602 169 636 203
rect 602 67 636 101
rect 691 89 725 123
rect 777 169 811 203
rect 777 67 811 101
rect 863 59 965 161
rect 1017 141 1051 175
rect 1017 59 1051 93
rect 1103 135 1137 169
rect 1189 169 1223 203
rect 1189 58 1223 92
rect 1275 169 1309 203
rect 1275 59 1309 93
<< pdiffc >>
rect 58 573 92 607
rect 58 497 92 531
rect 58 419 92 453
rect 144 565 178 599
rect 144 476 178 510
rect 144 379 178 413
rect 230 573 264 607
rect 230 497 264 531
rect 230 421 264 455
rect 316 565 350 599
rect 316 476 350 510
rect 316 379 350 413
rect 402 573 436 607
rect 402 476 436 510
rect 402 379 436 413
rect 535 565 569 599
rect 535 491 569 525
rect 621 561 655 595
rect 707 413 741 447
rect 793 561 827 595
rect 896 565 930 599
rect 896 485 930 519
rect 896 407 930 441
rect 995 537 1029 571
rect 1103 565 1137 599
rect 1103 476 1137 510
rect 1189 540 1223 574
rect 1275 565 1309 599
rect 1275 468 1309 502
rect 1275 379 1309 413
<< poly >>
rect 103 619 133 645
rect 189 619 219 645
rect 275 619 305 645
rect 361 619 391 645
rect 580 619 610 645
rect 666 619 696 645
rect 752 619 782 645
rect 846 619 876 645
rect 954 619 984 645
rect 1062 619 1092 645
rect 1148 619 1178 645
rect 1234 619 1264 645
rect 103 329 133 367
rect 189 329 219 367
rect 275 329 305 367
rect 361 329 391 367
rect 580 335 610 367
rect 103 313 505 329
rect 103 279 119 313
rect 153 279 187 313
rect 221 279 255 313
rect 289 279 323 313
rect 357 279 391 313
rect 425 279 505 313
rect 103 263 505 279
rect 547 319 613 335
rect 547 285 563 319
rect 597 285 613 319
rect 666 303 696 367
rect 752 303 782 367
rect 846 333 876 367
rect 954 345 984 367
rect 547 269 613 285
rect 655 291 782 303
rect 824 317 890 333
rect 655 288 780 291
rect 655 287 779 288
rect 214 215 244 263
rect 300 215 330 263
rect 386 215 416 263
rect 475 215 505 263
rect 561 215 591 269
rect 655 253 707 287
rect 741 281 779 287
rect 824 283 840 317
rect 874 283 890 317
rect 741 276 773 281
rect 824 278 890 283
rect 741 253 766 276
rect 655 251 766 253
rect 652 248 766 251
rect 650 230 766 248
rect 650 215 680 230
rect 736 215 766 230
rect 822 267 890 278
rect 954 319 1020 345
rect 954 285 970 319
rect 1004 285 1020 319
rect 954 269 1020 285
rect 1062 335 1092 367
rect 1148 335 1178 367
rect 1062 319 1178 335
rect 1062 285 1078 319
rect 1112 285 1178 319
rect 1062 269 1178 285
rect 822 215 852 267
rect 976 215 1006 269
rect 1062 215 1092 269
rect 1148 215 1178 269
rect 1234 335 1264 367
rect 1234 319 1300 335
rect 1234 285 1250 319
rect 1284 285 1300 319
rect 1234 269 1300 285
rect 1234 215 1264 269
rect 214 21 244 47
rect 300 21 330 47
rect 386 21 416 47
rect 475 21 505 47
rect 561 21 591 47
rect 650 21 680 47
rect 736 21 766 47
rect 822 21 852 47
rect 976 21 1006 47
rect 1062 21 1092 47
rect 1148 21 1178 47
rect 1234 21 1264 47
<< polycont >>
rect 119 279 153 313
rect 187 279 221 313
rect 255 279 289 313
rect 323 279 357 313
rect 391 279 425 313
rect 563 285 597 319
rect 707 253 741 287
rect 840 283 874 317
rect 970 285 1004 319
rect 1078 285 1112 319
rect 1250 285 1284 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 42 607 108 649
rect 42 573 58 607
rect 92 573 108 607
rect 42 531 108 573
rect 42 497 58 531
rect 92 497 108 531
rect 42 453 108 497
rect 42 419 58 453
rect 92 419 108 453
rect 142 599 180 615
rect 142 565 144 599
rect 178 565 180 599
rect 142 510 180 565
rect 142 476 144 510
rect 178 476 180 510
rect 142 413 180 476
rect 214 607 280 649
rect 214 573 230 607
rect 264 573 280 607
rect 214 531 280 573
rect 214 497 230 531
rect 264 497 280 531
rect 214 455 280 497
rect 214 421 230 455
rect 264 421 280 455
rect 314 599 352 615
rect 314 565 316 599
rect 350 565 352 599
rect 314 510 352 565
rect 314 476 316 510
rect 350 476 352 510
rect 142 385 144 413
rect 18 379 144 385
rect 178 385 180 413
rect 314 413 352 476
rect 314 385 316 413
rect 178 379 316 385
rect 350 379 352 413
rect 18 351 352 379
rect 386 607 452 649
rect 386 573 402 607
rect 436 573 452 607
rect 386 510 452 573
rect 386 476 402 510
rect 436 476 452 510
rect 386 413 452 476
rect 519 599 571 615
rect 519 565 535 599
rect 569 565 571 599
rect 519 525 571 565
rect 605 595 843 611
rect 605 561 621 595
rect 655 561 793 595
rect 827 561 843 595
rect 605 553 843 561
rect 877 599 945 615
rect 877 565 896 599
rect 930 565 945 599
rect 519 491 535 525
rect 569 519 571 525
rect 877 519 945 565
rect 979 571 1045 649
rect 979 537 995 571
rect 1029 537 1045 571
rect 979 526 1045 537
rect 1087 599 1139 615
rect 1087 565 1103 599
rect 1137 565 1139 599
rect 569 491 896 519
rect 519 485 896 491
rect 930 492 945 519
rect 1087 510 1139 565
rect 1173 574 1239 649
rect 1173 540 1189 574
rect 1223 540 1239 574
rect 1173 526 1239 540
rect 1273 599 1325 615
rect 1273 565 1275 599
rect 1309 565 1325 599
rect 1087 492 1103 510
rect 930 485 1103 492
rect 519 475 585 485
rect 871 476 1103 485
rect 1137 492 1139 510
rect 1273 502 1325 565
rect 1273 492 1275 502
rect 1137 476 1275 492
rect 871 468 1275 476
rect 1309 468 1325 502
rect 871 458 1325 468
rect 691 447 757 451
rect 691 441 707 447
rect 386 379 402 413
rect 436 379 452 413
rect 386 363 452 379
rect 495 413 707 441
rect 741 413 757 447
rect 495 407 757 413
rect 871 441 946 458
rect 871 407 896 441
rect 930 407 946 441
rect 18 245 69 351
rect 495 317 529 407
rect 980 390 1225 424
rect 103 313 529 317
rect 103 279 119 313
rect 153 279 187 313
rect 221 279 255 313
rect 289 279 323 313
rect 357 279 391 313
rect 425 279 529 313
rect 18 211 461 245
rect 18 78 81 211
rect 253 209 461 211
rect 253 203 291 209
rect 153 176 219 177
rect 153 142 169 176
rect 203 142 219 176
rect 153 93 219 142
rect 153 59 169 93
rect 203 59 219 93
rect 153 17 219 59
rect 253 169 255 203
rect 289 169 291 203
rect 425 203 461 209
rect 253 101 291 169
rect 253 67 255 101
rect 289 67 291 101
rect 253 51 291 67
rect 325 174 391 175
rect 325 140 341 174
rect 375 140 391 174
rect 325 89 391 140
rect 325 55 341 89
rect 375 55 391 89
rect 325 17 391 55
rect 425 169 427 203
rect 495 231 529 279
rect 563 339 890 373
rect 980 364 1020 390
rect 563 319 641 339
rect 597 285 641 319
rect 824 317 890 339
rect 563 269 641 285
rect 675 287 742 303
rect 675 253 707 287
rect 741 253 742 287
rect 824 283 840 317
rect 874 283 890 317
rect 954 319 1020 364
rect 954 285 970 319
rect 1004 285 1020 319
rect 1062 319 1128 356
rect 1062 285 1078 319
rect 1112 285 1128 319
rect 1183 329 1225 390
rect 1259 413 1325 458
rect 1259 379 1275 413
rect 1309 379 1325 413
rect 1259 363 1325 379
rect 1183 319 1300 329
rect 1183 285 1250 319
rect 1284 285 1300 319
rect 1183 269 1300 285
rect 675 237 742 253
rect 495 203 641 231
rect 777 213 1139 247
rect 777 203 822 213
rect 495 197 602 203
rect 425 101 461 169
rect 600 169 602 197
rect 636 169 777 203
rect 811 169 822 203
rect 425 67 427 101
rect 425 51 461 67
rect 500 160 566 161
rect 500 126 516 160
rect 550 126 566 160
rect 500 89 566 126
rect 500 55 516 89
rect 550 55 566 89
rect 500 17 566 55
rect 600 101 641 169
rect 600 67 602 101
rect 636 67 641 101
rect 600 51 641 67
rect 675 123 741 135
rect 675 89 691 123
rect 725 89 741 123
rect 675 17 741 89
rect 775 101 822 169
rect 775 67 777 101
rect 811 67 822 101
rect 775 51 822 67
rect 856 161 967 177
rect 856 59 863 161
rect 965 59 967 161
rect 856 17 967 59
rect 1001 175 1067 179
rect 1001 141 1017 175
rect 1051 141 1067 175
rect 1001 93 1067 141
rect 1101 169 1139 213
rect 1101 135 1103 169
rect 1137 135 1139 169
rect 1101 119 1139 135
rect 1173 203 1239 219
rect 1173 169 1189 203
rect 1223 169 1239 203
rect 1001 59 1017 93
rect 1051 85 1067 93
rect 1173 92 1239 169
rect 1173 85 1189 92
rect 1051 59 1189 85
rect 1001 58 1189 59
rect 1223 58 1239 92
rect 1001 51 1239 58
rect 1273 203 1325 219
rect 1273 169 1275 203
rect 1309 169 1325 203
rect 1273 93 1325 169
rect 1273 59 1275 93
rect 1309 59 1325 93
rect 1273 17 1325 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a211o_4
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1087 390 1121 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1183 390 1217 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1947050
string GDS_START 1935408
<< end >>
