magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2310 1852
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 35 67 997 203
rect 35 21 859 67
rect 35 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 132 47 162 177
rect 247 47 277 177
rect 333 47 363 177
rect 448 47 478 177
rect 544 47 574 177
rect 640 47 670 177
rect 746 47 776 177
rect 858 93 888 177
<< scpmoshvt >>
rect 124 297 160 497
rect 239 297 275 497
rect 339 297 375 497
rect 450 297 486 497
rect 548 297 584 497
rect 642 297 678 497
rect 738 297 774 497
rect 850 345 886 429
<< ndiff >>
rect 61 161 132 177
rect 61 127 77 161
rect 111 127 132 161
rect 61 93 132 127
rect 61 59 77 93
rect 111 59 132 93
rect 61 47 132 59
rect 162 47 247 177
rect 277 47 333 177
rect 363 89 448 177
rect 363 55 402 89
rect 436 55 448 89
rect 363 47 448 55
rect 478 153 544 177
rect 478 119 499 153
rect 533 119 544 153
rect 478 47 544 119
rect 574 89 640 177
rect 574 55 589 89
rect 623 55 640 89
rect 574 47 640 55
rect 670 169 746 177
rect 670 135 691 169
rect 725 135 746 169
rect 670 101 746 135
rect 670 67 691 101
rect 725 67 746 101
rect 670 47 746 67
rect 776 93 858 177
rect 888 135 971 177
rect 888 101 925 135
rect 959 101 971 135
rect 888 93 971 101
rect 776 89 833 93
rect 776 55 787 89
rect 821 55 833 89
rect 776 47 833 55
<< pdiff >>
rect 56 417 124 497
rect 56 383 68 417
rect 102 383 124 417
rect 56 349 124 383
rect 56 315 68 349
rect 102 315 124 349
rect 56 297 124 315
rect 160 489 239 497
rect 160 455 186 489
rect 220 455 239 489
rect 160 297 239 455
rect 275 339 339 497
rect 275 305 292 339
rect 326 305 339 339
rect 275 297 339 305
rect 375 489 450 497
rect 375 455 395 489
rect 429 455 450 489
rect 375 297 450 455
rect 486 341 548 497
rect 486 307 501 341
rect 535 307 548 341
rect 486 297 548 307
rect 584 489 642 497
rect 584 455 596 489
rect 630 455 642 489
rect 584 297 642 455
rect 678 341 738 497
rect 678 307 691 341
rect 725 307 738 341
rect 678 297 738 307
rect 774 489 833 497
rect 774 455 787 489
rect 821 455 833 489
rect 774 429 833 455
rect 774 345 850 429
rect 886 421 945 429
rect 886 387 899 421
rect 933 387 945 421
rect 886 345 945 387
rect 774 297 833 345
<< ndiffc >>
rect 77 127 111 161
rect 77 59 111 93
rect 402 55 436 89
rect 499 119 533 153
rect 589 55 623 89
rect 691 135 725 169
rect 691 67 725 101
rect 925 101 959 135
rect 787 55 821 89
<< pdiffc >>
rect 68 383 102 417
rect 68 315 102 349
rect 186 455 220 489
rect 292 305 326 339
rect 395 455 429 489
rect 501 307 535 341
rect 596 455 630 489
rect 691 307 725 341
rect 787 455 821 489
rect 899 387 933 421
<< poly >>
rect 124 497 160 523
rect 239 497 275 523
rect 339 497 375 523
rect 450 497 486 523
rect 548 497 584 523
rect 642 497 678 523
rect 738 497 774 523
rect 848 455 888 523
rect 850 429 886 455
rect 850 330 886 345
rect 124 282 160 297
rect 239 282 275 297
rect 339 282 375 297
rect 450 282 486 297
rect 548 282 584 297
rect 642 282 678 297
rect 738 282 774 297
rect 122 265 162 282
rect 237 265 277 282
rect 337 265 377 282
rect 448 265 488 282
rect 546 265 586 282
rect 640 265 680 282
rect 736 265 776 282
rect 848 265 888 330
rect 98 249 162 265
rect 98 215 108 249
rect 142 215 162 249
rect 98 199 162 215
rect 204 249 277 265
rect 204 215 214 249
rect 248 215 277 249
rect 204 199 277 215
rect 319 249 383 265
rect 319 215 329 249
rect 363 215 383 249
rect 319 199 383 215
rect 448 249 776 265
rect 448 215 464 249
rect 498 215 542 249
rect 576 215 620 249
rect 654 215 776 249
rect 448 199 776 215
rect 823 249 888 265
rect 823 215 833 249
rect 867 215 888 249
rect 823 199 888 215
rect 132 177 162 199
rect 247 177 277 199
rect 333 177 363 199
rect 448 177 478 199
rect 544 177 574 199
rect 640 177 670 199
rect 746 177 776 199
rect 858 177 888 199
rect 132 21 162 47
rect 247 21 277 47
rect 333 21 363 47
rect 448 21 478 47
rect 544 21 574 47
rect 640 21 670 47
rect 746 21 776 47
rect 858 27 888 93
<< polycont >>
rect 108 215 142 249
rect 214 215 248 249
rect 329 215 363 249
rect 464 215 498 249
rect 542 215 576 249
rect 620 215 654 249
rect 833 215 867 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 146 489 246 527
rect 146 455 186 489
rect 220 455 246 489
rect 379 489 445 527
rect 379 455 395 489
rect 429 455 445 489
rect 569 489 646 527
rect 569 455 596 489
rect 630 455 646 489
rect 761 489 837 527
rect 761 455 787 489
rect 821 455 837 489
rect 30 417 102 433
rect 30 383 68 417
rect 30 349 102 383
rect 30 315 68 349
rect 30 299 102 315
rect 136 387 899 421
rect 933 387 981 421
rect 136 375 981 387
rect 30 161 74 299
rect 136 265 173 375
rect 266 305 292 339
rect 326 305 441 339
rect 475 307 501 341
rect 535 307 691 341
rect 725 307 799 341
rect 407 271 441 305
rect 108 249 173 265
rect 142 215 173 249
rect 108 199 173 215
rect 207 249 257 268
rect 207 215 214 249
rect 248 215 257 249
rect 30 127 77 161
rect 111 127 127 161
rect 207 145 257 215
rect 298 249 373 268
rect 298 215 329 249
rect 363 215 373 249
rect 298 199 373 215
rect 407 249 680 271
rect 407 215 464 249
rect 498 215 542 249
rect 576 215 620 249
rect 654 215 680 249
rect 407 204 680 215
rect 407 161 453 204
rect 714 169 799 307
rect 30 109 127 127
rect 304 123 453 161
rect 497 153 691 169
rect 304 109 340 123
rect 30 93 340 109
rect 497 119 499 153
rect 533 135 691 153
rect 725 135 799 169
rect 533 123 799 135
rect 833 249 891 341
rect 867 215 891 249
rect 833 123 891 215
rect 925 135 981 375
rect 533 119 535 123
rect 497 103 535 119
rect 30 59 77 93
rect 111 71 340 93
rect 673 101 727 123
rect 111 59 127 71
rect 30 51 127 59
rect 386 55 402 89
rect 436 55 452 89
rect 386 17 452 55
rect 569 55 589 89
rect 623 55 639 89
rect 569 17 639 55
rect 673 67 691 101
rect 725 67 727 101
rect 959 101 981 135
rect 673 51 727 67
rect 761 55 787 89
rect 821 55 837 89
rect 925 85 981 101
rect 761 17 837 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel locali s 855 221 889 255 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 743 153 777 187 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 298 199 373 268 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 221 257 255 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and3b_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1012 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1825788
string GDS_START 1818756
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
