magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 331 1478 704
<< pwell >>
rect 61 49 1439 243
rect 0 0 1440 49
<< scnmos >>
rect 140 49 170 217
rect 226 49 256 217
rect 312 49 342 217
rect 398 49 428 217
rect 484 49 514 217
rect 570 49 600 217
rect 656 49 686 217
rect 742 49 772 217
rect 837 49 867 217
rect 923 49 953 217
rect 1009 49 1039 217
rect 1217 49 1247 217
rect 1330 133 1360 217
<< scpmoshvt >>
rect 140 367 170 619
rect 226 367 256 619
rect 312 367 342 619
rect 398 367 428 619
rect 484 367 514 619
rect 570 367 600 619
rect 656 367 686 619
rect 742 367 772 619
rect 837 367 867 619
rect 923 367 953 619
rect 1009 367 1039 619
rect 1225 367 1255 619
rect 1330 367 1360 495
<< ndiff >>
rect 87 168 140 217
rect 87 134 95 168
rect 129 134 140 168
rect 87 100 140 134
rect 87 66 95 100
rect 129 66 140 100
rect 87 49 140 66
rect 170 192 226 217
rect 170 158 181 192
rect 215 158 226 192
rect 170 108 226 158
rect 170 74 181 108
rect 215 74 226 108
rect 170 49 226 74
rect 256 168 312 217
rect 256 134 267 168
rect 301 134 312 168
rect 256 100 312 134
rect 256 66 267 100
rect 301 66 312 100
rect 256 49 312 66
rect 342 192 398 217
rect 342 158 353 192
rect 387 158 398 192
rect 342 108 398 158
rect 342 74 353 108
rect 387 74 398 108
rect 342 49 398 74
rect 428 168 484 217
rect 428 134 439 168
rect 473 134 484 168
rect 428 100 484 134
rect 428 66 439 100
rect 473 66 484 100
rect 428 49 484 66
rect 514 192 570 217
rect 514 158 525 192
rect 559 158 570 192
rect 514 108 570 158
rect 514 74 525 108
rect 559 74 570 108
rect 514 49 570 74
rect 600 168 656 217
rect 600 134 611 168
rect 645 134 656 168
rect 600 100 656 134
rect 600 66 611 100
rect 645 66 656 100
rect 600 49 656 66
rect 686 192 742 217
rect 686 158 697 192
rect 731 158 742 192
rect 686 108 742 158
rect 686 74 697 108
rect 731 74 742 108
rect 686 49 742 74
rect 772 168 837 217
rect 772 134 788 168
rect 822 134 837 168
rect 772 100 837 134
rect 772 66 788 100
rect 822 66 837 100
rect 772 49 837 66
rect 867 192 923 217
rect 867 158 878 192
rect 912 158 923 192
rect 867 108 923 158
rect 867 74 878 108
rect 912 74 923 108
rect 867 49 923 74
rect 953 168 1009 217
rect 953 134 964 168
rect 998 134 1009 168
rect 953 100 1009 134
rect 953 66 964 100
rect 998 66 1009 100
rect 953 49 1009 66
rect 1039 192 1092 217
rect 1039 158 1050 192
rect 1084 158 1092 192
rect 1039 108 1092 158
rect 1039 74 1050 108
rect 1084 74 1092 108
rect 1039 49 1092 74
rect 1160 205 1217 217
rect 1160 171 1168 205
rect 1202 171 1217 205
rect 1160 137 1217 171
rect 1160 103 1168 137
rect 1202 103 1217 137
rect 1160 49 1217 103
rect 1247 174 1330 217
rect 1247 140 1258 174
rect 1292 140 1330 174
rect 1247 133 1330 140
rect 1360 192 1413 217
rect 1360 158 1371 192
rect 1405 158 1413 192
rect 1360 133 1413 158
rect 1247 95 1300 133
rect 1247 61 1258 95
rect 1292 61 1300 95
rect 1247 49 1300 61
<< pdiff >>
rect 83 607 140 619
rect 83 573 95 607
rect 129 573 140 607
rect 83 539 140 573
rect 83 505 95 539
rect 129 505 140 539
rect 83 471 140 505
rect 83 437 95 471
rect 129 437 140 471
rect 83 367 140 437
rect 170 585 226 619
rect 170 551 181 585
rect 215 551 226 585
rect 170 506 226 551
rect 170 472 181 506
rect 215 472 226 506
rect 170 427 226 472
rect 170 393 181 427
rect 215 393 226 427
rect 170 367 226 393
rect 256 607 312 619
rect 256 573 267 607
rect 301 573 312 607
rect 256 539 312 573
rect 256 505 267 539
rect 301 505 312 539
rect 256 471 312 505
rect 256 437 267 471
rect 301 437 312 471
rect 256 367 312 437
rect 342 585 398 619
rect 342 551 353 585
rect 387 551 398 585
rect 342 506 398 551
rect 342 472 353 506
rect 387 472 398 506
rect 342 427 398 472
rect 342 393 353 427
rect 387 393 398 427
rect 342 367 398 393
rect 428 607 484 619
rect 428 573 439 607
rect 473 573 484 607
rect 428 539 484 573
rect 428 505 439 539
rect 473 505 484 539
rect 428 471 484 505
rect 428 437 439 471
rect 473 437 484 471
rect 428 367 484 437
rect 514 585 570 619
rect 514 551 525 585
rect 559 551 570 585
rect 514 506 570 551
rect 514 472 525 506
rect 559 472 570 506
rect 514 427 570 472
rect 514 393 525 427
rect 559 393 570 427
rect 514 367 570 393
rect 600 607 656 619
rect 600 573 611 607
rect 645 573 656 607
rect 600 539 656 573
rect 600 505 611 539
rect 645 505 656 539
rect 600 471 656 505
rect 600 437 611 471
rect 645 437 656 471
rect 600 367 656 437
rect 686 585 742 619
rect 686 551 697 585
rect 731 551 742 585
rect 686 506 742 551
rect 686 472 697 506
rect 731 472 742 506
rect 686 427 742 472
rect 686 393 697 427
rect 731 393 742 427
rect 686 367 742 393
rect 772 599 837 619
rect 772 565 783 599
rect 817 565 837 599
rect 772 531 837 565
rect 772 497 783 531
rect 817 497 837 531
rect 772 463 837 497
rect 772 429 783 463
rect 817 429 837 463
rect 772 367 837 429
rect 867 585 923 619
rect 867 551 878 585
rect 912 551 923 585
rect 867 506 923 551
rect 867 472 878 506
rect 912 472 923 506
rect 867 427 923 472
rect 867 393 878 427
rect 912 393 923 427
rect 867 367 923 393
rect 953 605 1009 619
rect 953 571 964 605
rect 998 571 1009 605
rect 953 537 1009 571
rect 953 503 964 537
rect 998 503 1009 537
rect 953 469 1009 503
rect 953 435 964 469
rect 998 435 1009 469
rect 953 367 1009 435
rect 1039 585 1092 619
rect 1039 551 1050 585
rect 1084 551 1092 585
rect 1039 506 1092 551
rect 1039 472 1050 506
rect 1084 472 1092 506
rect 1039 427 1092 472
rect 1039 393 1050 427
rect 1084 393 1092 427
rect 1039 367 1092 393
rect 1172 549 1225 619
rect 1172 515 1180 549
rect 1214 515 1225 549
rect 1172 481 1225 515
rect 1172 447 1180 481
rect 1214 447 1225 481
rect 1172 413 1225 447
rect 1172 379 1180 413
rect 1214 379 1225 413
rect 1172 367 1225 379
rect 1255 588 1308 619
rect 1255 554 1266 588
rect 1300 554 1308 588
rect 1255 512 1308 554
rect 1255 478 1266 512
rect 1300 495 1308 512
rect 1300 478 1330 495
rect 1255 367 1330 478
rect 1360 429 1413 495
rect 1360 395 1371 429
rect 1405 395 1413 429
rect 1360 367 1413 395
<< ndiffc >>
rect 95 134 129 168
rect 95 66 129 100
rect 181 158 215 192
rect 181 74 215 108
rect 267 134 301 168
rect 267 66 301 100
rect 353 158 387 192
rect 353 74 387 108
rect 439 134 473 168
rect 439 66 473 100
rect 525 158 559 192
rect 525 74 559 108
rect 611 134 645 168
rect 611 66 645 100
rect 697 158 731 192
rect 697 74 731 108
rect 788 134 822 168
rect 788 66 822 100
rect 878 158 912 192
rect 878 74 912 108
rect 964 134 998 168
rect 964 66 998 100
rect 1050 158 1084 192
rect 1050 74 1084 108
rect 1168 171 1202 205
rect 1168 103 1202 137
rect 1258 140 1292 174
rect 1371 158 1405 192
rect 1258 61 1292 95
<< pdiffc >>
rect 95 573 129 607
rect 95 505 129 539
rect 95 437 129 471
rect 181 551 215 585
rect 181 472 215 506
rect 181 393 215 427
rect 267 573 301 607
rect 267 505 301 539
rect 267 437 301 471
rect 353 551 387 585
rect 353 472 387 506
rect 353 393 387 427
rect 439 573 473 607
rect 439 505 473 539
rect 439 437 473 471
rect 525 551 559 585
rect 525 472 559 506
rect 525 393 559 427
rect 611 573 645 607
rect 611 505 645 539
rect 611 437 645 471
rect 697 551 731 585
rect 697 472 731 506
rect 697 393 731 427
rect 783 565 817 599
rect 783 497 817 531
rect 783 429 817 463
rect 878 551 912 585
rect 878 472 912 506
rect 878 393 912 427
rect 964 571 998 605
rect 964 503 998 537
rect 964 435 998 469
rect 1050 551 1084 585
rect 1050 472 1084 506
rect 1050 393 1084 427
rect 1180 515 1214 549
rect 1180 447 1214 481
rect 1180 379 1214 413
rect 1266 554 1300 588
rect 1266 478 1300 512
rect 1371 395 1405 429
<< poly >>
rect 140 619 170 645
rect 226 619 256 645
rect 312 619 342 645
rect 398 619 428 645
rect 484 619 514 645
rect 570 619 600 645
rect 656 619 686 645
rect 742 619 772 645
rect 837 619 867 645
rect 923 619 953 645
rect 1009 619 1039 645
rect 1225 619 1255 645
rect 1330 495 1360 521
rect 140 331 170 367
rect 226 331 256 367
rect 312 331 342 367
rect 398 331 428 367
rect 484 331 514 367
rect 570 331 600 367
rect 656 331 686 367
rect 742 331 772 367
rect 837 331 867 367
rect 923 331 953 367
rect 1009 331 1039 367
rect 117 315 795 331
rect 117 281 133 315
rect 167 281 201 315
rect 235 281 269 315
rect 303 281 337 315
rect 371 281 405 315
rect 439 281 473 315
rect 507 281 541 315
rect 575 281 609 315
rect 643 281 677 315
rect 711 281 745 315
rect 779 281 795 315
rect 117 265 795 281
rect 837 315 1175 331
rect 837 281 853 315
rect 887 281 921 315
rect 955 281 989 315
rect 1023 281 1057 315
rect 1091 281 1125 315
rect 1159 281 1175 315
rect 1225 305 1255 367
rect 1330 335 1360 367
rect 1330 315 1396 335
rect 837 265 1175 281
rect 1217 289 1288 305
rect 140 217 170 265
rect 226 217 256 265
rect 312 217 342 265
rect 398 217 428 265
rect 484 217 514 265
rect 570 217 600 265
rect 656 217 686 265
rect 742 217 772 265
rect 837 217 867 265
rect 923 217 953 265
rect 1009 217 1039 265
rect 1217 255 1238 289
rect 1272 255 1288 289
rect 1217 239 1288 255
rect 1330 281 1346 315
rect 1380 281 1396 315
rect 1330 265 1396 281
rect 1217 217 1247 239
rect 1330 217 1360 265
rect 1330 107 1360 133
rect 140 23 170 49
rect 226 23 256 49
rect 312 23 342 49
rect 398 23 428 49
rect 484 23 514 49
rect 570 23 600 49
rect 656 23 686 49
rect 742 23 772 49
rect 837 23 867 49
rect 923 23 953 49
rect 1009 23 1039 49
rect 1217 23 1247 49
<< polycont >>
rect 133 281 167 315
rect 201 281 235 315
rect 269 281 303 315
rect 337 281 371 315
rect 405 281 439 315
rect 473 281 507 315
rect 541 281 575 315
rect 609 281 643 315
rect 677 281 711 315
rect 745 281 779 315
rect 853 281 887 315
rect 921 281 955 315
rect 989 281 1023 315
rect 1057 281 1091 315
rect 1125 281 1159 315
rect 1238 255 1272 289
rect 1346 281 1380 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 79 607 138 649
rect 79 573 95 607
rect 129 573 138 607
rect 79 539 138 573
rect 79 505 95 539
rect 129 505 138 539
rect 79 471 138 505
rect 79 437 95 471
rect 129 437 138 471
rect 79 421 138 437
rect 172 585 224 615
rect 172 551 181 585
rect 215 551 224 585
rect 172 506 224 551
rect 172 472 181 506
rect 215 472 224 506
rect 172 427 224 472
rect 172 393 181 427
rect 215 393 224 427
rect 258 607 310 649
rect 258 573 267 607
rect 301 573 310 607
rect 258 539 310 573
rect 258 505 267 539
rect 301 505 310 539
rect 258 471 310 505
rect 258 437 267 471
rect 301 437 310 471
rect 258 421 310 437
rect 344 585 396 615
rect 344 551 353 585
rect 387 551 396 585
rect 344 506 396 551
rect 344 472 353 506
rect 387 472 396 506
rect 344 427 396 472
rect 172 385 224 393
rect 344 393 353 427
rect 387 393 396 427
rect 430 607 482 649
rect 430 573 439 607
rect 473 573 482 607
rect 430 539 482 573
rect 430 505 439 539
rect 473 505 482 539
rect 430 471 482 505
rect 430 437 439 471
rect 473 437 482 471
rect 430 421 482 437
rect 516 585 568 615
rect 516 551 525 585
rect 559 551 568 585
rect 516 506 568 551
rect 516 472 525 506
rect 559 472 568 506
rect 516 427 568 472
rect 344 385 396 393
rect 516 393 525 427
rect 559 393 568 427
rect 602 607 654 649
rect 602 573 611 607
rect 645 573 654 607
rect 602 539 654 573
rect 602 505 611 539
rect 645 505 654 539
rect 602 471 654 505
rect 602 437 611 471
rect 645 437 654 471
rect 602 421 654 437
rect 688 585 733 615
rect 688 551 697 585
rect 731 551 733 585
rect 688 506 733 551
rect 688 472 697 506
rect 731 472 733 506
rect 688 427 733 472
rect 516 385 568 393
rect 688 393 697 427
rect 731 393 733 427
rect 767 599 833 649
rect 767 565 783 599
rect 817 565 833 599
rect 767 531 833 565
rect 767 497 783 531
rect 817 497 833 531
rect 767 463 833 497
rect 767 429 783 463
rect 817 429 833 463
rect 767 419 833 429
rect 867 585 922 615
rect 867 551 878 585
rect 912 551 922 585
rect 867 506 922 551
rect 867 472 878 506
rect 912 472 922 506
rect 867 427 922 472
rect 688 385 733 393
rect 867 393 878 427
rect 912 393 922 427
rect 956 605 1008 649
rect 956 571 964 605
rect 998 571 1008 605
rect 956 537 1008 571
rect 956 503 964 537
rect 998 503 1008 537
rect 956 469 1008 503
rect 956 435 964 469
rect 998 435 1008 469
rect 956 419 1008 435
rect 1042 585 1100 615
rect 1042 551 1050 585
rect 1084 551 1100 585
rect 1250 588 1316 649
rect 1042 506 1100 551
rect 1042 472 1050 506
rect 1084 472 1100 506
rect 1042 427 1100 472
rect 867 385 922 393
rect 1042 393 1050 427
rect 1084 393 1100 427
rect 1042 385 1100 393
rect 17 351 733 385
rect 767 351 1100 385
rect 1168 549 1214 565
rect 1168 515 1180 549
rect 1168 481 1214 515
rect 1168 447 1180 481
rect 1250 554 1266 588
rect 1300 554 1316 588
rect 1250 512 1316 554
rect 1250 478 1266 512
rect 1300 478 1316 512
rect 1250 474 1316 478
rect 1168 413 1214 447
rect 1168 379 1180 413
rect 1168 363 1214 379
rect 1248 429 1421 440
rect 1248 395 1371 429
rect 1405 395 1421 429
rect 1248 385 1421 395
rect 17 245 81 351
rect 767 317 801 351
rect 1168 317 1204 363
rect 117 315 801 317
rect 117 281 133 315
rect 167 281 201 315
rect 235 281 269 315
rect 303 281 337 315
rect 371 281 405 315
rect 439 281 473 315
rect 507 281 541 315
rect 575 281 609 315
rect 643 281 677 315
rect 711 281 745 315
rect 779 281 801 315
rect 117 279 801 281
rect 837 315 1204 317
rect 837 281 853 315
rect 887 281 921 315
rect 955 281 989 315
rect 1023 281 1057 315
rect 1091 281 1125 315
rect 1159 281 1204 315
rect 1248 305 1288 385
rect 837 279 1204 281
rect 767 245 801 279
rect 17 211 733 245
rect 767 211 1100 245
rect 179 192 217 211
rect 79 168 145 177
rect 79 134 95 168
rect 129 134 145 168
rect 79 100 145 134
rect 79 66 95 100
rect 129 66 145 100
rect 79 17 145 66
rect 179 158 181 192
rect 215 158 217 192
rect 351 192 389 211
rect 179 108 217 158
rect 179 74 181 108
rect 215 74 217 108
rect 179 58 217 74
rect 251 168 317 177
rect 251 134 267 168
rect 301 134 317 168
rect 251 100 317 134
rect 251 66 267 100
rect 301 66 317 100
rect 251 17 317 66
rect 351 158 353 192
rect 387 158 389 192
rect 523 192 561 211
rect 351 108 389 158
rect 351 74 353 108
rect 387 74 389 108
rect 351 58 389 74
rect 423 168 489 177
rect 423 134 439 168
rect 473 134 489 168
rect 423 100 489 134
rect 423 66 439 100
rect 473 66 489 100
rect 423 17 489 66
rect 523 158 525 192
rect 559 158 561 192
rect 695 192 733 211
rect 523 108 561 158
rect 523 74 525 108
rect 559 74 561 108
rect 523 58 561 74
rect 595 168 661 177
rect 595 134 611 168
rect 645 134 661 168
rect 595 100 661 134
rect 595 66 611 100
rect 645 66 661 100
rect 595 17 661 66
rect 695 158 697 192
rect 731 158 733 192
rect 872 192 914 211
rect 695 108 733 158
rect 695 74 697 108
rect 731 74 733 108
rect 695 58 733 74
rect 767 168 838 177
rect 767 134 788 168
rect 822 134 838 168
rect 767 100 838 134
rect 767 66 788 100
rect 822 66 838 100
rect 767 17 838 66
rect 872 158 878 192
rect 912 158 914 192
rect 1048 192 1100 211
rect 872 108 914 158
rect 872 74 878 108
rect 912 74 914 108
rect 872 58 914 74
rect 948 168 1014 177
rect 948 134 964 168
rect 998 134 1014 168
rect 948 100 1014 134
rect 948 66 964 100
rect 998 66 1014 100
rect 948 17 1014 66
rect 1048 158 1050 192
rect 1084 158 1100 192
rect 1048 108 1100 158
rect 1048 74 1050 108
rect 1084 74 1100 108
rect 1152 205 1204 279
rect 1238 289 1288 305
rect 1272 255 1288 289
rect 1330 315 1423 351
rect 1330 281 1346 315
rect 1380 281 1423 315
rect 1238 247 1288 255
rect 1238 213 1421 247
rect 1152 171 1168 205
rect 1202 171 1204 205
rect 1355 192 1421 213
rect 1152 137 1204 171
rect 1152 103 1168 137
rect 1202 103 1204 137
rect 1152 87 1204 103
rect 1242 174 1308 179
rect 1242 140 1258 174
rect 1292 140 1308 174
rect 1242 95 1308 140
rect 1355 158 1371 192
rect 1405 158 1421 192
rect 1355 133 1421 158
rect 1048 58 1100 74
rect 1242 61 1258 95
rect 1292 61 1308 95
rect 1242 17 1308 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 bufbuf_8
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6817232
string GDS_START 6805032
<< end >>
