magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2126 1852
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 16 21 787 203
rect 29 -17 63 21
<< scnmos >>
rect 94 47 124 177
rect 200 47 230 177
rect 289 47 319 177
rect 487 47 517 177
rect 581 47 611 177
rect 665 47 695 177
<< scpmoshvt >>
rect 86 297 122 497
rect 192 297 228 497
rect 274 297 310 497
rect 479 297 515 497
rect 561 297 597 497
rect 667 297 703 497
<< ndiff >>
rect 42 163 94 177
rect 42 129 50 163
rect 84 129 94 163
rect 42 95 94 129
rect 42 61 50 95
rect 84 61 94 95
rect 42 47 94 61
rect 124 95 200 177
rect 124 61 156 95
rect 190 61 200 95
rect 124 47 200 61
rect 230 163 289 177
rect 230 129 240 163
rect 274 129 289 163
rect 230 47 289 129
rect 319 95 371 177
rect 319 61 329 95
rect 363 61 371 95
rect 319 47 371 61
rect 425 95 487 177
rect 425 61 433 95
rect 467 61 487 95
rect 425 47 487 61
rect 517 163 581 177
rect 517 129 537 163
rect 571 129 581 163
rect 517 95 581 129
rect 517 61 537 95
rect 571 61 581 95
rect 517 47 581 61
rect 611 95 665 177
rect 611 61 621 95
rect 655 61 665 95
rect 611 47 665 61
rect 695 163 761 177
rect 695 129 715 163
rect 749 129 761 163
rect 695 95 761 129
rect 695 61 715 95
rect 749 61 761 95
rect 695 47 761 61
<< pdiff >>
rect 27 477 86 497
rect 27 443 39 477
rect 73 443 86 477
rect 27 409 86 443
rect 27 375 39 409
rect 73 375 86 409
rect 27 341 86 375
rect 27 307 39 341
rect 73 307 86 341
rect 27 297 86 307
rect 122 477 192 497
rect 122 443 138 477
rect 172 443 192 477
rect 122 297 192 443
rect 228 297 274 497
rect 310 477 479 497
rect 310 443 322 477
rect 356 443 433 477
rect 467 443 479 477
rect 310 409 479 443
rect 310 375 322 409
rect 356 375 433 409
rect 467 375 479 409
rect 310 297 479 375
rect 515 297 561 497
rect 597 477 667 497
rect 597 443 609 477
rect 643 443 667 477
rect 597 409 667 443
rect 597 375 609 409
rect 643 375 667 409
rect 597 297 667 375
rect 703 477 761 497
rect 703 443 719 477
rect 753 443 761 477
rect 703 409 761 443
rect 703 375 719 409
rect 753 375 761 409
rect 703 297 761 375
<< ndiffc >>
rect 50 129 84 163
rect 50 61 84 95
rect 156 61 190 95
rect 240 129 274 163
rect 329 61 363 95
rect 433 61 467 95
rect 537 129 571 163
rect 537 61 571 95
rect 621 61 655 95
rect 715 129 749 163
rect 715 61 749 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 138 443 172 477
rect 322 443 356 477
rect 433 443 467 477
rect 322 375 356 409
rect 433 375 467 409
rect 609 443 643 477
rect 609 375 643 409
rect 719 443 753 477
rect 719 375 753 409
<< poly >>
rect 86 497 122 523
rect 192 497 228 523
rect 274 497 310 523
rect 479 497 515 523
rect 561 497 597 523
rect 667 497 703 523
rect 86 282 122 297
rect 192 282 228 297
rect 274 282 310 297
rect 479 282 515 297
rect 561 282 597 297
rect 667 282 703 297
rect 84 265 124 282
rect 190 265 230 282
rect 23 249 124 265
rect 23 215 33 249
rect 67 215 124 249
rect 23 199 124 215
rect 94 177 124 199
rect 176 249 230 265
rect 176 215 186 249
rect 220 215 230 249
rect 176 197 230 215
rect 272 265 312 282
rect 477 265 517 282
rect 272 249 326 265
rect 272 215 282 249
rect 316 215 326 249
rect 272 199 326 215
rect 463 249 517 265
rect 463 215 473 249
rect 507 215 517 249
rect 463 199 517 215
rect 559 265 599 282
rect 665 265 705 282
rect 559 249 623 265
rect 559 215 579 249
rect 613 215 623 249
rect 559 199 623 215
rect 665 249 719 265
rect 665 215 675 249
rect 709 215 719 249
rect 665 199 719 215
rect 200 177 230 197
rect 289 177 319 199
rect 487 177 517 199
rect 581 177 611 199
rect 665 177 695 199
rect 94 21 124 47
rect 200 21 230 47
rect 289 21 319 47
rect 487 21 517 47
rect 581 21 611 47
rect 665 21 695 47
<< polycont >>
rect 33 215 67 249
rect 186 215 220 249
rect 282 215 316 249
rect 473 215 507 249
rect 579 215 613 249
rect 675 215 709 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 477 73 493
rect 17 443 39 477
rect 17 409 73 443
rect 112 477 172 527
rect 112 443 138 477
rect 112 417 172 443
rect 300 477 471 493
rect 300 443 322 477
rect 356 443 433 477
rect 467 443 471 477
rect 300 409 471 443
rect 583 477 659 527
rect 583 443 609 477
rect 643 443 659 477
rect 583 409 659 443
rect 17 375 39 409
rect 17 344 73 375
rect 206 375 322 409
rect 356 375 433 409
rect 467 375 549 409
rect 206 344 247 375
rect 17 341 247 344
rect 17 307 39 341
rect 73 307 247 341
rect 17 299 247 307
rect 17 291 151 299
rect 17 249 83 257
rect 17 215 33 249
rect 67 215 83 249
rect 17 199 83 215
rect 117 165 151 291
rect 185 249 247 265
rect 185 215 186 249
rect 220 215 247 249
rect 185 197 247 215
rect 281 249 358 341
rect 281 215 282 249
rect 316 215 358 249
rect 281 197 358 215
rect 396 251 463 341
rect 515 325 549 375
rect 583 375 609 409
rect 643 375 659 409
rect 693 477 806 493
rect 693 443 719 477
rect 753 443 806 477
rect 693 409 806 443
rect 693 375 719 409
rect 753 375 806 409
rect 583 359 659 375
rect 515 291 709 325
rect 396 249 523 251
rect 396 215 473 249
rect 507 215 523 249
rect 563 249 629 257
rect 563 215 579 249
rect 613 215 629 249
rect 675 249 709 291
rect 396 197 523 215
rect 675 199 709 215
rect 743 165 806 375
rect 34 163 151 165
rect 689 163 806 165
rect 34 129 50 163
rect 84 129 151 163
rect 207 129 240 163
rect 274 129 537 163
rect 571 129 587 163
rect 34 95 100 129
rect 521 95 587 129
rect 689 129 715 163
rect 749 129 806 163
rect 34 61 50 95
rect 84 61 100 95
rect 140 61 156 95
rect 190 61 329 95
rect 363 61 381 95
rect 417 61 433 95
rect 467 61 485 95
rect 34 51 100 61
rect 417 17 485 61
rect 521 61 537 95
rect 571 61 587 95
rect 521 54 587 61
rect 621 95 655 128
rect 621 17 655 61
rect 689 95 806 129
rect 689 61 715 95
rect 749 61 806 95
rect 689 53 806 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 396 251 463 341 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 759 357 793 391 0 FreeSans 400 0 0 0 X
port 10 nsew signal output
flabel locali s 188 221 232 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 C1
port 5 nsew signal input
flabel locali s 570 221 604 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 432 306 432 306 0 FreeSans 400 0 0 0 A2
port 2 nsew
flabel locali s 290 221 324 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 290 293 324 327 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221a_1
rlabel locali s 396 197 523 251 1 A2
port 2 nsew signal input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2484088
string GDS_START 2476826
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
