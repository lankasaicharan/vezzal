magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3322 1852
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 2 21 2019 203
rect 30 -17 64 21
<< scnmos >>
rect 93 47 123 177
rect 177 47 207 177
rect 383 47 413 177
rect 477 47 507 177
rect 571 47 601 177
rect 675 47 705 177
rect 759 47 789 177
rect 853 47 883 177
rect 947 47 977 177
rect 1051 47 1081 177
rect 1239 47 1269 177
rect 1333 47 1363 177
rect 1427 47 1457 177
rect 1531 47 1561 177
rect 1615 47 1645 177
rect 1709 47 1739 177
rect 1803 47 1833 177
rect 1907 47 1937 177
<< scpmoshvt >>
rect 85 297 121 497
rect 179 297 215 497
rect 385 297 421 497
rect 479 297 515 497
rect 573 297 609 497
rect 667 297 703 497
rect 761 297 797 497
rect 855 297 891 497
rect 949 297 985 497
rect 1043 297 1079 497
rect 1241 297 1277 497
rect 1335 297 1371 497
rect 1429 297 1465 497
rect 1523 297 1559 497
rect 1617 297 1653 497
rect 1711 297 1747 497
rect 1805 297 1841 497
rect 1899 297 1935 497
<< ndiff >>
rect 28 163 93 177
rect 28 129 39 163
rect 73 129 93 163
rect 28 95 93 129
rect 28 61 39 95
rect 73 61 93 95
rect 28 47 93 61
rect 123 95 177 177
rect 123 61 133 95
rect 167 61 177 95
rect 123 47 177 61
rect 207 163 269 177
rect 207 129 227 163
rect 261 129 269 163
rect 207 95 269 129
rect 207 61 227 95
rect 261 61 269 95
rect 207 47 269 61
rect 331 95 383 177
rect 331 61 339 95
rect 373 61 383 95
rect 331 47 383 61
rect 413 163 477 177
rect 413 129 433 163
rect 467 129 477 163
rect 413 95 477 129
rect 413 61 433 95
rect 467 61 477 95
rect 413 47 477 61
rect 507 95 571 177
rect 507 61 527 95
rect 561 61 571 95
rect 507 47 571 61
rect 601 163 675 177
rect 601 129 621 163
rect 655 129 675 163
rect 601 95 675 129
rect 601 61 621 95
rect 655 61 675 95
rect 601 47 675 61
rect 705 95 759 177
rect 705 61 715 95
rect 749 61 759 95
rect 705 47 759 61
rect 789 163 853 177
rect 789 129 809 163
rect 843 129 853 163
rect 789 95 853 129
rect 789 61 809 95
rect 843 61 853 95
rect 789 47 853 61
rect 883 95 947 177
rect 883 61 903 95
rect 937 61 947 95
rect 883 47 947 61
rect 977 163 1051 177
rect 977 129 997 163
rect 1031 129 1051 163
rect 977 95 1051 129
rect 977 61 997 95
rect 1031 61 1051 95
rect 977 47 1051 61
rect 1081 95 1239 177
rect 1081 61 1091 95
rect 1125 61 1195 95
rect 1229 61 1239 95
rect 1081 47 1239 61
rect 1269 163 1333 177
rect 1269 129 1289 163
rect 1323 129 1333 163
rect 1269 95 1333 129
rect 1269 61 1289 95
rect 1323 61 1333 95
rect 1269 47 1333 61
rect 1363 95 1427 177
rect 1363 61 1383 95
rect 1417 61 1427 95
rect 1363 47 1427 61
rect 1457 163 1531 177
rect 1457 129 1477 163
rect 1511 129 1531 163
rect 1457 95 1531 129
rect 1457 61 1477 95
rect 1511 61 1531 95
rect 1457 47 1531 61
rect 1561 95 1615 177
rect 1561 61 1571 95
rect 1605 61 1615 95
rect 1561 47 1615 61
rect 1645 163 1709 177
rect 1645 129 1665 163
rect 1699 129 1709 163
rect 1645 95 1709 129
rect 1645 61 1665 95
rect 1699 61 1709 95
rect 1645 47 1709 61
rect 1739 95 1803 177
rect 1739 61 1759 95
rect 1793 61 1803 95
rect 1739 47 1803 61
rect 1833 163 1907 177
rect 1833 129 1853 163
rect 1887 129 1907 163
rect 1833 95 1907 129
rect 1833 61 1853 95
rect 1887 61 1907 95
rect 1833 47 1907 61
rect 1937 163 1993 177
rect 1937 129 1947 163
rect 1981 129 1993 163
rect 1937 95 1993 129
rect 1937 61 1947 95
rect 1981 61 1993 95
rect 1937 47 1993 61
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 179 497
rect 121 443 133 477
rect 167 443 179 477
rect 121 297 179 443
rect 215 341 273 497
rect 215 307 227 341
rect 261 307 273 341
rect 215 297 273 307
rect 331 477 385 497
rect 331 443 339 477
rect 373 443 385 477
rect 331 297 385 443
rect 421 341 479 497
rect 421 307 433 341
rect 467 307 479 341
rect 421 297 479 307
rect 515 477 573 497
rect 515 443 527 477
rect 561 443 573 477
rect 515 297 573 443
rect 609 341 667 497
rect 609 307 621 341
rect 655 307 667 341
rect 609 297 667 307
rect 703 477 761 497
rect 703 443 715 477
rect 749 443 761 477
rect 703 297 761 443
rect 797 409 855 497
rect 797 375 809 409
rect 843 375 855 409
rect 797 341 855 375
rect 797 307 809 341
rect 843 307 855 341
rect 797 297 855 307
rect 891 477 949 497
rect 891 443 903 477
rect 937 443 949 477
rect 891 409 949 443
rect 891 375 903 409
rect 937 375 949 409
rect 891 297 949 375
rect 985 409 1043 497
rect 985 375 997 409
rect 1031 375 1043 409
rect 985 341 1043 375
rect 985 307 997 341
rect 1031 307 1043 341
rect 985 297 1043 307
rect 1079 477 1133 497
rect 1079 443 1091 477
rect 1125 443 1133 477
rect 1079 409 1133 443
rect 1079 375 1091 409
rect 1125 375 1133 409
rect 1079 297 1133 375
rect 1187 477 1241 497
rect 1187 443 1195 477
rect 1229 443 1241 477
rect 1187 409 1241 443
rect 1187 375 1195 409
rect 1229 375 1241 409
rect 1187 297 1241 375
rect 1277 409 1335 497
rect 1277 375 1289 409
rect 1323 375 1335 409
rect 1277 341 1335 375
rect 1277 307 1289 341
rect 1323 307 1335 341
rect 1277 297 1335 307
rect 1371 477 1429 497
rect 1371 443 1383 477
rect 1417 443 1429 477
rect 1371 409 1429 443
rect 1371 375 1383 409
rect 1417 375 1429 409
rect 1371 297 1429 375
rect 1465 409 1523 497
rect 1465 375 1477 409
rect 1511 375 1523 409
rect 1465 341 1523 375
rect 1465 307 1477 341
rect 1511 307 1523 341
rect 1465 297 1523 307
rect 1559 477 1617 497
rect 1559 443 1571 477
rect 1605 443 1617 477
rect 1559 409 1617 443
rect 1559 375 1571 409
rect 1605 375 1617 409
rect 1559 341 1617 375
rect 1559 307 1571 341
rect 1605 307 1617 341
rect 1559 297 1617 307
rect 1653 477 1711 497
rect 1653 443 1665 477
rect 1699 443 1711 477
rect 1653 409 1711 443
rect 1653 375 1665 409
rect 1699 375 1711 409
rect 1653 297 1711 375
rect 1747 477 1805 497
rect 1747 443 1759 477
rect 1793 443 1805 477
rect 1747 409 1805 443
rect 1747 375 1759 409
rect 1793 375 1805 409
rect 1747 341 1805 375
rect 1747 307 1759 341
rect 1793 307 1805 341
rect 1747 297 1805 307
rect 1841 477 1899 497
rect 1841 443 1853 477
rect 1887 443 1899 477
rect 1841 409 1899 443
rect 1841 375 1853 409
rect 1887 375 1899 409
rect 1841 297 1899 375
rect 1935 477 1993 497
rect 1935 443 1947 477
rect 1981 443 1993 477
rect 1935 409 1993 443
rect 1935 375 1947 409
rect 1981 375 1993 409
rect 1935 341 1993 375
rect 1935 307 1947 341
rect 1981 307 1993 341
rect 1935 297 1993 307
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 133 61 167 95
rect 227 129 261 163
rect 227 61 261 95
rect 339 61 373 95
rect 433 129 467 163
rect 433 61 467 95
rect 527 61 561 95
rect 621 129 655 163
rect 621 61 655 95
rect 715 61 749 95
rect 809 129 843 163
rect 809 61 843 95
rect 903 61 937 95
rect 997 129 1031 163
rect 997 61 1031 95
rect 1091 61 1125 95
rect 1195 61 1229 95
rect 1289 129 1323 163
rect 1289 61 1323 95
rect 1383 61 1417 95
rect 1477 129 1511 163
rect 1477 61 1511 95
rect 1571 61 1605 95
rect 1665 129 1699 163
rect 1665 61 1699 95
rect 1759 61 1793 95
rect 1853 129 1887 163
rect 1853 61 1887 95
rect 1947 129 1981 163
rect 1947 61 1981 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 133 443 167 477
rect 227 307 261 341
rect 339 443 373 477
rect 433 307 467 341
rect 527 443 561 477
rect 621 307 655 341
rect 715 443 749 477
rect 809 375 843 409
rect 809 307 843 341
rect 903 443 937 477
rect 903 375 937 409
rect 997 375 1031 409
rect 997 307 1031 341
rect 1091 443 1125 477
rect 1091 375 1125 409
rect 1195 443 1229 477
rect 1195 375 1229 409
rect 1289 375 1323 409
rect 1289 307 1323 341
rect 1383 443 1417 477
rect 1383 375 1417 409
rect 1477 375 1511 409
rect 1477 307 1511 341
rect 1571 443 1605 477
rect 1571 375 1605 409
rect 1571 307 1605 341
rect 1665 443 1699 477
rect 1665 375 1699 409
rect 1759 443 1793 477
rect 1759 375 1793 409
rect 1759 307 1793 341
rect 1853 443 1887 477
rect 1853 375 1887 409
rect 1947 443 1981 477
rect 1947 375 1981 409
rect 1947 307 1981 341
<< poly >>
rect 85 497 121 523
rect 179 497 215 523
rect 385 497 421 523
rect 479 497 515 523
rect 573 497 609 523
rect 667 497 703 523
rect 761 497 797 523
rect 855 497 891 523
rect 949 497 985 523
rect 1043 497 1079 523
rect 1241 497 1277 523
rect 1335 497 1371 523
rect 1429 497 1465 523
rect 1523 497 1559 523
rect 1617 497 1653 523
rect 1711 497 1747 523
rect 1805 497 1841 523
rect 1899 497 1935 523
rect 85 282 121 297
rect 179 282 215 297
rect 385 282 421 297
rect 479 282 515 297
rect 573 282 609 297
rect 667 282 703 297
rect 761 282 797 297
rect 855 282 891 297
rect 949 282 985 297
rect 1043 282 1079 297
rect 1241 282 1277 297
rect 1335 282 1371 297
rect 1429 282 1465 297
rect 1523 282 1559 297
rect 1617 282 1653 297
rect 1711 282 1747 297
rect 1805 282 1841 297
rect 1899 282 1935 297
rect 83 265 123 282
rect 29 249 123 265
rect 29 215 39 249
rect 73 215 123 249
rect 29 199 123 215
rect 93 177 123 199
rect 177 265 217 282
rect 383 265 423 282
rect 477 265 517 282
rect 571 265 611 282
rect 665 265 705 282
rect 177 249 277 265
rect 177 215 227 249
rect 261 215 277 249
rect 177 199 277 215
rect 383 249 705 265
rect 383 215 403 249
rect 437 215 481 249
rect 515 215 559 249
rect 593 215 705 249
rect 383 199 705 215
rect 177 177 207 199
rect 383 177 413 199
rect 477 177 507 199
rect 571 177 601 199
rect 675 177 705 199
rect 759 265 799 282
rect 853 265 893 282
rect 947 265 987 282
rect 1041 265 1081 282
rect 759 249 1081 265
rect 759 215 787 249
rect 821 215 865 249
rect 899 215 943 249
rect 977 215 1021 249
rect 1055 215 1081 249
rect 759 199 1081 215
rect 759 177 789 199
rect 853 177 883 199
rect 947 177 977 199
rect 1051 177 1081 199
rect 1239 265 1279 282
rect 1333 265 1373 282
rect 1427 265 1467 282
rect 1521 265 1561 282
rect 1239 249 1561 265
rect 1239 215 1267 249
rect 1301 215 1345 249
rect 1379 215 1423 249
rect 1457 215 1501 249
rect 1535 215 1561 249
rect 1239 199 1561 215
rect 1239 177 1269 199
rect 1333 177 1363 199
rect 1427 177 1457 199
rect 1531 177 1561 199
rect 1615 265 1655 282
rect 1709 265 1749 282
rect 1803 265 1843 282
rect 1897 265 1937 282
rect 1615 249 1937 265
rect 1615 215 1643 249
rect 1677 215 1721 249
rect 1755 215 1799 249
rect 1833 215 1877 249
rect 1911 215 1937 249
rect 1615 199 1937 215
rect 1615 177 1645 199
rect 1709 177 1739 199
rect 1803 177 1833 199
rect 1907 177 1937 199
rect 93 21 123 47
rect 177 21 207 47
rect 383 21 413 47
rect 477 21 507 47
rect 571 21 601 47
rect 675 21 705 47
rect 759 21 789 47
rect 853 21 883 47
rect 947 21 977 47
rect 1051 21 1081 47
rect 1239 21 1269 47
rect 1333 21 1363 47
rect 1427 21 1457 47
rect 1531 21 1561 47
rect 1615 21 1645 47
rect 1709 21 1739 47
rect 1803 21 1833 47
rect 1907 21 1937 47
<< polycont >>
rect 39 215 73 249
rect 227 215 261 249
rect 403 215 437 249
rect 481 215 515 249
rect 559 215 593 249
rect 787 215 821 249
rect 865 215 899 249
rect 943 215 977 249
rect 1021 215 1055 249
rect 1267 215 1301 249
rect 1345 215 1379 249
rect 1423 215 1457 249
rect 1501 215 1535 249
rect 1643 215 1677 249
rect 1721 215 1755 249
rect 1799 215 1833 249
rect 1877 215 1911 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 17 477 73 493
rect 17 443 39 477
rect 107 477 183 527
rect 107 443 133 477
rect 167 443 183 477
rect 323 477 1139 493
rect 323 443 339 477
rect 373 443 527 477
rect 561 443 715 477
rect 749 459 903 477
rect 749 443 765 459
rect 895 443 903 459
rect 937 459 1091 477
rect 937 443 945 459
rect 17 409 73 443
rect 809 409 851 425
rect 17 375 39 409
rect 73 375 765 409
rect 17 341 167 375
rect 17 307 39 341
rect 73 307 167 341
rect 201 307 227 341
rect 261 307 347 341
rect 22 249 89 273
rect 22 215 39 249
rect 73 215 89 249
rect 133 179 167 307
rect 201 249 279 265
rect 201 215 227 249
rect 261 215 279 249
rect 313 249 347 307
rect 388 307 433 341
rect 467 307 621 341
rect 655 307 687 341
rect 388 283 687 307
rect 313 215 403 249
rect 437 215 481 249
rect 515 215 559 249
rect 593 215 619 249
rect 313 181 347 215
rect 653 181 687 283
rect 731 257 765 375
rect 843 375 851 409
rect 809 341 851 375
rect 895 409 945 443
rect 1083 443 1091 459
rect 1125 443 1139 477
rect 895 375 903 409
rect 937 375 945 409
rect 895 359 945 375
rect 989 409 1039 425
rect 989 375 997 409
rect 1031 375 1039 409
rect 843 325 851 341
rect 989 341 1039 375
rect 1083 409 1139 443
rect 1083 375 1091 409
rect 1125 375 1139 409
rect 1083 359 1139 375
rect 1176 477 1613 493
rect 1176 443 1195 477
rect 1229 459 1383 477
rect 1229 443 1237 459
rect 1176 409 1237 443
rect 1375 443 1383 459
rect 1417 459 1571 477
rect 1417 443 1425 459
rect 1176 375 1195 409
rect 1229 375 1237 409
rect 1176 359 1237 375
rect 1281 409 1331 425
rect 1281 375 1289 409
rect 1323 375 1331 409
rect 989 325 997 341
rect 843 307 997 325
rect 1031 325 1039 341
rect 1281 341 1331 375
rect 1375 409 1425 443
rect 1563 443 1571 459
rect 1605 443 1613 477
rect 1375 375 1383 409
rect 1417 375 1425 409
rect 1375 359 1425 375
rect 1469 409 1519 425
rect 1469 375 1477 409
rect 1511 375 1519 409
rect 1281 325 1289 341
rect 1031 307 1289 325
rect 1323 325 1331 341
rect 1469 341 1519 375
rect 1469 325 1477 341
rect 1323 307 1477 325
rect 1511 307 1519 341
rect 809 291 1519 307
rect 1563 409 1613 443
rect 1563 375 1571 409
rect 1605 375 1613 409
rect 1563 341 1613 375
rect 1657 477 1707 527
rect 1657 443 1665 477
rect 1699 443 1707 477
rect 1657 409 1707 443
rect 1657 375 1665 409
rect 1699 375 1707 409
rect 1657 359 1707 375
rect 1751 477 1801 493
rect 1751 443 1759 477
rect 1793 443 1801 477
rect 1751 409 1801 443
rect 1751 375 1759 409
rect 1793 375 1801 409
rect 1563 307 1571 341
rect 1605 325 1613 341
rect 1751 341 1801 375
rect 1845 477 1895 527
rect 1845 443 1853 477
rect 1887 443 1895 477
rect 1845 409 1895 443
rect 1845 375 1853 409
rect 1887 375 1895 409
rect 1845 359 1895 375
rect 1939 477 2002 493
rect 1939 443 1947 477
rect 1981 443 2002 477
rect 1939 409 2002 443
rect 1939 375 1947 409
rect 1981 375 2002 409
rect 1751 325 1759 341
rect 1605 307 1759 325
rect 1793 325 1801 341
rect 1939 341 2002 375
rect 1939 325 1947 341
rect 1793 307 1947 325
rect 1981 307 2002 341
rect 1563 291 2002 307
rect 731 249 1081 257
rect 731 215 787 249
rect 821 215 865 249
rect 899 215 943 249
rect 977 215 1021 249
rect 1055 215 1081 249
rect 1130 249 1561 257
rect 1130 215 1267 249
rect 1301 215 1345 249
rect 1379 215 1423 249
rect 1457 215 1501 249
rect 1535 215 1561 249
rect 1615 249 2002 257
rect 1615 215 1643 249
rect 1677 215 1721 249
rect 1755 215 1799 249
rect 1833 215 1877 249
rect 1911 215 2002 249
rect 17 163 167 179
rect 17 129 39 163
rect 73 145 167 163
rect 201 163 347 181
rect 73 129 89 145
rect 17 95 89 129
rect 201 129 227 163
rect 261 147 347 163
rect 407 163 1903 181
rect 261 129 277 147
rect 17 61 39 95
rect 73 61 89 95
rect 17 51 89 61
rect 133 95 167 111
rect 133 17 167 61
rect 201 95 277 129
rect 407 129 433 163
rect 467 145 621 163
rect 467 129 483 145
rect 201 61 227 95
rect 261 61 277 95
rect 201 51 277 61
rect 339 95 373 111
rect 339 17 373 61
rect 407 95 483 129
rect 595 129 621 145
rect 655 145 809 163
rect 655 129 671 145
rect 407 61 433 95
rect 467 61 483 95
rect 407 51 483 61
rect 527 95 561 111
rect 527 17 561 61
rect 595 95 671 129
rect 783 129 809 145
rect 843 145 997 163
rect 843 129 859 145
rect 595 61 621 95
rect 655 61 671 95
rect 595 51 671 61
rect 715 95 749 111
rect 715 17 749 61
rect 783 95 859 129
rect 971 129 997 145
rect 1031 145 1289 163
rect 1031 129 1047 145
rect 783 61 809 95
rect 843 61 859 95
rect 783 51 859 61
rect 903 95 937 111
rect 903 17 937 61
rect 971 95 1047 129
rect 1263 129 1289 145
rect 1323 145 1477 163
rect 1323 129 1339 145
rect 971 61 997 95
rect 1031 61 1047 95
rect 971 51 1047 61
rect 1091 95 1229 111
rect 1125 61 1195 95
rect 1091 17 1229 61
rect 1263 95 1339 129
rect 1451 129 1477 145
rect 1511 145 1665 163
rect 1511 129 1527 145
rect 1263 61 1289 95
rect 1323 61 1339 95
rect 1263 51 1339 61
rect 1383 95 1417 111
rect 1383 17 1417 61
rect 1451 95 1527 129
rect 1639 129 1665 145
rect 1699 145 1853 163
rect 1699 129 1715 145
rect 1451 61 1477 95
rect 1511 61 1527 95
rect 1451 51 1527 61
rect 1571 95 1605 111
rect 1571 17 1605 61
rect 1639 95 1715 129
rect 1827 129 1853 145
rect 1887 129 1903 163
rect 1639 61 1665 95
rect 1699 61 1715 95
rect 1639 51 1715 61
rect 1759 95 1793 111
rect 1759 17 1793 61
rect 1827 95 1903 129
rect 1827 61 1853 95
rect 1887 61 1903 95
rect 1827 51 1903 61
rect 1947 163 2002 181
rect 1981 129 2002 163
rect 1947 95 2002 129
rect 1981 61 2002 95
rect 1947 17 2002 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 215 221 249 255 0 FreeSans 400 180 0 0 D_N
port 4 nsew signal input
flabel locali s 582 289 616 323 0 FreeSans 400 180 0 0 Y
port 9 nsew signal output
flabel locali s 1615 215 2002 257 0 FreeSans 400 180 0 0 A
port 1 nsew signal input
flabel locali s 1130 215 1561 257 0 FreeSans 400 180 0 0 B
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4bb_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2024 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1516110
string GDS_START 1501766
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
