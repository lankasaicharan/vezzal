magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 3506 1975
<< nwell >>
rect -38 388 2246 704
rect -38 332 740 388
rect 1041 332 2246 388
<< pwell >>
rect 232 248 342 286
rect 1 229 342 248
rect 889 238 999 312
rect 1421 248 1812 252
rect 1421 238 2207 248
rect 1 212 698 229
rect 889 212 2207 238
rect 1 49 2207 212
rect 0 0 2208 49
<< scpmos >>
rect 86 368 116 592
rect 176 368 206 592
rect 421 503 451 587
rect 528 445 558 529
rect 672 445 702 529
rect 756 445 786 529
rect 880 424 910 592
rect 970 424 1000 592
rect 1178 479 1208 563
rect 1293 479 1323 563
rect 1405 424 1435 592
rect 1495 424 1525 592
rect 1602 368 1632 592
rect 1692 368 1722 592
rect 1894 368 1924 568
rect 2001 368 2031 592
rect 2091 368 2121 592
<< nmoslvt >>
rect 84 74 114 222
rect 213 74 243 222
rect 499 119 529 203
rect 585 119 615 203
rect 687 102 717 186
rect 765 102 795 186
rect 870 76 900 186
rect 988 76 1018 186
rect 1218 128 1248 212
rect 1290 128 1320 212
rect 1504 78 1534 226
rect 1599 78 1629 226
rect 1685 78 1715 226
rect 1897 94 1927 222
rect 2008 74 2038 222
rect 2094 74 2124 222
<< ndiff >>
rect 258 248 316 260
rect 258 222 270 248
rect 27 202 84 222
rect 27 168 39 202
rect 73 168 84 202
rect 27 120 84 168
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 96 213 222
rect 114 74 146 96
rect 129 62 146 74
rect 180 74 213 96
rect 243 214 270 222
rect 304 214 316 248
rect 243 74 316 214
rect 180 62 198 74
rect 129 50 198 62
rect 376 119 499 203
rect 529 180 585 203
rect 529 146 540 180
rect 574 146 585 180
rect 529 119 585 146
rect 615 186 672 203
rect 915 274 973 286
rect 915 240 927 274
rect 961 240 973 274
rect 915 186 973 240
rect 1447 214 1504 226
rect 1161 186 1218 212
rect 615 180 687 186
rect 615 146 626 180
rect 660 146 687 180
rect 615 119 687 146
rect 376 112 450 119
rect 376 78 388 112
rect 422 78 450 112
rect 637 102 687 119
rect 717 102 765 186
rect 795 122 870 186
rect 795 102 823 122
rect 376 66 450 78
rect 810 88 823 102
rect 857 88 870 122
rect 810 76 870 88
rect 900 76 988 186
rect 1018 174 1218 186
rect 1018 140 1173 174
rect 1207 140 1218 174
rect 1018 128 1218 140
rect 1248 128 1290 212
rect 1320 179 1393 212
rect 1320 145 1347 179
rect 1381 145 1393 179
rect 1320 128 1393 145
rect 1447 180 1459 214
rect 1493 180 1504 214
rect 1018 76 1068 128
rect 1447 124 1504 180
rect 1447 90 1459 124
rect 1493 90 1504 124
rect 1447 78 1504 90
rect 1534 214 1599 226
rect 1534 180 1545 214
rect 1579 180 1599 214
rect 1534 124 1599 180
rect 1534 90 1545 124
rect 1579 90 1599 124
rect 1534 78 1599 90
rect 1629 214 1685 226
rect 1629 180 1640 214
rect 1674 180 1685 214
rect 1629 124 1685 180
rect 1629 90 1640 124
rect 1674 90 1685 124
rect 1629 78 1685 90
rect 1715 214 1786 226
rect 1715 180 1740 214
rect 1774 180 1786 214
rect 1715 124 1786 180
rect 1715 90 1740 124
rect 1774 90 1786 124
rect 1840 184 1897 222
rect 1840 150 1852 184
rect 1886 150 1897 184
rect 1840 94 1897 150
rect 1927 210 2008 222
rect 1927 176 1963 210
rect 1997 176 2008 210
rect 1927 120 2008 176
rect 1927 94 1963 120
rect 1715 78 1786 90
rect 1951 86 1963 94
rect 1997 86 2008 120
rect 1951 74 2008 86
rect 2038 210 2094 222
rect 2038 176 2049 210
rect 2083 176 2094 210
rect 2038 120 2094 176
rect 2038 86 2049 120
rect 2083 86 2094 120
rect 2038 74 2094 86
rect 2124 210 2181 222
rect 2124 176 2135 210
rect 2169 176 2181 210
rect 2124 120 2181 176
rect 2124 86 2135 120
rect 2169 86 2181 120
rect 2124 74 2181 86
<< pdiff >>
rect 319 627 403 639
rect 319 593 344 627
rect 378 593 403 627
rect 804 627 862 639
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 462 176 546
rect 116 428 129 462
rect 163 428 176 462
rect 116 368 176 428
rect 206 580 265 592
rect 206 546 219 580
rect 253 546 265 580
rect 206 497 265 546
rect 319 587 403 593
rect 804 593 816 627
rect 850 593 862 627
rect 804 592 862 593
rect 319 503 421 587
rect 451 529 504 587
rect 804 529 880 592
rect 451 503 528 529
rect 206 463 219 497
rect 253 463 265 497
rect 469 491 528 503
rect 206 414 265 463
rect 206 380 219 414
rect 253 380 265 414
rect 469 457 481 491
rect 515 457 528 491
rect 469 445 528 457
rect 558 491 672 529
rect 558 457 600 491
rect 634 457 672 491
rect 558 445 672 457
rect 702 445 756 529
rect 786 445 880 529
rect 206 368 265 380
rect 827 424 880 445
rect 910 472 970 592
rect 910 438 923 472
rect 957 438 970 472
rect 910 424 970 438
rect 1000 563 1053 592
rect 1352 563 1405 592
rect 1000 525 1178 563
rect 1000 491 1091 525
rect 1125 491 1178 525
rect 1000 479 1178 491
rect 1208 479 1293 563
rect 1323 538 1405 563
rect 1323 504 1336 538
rect 1370 504 1405 538
rect 1323 479 1405 504
rect 1000 424 1053 479
rect 1352 424 1405 479
rect 1435 580 1495 592
rect 1435 546 1448 580
rect 1482 546 1495 580
rect 1435 476 1495 546
rect 1435 442 1448 476
rect 1482 442 1495 476
rect 1435 424 1495 442
rect 1525 573 1602 592
rect 1525 539 1555 573
rect 1589 539 1602 573
rect 1525 424 1602 539
rect 1549 368 1602 424
rect 1632 414 1692 592
rect 1632 380 1645 414
rect 1679 380 1692 414
rect 1632 368 1692 380
rect 1722 573 1781 592
rect 1722 539 1735 573
rect 1769 539 1781 573
rect 1942 580 2001 592
rect 1942 568 1954 580
rect 1722 368 1781 539
rect 1835 556 1894 568
rect 1835 522 1847 556
rect 1881 522 1894 556
rect 1835 485 1894 522
rect 1835 451 1847 485
rect 1881 451 1894 485
rect 1835 414 1894 451
rect 1835 380 1847 414
rect 1881 380 1894 414
rect 1835 368 1894 380
rect 1924 546 1954 568
rect 1988 546 2001 580
rect 1924 497 2001 546
rect 1924 463 1954 497
rect 1988 463 2001 497
rect 1924 414 2001 463
rect 1924 380 1954 414
rect 1988 380 2001 414
rect 1924 368 2001 380
rect 2031 580 2091 592
rect 2031 546 2044 580
rect 2078 546 2091 580
rect 2031 497 2091 546
rect 2031 463 2044 497
rect 2078 463 2091 497
rect 2031 414 2091 463
rect 2031 380 2044 414
rect 2078 380 2091 414
rect 2031 368 2091 380
rect 2121 580 2181 592
rect 2121 546 2135 580
rect 2169 546 2181 580
rect 2121 497 2181 546
rect 2121 463 2135 497
rect 2169 463 2181 497
rect 2121 414 2181 463
rect 2121 380 2135 414
rect 2169 380 2181 414
rect 2121 368 2181 380
<< ndiffc >>
rect 39 168 73 202
rect 39 86 73 120
rect 146 62 180 96
rect 270 214 304 248
rect 540 146 574 180
rect 927 240 961 274
rect 626 146 660 180
rect 388 78 422 112
rect 823 88 857 122
rect 1173 140 1207 174
rect 1347 145 1381 179
rect 1459 180 1493 214
rect 1459 90 1493 124
rect 1545 180 1579 214
rect 1545 90 1579 124
rect 1640 180 1674 214
rect 1640 90 1674 124
rect 1740 180 1774 214
rect 1740 90 1774 124
rect 1852 150 1886 184
rect 1963 176 1997 210
rect 1963 86 1997 120
rect 2049 176 2083 210
rect 2049 86 2083 120
rect 2135 176 2169 210
rect 2135 86 2169 120
<< pdiffc >>
rect 344 593 378 627
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 428 163 462
rect 219 546 253 580
rect 816 593 850 627
rect 219 463 253 497
rect 219 380 253 414
rect 481 457 515 491
rect 600 457 634 491
rect 923 438 957 472
rect 1091 491 1125 525
rect 1336 504 1370 538
rect 1448 546 1482 580
rect 1448 442 1482 476
rect 1555 539 1589 573
rect 1645 380 1679 414
rect 1735 539 1769 573
rect 1847 522 1881 556
rect 1847 451 1881 485
rect 1847 380 1881 414
rect 1954 546 1988 580
rect 1954 463 1988 497
rect 1954 380 1988 414
rect 2044 546 2078 580
rect 2044 463 2078 497
rect 2044 380 2078 414
rect 2135 546 2169 580
rect 2135 463 2169 497
rect 2135 380 2169 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 421 587 451 613
rect 880 592 910 618
rect 970 592 1000 618
rect 1405 592 1435 618
rect 1495 592 1525 618
rect 1602 592 1632 618
rect 1692 592 1722 618
rect 528 529 558 555
rect 672 529 702 555
rect 756 529 786 555
rect 421 488 451 503
rect 418 471 454 488
rect 365 455 454 471
rect 365 421 381 455
rect 415 421 454 455
rect 528 430 558 445
rect 672 430 702 445
rect 756 430 786 445
rect 365 405 454 421
rect 86 353 116 368
rect 176 353 206 368
rect 525 363 561 430
rect 669 413 705 430
rect 83 310 119 353
rect 173 310 209 353
rect 297 347 561 363
rect 297 313 313 347
rect 347 333 561 347
rect 609 397 711 413
rect 609 363 661 397
rect 695 363 711 397
rect 609 347 711 363
rect 347 313 363 333
rect 51 294 119 310
rect 51 260 67 294
rect 101 260 119 294
rect 51 244 119 260
rect 161 294 243 310
rect 297 297 363 313
rect 161 260 177 294
rect 211 260 243 294
rect 161 244 243 260
rect 84 222 114 244
rect 213 222 243 244
rect 84 48 114 74
rect 213 48 243 74
rect 331 51 361 297
rect 409 275 475 291
rect 409 241 425 275
rect 459 255 475 275
rect 459 241 529 255
rect 609 248 639 347
rect 753 284 789 430
rect 1178 563 1208 589
rect 1293 563 1323 589
rect 1178 464 1208 479
rect 1293 464 1323 479
rect 1175 447 1211 464
rect 1175 431 1241 447
rect 880 409 910 424
rect 970 409 1000 424
rect 877 392 913 409
rect 831 376 913 392
rect 831 342 847 376
rect 881 342 913 376
rect 831 326 913 342
rect 967 368 1003 409
rect 1175 397 1191 431
rect 1225 397 1241 431
rect 1175 381 1241 397
rect 967 338 1133 368
rect 409 225 529 241
rect 499 203 529 225
rect 585 218 639 248
rect 759 268 828 284
rect 759 234 778 268
rect 812 234 828 268
rect 759 218 828 234
rect 585 203 615 218
rect 687 186 717 212
rect 765 186 795 218
rect 870 186 900 326
rect 1103 300 1133 338
rect 1290 348 1326 464
rect 1405 409 1435 424
rect 1495 409 1525 424
rect 1402 392 1438 409
rect 1492 392 1528 409
rect 1402 376 1534 392
rect 1402 362 1467 376
rect 1290 300 1320 348
rect 1451 342 1467 362
rect 1501 342 1534 376
rect 1894 568 1924 594
rect 2001 592 2031 618
rect 2091 592 2121 618
rect 1602 353 1632 368
rect 1692 353 1722 368
rect 1894 353 1924 368
rect 2001 353 2031 368
rect 2091 353 2121 368
rect 1451 326 1534 342
rect 988 274 1061 290
rect 988 240 1011 274
rect 1045 240 1061 274
rect 988 224 1061 240
rect 1103 284 1169 300
rect 1103 250 1119 284
rect 1153 264 1169 284
rect 1290 284 1409 300
rect 1153 250 1248 264
rect 1103 234 1248 250
rect 988 186 1018 224
rect 1218 212 1248 234
rect 1290 250 1359 284
rect 1393 250 1409 284
rect 1290 234 1409 250
rect 1290 212 1320 234
rect 1504 226 1534 326
rect 1599 294 1635 353
rect 1689 330 1725 353
rect 1891 330 1927 353
rect 1685 314 1927 330
rect 1998 326 2034 353
rect 2088 326 2124 353
rect 1685 294 1753 314
rect 1599 280 1753 294
rect 1787 280 1927 314
rect 1599 264 1927 280
rect 1599 226 1629 264
rect 1685 226 1715 264
rect 499 93 529 119
rect 585 93 615 119
rect 687 51 717 102
rect 765 76 795 102
rect 1218 106 1248 128
rect 1114 90 1248 106
rect 1290 102 1320 128
rect 331 21 717 51
rect 870 50 900 76
rect 988 50 1018 76
rect 1114 56 1130 90
rect 1164 56 1198 90
rect 1232 56 1248 90
rect 1897 222 1927 264
rect 1969 310 2124 326
rect 1969 276 1985 310
rect 2019 276 2124 310
rect 1969 260 2124 276
rect 2008 222 2038 260
rect 2094 222 2124 260
rect 1114 40 1248 56
rect 1504 52 1534 78
rect 1599 52 1629 78
rect 1685 52 1715 78
rect 1897 68 1927 94
rect 2008 48 2038 74
rect 2094 48 2124 74
<< polycont >>
rect 381 421 415 455
rect 313 313 347 347
rect 661 363 695 397
rect 67 260 101 294
rect 177 260 211 294
rect 425 241 459 275
rect 847 342 881 376
rect 1191 397 1225 431
rect 778 234 812 268
rect 1467 342 1501 376
rect 1011 240 1045 274
rect 1119 250 1153 284
rect 1359 250 1393 284
rect 1753 280 1787 314
rect 1130 56 1164 90
rect 1198 56 1232 90
rect 1985 276 2019 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 497 89 546
rect 23 463 39 497
rect 73 463 89 497
rect 23 414 89 463
rect 23 380 39 414
rect 73 380 89 414
rect 129 580 179 649
rect 315 627 407 649
rect 163 546 179 580
rect 129 462 179 546
rect 163 428 179 462
rect 129 412 179 428
rect 219 580 269 596
rect 315 593 344 627
rect 378 593 407 627
rect 800 627 866 649
rect 800 593 816 627
rect 850 593 866 627
rect 253 559 269 580
rect 1007 559 1241 593
rect 253 546 1041 559
rect 219 525 1041 546
rect 219 497 288 525
rect 253 463 288 497
rect 219 414 288 463
rect 23 378 89 380
rect 253 380 288 414
rect 365 455 431 471
rect 365 421 381 455
rect 415 421 431 455
rect 465 457 481 491
rect 515 457 543 491
rect 465 441 543 457
rect 365 405 431 421
rect 23 344 185 378
rect 219 363 288 380
rect 151 310 185 344
rect 254 347 363 363
rect 254 313 313 347
rect 347 313 363 347
rect 25 294 117 310
rect 25 260 67 294
rect 101 260 117 294
rect 25 236 117 260
rect 151 294 220 310
rect 151 260 177 294
rect 211 260 220 294
rect 151 202 220 260
rect 254 297 363 313
rect 397 356 431 405
rect 254 248 320 297
rect 254 214 270 248
rect 304 214 320 248
rect 397 275 475 356
rect 397 241 425 275
rect 459 241 475 275
rect 397 225 475 241
rect 509 248 543 441
rect 577 457 600 491
rect 634 457 865 491
rect 577 316 611 457
rect 645 397 728 413
rect 645 363 661 397
rect 695 363 728 397
rect 645 350 728 363
rect 577 282 660 316
rect 509 214 574 248
rect 23 168 39 202
rect 73 180 220 202
rect 540 180 574 214
rect 73 168 506 180
rect 23 146 506 168
rect 23 120 89 146
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 125 96 202 112
rect 125 62 146 96
rect 180 62 202 96
rect 125 17 202 62
rect 372 78 388 112
rect 422 78 438 112
rect 372 17 438 78
rect 472 85 506 146
rect 540 119 574 146
rect 610 180 660 282
rect 610 146 626 180
rect 610 119 660 146
rect 694 190 728 350
rect 831 392 865 457
rect 907 472 973 491
rect 907 438 923 472
rect 957 438 973 472
rect 907 436 973 438
rect 831 376 895 392
rect 831 342 847 376
rect 881 342 895 376
rect 831 326 895 342
rect 929 290 963 436
rect 1007 290 1041 525
rect 1075 491 1091 525
rect 1125 491 1141 525
rect 1075 358 1141 491
rect 1175 431 1241 559
rect 1320 538 1386 649
rect 1320 504 1336 538
rect 1370 504 1386 538
rect 1320 475 1386 504
rect 1432 580 1498 596
rect 1432 546 1448 580
rect 1482 546 1498 580
rect 1432 482 1498 546
rect 1539 573 1605 649
rect 1539 539 1555 573
rect 1589 539 1605 573
rect 1539 516 1605 539
rect 1719 573 1785 649
rect 1719 539 1735 573
rect 1769 539 1785 573
rect 1938 580 1988 649
rect 1719 516 1785 539
rect 1847 556 1897 572
rect 1881 522 1897 556
rect 1847 485 1897 522
rect 1432 476 1803 482
rect 1175 397 1191 431
rect 1225 397 1241 431
rect 1432 442 1448 476
rect 1482 448 1803 476
rect 1482 442 1585 448
rect 1432 426 1585 442
rect 1175 392 1241 397
rect 1275 376 1517 392
rect 1275 358 1467 376
rect 1075 342 1467 358
rect 1501 342 1517 376
rect 1075 334 1517 342
rect 1075 324 1309 334
rect 762 274 963 290
rect 762 268 927 274
rect 762 234 778 268
rect 812 240 927 268
rect 961 240 963 274
rect 812 234 963 240
rect 762 224 963 234
rect 997 274 1055 290
rect 997 240 1011 274
rect 1045 240 1055 274
rect 997 224 1055 240
rect 1089 284 1169 290
rect 1089 250 1119 284
rect 1153 250 1169 284
rect 1089 234 1169 250
rect 694 156 963 190
rect 694 85 728 156
rect 472 51 728 85
rect 806 88 823 122
rect 857 88 874 122
rect 806 17 874 88
rect 929 106 963 156
rect 1089 106 1123 234
rect 1203 190 1237 324
rect 1551 300 1585 426
rect 1343 284 1585 300
rect 1343 250 1359 284
rect 1393 266 1585 284
rect 1629 380 1645 414
rect 1679 380 1703 414
rect 1629 310 1703 380
rect 1737 314 1803 448
rect 1393 250 1493 266
rect 1343 234 1493 250
rect 1443 214 1493 234
rect 1157 174 1237 190
rect 1157 140 1173 174
rect 1207 140 1237 174
rect 1331 179 1397 200
rect 1331 145 1347 179
rect 1381 145 1397 179
rect 929 90 1248 106
rect 929 56 1130 90
rect 1164 56 1198 90
rect 1232 56 1248 90
rect 929 51 1248 56
rect 1331 17 1397 145
rect 1443 180 1459 214
rect 1443 124 1493 180
rect 1443 90 1459 124
rect 1443 74 1493 90
rect 1529 214 1595 230
rect 1529 180 1545 214
rect 1579 180 1595 214
rect 1529 124 1595 180
rect 1529 90 1545 124
rect 1579 90 1595 124
rect 1529 17 1595 90
rect 1629 214 1690 310
rect 1737 280 1753 314
rect 1787 280 1803 314
rect 1737 264 1803 280
rect 1881 451 1897 485
rect 1847 414 1897 451
rect 1881 380 1897 414
rect 1847 326 1897 380
rect 1938 546 1954 580
rect 1938 497 1988 546
rect 1938 463 1954 497
rect 1938 414 1988 463
rect 1938 380 1954 414
rect 1938 364 1988 380
rect 2028 580 2101 596
rect 2028 546 2044 580
rect 2078 546 2101 580
rect 2028 497 2101 546
rect 2028 463 2044 497
rect 2078 463 2101 497
rect 2028 414 2101 463
rect 2028 380 2044 414
rect 2078 380 2101 414
rect 2028 364 2101 380
rect 2135 580 2185 649
rect 2169 546 2185 580
rect 2135 497 2185 546
rect 2169 463 2185 497
rect 2135 414 2185 463
rect 2169 380 2185 414
rect 2135 364 2185 380
rect 1847 310 2033 326
rect 1847 276 1985 310
rect 2019 276 2033 310
rect 1847 260 2033 276
rect 1629 180 1640 214
rect 1674 180 1690 214
rect 1629 124 1690 180
rect 1629 90 1640 124
rect 1674 90 1690 124
rect 1629 74 1690 90
rect 1724 214 1790 230
rect 1724 180 1740 214
rect 1774 180 1790 214
rect 1724 124 1790 180
rect 1724 90 1740 124
rect 1774 90 1790 124
rect 1847 184 1902 260
rect 2067 226 2101 364
rect 1847 150 1852 184
rect 1886 150 1902 184
rect 1847 90 1902 150
rect 1947 210 1997 226
rect 1947 176 1963 210
rect 1947 120 1997 176
rect 1724 17 1790 90
rect 1947 86 1963 120
rect 1947 17 1997 86
rect 2033 210 2101 226
rect 2033 176 2049 210
rect 2083 176 2101 210
rect 2033 120 2101 176
rect 2033 86 2049 120
rect 2083 86 2101 120
rect 2033 70 2101 86
rect 2135 210 2185 226
rect 2169 176 2185 210
rect 2135 120 2185 176
rect 2169 86 2185 120
rect 2135 17 2185 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfxbp_2
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2047 464 2081 498 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 2047 538 2081 572 0 FreeSans 340 0 0 0 Q_N
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 1471318
string GDS_START 1455038
<< end >>
