magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 464 232 652 251
rect 464 157 843 232
rect 1 49 843 157
rect 0 0 864 49
<< scnmos >>
rect 84 47 114 131
rect 156 47 186 131
rect 242 47 272 131
rect 328 47 358 131
rect 546 141 576 225
rect 648 122 678 206
rect 734 122 764 206
<< scpmoshvt >>
rect 93 419 143 619
rect 220 419 270 619
rect 318 419 368 619
rect 432 419 482 619
rect 530 419 580 619
rect 636 419 686 619
<< ndiff >>
rect 27 111 84 131
rect 27 77 39 111
rect 73 77 84 111
rect 27 47 84 77
rect 114 47 156 131
rect 186 106 242 131
rect 186 72 197 106
rect 231 72 242 106
rect 186 47 242 72
rect 272 111 328 131
rect 272 77 283 111
rect 317 77 328 111
rect 272 47 328 77
rect 358 73 430 131
rect 490 213 546 225
rect 490 179 501 213
rect 535 179 546 213
rect 490 141 546 179
rect 576 206 626 225
rect 576 164 648 206
rect 576 141 603 164
rect 591 130 603 141
rect 637 130 648 164
rect 591 122 648 130
rect 678 187 734 206
rect 678 153 689 187
rect 723 153 734 187
rect 678 122 734 153
rect 764 187 817 206
rect 764 153 775 187
rect 809 153 817 187
rect 764 122 817 153
rect 358 47 385 73
rect 373 39 385 47
rect 419 39 430 73
rect 373 27 430 39
<< pdiff >>
rect 36 597 93 619
rect 36 563 48 597
rect 82 563 93 597
rect 36 465 93 563
rect 36 431 48 465
rect 82 431 93 465
rect 36 419 93 431
rect 143 607 220 619
rect 143 573 154 607
rect 188 573 220 607
rect 143 514 220 573
rect 143 480 154 514
rect 188 480 220 514
rect 143 419 220 480
rect 270 419 318 619
rect 368 597 432 619
rect 368 563 379 597
rect 413 563 432 597
rect 368 465 432 563
rect 368 431 379 465
rect 413 431 432 465
rect 368 419 432 431
rect 482 419 530 619
rect 580 607 636 619
rect 580 573 591 607
rect 625 573 636 607
rect 580 514 636 573
rect 580 480 591 514
rect 625 480 636 514
rect 580 419 636 480
rect 686 597 743 619
rect 686 563 697 597
rect 731 563 743 597
rect 686 465 743 563
rect 686 431 697 465
rect 731 431 743 465
rect 686 419 743 431
<< ndiffc >>
rect 39 77 73 111
rect 197 72 231 106
rect 283 77 317 111
rect 501 179 535 213
rect 603 130 637 164
rect 689 153 723 187
rect 775 153 809 187
rect 385 39 419 73
<< pdiffc >>
rect 48 563 82 597
rect 48 431 82 465
rect 154 573 188 607
rect 154 480 188 514
rect 379 563 413 597
rect 379 431 413 465
rect 591 573 625 607
rect 591 480 625 514
rect 697 563 731 597
rect 697 431 731 465
<< poly >>
rect 93 619 143 645
rect 220 619 270 645
rect 318 619 368 645
rect 432 619 482 645
rect 530 619 580 645
rect 636 619 686 645
rect 93 379 143 419
rect 84 363 156 379
rect 84 329 106 363
rect 140 329 156 363
rect 220 358 270 419
rect 84 295 156 329
rect 84 261 106 295
rect 140 261 156 295
rect 84 245 156 261
rect 204 342 270 358
rect 204 308 220 342
rect 254 308 270 342
rect 204 274 270 308
rect 84 176 114 245
rect 204 240 220 274
rect 254 240 270 274
rect 204 224 270 240
rect 318 358 368 419
rect 318 342 384 358
rect 318 308 334 342
rect 368 308 384 342
rect 318 274 384 308
rect 432 345 482 419
rect 530 393 580 419
rect 432 329 498 345
rect 432 295 448 329
rect 482 295 498 329
rect 550 332 580 393
rect 636 404 686 419
rect 636 374 764 404
rect 734 332 764 374
rect 550 316 682 332
rect 550 302 632 316
rect 432 279 498 295
rect 616 282 632 302
rect 666 282 682 316
rect 318 240 334 274
rect 368 240 384 274
rect 318 224 384 240
rect 240 176 270 224
rect 84 146 186 176
rect 240 146 272 176
rect 84 131 114 146
rect 156 131 186 146
rect 242 131 272 146
rect 328 131 358 224
rect 445 126 475 279
rect 616 266 682 282
rect 724 316 790 332
rect 724 282 740 316
rect 774 282 790 316
rect 724 266 790 282
rect 546 225 576 251
rect 648 206 678 266
rect 734 206 764 266
rect 546 126 576 141
rect 445 96 576 126
rect 648 96 678 122
rect 734 96 764 122
rect 84 21 114 47
rect 156 21 186 47
rect 242 21 272 47
rect 328 21 358 47
<< polycont >>
rect 106 329 140 363
rect 106 261 140 295
rect 220 308 254 342
rect 220 240 254 274
rect 334 308 368 342
rect 448 295 482 329
rect 632 282 666 316
rect 334 240 368 274
rect 740 282 774 316
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 20 597 98 613
rect 20 563 48 597
rect 82 563 98 597
rect 20 465 98 563
rect 20 431 48 465
rect 82 431 98 465
rect 138 607 204 649
rect 138 573 154 607
rect 188 573 204 607
rect 138 514 204 573
rect 138 480 154 514
rect 188 480 204 514
rect 138 464 204 480
rect 363 597 429 613
rect 363 563 379 597
rect 413 563 429 597
rect 363 465 429 563
rect 20 415 98 431
rect 363 431 379 465
rect 413 431 429 465
rect 575 607 641 649
rect 575 573 591 607
rect 625 573 641 607
rect 575 514 641 573
rect 575 480 591 514
rect 625 480 641 514
rect 575 464 641 480
rect 681 597 847 613
rect 681 563 697 597
rect 731 563 847 597
rect 681 465 847 563
rect 363 428 429 431
rect 681 431 697 465
rect 731 431 847 465
rect 681 428 847 431
rect 20 208 54 415
rect 134 394 847 428
rect 134 379 168 394
rect 90 363 168 379
rect 90 329 106 363
rect 140 329 168 363
rect 90 295 168 329
rect 90 261 106 295
rect 140 261 168 295
rect 90 245 168 261
rect 204 342 270 358
rect 204 308 220 342
rect 254 308 270 342
rect 204 274 270 308
rect 204 240 220 274
rect 254 240 270 274
rect 204 224 270 240
rect 313 342 374 358
rect 313 308 334 342
rect 368 308 374 342
rect 313 274 374 308
rect 408 329 553 356
rect 408 295 448 329
rect 482 295 553 329
rect 408 279 553 295
rect 601 316 666 356
rect 601 282 632 316
rect 313 240 334 274
rect 368 240 374 274
rect 601 266 666 282
rect 700 316 779 358
rect 700 282 740 316
rect 774 282 779 316
rect 700 266 779 282
rect 313 224 374 240
rect 485 213 739 232
rect 20 111 89 208
rect 485 179 501 213
rect 535 198 739 213
rect 813 203 847 394
rect 535 179 551 198
rect 689 187 739 198
rect 587 143 603 164
rect 20 77 39 111
rect 73 77 89 111
rect 20 53 89 77
rect 181 106 231 135
rect 181 72 197 106
rect 181 17 231 72
rect 267 130 603 143
rect 637 130 653 164
rect 723 153 739 187
rect 689 137 739 153
rect 773 187 847 203
rect 773 153 775 187
rect 809 153 847 187
rect 773 137 847 153
rect 267 111 653 130
rect 267 77 283 111
rect 317 109 653 111
rect 317 77 333 109
rect 267 53 333 77
rect 369 39 385 73
rect 419 39 435 73
rect 369 17 435 39
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221a_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4801028
string GDS_START 4793146
<< end >>
