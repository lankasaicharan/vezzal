magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
rect 691 299 971 331
<< pwell >>
rect 963 241 1151 257
rect 762 235 1151 241
rect 335 159 1151 235
rect 29 49 1151 159
rect 0 0 1152 49
<< scnmos >>
rect 108 49 138 133
rect 194 49 224 133
rect 414 125 444 209
rect 500 125 530 209
rect 572 125 602 209
rect 661 125 691 209
rect 733 125 763 209
rect 841 47 871 215
rect 1042 63 1072 231
<< scpmoshvt >>
rect 80 425 110 553
rect 166 425 196 553
rect 370 461 400 589
rect 494 419 524 547
rect 566 419 596 547
rect 671 419 701 503
rect 743 419 773 503
rect 852 335 882 587
rect 1042 367 1072 619
<< ndiff >>
rect 55 105 108 133
rect 55 71 63 105
rect 97 71 108 105
rect 55 49 108 71
rect 138 105 194 133
rect 138 71 149 105
rect 183 71 194 105
rect 138 49 194 71
rect 224 105 277 133
rect 224 71 235 105
rect 269 71 277 105
rect 788 209 841 215
rect 361 185 414 209
rect 361 151 369 185
rect 403 151 414 185
rect 361 125 414 151
rect 444 167 500 209
rect 444 133 455 167
rect 489 133 500 167
rect 444 125 500 133
rect 530 125 572 209
rect 602 197 661 209
rect 602 163 616 197
rect 650 163 661 197
rect 602 125 661 163
rect 691 125 733 209
rect 763 125 841 209
rect 224 49 277 71
rect 788 117 841 125
rect 788 83 796 117
rect 830 83 841 117
rect 788 47 841 83
rect 871 109 924 215
rect 871 75 882 109
rect 916 75 924 109
rect 871 47 924 75
rect 989 203 1042 231
rect 989 169 997 203
rect 1031 169 1042 203
rect 989 109 1042 169
rect 989 75 997 109
rect 1031 75 1042 109
rect 989 63 1042 75
rect 1072 212 1125 231
rect 1072 178 1083 212
rect 1117 178 1125 212
rect 1072 109 1125 178
rect 1072 75 1083 109
rect 1117 75 1125 109
rect 1072 63 1125 75
<< pdiff >>
rect 27 539 80 553
rect 27 505 35 539
rect 69 505 80 539
rect 27 471 80 505
rect 27 437 35 471
rect 69 437 80 471
rect 27 425 80 437
rect 110 545 166 553
rect 110 511 121 545
rect 155 511 166 545
rect 110 477 166 511
rect 110 443 121 477
rect 155 443 166 477
rect 110 425 166 443
rect 196 539 249 553
rect 196 505 207 539
rect 241 505 249 539
rect 196 471 249 505
rect 196 437 207 471
rect 241 437 249 471
rect 196 425 249 437
rect 317 577 370 589
rect 317 543 325 577
rect 359 543 370 577
rect 317 507 370 543
rect 317 473 325 507
rect 359 473 370 507
rect 317 461 370 473
rect 400 567 472 589
rect 400 533 430 567
rect 464 547 472 567
rect 989 607 1042 619
rect 795 579 852 587
rect 464 533 494 547
rect 400 461 494 533
rect 422 419 494 461
rect 524 419 566 547
rect 596 533 649 547
rect 596 499 607 533
rect 641 503 649 533
rect 795 545 807 579
rect 841 545 852 579
rect 795 511 852 545
rect 795 503 807 511
rect 641 499 671 503
rect 596 465 671 499
rect 596 431 619 465
rect 653 431 671 465
rect 596 419 671 431
rect 701 419 743 503
rect 773 477 807 503
rect 841 477 852 511
rect 773 441 852 477
rect 773 419 807 441
rect 795 407 807 419
rect 841 407 852 441
rect 795 335 852 407
rect 882 574 935 587
rect 882 540 893 574
rect 927 540 935 574
rect 882 482 935 540
rect 882 448 893 482
rect 927 448 935 482
rect 882 389 935 448
rect 882 355 893 389
rect 927 355 935 389
rect 989 573 997 607
rect 1031 573 1042 607
rect 989 507 1042 573
rect 989 473 997 507
rect 1031 473 1042 507
rect 989 413 1042 473
rect 989 379 997 413
rect 1031 379 1042 413
rect 989 367 1042 379
rect 1072 599 1125 619
rect 1072 565 1083 599
rect 1117 565 1125 599
rect 1072 508 1125 565
rect 1072 474 1083 508
rect 1117 474 1125 508
rect 1072 413 1125 474
rect 1072 379 1083 413
rect 1117 379 1125 413
rect 1072 367 1125 379
rect 882 335 935 355
<< ndiffc >>
rect 63 71 97 105
rect 149 71 183 105
rect 235 71 269 105
rect 369 151 403 185
rect 455 133 489 167
rect 616 163 650 197
rect 796 83 830 117
rect 882 75 916 109
rect 997 169 1031 203
rect 997 75 1031 109
rect 1083 178 1117 212
rect 1083 75 1117 109
<< pdiffc >>
rect 35 505 69 539
rect 35 437 69 471
rect 121 511 155 545
rect 121 443 155 477
rect 207 505 241 539
rect 207 437 241 471
rect 325 543 359 577
rect 325 473 359 507
rect 430 533 464 567
rect 607 499 641 533
rect 807 545 841 579
rect 619 431 653 465
rect 807 477 841 511
rect 807 407 841 441
rect 893 540 927 574
rect 893 448 927 482
rect 893 355 927 389
rect 997 573 1031 607
rect 997 473 1031 507
rect 997 379 1031 413
rect 1083 565 1117 599
rect 1083 474 1117 508
rect 1083 379 1117 413
<< poly >>
rect 272 615 596 645
rect 1042 619 1072 645
rect 80 553 110 579
rect 166 553 196 579
rect 80 289 110 425
rect 166 367 196 425
rect 272 393 302 615
rect 370 589 400 615
rect 494 547 524 573
rect 566 547 596 615
rect 852 587 882 613
rect 370 435 400 461
rect 671 503 701 529
rect 743 503 773 529
rect 272 377 338 393
rect 166 337 224 367
rect 80 273 146 289
rect 80 239 96 273
rect 130 239 146 273
rect 80 205 146 239
rect 80 171 96 205
rect 130 171 146 205
rect 80 155 146 171
rect 194 221 224 337
rect 272 343 288 377
rect 322 343 338 377
rect 494 349 524 419
rect 566 393 596 419
rect 671 381 701 419
rect 272 327 338 343
rect 194 205 260 221
rect 194 171 210 205
rect 244 171 260 205
rect 194 155 260 171
rect 108 133 138 155
rect 194 133 224 155
rect 308 103 338 327
rect 444 333 524 349
rect 644 351 701 381
rect 644 345 674 351
rect 444 299 460 333
rect 494 313 524 333
rect 572 329 674 345
rect 494 299 530 313
rect 444 283 530 299
rect 414 209 444 235
rect 500 209 530 283
rect 572 295 588 329
rect 622 315 674 329
rect 622 295 638 315
rect 743 303 773 419
rect 852 303 882 335
rect 1042 319 1072 367
rect 993 303 1072 319
rect 572 279 638 295
rect 733 287 799 303
rect 572 209 602 279
rect 733 253 749 287
rect 783 253 799 287
rect 733 237 799 253
rect 841 287 907 303
rect 841 253 857 287
rect 891 253 907 287
rect 993 269 1009 303
rect 1043 269 1072 303
rect 993 253 1072 269
rect 841 237 907 253
rect 661 209 691 235
rect 733 209 763 237
rect 841 215 871 237
rect 1042 231 1072 253
rect 414 103 444 125
rect 308 87 444 103
rect 500 99 530 125
rect 572 99 602 125
rect 308 73 394 87
rect 378 53 394 73
rect 428 53 444 87
rect 378 51 444 53
rect 661 51 691 125
rect 733 99 763 125
rect 108 23 138 49
rect 194 23 224 49
rect 378 21 691 51
rect 841 21 871 47
rect 1042 37 1072 63
<< polycont >>
rect 96 239 130 273
rect 96 171 130 205
rect 288 343 322 377
rect 210 171 244 205
rect 460 299 494 333
rect 588 295 622 329
rect 749 253 783 287
rect 857 253 891 287
rect 1009 269 1043 303
rect 394 53 428 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 17 539 73 555
rect 17 505 35 539
rect 69 505 73 539
rect 17 471 73 505
rect 17 437 35 471
rect 69 437 73 471
rect 17 359 73 437
rect 117 545 159 649
rect 309 577 375 593
rect 117 511 121 545
rect 155 511 159 545
rect 117 477 159 511
rect 117 443 121 477
rect 155 443 159 477
rect 117 427 159 443
rect 203 539 267 555
rect 203 505 207 539
rect 241 505 267 539
rect 203 471 267 505
rect 203 437 207 471
rect 241 437 267 471
rect 309 543 325 577
rect 359 543 375 577
rect 309 507 375 543
rect 414 567 480 649
rect 414 533 430 567
rect 464 533 480 567
rect 791 579 857 649
rect 981 607 1043 649
rect 414 529 480 533
rect 603 533 692 549
rect 309 473 325 507
rect 359 495 375 507
rect 603 499 607 533
rect 641 499 692 533
rect 359 473 564 495
rect 309 461 564 473
rect 203 427 267 437
rect 203 393 338 427
rect 267 377 338 393
rect 17 325 231 359
rect 267 343 288 377
rect 322 343 338 377
rect 267 341 338 343
rect 17 121 60 325
rect 197 307 231 325
rect 444 333 496 349
rect 444 307 460 333
rect 197 299 460 307
rect 494 299 496 333
rect 94 273 163 289
rect 197 273 496 299
rect 530 345 564 461
rect 603 465 692 499
rect 603 431 619 465
rect 653 431 692 465
rect 603 415 692 431
rect 530 329 624 345
rect 530 295 588 329
rect 622 295 624 329
rect 530 279 624 295
rect 94 239 96 273
rect 130 239 163 273
rect 94 205 163 239
rect 530 237 564 279
rect 94 171 96 205
rect 130 171 163 205
rect 94 155 163 171
rect 210 205 257 221
rect 244 171 257 205
rect 210 155 257 171
rect 353 203 564 237
rect 353 185 405 203
rect 658 201 692 415
rect 791 545 807 579
rect 841 545 857 579
rect 791 511 857 545
rect 791 477 807 511
rect 841 477 857 511
rect 791 441 857 477
rect 791 407 807 441
rect 841 407 857 441
rect 891 574 943 590
rect 891 540 893 574
rect 927 540 943 574
rect 891 482 943 540
rect 891 448 893 482
rect 927 448 943 482
rect 891 389 943 448
rect 981 573 997 607
rect 1031 573 1043 607
rect 981 507 1043 573
rect 981 473 997 507
rect 1031 473 1043 507
rect 981 413 1043 473
rect 981 407 997 413
rect 891 373 893 389
rect 733 355 893 373
rect 927 373 943 389
rect 995 379 997 407
rect 1031 379 1043 413
rect 927 355 961 373
rect 995 363 1043 379
rect 1077 599 1135 615
rect 1077 565 1083 599
rect 1117 565 1135 599
rect 1077 508 1135 565
rect 1077 474 1083 508
rect 1117 474 1135 508
rect 1077 413 1135 474
rect 1077 379 1083 413
rect 1117 379 1135 413
rect 733 339 961 355
rect 733 287 799 339
rect 927 319 961 339
rect 927 303 1043 319
rect 733 253 749 287
rect 783 253 799 287
rect 733 237 799 253
rect 841 287 893 303
rect 841 253 857 287
rect 891 253 893 287
rect 841 201 893 253
rect 353 151 369 185
rect 403 151 405 185
rect 600 197 893 201
rect 353 135 405 151
rect 439 167 514 169
rect 439 133 455 167
rect 489 133 514 167
rect 600 163 616 197
rect 650 163 893 197
rect 600 159 893 163
rect 927 269 1009 303
rect 927 253 1043 269
rect 439 121 514 133
rect 927 125 961 253
rect 17 105 107 121
rect 17 71 63 105
rect 97 71 107 105
rect 17 53 107 71
rect 141 105 190 121
rect 141 71 149 105
rect 183 71 190 105
rect 141 17 190 71
rect 224 105 285 121
rect 224 71 235 105
rect 269 87 285 105
rect 269 71 394 87
rect 224 53 394 71
rect 428 53 444 87
rect 224 51 444 53
rect 480 17 514 121
rect 780 117 846 125
rect 780 83 796 117
rect 830 83 846 117
rect 780 17 846 83
rect 880 109 961 125
rect 880 75 882 109
rect 916 75 961 109
rect 880 57 961 75
rect 995 203 1043 219
rect 995 169 997 203
rect 1031 169 1043 203
rect 995 109 1043 169
rect 995 75 997 109
rect 1031 75 1043 109
rect 995 17 1043 75
rect 1077 212 1135 379
rect 1077 178 1083 212
rect 1117 178 1135 212
rect 1077 109 1135 178
rect 1077 75 1083 109
rect 1117 75 1135 109
rect 1077 59 1135 75
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlxtp_1
flabel comment s 318 204 318 204 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1087 94 1121 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1087 390 1121 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1087 464 1121 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1087 538 1121 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 37514
string GDS_START 27110
<< end >>
