magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 29 49 767 243
rect 0 0 768 49
<< scnmos >>
rect 108 133 138 217
rect 213 49 243 217
rect 299 49 329 217
rect 385 49 415 217
rect 471 49 501 217
rect 586 49 616 217
rect 658 49 688 217
<< scpmoshvt >>
rect 96 367 126 451
rect 213 367 243 619
rect 299 367 329 619
rect 385 367 415 619
rect 471 367 501 619
rect 572 367 602 619
rect 658 367 688 619
<< ndiff >>
rect 55 192 108 217
rect 55 158 63 192
rect 97 158 108 192
rect 55 133 108 158
rect 138 165 213 217
rect 138 133 168 165
rect 160 131 168 133
rect 202 131 213 165
rect 160 95 213 131
rect 160 61 168 95
rect 202 61 213 95
rect 160 49 213 61
rect 243 205 299 217
rect 243 171 254 205
rect 288 171 299 205
rect 243 101 299 171
rect 243 67 254 101
rect 288 67 299 101
rect 243 49 299 67
rect 329 176 385 217
rect 329 142 340 176
rect 374 142 385 176
rect 329 95 385 142
rect 329 61 340 95
rect 374 61 385 95
rect 329 49 385 61
rect 415 205 471 217
rect 415 171 426 205
rect 460 171 471 205
rect 415 101 471 171
rect 415 67 426 101
rect 460 67 471 101
rect 415 49 471 67
rect 501 159 586 217
rect 501 125 526 159
rect 560 125 586 159
rect 501 91 586 125
rect 501 57 526 91
rect 560 57 586 91
rect 501 49 586 57
rect 616 49 658 217
rect 688 205 741 217
rect 688 171 699 205
rect 733 171 741 205
rect 688 95 741 171
rect 688 61 699 95
rect 733 61 741 95
rect 688 49 741 61
<< pdiff >>
rect 160 600 213 619
rect 160 566 168 600
rect 202 566 213 600
rect 160 451 213 566
rect 43 439 96 451
rect 43 405 51 439
rect 85 405 96 439
rect 43 367 96 405
rect 126 367 213 451
rect 243 413 299 619
rect 243 379 254 413
rect 288 379 299 413
rect 243 367 299 379
rect 329 600 385 619
rect 329 566 340 600
rect 374 566 385 600
rect 329 367 385 566
rect 415 413 471 619
rect 415 379 426 413
rect 460 379 471 413
rect 415 367 471 379
rect 501 600 572 619
rect 501 566 519 600
rect 553 566 572 600
rect 501 367 572 566
rect 602 436 658 619
rect 602 402 613 436
rect 647 402 658 436
rect 602 367 658 402
rect 688 600 741 619
rect 688 566 699 600
rect 733 566 741 600
rect 688 367 741 566
<< ndiffc >>
rect 63 158 97 192
rect 168 131 202 165
rect 168 61 202 95
rect 254 171 288 205
rect 254 67 288 101
rect 340 142 374 176
rect 340 61 374 95
rect 426 171 460 205
rect 426 67 460 101
rect 526 125 560 159
rect 526 57 560 91
rect 699 171 733 205
rect 699 61 733 95
<< pdiffc >>
rect 168 566 202 600
rect 51 405 85 439
rect 254 379 288 413
rect 340 566 374 600
rect 426 379 460 413
rect 519 566 553 600
rect 613 402 647 436
rect 699 566 733 600
<< poly >>
rect 213 619 243 645
rect 299 619 329 645
rect 385 619 415 645
rect 471 619 501 645
rect 572 619 602 645
rect 658 619 688 645
rect 96 451 126 477
rect 96 308 126 367
rect 213 335 243 367
rect 299 335 329 367
rect 385 335 415 367
rect 471 335 501 367
rect 572 335 602 367
rect 213 319 501 335
rect 96 292 171 308
rect 96 258 121 292
rect 155 258 171 292
rect 96 242 171 258
rect 213 285 315 319
rect 349 285 383 319
rect 417 285 451 319
rect 485 285 501 319
rect 213 269 501 285
rect 550 319 616 335
rect 550 285 566 319
rect 600 285 616 319
rect 550 269 616 285
rect 108 217 138 242
rect 213 217 243 269
rect 299 217 329 269
rect 385 217 415 269
rect 471 217 501 269
rect 586 217 616 269
rect 658 325 688 367
rect 658 309 743 325
rect 658 275 693 309
rect 727 275 743 309
rect 658 259 743 275
rect 658 217 688 259
rect 108 107 138 133
rect 213 23 243 49
rect 299 23 329 49
rect 385 23 415 49
rect 471 23 501 49
rect 586 23 616 49
rect 658 23 688 49
<< polycont >>
rect 121 258 155 292
rect 315 285 349 319
rect 383 285 417 319
rect 451 285 485 319
rect 566 285 600 319
rect 693 275 727 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 152 600 218 649
rect 152 566 168 600
rect 202 566 218 600
rect 152 556 218 566
rect 324 600 390 649
rect 324 566 340 600
rect 374 566 390 600
rect 324 556 390 566
rect 503 600 569 649
rect 503 566 519 600
rect 553 566 569 600
rect 503 556 569 566
rect 683 600 749 649
rect 683 566 699 600
rect 733 566 749 600
rect 683 556 749 566
rect 35 486 743 522
rect 35 439 85 486
rect 35 405 51 439
rect 35 204 85 405
rect 121 292 176 441
rect 496 436 651 452
rect 155 258 176 292
rect 121 238 176 258
rect 210 413 460 429
rect 210 379 254 413
rect 288 379 426 413
rect 210 363 460 379
rect 496 402 613 436
rect 647 402 651 436
rect 496 386 651 402
rect 210 249 257 363
rect 496 329 532 386
rect 299 319 532 329
rect 299 285 315 319
rect 349 285 383 319
rect 417 285 451 319
rect 485 285 532 319
rect 299 283 532 285
rect 210 215 462 249
rect 246 205 290 215
rect 35 192 113 204
rect 35 158 63 192
rect 97 158 113 192
rect 35 144 113 158
rect 152 165 212 181
rect 152 131 168 165
rect 202 131 212 165
rect 152 95 212 131
rect 152 61 168 95
rect 202 61 212 95
rect 152 17 212 61
rect 246 171 254 205
rect 288 171 290 205
rect 424 205 462 215
rect 246 101 290 171
rect 246 67 254 101
rect 288 67 290 101
rect 246 51 290 67
rect 324 176 390 179
rect 324 142 340 176
rect 374 142 390 176
rect 324 95 390 142
rect 324 61 340 95
rect 374 61 390 95
rect 324 17 390 61
rect 424 171 426 205
rect 460 171 462 205
rect 496 233 532 283
rect 566 319 643 352
rect 600 285 643 319
rect 709 309 743 486
rect 566 269 643 285
rect 677 275 693 309
rect 727 275 743 309
rect 496 205 749 233
rect 496 199 699 205
rect 424 101 462 171
rect 683 171 699 199
rect 733 171 749 205
rect 424 67 426 101
rect 460 67 462 101
rect 424 51 462 67
rect 510 159 576 163
rect 510 125 526 159
rect 560 125 576 159
rect 510 91 576 125
rect 510 57 526 91
rect 560 57 576 91
rect 510 17 576 57
rect 683 95 749 171
rect 683 61 699 95
rect 733 61 749 95
rect 683 51 749 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and2b_4
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5133220
string GDS_START 5126718
<< end >>
