magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 198 179 575 241
rect 1 49 575 179
rect 0 0 576 49
<< scnmos >>
rect 80 69 110 153
rect 280 47 310 215
rect 367 47 397 215
rect 466 47 496 215
<< scpmoshvt >>
rect 175 403 205 487
rect 280 367 310 619
rect 394 367 424 619
rect 466 367 496 619
<< ndiff >>
rect 224 203 280 215
rect 224 169 232 203
rect 266 169 280 203
rect 27 127 80 153
rect 27 93 35 127
rect 69 93 80 127
rect 27 69 80 93
rect 110 127 163 153
rect 110 93 121 127
rect 155 93 163 127
rect 110 69 163 93
rect 224 93 280 169
rect 224 59 232 93
rect 266 59 280 93
rect 224 47 280 59
rect 310 203 367 215
rect 310 169 322 203
rect 356 169 367 203
rect 310 101 367 169
rect 310 67 322 101
rect 356 67 367 101
rect 310 47 367 67
rect 397 173 466 215
rect 397 139 412 173
rect 446 139 466 173
rect 397 93 466 139
rect 397 59 412 93
rect 446 59 466 93
rect 397 47 466 59
rect 496 203 549 215
rect 496 169 507 203
rect 541 169 549 203
rect 496 101 549 169
rect 496 67 507 101
rect 541 67 549 101
rect 496 47 549 67
<< pdiff >>
rect 227 607 280 619
rect 227 573 235 607
rect 269 573 280 607
rect 227 493 280 573
rect 227 487 235 493
rect 122 462 175 487
rect 122 428 130 462
rect 164 428 175 462
rect 122 403 175 428
rect 205 459 235 487
rect 269 459 280 493
rect 205 403 280 459
rect 227 367 280 403
rect 310 599 394 619
rect 310 565 335 599
rect 369 565 394 599
rect 310 510 394 565
rect 310 476 335 510
rect 369 476 394 510
rect 310 420 394 476
rect 310 386 335 420
rect 369 386 394 420
rect 310 367 394 386
rect 424 367 466 619
rect 496 607 549 619
rect 496 573 507 607
rect 541 573 549 607
rect 496 510 549 573
rect 496 476 507 510
rect 541 476 549 510
rect 496 418 549 476
rect 496 384 507 418
rect 541 384 549 418
rect 496 367 549 384
<< ndiffc >>
rect 232 169 266 203
rect 35 93 69 127
rect 121 93 155 127
rect 232 59 266 93
rect 322 169 356 203
rect 322 67 356 101
rect 412 139 446 173
rect 412 59 446 93
rect 507 169 541 203
rect 507 67 541 101
<< pdiffc >>
rect 235 573 269 607
rect 130 428 164 462
rect 235 459 269 493
rect 335 565 369 599
rect 335 476 369 510
rect 335 386 369 420
rect 507 573 541 607
rect 507 476 541 510
rect 507 384 541 418
<< poly >>
rect 280 619 310 645
rect 394 619 424 645
rect 466 619 496 645
rect 175 487 205 513
rect 175 381 205 403
rect 44 355 205 381
rect 44 321 60 355
rect 94 351 205 355
rect 94 321 110 351
rect 44 287 110 321
rect 280 303 310 367
rect 394 335 424 367
rect 44 253 60 287
rect 94 253 110 287
rect 44 237 110 253
rect 158 287 310 303
rect 158 253 174 287
rect 208 253 310 287
rect 352 319 424 335
rect 352 285 368 319
rect 402 285 424 319
rect 352 269 424 285
rect 466 325 496 367
rect 466 309 551 325
rect 466 275 501 309
rect 535 275 551 309
rect 158 237 310 253
rect 80 153 110 237
rect 280 215 310 237
rect 367 215 397 269
rect 466 259 551 275
rect 466 215 496 259
rect 80 43 110 69
rect 280 21 310 47
rect 367 21 397 47
rect 466 21 496 47
<< polycont >>
rect 60 321 94 355
rect 60 253 94 287
rect 174 253 208 287
rect 368 285 402 319
rect 501 275 535 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 214 607 285 649
rect 214 573 235 607
rect 269 573 285 607
rect 214 493 285 573
rect 114 462 180 478
rect 114 428 130 462
rect 164 428 180 462
rect 214 459 235 493
rect 269 459 285 493
rect 214 454 285 459
rect 319 599 385 615
rect 319 565 335 599
rect 369 565 385 599
rect 319 510 385 565
rect 319 476 335 510
rect 369 476 385 510
rect 114 412 180 428
rect 319 420 385 476
rect 17 355 103 378
rect 17 321 60 355
rect 94 321 103 355
rect 17 287 103 321
rect 17 253 60 287
rect 94 253 103 287
rect 17 237 103 253
rect 137 303 180 412
rect 248 386 335 420
rect 369 386 385 420
rect 491 607 557 649
rect 491 573 507 607
rect 541 573 557 607
rect 491 510 557 573
rect 491 476 507 510
rect 541 476 557 510
rect 491 418 557 476
rect 137 287 214 303
rect 137 253 174 287
rect 208 253 214 287
rect 137 237 214 253
rect 137 203 182 237
rect 248 203 282 386
rect 491 384 507 418
rect 541 384 557 418
rect 316 319 451 350
rect 316 285 368 319
rect 402 285 451 319
rect 316 275 451 285
rect 485 309 559 350
rect 485 275 501 309
rect 535 275 559 309
rect 19 169 182 203
rect 216 169 232 203
rect 266 169 282 203
rect 19 127 71 169
rect 19 93 35 127
rect 69 93 71 127
rect 19 77 71 93
rect 105 127 171 135
rect 105 93 121 127
rect 155 93 171 127
rect 105 17 171 93
rect 216 93 282 169
rect 216 59 232 93
rect 266 59 282 93
rect 216 51 282 59
rect 316 207 557 241
rect 316 203 362 207
rect 316 169 322 203
rect 356 169 362 203
rect 496 203 557 207
rect 316 101 362 169
rect 316 67 322 101
rect 356 67 362 101
rect 316 51 362 67
rect 396 139 412 173
rect 446 139 462 173
rect 396 93 462 139
rect 396 59 412 93
rect 446 59 462 93
rect 396 17 462 59
rect 496 169 507 203
rect 541 169 557 203
rect 496 101 557 169
rect 496 67 507 101
rect 541 67 557 101
rect 496 51 557 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21bai_1
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5208990
string GDS_START 5202940
<< end >>
