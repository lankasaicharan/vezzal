magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 284 228 666 248
rect 1 49 666 228
rect 0 0 672 49
<< scpmos >>
rect 101 383 131 551
rect 191 383 221 551
rect 370 368 400 592
rect 460 368 490 592
rect 556 368 586 592
<< nmoslvt >>
rect 84 74 114 202
rect 162 74 192 202
rect 367 74 397 222
rect 467 74 497 222
rect 553 74 583 222
<< ndiff >>
rect 310 210 367 222
rect 27 188 84 202
rect 27 154 39 188
rect 73 154 84 188
rect 27 120 84 154
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 74 162 202
rect 192 188 249 202
rect 192 154 203 188
rect 237 154 249 188
rect 192 120 249 154
rect 192 86 203 120
rect 237 86 249 120
rect 192 74 249 86
rect 310 176 322 210
rect 356 176 367 210
rect 310 120 367 176
rect 310 86 322 120
rect 356 86 367 120
rect 310 74 367 86
rect 397 139 467 222
rect 397 105 422 139
rect 456 105 467 139
rect 397 74 467 105
rect 497 131 553 222
rect 497 97 508 131
rect 542 97 553 131
rect 497 74 553 97
rect 583 210 640 222
rect 583 176 594 210
rect 628 176 640 210
rect 583 120 640 176
rect 583 86 594 120
rect 628 86 640 120
rect 583 74 640 86
<< pdiff >>
rect 276 580 370 592
rect 276 551 304 580
rect 32 539 101 551
rect 32 505 44 539
rect 78 505 101 539
rect 32 429 101 505
rect 32 395 44 429
rect 78 395 101 429
rect 32 383 101 395
rect 131 539 191 551
rect 131 505 144 539
rect 178 505 191 539
rect 131 429 191 505
rect 131 395 144 429
rect 178 395 191 429
rect 131 383 191 395
rect 221 546 304 551
rect 338 546 370 580
rect 221 503 370 546
rect 221 469 234 503
rect 268 469 304 503
rect 338 469 370 503
rect 221 429 370 469
rect 221 395 266 429
rect 300 395 370 429
rect 221 383 370 395
rect 317 368 370 383
rect 400 580 460 592
rect 400 546 413 580
rect 447 546 460 580
rect 400 510 460 546
rect 400 476 413 510
rect 447 476 460 510
rect 400 440 460 476
rect 400 406 413 440
rect 447 406 460 440
rect 400 368 460 406
rect 490 368 556 592
rect 586 580 645 592
rect 586 546 599 580
rect 633 546 645 580
rect 586 510 645 546
rect 586 476 599 510
rect 633 476 645 510
rect 586 440 645 476
rect 586 406 599 440
rect 633 406 645 440
rect 586 368 645 406
<< ndiffc >>
rect 39 154 73 188
rect 39 86 73 120
rect 203 154 237 188
rect 203 86 237 120
rect 322 176 356 210
rect 322 86 356 120
rect 422 105 456 139
rect 508 97 542 131
rect 594 176 628 210
rect 594 86 628 120
<< pdiffc >>
rect 44 505 78 539
rect 44 395 78 429
rect 144 505 178 539
rect 144 395 178 429
rect 304 546 338 580
rect 234 469 268 503
rect 304 469 338 503
rect 266 395 300 429
rect 413 546 447 580
rect 413 476 447 510
rect 413 406 447 440
rect 599 546 633 580
rect 599 476 633 510
rect 599 406 633 440
<< poly >>
rect 370 592 400 618
rect 460 592 490 618
rect 556 592 586 618
rect 101 551 131 577
rect 191 551 221 577
rect 101 368 131 383
rect 191 368 221 383
rect 84 338 134 368
rect 84 302 114 338
rect 21 286 114 302
rect 188 290 224 368
rect 370 353 400 368
rect 460 353 490 368
rect 556 353 586 368
rect 367 336 403 353
rect 21 252 37 286
rect 71 252 114 286
rect 21 236 114 252
rect 84 202 114 236
rect 156 274 224 290
rect 156 240 172 274
rect 206 260 224 274
rect 272 320 403 336
rect 457 326 493 353
rect 553 326 589 353
rect 272 286 288 320
rect 322 286 403 320
rect 272 270 403 286
rect 445 310 511 326
rect 445 276 461 310
rect 495 276 511 310
rect 206 240 222 260
rect 156 224 222 240
rect 162 202 192 224
rect 367 222 397 270
rect 445 260 511 276
rect 553 310 651 326
rect 553 276 601 310
rect 635 276 651 310
rect 553 260 651 276
rect 467 222 497 260
rect 553 222 583 260
rect 84 48 114 74
rect 162 48 192 74
rect 367 48 397 74
rect 467 48 497 74
rect 553 48 583 74
<< polycont >>
rect 37 252 71 286
rect 172 240 206 274
rect 288 286 322 320
rect 461 276 495 310
rect 601 276 635 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 28 539 94 649
rect 228 580 338 649
rect 28 505 44 539
rect 78 505 94 539
rect 28 429 94 505
rect 28 395 44 429
rect 78 395 94 429
rect 28 379 94 395
rect 128 539 194 555
rect 128 505 144 539
rect 178 505 194 539
rect 128 429 194 505
rect 128 395 144 429
rect 178 395 194 429
rect 228 546 304 580
rect 228 503 338 546
rect 228 469 234 503
rect 268 469 304 503
rect 228 429 338 469
rect 228 395 266 429
rect 300 395 338 429
rect 372 580 463 596
rect 372 546 413 580
rect 447 546 463 580
rect 372 510 463 546
rect 372 476 413 510
rect 447 476 463 510
rect 372 440 463 476
rect 372 406 413 440
rect 447 406 463 440
rect 128 358 194 395
rect 372 390 463 406
rect 599 580 649 649
rect 633 546 649 580
rect 599 510 649 546
rect 633 476 649 510
rect 599 440 649 476
rect 633 406 649 440
rect 599 390 649 406
rect 128 324 338 358
rect 254 320 338 324
rect 21 286 87 302
rect 21 252 37 286
rect 71 252 87 286
rect 21 236 87 252
rect 121 274 220 290
rect 121 240 172 274
rect 206 240 220 274
rect 121 224 220 240
rect 254 286 288 320
rect 322 286 338 320
rect 254 270 338 286
rect 254 190 288 270
rect 372 236 406 390
rect 445 310 551 356
rect 445 276 461 310
rect 495 276 551 310
rect 445 260 551 276
rect 585 310 651 356
rect 585 276 601 310
rect 635 276 651 310
rect 585 260 651 276
rect 23 188 89 190
rect 23 154 39 188
rect 73 154 89 188
rect 23 120 89 154
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 187 188 288 190
rect 187 154 203 188
rect 237 154 288 188
rect 187 120 288 154
rect 187 86 203 120
rect 237 86 288 120
rect 187 70 288 86
rect 322 210 406 236
rect 356 202 406 210
rect 440 210 644 226
rect 356 176 372 202
rect 322 120 372 176
rect 440 192 594 210
rect 440 168 474 192
rect 356 86 372 120
rect 406 139 474 168
rect 578 176 594 192
rect 628 176 644 210
rect 406 105 422 139
rect 456 105 474 139
rect 406 89 474 105
rect 508 131 542 158
rect 322 70 372 86
rect 508 17 542 97
rect 578 120 644 176
rect 578 86 594 120
rect 628 86 644 120
rect 578 70 644 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o2bb2ai_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 2990482
string GDS_START 2983882
<< end >>
