magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 1 49 855 247
rect 0 0 864 49
<< scnmos >>
rect 84 53 114 221
rect 170 53 200 221
rect 284 53 314 221
rect 370 53 400 221
rect 456 53 486 221
rect 542 53 572 221
rect 642 53 672 221
rect 742 53 772 221
<< scpmoshvt >>
rect 88 367 118 619
rect 174 367 204 619
rect 260 367 290 619
rect 346 367 376 619
rect 446 367 476 619
rect 546 367 576 619
rect 646 367 676 619
rect 732 367 762 619
<< ndiff >>
rect 27 209 84 221
rect 27 175 39 209
rect 73 175 84 209
rect 27 99 84 175
rect 27 65 39 99
rect 73 65 84 99
rect 27 53 84 65
rect 114 186 170 221
rect 114 152 125 186
rect 159 152 170 186
rect 114 101 170 152
rect 114 67 125 101
rect 159 67 170 101
rect 114 53 170 67
rect 200 99 284 221
rect 200 65 225 99
rect 259 65 284 99
rect 200 53 284 65
rect 314 126 370 221
rect 314 92 325 126
rect 359 92 370 126
rect 314 53 370 92
rect 400 189 456 221
rect 400 155 411 189
rect 445 155 456 189
rect 400 53 456 155
rect 486 167 542 221
rect 486 133 497 167
rect 531 133 542 167
rect 486 99 542 133
rect 486 65 497 99
rect 531 65 542 99
rect 486 53 542 65
rect 572 189 642 221
rect 572 155 597 189
rect 631 155 642 189
rect 572 53 642 155
rect 672 209 742 221
rect 672 175 697 209
rect 731 175 742 209
rect 672 101 742 175
rect 672 67 697 101
rect 731 67 742 101
rect 672 53 742 67
rect 772 209 829 221
rect 772 175 783 209
rect 817 175 829 209
rect 772 99 829 175
rect 772 65 783 99
rect 817 65 829 99
rect 772 53 829 65
<< pdiff >>
rect 31 607 88 619
rect 31 573 43 607
rect 77 573 88 607
rect 31 510 88 573
rect 31 476 43 510
rect 77 476 88 510
rect 31 413 88 476
rect 31 379 43 413
rect 77 379 88 413
rect 31 367 88 379
rect 118 599 174 619
rect 118 565 129 599
rect 163 565 174 599
rect 118 506 174 565
rect 118 472 129 506
rect 163 472 174 506
rect 118 413 174 472
rect 118 379 129 413
rect 163 379 174 413
rect 118 367 174 379
rect 204 591 260 619
rect 204 557 215 591
rect 249 557 260 591
rect 204 367 260 557
rect 290 599 346 619
rect 290 565 301 599
rect 335 565 346 599
rect 290 508 346 565
rect 290 474 301 508
rect 335 474 346 508
rect 290 367 346 474
rect 376 531 446 619
rect 376 497 401 531
rect 435 497 446 531
rect 376 440 446 497
rect 376 406 401 440
rect 435 406 446 440
rect 376 367 446 406
rect 476 599 546 619
rect 476 565 501 599
rect 535 565 546 599
rect 476 508 546 565
rect 476 474 501 508
rect 535 474 546 508
rect 476 367 546 474
rect 576 531 646 619
rect 576 497 601 531
rect 635 497 646 531
rect 576 419 646 497
rect 576 385 601 419
rect 635 385 646 419
rect 576 367 646 385
rect 676 599 732 619
rect 676 565 687 599
rect 721 565 732 599
rect 676 509 732 565
rect 676 475 687 509
rect 721 475 732 509
rect 676 419 732 475
rect 676 385 687 419
rect 721 385 732 419
rect 676 367 732 385
rect 762 607 833 619
rect 762 573 787 607
rect 821 573 833 607
rect 762 513 833 573
rect 762 479 787 513
rect 821 479 833 513
rect 762 419 833 479
rect 762 385 787 419
rect 821 385 833 419
rect 762 367 833 385
<< ndiffc >>
rect 39 175 73 209
rect 39 65 73 99
rect 125 152 159 186
rect 125 67 159 101
rect 225 65 259 99
rect 325 92 359 126
rect 411 155 445 189
rect 497 133 531 167
rect 497 65 531 99
rect 597 155 631 189
rect 697 175 731 209
rect 697 67 731 101
rect 783 175 817 209
rect 783 65 817 99
<< pdiffc >>
rect 43 573 77 607
rect 43 476 77 510
rect 43 379 77 413
rect 129 565 163 599
rect 129 472 163 506
rect 129 379 163 413
rect 215 557 249 591
rect 301 565 335 599
rect 301 474 335 508
rect 401 497 435 531
rect 401 406 435 440
rect 501 565 535 599
rect 501 474 535 508
rect 601 497 635 531
rect 601 385 635 419
rect 687 565 721 599
rect 687 475 721 509
rect 687 385 721 419
rect 787 573 821 607
rect 787 479 821 513
rect 787 385 821 419
<< poly >>
rect 88 619 118 645
rect 174 619 204 645
rect 260 619 290 645
rect 346 619 376 645
rect 446 619 476 645
rect 546 619 576 645
rect 646 619 676 645
rect 732 619 762 645
rect 88 335 118 367
rect 174 335 204 367
rect 260 335 290 367
rect 346 335 376 367
rect 446 335 476 367
rect 546 335 576 367
rect 646 335 676 367
rect 732 335 762 367
rect 84 319 819 335
rect 84 285 293 319
rect 327 285 361 319
rect 395 285 429 319
rect 463 285 497 319
rect 531 285 565 319
rect 599 285 633 319
rect 667 285 701 319
rect 735 285 769 319
rect 803 285 819 319
rect 84 269 819 285
rect 84 221 114 269
rect 170 221 200 269
rect 284 221 314 269
rect 370 221 400 269
rect 456 221 486 269
rect 542 221 572 269
rect 642 221 672 269
rect 742 221 772 269
rect 84 27 114 53
rect 170 27 200 53
rect 284 27 314 53
rect 370 27 400 53
rect 456 27 486 53
rect 542 27 572 53
rect 642 27 672 53
rect 742 27 772 53
<< polycont >>
rect 293 285 327 319
rect 361 285 395 319
rect 429 285 463 319
rect 497 285 531 319
rect 565 285 599 319
rect 633 285 667 319
rect 701 285 735 319
rect 769 285 803 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 27 607 77 649
rect 27 573 43 607
rect 27 510 77 573
rect 27 476 43 510
rect 27 413 77 476
rect 27 379 43 413
rect 27 363 77 379
rect 113 599 163 615
rect 113 565 129 599
rect 113 506 163 565
rect 199 591 249 649
rect 199 557 215 591
rect 199 526 249 557
rect 285 599 737 615
rect 285 565 301 599
rect 335 581 501 599
rect 335 565 351 581
rect 113 472 129 506
rect 285 508 351 565
rect 485 565 501 581
rect 535 581 687 599
rect 535 565 551 581
rect 285 492 301 508
rect 163 474 301 492
rect 335 474 351 508
rect 163 472 351 474
rect 113 458 351 472
rect 385 531 451 547
rect 385 497 401 531
rect 435 497 451 531
rect 113 413 163 458
rect 385 440 451 497
rect 485 508 551 565
rect 721 565 737 599
rect 485 474 501 508
rect 535 474 551 508
rect 485 458 551 474
rect 585 531 651 547
rect 585 497 601 531
rect 635 497 651 531
rect 385 424 401 440
rect 113 379 129 413
rect 113 363 163 379
rect 209 406 401 424
rect 435 424 451 440
rect 585 424 651 497
rect 435 419 651 424
rect 435 406 601 419
rect 209 390 601 406
rect 209 282 243 390
rect 585 385 601 390
rect 635 385 651 419
rect 585 369 651 385
rect 687 509 737 565
rect 721 475 737 509
rect 687 419 737 475
rect 721 385 737 419
rect 687 369 737 385
rect 771 607 837 649
rect 771 573 787 607
rect 821 573 837 607
rect 771 513 837 573
rect 771 479 787 513
rect 821 479 837 513
rect 771 419 837 479
rect 771 385 787 419
rect 821 385 837 419
rect 771 369 837 385
rect 313 335 551 356
rect 121 236 243 282
rect 277 319 819 335
rect 277 285 293 319
rect 327 285 361 319
rect 395 285 429 319
rect 463 285 497 319
rect 531 285 565 319
rect 599 285 633 319
rect 667 285 701 319
rect 735 285 769 319
rect 803 285 819 319
rect 277 269 819 285
rect 209 235 243 236
rect 23 209 73 225
rect 23 175 39 209
rect 23 99 73 175
rect 23 65 39 99
rect 23 17 73 65
rect 109 186 175 202
rect 209 201 647 235
rect 109 152 125 186
rect 159 167 175 186
rect 411 189 445 201
rect 159 152 375 167
rect 109 133 375 152
rect 109 101 175 133
rect 109 67 125 101
rect 159 67 175 101
rect 309 126 375 133
rect 109 51 175 67
rect 209 65 225 99
rect 259 65 275 99
rect 209 17 275 65
rect 309 92 325 126
rect 359 92 375 126
rect 581 189 647 201
rect 411 119 445 155
rect 481 133 497 167
rect 531 133 547 167
rect 309 85 375 92
rect 481 99 547 133
rect 581 155 597 189
rect 631 155 647 189
rect 581 119 647 155
rect 681 209 747 225
rect 681 175 697 209
rect 731 175 747 209
rect 481 85 497 99
rect 309 65 497 85
rect 531 85 547 99
rect 681 101 747 175
rect 681 85 697 101
rect 531 67 697 85
rect 731 67 747 101
rect 531 65 747 67
rect 309 51 747 65
rect 783 209 833 225
rect 817 175 833 209
rect 783 99 833 175
rect 817 65 833 99
rect 783 17 833 65
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 invlp_4
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6824574
string GDS_START 6817288
<< end >>
