magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 331 1478 704
<< pwell >>
rect 126 183 386 235
rect 1168 203 1439 287
rect 724 183 1439 203
rect 10 49 1439 183
rect 0 0 1440 49
<< scnmos >>
rect 93 73 123 157
rect 202 125 232 209
rect 280 125 310 209
rect 1254 177 1284 261
rect 1326 177 1356 261
rect 389 73 419 157
rect 491 73 521 157
rect 569 73 599 157
rect 807 93 837 177
rect 879 93 909 177
rect 979 93 1009 177
rect 1051 93 1081 177
<< scpmoshvt >>
rect 87 535 117 619
rect 251 535 281 619
rect 360 419 410 619
rect 458 419 508 619
rect 564 419 614 619
rect 887 415 917 543
rect 1128 387 1178 587
rect 1234 387 1284 587
<< ndiff >>
rect 152 157 202 209
rect 36 132 93 157
rect 36 98 48 132
rect 82 98 93 132
rect 36 73 93 98
rect 123 126 202 157
rect 123 92 134 126
rect 168 125 202 126
rect 232 125 280 209
rect 310 157 360 209
rect 1194 249 1254 261
rect 1194 215 1206 249
rect 1240 215 1254 249
rect 1194 177 1254 215
rect 1284 177 1326 261
rect 1356 236 1413 261
rect 1356 202 1367 236
rect 1401 202 1413 236
rect 1356 177 1413 202
rect 750 169 807 177
rect 310 125 389 157
rect 168 92 180 125
rect 332 124 389 125
rect 123 73 180 92
rect 332 90 344 124
rect 378 90 389 124
rect 332 73 389 90
rect 419 73 491 157
rect 521 73 569 157
rect 599 129 656 157
rect 599 95 610 129
rect 644 95 656 129
rect 599 73 656 95
rect 750 135 762 169
rect 796 135 807 169
rect 750 93 807 135
rect 837 93 879 177
rect 909 152 979 177
rect 909 118 920 152
rect 954 118 979 152
rect 909 93 979 118
rect 1009 93 1051 177
rect 1081 139 1134 177
rect 1081 105 1092 139
rect 1126 105 1134 139
rect 1081 93 1134 105
<< pdiff >>
rect 30 597 87 619
rect 30 563 42 597
rect 76 563 87 597
rect 30 535 87 563
rect 117 535 251 619
rect 281 535 360 619
rect 303 519 360 535
rect 303 485 315 519
rect 349 485 360 519
rect 303 419 360 485
rect 410 419 458 619
rect 508 597 564 619
rect 508 563 519 597
rect 553 563 564 597
rect 508 529 564 563
rect 508 495 519 529
rect 553 495 564 529
rect 508 461 564 495
rect 508 427 519 461
rect 553 427 564 461
rect 508 419 564 427
rect 614 597 671 619
rect 614 563 625 597
rect 659 563 671 597
rect 1071 575 1128 587
rect 614 529 671 563
rect 614 495 625 529
rect 659 495 671 529
rect 614 461 671 495
rect 807 531 887 543
rect 807 497 819 531
rect 853 497 887 531
rect 614 427 625 461
rect 659 427 671 461
rect 614 419 671 427
rect 807 461 887 497
rect 807 427 819 461
rect 853 427 887 461
rect 807 415 887 427
rect 917 519 1017 543
rect 917 485 971 519
rect 1005 485 1017 519
rect 917 415 1017 485
rect 1071 541 1083 575
rect 1117 541 1128 575
rect 1071 504 1128 541
rect 1071 470 1083 504
rect 1117 470 1128 504
rect 1071 433 1128 470
rect 1071 399 1083 433
rect 1117 399 1128 433
rect 1071 387 1128 399
rect 1178 575 1234 587
rect 1178 541 1189 575
rect 1223 541 1234 575
rect 1178 504 1234 541
rect 1178 470 1189 504
rect 1223 470 1234 504
rect 1178 433 1234 470
rect 1178 399 1189 433
rect 1223 399 1234 433
rect 1178 387 1234 399
rect 1284 575 1352 587
rect 1284 541 1306 575
rect 1340 541 1352 575
rect 1284 504 1352 541
rect 1284 470 1306 504
rect 1340 470 1352 504
rect 1284 433 1352 470
rect 1284 399 1306 433
rect 1340 399 1352 433
rect 1284 387 1352 399
<< ndiffc >>
rect 48 98 82 132
rect 134 92 168 126
rect 1206 215 1240 249
rect 1367 202 1401 236
rect 344 90 378 124
rect 610 95 644 129
rect 762 135 796 169
rect 920 118 954 152
rect 1092 105 1126 139
<< pdiffc >>
rect 42 563 76 597
rect 315 485 349 519
rect 519 563 553 597
rect 519 495 553 529
rect 519 427 553 461
rect 625 563 659 597
rect 625 495 659 529
rect 819 497 853 531
rect 625 427 659 461
rect 819 427 853 461
rect 971 485 1005 519
rect 1083 541 1117 575
rect 1083 470 1117 504
rect 1083 399 1117 433
rect 1189 541 1223 575
rect 1189 470 1223 504
rect 1189 399 1223 433
rect 1306 541 1340 575
rect 1306 470 1340 504
rect 1306 399 1340 433
<< poly >>
rect 87 619 117 645
rect 251 619 281 645
rect 360 619 410 645
rect 458 619 508 645
rect 564 619 614 645
rect 87 503 117 535
rect 51 487 117 503
rect 51 453 67 487
rect 101 453 117 487
rect 251 465 281 535
rect 51 437 117 453
rect 159 435 281 465
rect 159 395 189 435
rect 1128 587 1178 613
rect 1234 587 1284 613
rect 887 543 917 569
rect 703 475 769 491
rect 703 441 719 475
rect 753 441 769 475
rect 21 365 189 395
rect 360 387 410 419
rect 237 371 410 387
rect 21 209 51 365
rect 237 337 253 371
rect 287 337 410 371
rect 237 321 410 337
rect 458 323 508 419
rect 564 323 614 419
rect 703 407 769 441
rect 703 373 719 407
rect 753 373 769 407
rect 703 357 769 373
rect 99 301 195 317
rect 99 267 115 301
rect 149 273 195 301
rect 149 267 232 273
rect 99 251 232 267
rect 165 243 232 251
rect 202 209 232 243
rect 280 209 310 321
rect 458 293 521 323
rect 383 229 449 245
rect 21 179 123 209
rect 93 157 123 179
rect 383 195 399 229
rect 433 195 449 229
rect 383 179 449 195
rect 491 209 521 293
rect 564 307 630 323
rect 564 273 580 307
rect 614 273 630 307
rect 564 257 630 273
rect 703 209 733 357
rect 887 356 917 415
rect 871 340 937 356
rect 871 306 887 340
rect 921 306 937 340
rect 871 290 937 306
rect 491 179 733 209
rect 807 274 937 290
rect 979 333 1045 349
rect 979 299 995 333
rect 1029 299 1045 333
rect 807 260 909 274
rect 389 157 419 179
rect 491 157 521 179
rect 569 157 599 179
rect 807 177 837 260
rect 879 177 909 260
rect 979 265 1045 299
rect 979 231 995 265
rect 1029 245 1045 265
rect 1128 315 1178 387
rect 1234 315 1284 387
rect 1128 285 1356 315
rect 1128 245 1158 285
rect 1254 261 1284 285
rect 1326 261 1356 285
rect 1029 231 1158 245
rect 979 215 1158 231
rect 979 177 1009 215
rect 1051 177 1081 215
rect 202 99 232 125
rect 280 99 310 125
rect 1254 151 1284 177
rect 1326 151 1356 177
rect 93 51 123 73
rect 389 51 419 73
rect 93 21 419 51
rect 491 47 521 73
rect 569 47 599 73
rect 807 67 837 93
rect 879 67 909 93
rect 979 67 1009 93
rect 1051 67 1081 93
<< polycont >>
rect 67 453 101 487
rect 719 441 753 475
rect 253 337 287 371
rect 719 373 753 407
rect 115 267 149 301
rect 399 195 433 229
rect 580 273 614 307
rect 887 306 921 340
rect 995 299 1029 333
rect 995 231 1029 265
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 26 597 92 649
rect 26 563 42 597
rect 76 563 92 597
rect 26 537 92 563
rect 231 581 469 615
rect 25 487 117 503
rect 25 453 67 487
rect 101 453 117 487
rect 25 437 117 453
rect 25 356 59 437
rect 231 424 265 581
rect 299 519 371 547
rect 299 485 315 519
rect 349 485 371 519
rect 299 458 371 485
rect 231 390 303 424
rect 237 371 303 390
rect 25 301 167 356
rect 25 267 115 301
rect 149 267 167 301
rect 25 251 167 267
rect 237 337 253 371
rect 287 337 303 371
rect 237 334 303 337
rect 237 217 271 334
rect 337 300 371 458
rect 435 391 469 581
rect 503 597 569 615
rect 503 581 519 597
rect 503 547 511 581
rect 553 563 569 597
rect 545 547 569 563
rect 503 529 569 547
rect 503 495 519 529
rect 553 495 569 529
rect 503 461 569 495
rect 503 427 519 461
rect 553 427 569 461
rect 503 425 569 427
rect 609 597 659 615
rect 609 563 625 597
rect 609 529 659 563
rect 609 495 625 529
rect 609 461 659 495
rect 609 427 625 461
rect 609 391 659 427
rect 435 357 659 391
rect 703 581 921 615
rect 703 475 769 581
rect 703 441 719 475
rect 753 441 769 475
rect 703 407 769 441
rect 703 373 719 407
rect 753 373 769 407
rect 703 357 769 373
rect 803 531 853 547
rect 803 497 819 531
rect 803 461 853 497
rect 803 427 819 461
rect 803 411 853 427
rect 887 424 921 581
rect 955 547 991 581
rect 1025 547 1031 581
rect 955 519 1031 547
rect 955 485 971 519
rect 1005 485 1031 519
rect 955 458 1031 485
rect 1067 575 1133 591
rect 1067 541 1083 575
rect 1117 541 1133 575
rect 1067 504 1133 541
rect 1067 470 1083 504
rect 1117 470 1133 504
rect 1067 433 1133 470
rect 1067 424 1083 433
rect 803 323 837 411
rect 887 399 1083 424
rect 1117 399 1133 433
rect 887 390 1133 399
rect 1067 383 1133 390
rect 1173 581 1239 591
rect 1173 547 1183 581
rect 1217 575 1239 581
rect 1173 541 1189 547
rect 1223 541 1239 575
rect 1173 504 1239 541
rect 1173 470 1189 504
rect 1223 470 1239 504
rect 1173 433 1239 470
rect 1173 399 1189 433
rect 1223 399 1239 433
rect 1173 383 1239 399
rect 1290 575 1417 591
rect 1290 541 1306 575
rect 1340 541 1417 575
rect 1290 504 1417 541
rect 1290 470 1306 504
rect 1340 470 1417 504
rect 1290 433 1417 470
rect 1290 399 1306 433
rect 1340 399 1417 433
rect 32 183 271 217
rect 315 266 371 300
rect 415 307 837 323
rect 415 273 580 307
rect 614 289 837 307
rect 871 340 937 356
rect 871 306 887 340
rect 921 306 937 340
rect 871 290 937 306
rect 979 333 1045 349
rect 979 299 995 333
rect 1029 299 1045 333
rect 614 273 796 289
rect 32 132 82 183
rect 32 98 48 132
rect 32 69 82 98
rect 118 126 184 149
rect 118 92 134 126
rect 168 92 184 126
rect 118 17 184 92
rect 315 145 349 266
rect 415 257 796 273
rect 415 232 449 257
rect 383 229 449 232
rect 383 195 399 229
rect 433 195 449 229
rect 383 179 449 195
rect 483 189 712 223
rect 483 145 517 189
rect 315 124 517 145
rect 315 90 344 124
rect 378 111 517 124
rect 594 129 644 155
rect 378 90 394 111
rect 315 69 394 90
rect 594 95 610 129
rect 594 17 644 95
rect 678 85 712 189
rect 746 169 796 257
rect 979 265 1045 299
rect 979 249 995 265
rect 746 135 762 169
rect 746 119 796 135
rect 830 231 995 249
rect 1029 231 1045 265
rect 830 215 1045 231
rect 830 85 864 215
rect 678 51 864 85
rect 920 152 970 181
rect 1099 155 1133 383
rect 954 118 970 152
rect 920 17 970 118
rect 1092 139 1133 155
rect 1126 105 1133 139
rect 1092 89 1133 105
rect 1190 249 1256 265
rect 1190 215 1206 249
rect 1240 215 1256 249
rect 1190 17 1256 215
rect 1290 236 1417 399
rect 1290 202 1367 236
rect 1401 202 1417 236
rect 1290 88 1417 202
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 511 563 519 581
rect 519 563 545 581
rect 511 547 545 563
rect 991 547 1025 581
rect 1183 575 1217 581
rect 1183 547 1189 575
rect 1189 547 1217 575
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 14 581 1426 589
rect 14 547 511 581
rect 545 547 991 581
rect 1025 547 1183 581
rect 1217 547 1426 581
rect 14 535 1426 547
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 isolatch_lp
flabel metal1 s 14 535 1426 589 0 FreeSans 340 0 0 0 KAPWR
port 3 nsew power bidirectional
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 SLEEP_B
port 2 nsew clock input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1375 94 1409 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1375 168 1409 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1375 390 1409 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5086618
string GDS_START 5076048
<< end >>
