magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 48 49 1991 241
rect 0 0 2016 49
<< scnmos >>
rect 127 47 157 215
rect 213 47 243 215
rect 299 47 329 215
rect 385 47 415 215
rect 471 47 501 215
rect 557 47 587 215
rect 643 47 673 215
rect 729 47 759 215
rect 832 47 862 215
rect 918 47 948 215
rect 1004 47 1034 215
rect 1090 47 1120 215
rect 1176 47 1206 215
rect 1262 47 1292 215
rect 1348 47 1378 215
rect 1434 47 1464 215
rect 1624 47 1654 215
rect 1710 47 1740 215
rect 1796 47 1826 215
rect 1882 47 1912 215
<< scpmoshvt >>
rect 126 367 156 619
rect 212 367 242 619
rect 298 367 328 619
rect 384 367 414 619
rect 470 367 500 619
rect 556 367 586 619
rect 642 367 672 619
rect 760 367 790 619
rect 846 367 876 619
rect 932 367 962 619
rect 1018 367 1048 619
rect 1104 367 1134 619
rect 1294 367 1324 619
rect 1380 367 1410 619
rect 1466 367 1496 619
rect 1552 367 1582 619
rect 1638 367 1668 619
rect 1724 367 1754 619
rect 1810 367 1840 619
rect 1896 367 1926 619
<< ndiff >>
rect 74 203 127 215
rect 74 169 82 203
rect 116 169 127 203
rect 74 93 127 169
rect 74 59 82 93
rect 116 59 127 93
rect 74 47 127 59
rect 157 207 213 215
rect 157 173 168 207
rect 202 173 213 207
rect 157 101 213 173
rect 157 67 168 101
rect 202 67 213 101
rect 157 47 213 67
rect 243 168 299 215
rect 243 134 254 168
rect 288 134 299 168
rect 243 89 299 134
rect 243 55 254 89
rect 288 55 299 89
rect 243 47 299 55
rect 329 207 385 215
rect 329 173 340 207
rect 374 173 385 207
rect 329 101 385 173
rect 329 67 340 101
rect 374 67 385 101
rect 329 47 385 67
rect 415 195 471 215
rect 415 161 426 195
rect 460 161 471 195
rect 415 47 471 161
rect 501 101 557 215
rect 501 67 512 101
rect 546 67 557 101
rect 501 47 557 67
rect 587 195 643 215
rect 587 161 598 195
rect 632 161 643 195
rect 587 47 643 161
rect 673 101 729 215
rect 673 67 684 101
rect 718 67 729 101
rect 673 47 729 67
rect 759 110 832 215
rect 759 76 778 110
rect 812 76 832 110
rect 759 47 832 76
rect 862 203 918 215
rect 862 169 873 203
rect 907 169 918 203
rect 862 101 918 169
rect 862 67 873 101
rect 907 67 918 101
rect 862 47 918 67
rect 948 173 1004 215
rect 948 139 959 173
rect 993 139 1004 173
rect 948 89 1004 139
rect 948 55 959 89
rect 993 55 1004 89
rect 948 47 1004 55
rect 1034 203 1090 215
rect 1034 169 1045 203
rect 1079 169 1090 203
rect 1034 101 1090 169
rect 1034 67 1045 101
rect 1079 67 1090 101
rect 1034 47 1090 67
rect 1120 175 1176 215
rect 1120 141 1131 175
rect 1165 141 1176 175
rect 1120 89 1176 141
rect 1120 55 1131 89
rect 1165 55 1176 89
rect 1120 47 1176 55
rect 1206 203 1262 215
rect 1206 169 1217 203
rect 1251 169 1262 203
rect 1206 135 1262 169
rect 1206 101 1217 135
rect 1251 101 1262 135
rect 1206 47 1262 101
rect 1292 161 1348 215
rect 1292 127 1303 161
rect 1337 127 1348 161
rect 1292 93 1348 127
rect 1292 59 1303 93
rect 1337 59 1348 93
rect 1292 47 1348 59
rect 1378 203 1434 215
rect 1378 169 1389 203
rect 1423 169 1434 203
rect 1378 101 1434 169
rect 1378 67 1389 101
rect 1423 67 1434 101
rect 1378 47 1434 67
rect 1464 174 1624 215
rect 1464 140 1475 174
rect 1509 140 1624 174
rect 1464 124 1624 140
rect 1464 90 1579 124
rect 1613 90 1624 124
rect 1464 89 1624 90
rect 1464 55 1475 89
rect 1509 55 1624 89
rect 1464 47 1624 55
rect 1654 192 1710 215
rect 1654 158 1665 192
rect 1699 158 1710 192
rect 1654 101 1710 158
rect 1654 67 1665 101
rect 1699 67 1710 101
rect 1654 47 1710 67
rect 1740 124 1796 215
rect 1740 90 1751 124
rect 1785 90 1796 124
rect 1740 47 1796 90
rect 1826 203 1882 215
rect 1826 169 1837 203
rect 1871 169 1882 203
rect 1826 101 1882 169
rect 1826 67 1837 101
rect 1871 67 1882 101
rect 1826 47 1882 67
rect 1912 167 1965 215
rect 1912 133 1923 167
rect 1957 133 1965 167
rect 1912 93 1965 133
rect 1912 59 1923 93
rect 1957 59 1965 93
rect 1912 47 1965 59
<< pdiff >>
rect 687 619 745 627
rect 73 599 126 619
rect 73 565 81 599
rect 115 565 126 599
rect 73 505 126 565
rect 73 471 81 505
rect 115 471 126 505
rect 73 413 126 471
rect 73 379 81 413
rect 115 379 126 413
rect 73 367 126 379
rect 156 607 212 619
rect 156 573 167 607
rect 201 573 212 607
rect 156 530 212 573
rect 156 496 167 530
rect 201 496 212 530
rect 156 447 212 496
rect 156 413 167 447
rect 201 413 212 447
rect 156 367 212 413
rect 242 599 298 619
rect 242 565 253 599
rect 287 565 298 599
rect 242 505 298 565
rect 242 471 253 505
rect 287 471 298 505
rect 242 413 298 471
rect 242 379 253 413
rect 287 379 298 413
rect 242 367 298 379
rect 328 607 384 619
rect 328 573 339 607
rect 373 573 384 607
rect 328 505 384 573
rect 328 471 339 505
rect 373 471 384 505
rect 328 367 384 471
rect 414 599 470 619
rect 414 565 425 599
rect 459 565 470 599
rect 414 526 470 565
rect 414 492 425 526
rect 459 492 470 526
rect 414 453 470 492
rect 414 419 425 453
rect 459 419 470 453
rect 414 367 470 419
rect 500 607 556 619
rect 500 573 511 607
rect 545 573 556 607
rect 500 505 556 573
rect 500 471 511 505
rect 545 471 556 505
rect 500 367 556 471
rect 586 599 642 619
rect 586 565 597 599
rect 631 565 642 599
rect 586 526 642 565
rect 586 492 597 526
rect 631 492 642 526
rect 586 453 642 492
rect 586 419 597 453
rect 631 419 642 453
rect 586 367 642 419
rect 672 585 699 619
rect 733 585 760 619
rect 672 551 760 585
rect 672 517 699 551
rect 733 517 760 551
rect 672 367 760 517
rect 790 599 846 619
rect 790 565 801 599
rect 835 565 846 599
rect 790 501 846 565
rect 790 467 801 501
rect 835 467 846 501
rect 790 367 846 467
rect 876 547 932 619
rect 876 513 887 547
rect 921 513 932 547
rect 876 479 932 513
rect 876 445 887 479
rect 921 445 932 479
rect 876 411 932 445
rect 876 377 887 411
rect 921 377 932 411
rect 876 367 932 377
rect 962 599 1018 619
rect 962 565 973 599
rect 1007 565 1018 599
rect 962 501 1018 565
rect 962 467 973 501
rect 1007 467 1018 501
rect 962 367 1018 467
rect 1048 547 1104 619
rect 1048 513 1059 547
rect 1093 513 1104 547
rect 1048 428 1104 513
rect 1048 394 1059 428
rect 1093 394 1104 428
rect 1048 367 1104 394
rect 1134 599 1187 619
rect 1134 565 1145 599
rect 1179 565 1187 599
rect 1134 513 1187 565
rect 1134 479 1145 513
rect 1179 479 1187 513
rect 1134 428 1187 479
rect 1134 394 1145 428
rect 1179 394 1187 428
rect 1134 367 1187 394
rect 1241 599 1294 619
rect 1241 565 1249 599
rect 1283 565 1294 599
rect 1241 517 1294 565
rect 1241 483 1249 517
rect 1283 483 1294 517
rect 1241 436 1294 483
rect 1241 402 1249 436
rect 1283 402 1294 436
rect 1241 367 1294 402
rect 1324 611 1380 619
rect 1324 577 1335 611
rect 1369 577 1380 611
rect 1324 492 1380 577
rect 1324 458 1335 492
rect 1369 458 1380 492
rect 1324 367 1380 458
rect 1410 599 1466 619
rect 1410 565 1421 599
rect 1455 565 1466 599
rect 1410 517 1466 565
rect 1410 483 1421 517
rect 1455 483 1466 517
rect 1410 436 1466 483
rect 1410 402 1421 436
rect 1455 402 1466 436
rect 1410 367 1466 402
rect 1496 607 1552 619
rect 1496 573 1507 607
rect 1541 573 1552 607
rect 1496 492 1552 573
rect 1496 458 1507 492
rect 1541 458 1552 492
rect 1496 367 1552 458
rect 1582 599 1638 619
rect 1582 565 1593 599
rect 1627 565 1638 599
rect 1582 517 1638 565
rect 1582 483 1593 517
rect 1627 483 1638 517
rect 1582 436 1638 483
rect 1582 402 1593 436
rect 1627 402 1638 436
rect 1582 367 1638 402
rect 1668 531 1724 619
rect 1668 497 1679 531
rect 1713 497 1724 531
rect 1668 413 1724 497
rect 1668 379 1679 413
rect 1713 379 1724 413
rect 1668 367 1724 379
rect 1754 599 1810 619
rect 1754 565 1765 599
rect 1799 565 1810 599
rect 1754 529 1810 565
rect 1754 495 1765 529
rect 1799 495 1810 529
rect 1754 459 1810 495
rect 1754 425 1765 459
rect 1799 425 1810 459
rect 1754 367 1810 425
rect 1840 531 1896 619
rect 1840 497 1851 531
rect 1885 497 1896 531
rect 1840 413 1896 497
rect 1840 379 1851 413
rect 1885 379 1896 413
rect 1840 367 1896 379
rect 1926 599 1979 619
rect 1926 565 1937 599
rect 1971 565 1979 599
rect 1926 529 1979 565
rect 1926 495 1937 529
rect 1971 495 1979 529
rect 1926 459 1979 495
rect 1926 425 1937 459
rect 1971 425 1979 459
rect 1926 367 1979 425
<< ndiffc >>
rect 82 169 116 203
rect 82 59 116 93
rect 168 173 202 207
rect 168 67 202 101
rect 254 134 288 168
rect 254 55 288 89
rect 340 173 374 207
rect 340 67 374 101
rect 426 161 460 195
rect 512 67 546 101
rect 598 161 632 195
rect 684 67 718 101
rect 778 76 812 110
rect 873 169 907 203
rect 873 67 907 101
rect 959 139 993 173
rect 959 55 993 89
rect 1045 169 1079 203
rect 1045 67 1079 101
rect 1131 141 1165 175
rect 1131 55 1165 89
rect 1217 169 1251 203
rect 1217 101 1251 135
rect 1303 127 1337 161
rect 1303 59 1337 93
rect 1389 169 1423 203
rect 1389 67 1423 101
rect 1475 140 1509 174
rect 1579 90 1613 124
rect 1475 55 1509 89
rect 1665 158 1699 192
rect 1665 67 1699 101
rect 1751 90 1785 124
rect 1837 169 1871 203
rect 1837 67 1871 101
rect 1923 133 1957 167
rect 1923 59 1957 93
<< pdiffc >>
rect 81 565 115 599
rect 81 471 115 505
rect 81 379 115 413
rect 167 573 201 607
rect 167 496 201 530
rect 167 413 201 447
rect 253 565 287 599
rect 253 471 287 505
rect 253 379 287 413
rect 339 573 373 607
rect 339 471 373 505
rect 425 565 459 599
rect 425 492 459 526
rect 425 419 459 453
rect 511 573 545 607
rect 511 471 545 505
rect 597 565 631 599
rect 597 492 631 526
rect 597 419 631 453
rect 699 585 733 619
rect 699 517 733 551
rect 801 565 835 599
rect 801 467 835 501
rect 887 513 921 547
rect 887 445 921 479
rect 887 377 921 411
rect 973 565 1007 599
rect 973 467 1007 501
rect 1059 513 1093 547
rect 1059 394 1093 428
rect 1145 565 1179 599
rect 1145 479 1179 513
rect 1145 394 1179 428
rect 1249 565 1283 599
rect 1249 483 1283 517
rect 1249 402 1283 436
rect 1335 577 1369 611
rect 1335 458 1369 492
rect 1421 565 1455 599
rect 1421 483 1455 517
rect 1421 402 1455 436
rect 1507 573 1541 607
rect 1507 458 1541 492
rect 1593 565 1627 599
rect 1593 483 1627 517
rect 1593 402 1627 436
rect 1679 497 1713 531
rect 1679 379 1713 413
rect 1765 565 1799 599
rect 1765 495 1799 529
rect 1765 425 1799 459
rect 1851 497 1885 531
rect 1851 379 1885 413
rect 1937 565 1971 599
rect 1937 495 1971 529
rect 1937 425 1971 459
<< poly >>
rect 126 619 156 645
rect 212 619 242 645
rect 298 619 328 645
rect 384 619 414 645
rect 470 619 500 645
rect 556 619 586 645
rect 642 619 672 645
rect 760 619 790 645
rect 846 619 876 645
rect 932 619 962 645
rect 1018 619 1048 645
rect 1104 619 1134 645
rect 1294 619 1324 645
rect 1380 619 1410 645
rect 1466 619 1496 645
rect 1552 619 1582 645
rect 1638 619 1668 645
rect 1724 619 1754 645
rect 1810 619 1840 645
rect 1896 619 1926 645
rect 126 325 156 367
rect 212 325 242 367
rect 298 325 328 367
rect 59 309 329 325
rect 59 275 75 309
rect 109 275 143 309
rect 177 275 211 309
rect 245 275 279 309
rect 313 275 329 309
rect 59 259 329 275
rect 127 215 157 259
rect 213 215 243 259
rect 299 215 329 259
rect 384 313 414 367
rect 470 313 500 367
rect 556 313 586 367
rect 642 313 672 367
rect 384 297 672 313
rect 760 308 790 367
rect 846 331 876 367
rect 932 331 962 367
rect 1018 331 1048 367
rect 1104 331 1134 367
rect 1294 335 1324 367
rect 1380 335 1410 367
rect 1466 335 1496 367
rect 1552 335 1582 367
rect 384 263 413 297
rect 447 263 481 297
rect 515 263 549 297
rect 583 263 617 297
rect 651 277 672 297
rect 715 292 790 308
rect 651 263 673 277
rect 384 247 673 263
rect 385 215 415 247
rect 471 215 501 247
rect 557 215 587 247
rect 643 215 673 247
rect 715 258 731 292
rect 765 278 790 292
rect 832 315 1134 331
rect 832 281 883 315
rect 917 281 987 315
rect 1021 281 1134 315
rect 765 258 781 278
rect 715 242 781 258
rect 832 265 1134 281
rect 1176 319 1582 335
rect 1638 321 1668 367
rect 1724 321 1754 367
rect 1810 321 1840 367
rect 1896 321 1926 367
rect 1176 285 1260 319
rect 1294 285 1328 319
rect 1362 285 1396 319
rect 1430 285 1464 319
rect 1498 285 1532 319
rect 1566 285 1582 319
rect 1176 269 1582 285
rect 1624 305 1926 321
rect 1624 271 1658 305
rect 1692 271 1726 305
rect 1760 271 1794 305
rect 1828 271 1862 305
rect 1896 271 1926 305
rect 729 215 759 242
rect 832 215 862 265
rect 918 215 948 265
rect 1004 215 1034 265
rect 1090 215 1120 265
rect 1176 215 1206 269
rect 1262 215 1292 269
rect 1348 215 1378 269
rect 1434 215 1464 269
rect 1624 255 1926 271
rect 1624 215 1654 255
rect 1710 215 1740 255
rect 1796 215 1826 255
rect 1882 215 1912 255
rect 127 21 157 47
rect 213 21 243 47
rect 299 21 329 47
rect 385 21 415 47
rect 471 21 501 47
rect 557 21 587 47
rect 643 21 673 47
rect 729 21 759 47
rect 832 21 862 47
rect 918 21 948 47
rect 1004 21 1034 47
rect 1090 21 1120 47
rect 1176 21 1206 47
rect 1262 21 1292 47
rect 1348 21 1378 47
rect 1434 21 1464 47
rect 1624 21 1654 47
rect 1710 21 1740 47
rect 1796 21 1826 47
rect 1882 21 1912 47
<< polycont >>
rect 75 275 109 309
rect 143 275 177 309
rect 211 275 245 309
rect 279 275 313 309
rect 413 263 447 297
rect 481 263 515 297
rect 549 263 583 297
rect 617 263 651 297
rect 731 258 765 292
rect 883 281 917 315
rect 987 281 1021 315
rect 1260 285 1294 319
rect 1328 285 1362 319
rect 1396 285 1430 319
rect 1464 285 1498 319
rect 1532 285 1566 319
rect 1658 271 1692 305
rect 1726 271 1760 305
rect 1794 271 1828 305
rect 1862 271 1896 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 65 599 117 615
rect 65 565 81 599
rect 115 565 117 599
rect 65 505 117 565
rect 65 471 81 505
rect 115 471 117 505
rect 65 413 117 471
rect 151 607 217 649
rect 151 573 167 607
rect 201 573 217 607
rect 151 530 217 573
rect 151 496 167 530
rect 201 496 217 530
rect 151 447 217 496
rect 151 413 167 447
rect 201 413 217 447
rect 251 599 289 615
rect 251 565 253 599
rect 287 565 289 599
rect 251 505 289 565
rect 251 471 253 505
rect 287 471 289 505
rect 323 607 389 649
rect 323 573 339 607
rect 373 573 389 607
rect 323 505 389 573
rect 323 471 339 505
rect 373 471 389 505
rect 423 599 461 615
rect 423 565 425 599
rect 459 565 461 599
rect 423 526 461 565
rect 423 492 425 526
rect 459 492 461 526
rect 251 437 289 471
rect 423 453 461 492
rect 495 607 561 649
rect 683 619 749 649
rect 495 573 511 607
rect 545 573 561 607
rect 495 505 561 573
rect 495 471 511 505
rect 545 471 561 505
rect 595 599 635 615
rect 595 565 597 599
rect 631 565 635 599
rect 595 526 635 565
rect 595 492 597 526
rect 631 492 635 526
rect 683 585 699 619
rect 733 585 749 619
rect 683 551 749 585
rect 683 517 699 551
rect 733 517 749 551
rect 783 599 1195 615
rect 783 565 801 599
rect 835 581 973 599
rect 835 565 837 581
rect 595 483 635 492
rect 783 501 837 565
rect 971 565 973 581
rect 1007 581 1145 599
rect 1007 565 1009 581
rect 783 485 801 501
rect 769 483 801 485
rect 423 437 425 453
rect 251 419 425 437
rect 459 437 461 453
rect 595 467 801 483
rect 835 467 837 501
rect 595 453 837 467
rect 595 437 597 453
rect 459 419 597 437
rect 631 451 837 453
rect 871 513 887 547
rect 921 513 937 547
rect 871 479 937 513
rect 631 449 781 451
rect 631 419 743 449
rect 251 413 743 419
rect 871 445 887 479
rect 921 445 937 479
rect 971 501 1009 565
rect 1143 565 1145 581
rect 1179 565 1195 599
rect 971 467 973 501
rect 1007 467 1009 501
rect 971 451 1009 467
rect 1043 513 1059 547
rect 1093 513 1109 547
rect 871 417 937 445
rect 1043 428 1109 513
rect 1043 417 1059 428
rect 65 379 81 413
rect 115 379 117 413
rect 251 379 253 413
rect 287 403 743 413
rect 799 411 1059 417
rect 287 379 293 403
rect 65 345 293 379
rect 799 377 887 411
rect 921 394 1059 411
rect 1093 394 1109 428
rect 921 378 1109 394
rect 1143 513 1195 565
rect 1143 479 1145 513
rect 1179 479 1195 513
rect 1143 428 1195 479
rect 1143 394 1145 428
rect 1179 394 1195 428
rect 1143 378 1195 394
rect 1233 599 1285 615
rect 1233 565 1249 599
rect 1283 565 1285 599
rect 1233 517 1285 565
rect 1233 483 1249 517
rect 1283 483 1285 517
rect 1233 436 1285 483
rect 1319 611 1385 649
rect 1319 577 1335 611
rect 1369 577 1385 611
rect 1319 492 1385 577
rect 1319 458 1335 492
rect 1369 458 1385 492
rect 1319 454 1385 458
rect 1419 599 1457 615
rect 1419 565 1421 599
rect 1455 565 1457 599
rect 1419 517 1457 565
rect 1419 483 1421 517
rect 1455 483 1457 517
rect 1233 402 1249 436
rect 1283 420 1285 436
rect 1419 436 1457 483
rect 1491 607 1557 649
rect 1491 573 1507 607
rect 1541 573 1557 607
rect 1491 492 1557 573
rect 1491 458 1507 492
rect 1541 458 1557 492
rect 1491 454 1557 458
rect 1591 599 1987 615
rect 1591 565 1593 599
rect 1627 581 1765 599
rect 1627 565 1634 581
rect 1591 517 1634 565
rect 1757 565 1765 581
rect 1799 581 1937 599
rect 1799 565 1809 581
rect 1591 483 1593 517
rect 1627 483 1634 517
rect 1419 420 1421 436
rect 1283 402 1421 420
rect 1455 420 1457 436
rect 1591 436 1634 483
rect 1591 420 1593 436
rect 1455 402 1593 420
rect 1627 402 1634 436
rect 1233 386 1634 402
rect 1668 531 1723 547
rect 1668 497 1679 531
rect 1713 497 1723 531
rect 1668 413 1723 497
rect 1668 379 1679 413
rect 1713 379 1723 413
rect 1757 529 1809 565
rect 1929 565 1937 581
rect 1971 565 1987 599
rect 1757 495 1765 529
rect 1799 495 1809 529
rect 1757 459 1809 495
rect 1757 425 1765 459
rect 1799 425 1809 459
rect 1757 409 1809 425
rect 1843 531 1895 547
rect 1843 497 1851 531
rect 1885 497 1895 531
rect 1843 413 1895 497
rect 921 377 954 378
rect 327 333 765 367
rect 327 311 361 333
rect 59 309 361 311
rect 59 275 75 309
rect 109 275 143 309
rect 177 275 211 309
rect 245 275 279 309
rect 313 275 361 309
rect 59 270 361 275
rect 397 263 413 297
rect 447 263 481 297
rect 515 263 549 297
rect 583 263 617 297
rect 651 263 667 297
rect 408 240 667 263
rect 701 292 765 333
rect 701 258 731 292
rect 701 240 765 258
rect 66 203 124 219
rect 66 169 82 203
rect 116 169 124 203
rect 66 93 124 169
rect 66 59 82 93
rect 116 59 124 93
rect 66 17 124 59
rect 158 207 374 236
rect 158 173 168 207
rect 202 202 340 207
rect 202 173 204 202
rect 158 101 204 173
rect 338 173 340 202
rect 799 206 833 377
rect 1668 375 1723 379
rect 1843 379 1851 413
rect 1885 379 1895 413
rect 1929 529 1987 565
rect 1929 495 1937 529
rect 1971 495 1987 529
rect 1929 459 1987 495
rect 1929 425 1937 459
rect 1971 425 1987 459
rect 1929 409 1987 425
rect 1843 375 1895 379
rect 988 343 1210 344
rect 867 315 1210 343
rect 867 281 883 315
rect 917 281 987 315
rect 1021 310 1210 315
rect 1021 281 1037 310
rect 867 277 1037 281
rect 1071 243 1140 276
rect 869 209 1140 243
rect 1176 247 1210 310
rect 1244 319 1608 351
rect 1668 339 1987 375
rect 1244 285 1260 319
rect 1294 285 1328 319
rect 1362 285 1396 319
rect 1430 285 1464 319
rect 1498 285 1532 319
rect 1566 285 1608 319
rect 1244 281 1608 285
rect 1642 271 1658 305
rect 1692 271 1726 305
rect 1760 271 1794 305
rect 1828 271 1862 305
rect 1896 271 1912 305
rect 1642 269 1912 271
rect 1176 213 1608 247
rect 1642 242 1793 269
rect 1946 235 1987 339
rect 869 206 909 209
rect 158 67 168 101
rect 202 67 204 101
rect 158 51 204 67
rect 238 134 254 168
rect 288 134 304 168
rect 238 89 304 134
rect 238 55 254 89
rect 288 55 304 89
rect 238 17 304 55
rect 338 117 374 173
rect 410 203 909 206
rect 410 195 873 203
rect 410 161 426 195
rect 460 161 598 195
rect 632 169 873 195
rect 907 169 909 203
rect 1043 203 1081 209
rect 632 161 909 169
rect 410 151 909 161
rect 338 101 728 117
rect 338 67 340 101
rect 374 67 512 101
rect 546 67 684 101
rect 718 67 728 101
rect 338 51 728 67
rect 762 110 828 117
rect 762 76 778 110
rect 812 76 828 110
rect 762 17 828 76
rect 862 101 909 151
rect 862 67 873 101
rect 907 67 909 101
rect 862 51 909 67
rect 943 139 959 173
rect 993 139 1009 173
rect 943 89 1009 139
rect 943 55 959 89
rect 993 55 1009 89
rect 943 17 1009 55
rect 1043 169 1045 203
rect 1079 169 1081 203
rect 1215 203 1253 213
rect 1043 101 1081 169
rect 1043 67 1045 101
rect 1079 67 1081 101
rect 1043 51 1081 67
rect 1115 141 1131 175
rect 1165 141 1181 175
rect 1115 89 1181 141
rect 1115 55 1131 89
rect 1165 55 1181 89
rect 1115 17 1181 55
rect 1215 169 1217 203
rect 1251 169 1253 203
rect 1387 208 1608 213
rect 1833 208 1987 235
rect 1387 203 1425 208
rect 1215 135 1253 169
rect 1215 101 1217 135
rect 1251 101 1253 135
rect 1215 51 1253 101
rect 1287 161 1353 179
rect 1287 127 1303 161
rect 1337 127 1353 161
rect 1287 93 1353 127
rect 1287 59 1303 93
rect 1337 59 1353 93
rect 1287 17 1353 59
rect 1387 169 1389 203
rect 1423 169 1425 203
rect 1574 203 1987 208
rect 1574 192 1837 203
rect 1574 174 1665 192
rect 1387 101 1425 169
rect 1387 67 1389 101
rect 1423 67 1425 101
rect 1387 51 1425 67
rect 1459 140 1475 174
rect 1509 140 1525 174
rect 1661 158 1665 174
rect 1699 174 1837 192
rect 1699 158 1701 174
rect 1459 124 1627 140
rect 1459 90 1579 124
rect 1613 90 1627 124
rect 1459 89 1627 90
rect 1459 55 1475 89
rect 1509 55 1627 89
rect 1459 17 1627 55
rect 1661 101 1701 158
rect 1835 169 1837 174
rect 1871 201 1987 203
rect 1871 169 1873 201
rect 1661 67 1665 101
rect 1699 67 1701 101
rect 1661 51 1701 67
rect 1735 124 1801 140
rect 1735 90 1751 124
rect 1785 90 1801 124
rect 1735 17 1801 90
rect 1835 101 1873 169
rect 1835 67 1837 101
rect 1871 67 1873 101
rect 1835 51 1873 67
rect 1907 133 1923 167
rect 1957 133 1973 167
rect 1907 93 1973 133
rect 1907 59 1923 93
rect 1957 59 1973 93
rect 1907 17 1973 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2bb2oi_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3104868
string GDS_START 3088112
<< end >>
