magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 332 1670 704
<< pwell >>
rect 871 274 1631 275
rect 1 228 333 272
rect 657 228 1631 274
rect 1 49 1631 228
rect 0 0 1632 49
<< scpmos >>
rect 81 368 117 592
rect 217 368 253 496
rect 419 394 455 562
rect 540 394 576 562
rect 754 368 790 592
rect 973 373 1009 541
rect 1080 383 1116 511
rect 1170 383 1206 511
rect 1297 383 1333 551
rect 1405 383 1441 583
rect 1512 383 1548 583
<< nmoslvt >>
rect 84 98 114 246
rect 202 162 232 246
rect 428 74 458 202
rect 528 74 558 202
rect 756 100 786 248
rect 979 121 1009 249
rect 1092 121 1122 249
rect 1204 165 1234 249
rect 1303 121 1333 249
rect 1402 121 1432 249
rect 1518 121 1548 249
<< ndiff >>
rect 27 218 84 246
rect 27 184 39 218
rect 73 184 84 218
rect 27 144 84 184
rect 27 110 39 144
rect 73 110 84 144
rect 27 98 84 110
rect 114 162 202 246
rect 232 234 307 246
rect 232 200 243 234
rect 277 200 307 234
rect 232 162 307 200
rect 371 179 428 202
rect 114 98 187 162
rect 371 145 383 179
rect 417 145 428 179
rect 129 82 187 98
rect 129 48 141 82
rect 175 48 187 82
rect 371 74 428 145
rect 458 194 528 202
rect 458 160 483 194
rect 517 160 528 194
rect 458 126 528 160
rect 458 92 483 126
rect 517 92 528 126
rect 458 74 528 92
rect 558 188 629 202
rect 558 154 583 188
rect 617 154 629 188
rect 558 120 629 154
rect 558 86 569 120
rect 603 86 629 120
rect 558 74 629 86
rect 683 100 756 248
rect 786 236 843 248
rect 786 202 797 236
rect 831 202 843 236
rect 786 100 843 202
rect 897 121 979 249
rect 1009 237 1092 249
rect 1009 203 1033 237
rect 1067 203 1092 237
rect 1009 121 1092 203
rect 1122 237 1204 249
rect 1122 203 1155 237
rect 1189 203 1204 237
rect 1122 165 1204 203
rect 1234 226 1303 249
rect 1234 192 1258 226
rect 1292 192 1303 226
rect 1234 165 1303 192
rect 1122 121 1172 165
rect 897 100 964 121
rect 683 84 741 100
rect 683 50 695 84
rect 729 50 741 84
rect 897 66 913 100
rect 947 66 964 100
rect 897 54 964 66
rect 129 36 187 48
rect 683 38 741 50
rect 1253 121 1303 165
rect 1333 235 1402 249
rect 1333 201 1357 235
rect 1391 201 1402 235
rect 1333 167 1402 201
rect 1333 133 1357 167
rect 1391 133 1402 167
rect 1333 121 1402 133
rect 1432 167 1518 249
rect 1432 133 1465 167
rect 1499 133 1518 167
rect 1432 121 1518 133
rect 1548 235 1605 249
rect 1548 201 1559 235
rect 1593 201 1605 235
rect 1548 167 1605 201
rect 1548 133 1559 167
rect 1593 133 1605 167
rect 1548 121 1605 133
<< pdiff >>
rect 685 592 739 604
rect 27 580 81 592
rect 27 546 37 580
rect 71 546 81 580
rect 27 499 81 546
rect 27 465 37 499
rect 71 465 81 499
rect 27 418 81 465
rect 27 384 37 418
rect 71 384 81 418
rect 27 368 81 384
rect 117 580 173 592
rect 117 546 127 580
rect 161 546 173 580
rect 470 576 525 588
rect 470 562 481 576
rect 117 508 173 546
rect 363 531 419 562
rect 117 474 127 508
rect 161 496 173 508
rect 363 497 375 531
rect 409 497 419 531
rect 161 474 217 496
rect 117 368 217 474
rect 253 462 309 496
rect 253 428 263 462
rect 297 428 309 462
rect 253 368 309 428
rect 363 440 419 497
rect 363 406 375 440
rect 409 406 419 440
rect 363 394 419 406
rect 455 542 481 562
rect 515 562 525 576
rect 515 542 540 562
rect 455 394 540 542
rect 576 440 631 562
rect 576 406 586 440
rect 620 406 631 440
rect 576 394 631 406
rect 685 558 695 592
rect 729 558 754 592
rect 685 368 754 558
rect 790 440 844 592
rect 790 406 800 440
rect 834 406 844 440
rect 790 368 844 406
rect 904 576 958 588
rect 904 542 914 576
rect 948 542 958 576
rect 904 541 958 542
rect 904 373 973 541
rect 1009 511 1065 541
rect 1353 551 1405 583
rect 1240 511 1297 551
rect 1009 499 1080 511
rect 1009 465 1019 499
rect 1053 465 1080 499
rect 1009 421 1080 465
rect 1009 387 1019 421
rect 1053 387 1080 421
rect 1009 383 1080 387
rect 1116 471 1170 511
rect 1116 437 1126 471
rect 1160 437 1170 471
rect 1116 383 1170 437
rect 1206 456 1297 511
rect 1206 422 1216 456
rect 1250 422 1297 456
rect 1206 383 1297 422
rect 1333 539 1405 551
rect 1333 505 1360 539
rect 1394 505 1405 539
rect 1333 440 1405 505
rect 1333 406 1360 440
rect 1394 406 1405 440
rect 1333 383 1405 406
rect 1441 569 1512 583
rect 1441 535 1468 569
rect 1502 535 1512 569
rect 1441 492 1512 535
rect 1441 458 1468 492
rect 1502 458 1512 492
rect 1441 383 1512 458
rect 1548 570 1605 583
rect 1548 536 1558 570
rect 1592 536 1605 570
rect 1548 488 1605 536
rect 1548 454 1558 488
rect 1592 454 1605 488
rect 1548 383 1605 454
rect 1009 373 1065 383
<< ndiffc >>
rect 39 184 73 218
rect 39 110 73 144
rect 243 200 277 234
rect 383 145 417 179
rect 141 48 175 82
rect 483 160 517 194
rect 483 92 517 126
rect 583 154 617 188
rect 569 86 603 120
rect 797 202 831 236
rect 1033 203 1067 237
rect 1155 203 1189 237
rect 1258 192 1292 226
rect 695 50 729 84
rect 913 66 947 100
rect 1357 201 1391 235
rect 1357 133 1391 167
rect 1465 133 1499 167
rect 1559 201 1593 235
rect 1559 133 1593 167
<< pdiffc >>
rect 37 546 71 580
rect 37 465 71 499
rect 37 384 71 418
rect 127 546 161 580
rect 127 474 161 508
rect 375 497 409 531
rect 263 428 297 462
rect 375 406 409 440
rect 481 542 515 576
rect 586 406 620 440
rect 695 558 729 592
rect 800 406 834 440
rect 914 542 948 576
rect 1019 465 1053 499
rect 1019 387 1053 421
rect 1126 437 1160 471
rect 1216 422 1250 456
rect 1360 505 1394 539
rect 1360 406 1394 440
rect 1468 535 1502 569
rect 1468 458 1502 492
rect 1558 536 1592 570
rect 1558 454 1592 488
<< poly >>
rect 81 592 117 618
rect 754 592 790 618
rect 859 615 1333 645
rect 419 562 455 588
rect 217 496 253 522
rect 540 562 576 588
rect 81 334 117 368
rect 217 336 253 368
rect 81 318 151 334
rect 81 284 101 318
rect 135 284 151 318
rect 81 268 151 284
rect 199 320 265 336
rect 199 286 215 320
rect 249 300 265 320
rect 419 300 455 394
rect 540 362 576 394
rect 503 346 576 362
rect 503 312 519 346
rect 553 312 576 346
rect 754 336 790 368
rect 859 336 889 615
rect 973 541 1009 567
rect 1080 511 1116 615
rect 1297 551 1333 615
rect 1405 583 1441 609
rect 1512 583 1548 609
rect 1170 511 1206 537
rect 973 337 1009 373
rect 1080 368 1116 383
rect 1080 338 1122 368
rect 249 286 449 300
rect 503 296 576 312
rect 741 320 889 336
rect 199 270 449 286
rect 84 246 114 268
rect 202 246 232 270
rect 419 247 449 270
rect 419 217 458 247
rect 428 202 458 217
rect 528 202 558 296
rect 741 286 757 320
rect 791 286 825 320
rect 859 286 889 320
rect 741 270 889 286
rect 943 321 1009 337
rect 943 287 959 321
rect 993 287 1009 321
rect 943 271 1009 287
rect 756 248 786 270
rect 979 249 1009 271
rect 1092 249 1122 338
rect 1170 294 1206 383
rect 1297 338 1333 383
rect 1405 351 1441 383
rect 1512 351 1548 383
rect 1170 264 1234 294
rect 1204 249 1234 264
rect 1303 249 1333 338
rect 1375 335 1441 351
rect 1375 301 1391 335
rect 1425 301 1441 335
rect 1375 285 1441 301
rect 1483 335 1549 351
rect 1483 301 1499 335
rect 1533 301 1549 335
rect 1483 285 1549 301
rect 1402 249 1432 285
rect 1518 249 1548 285
rect 202 136 232 162
rect 84 72 114 98
rect 428 48 458 74
rect 528 48 558 74
rect 756 74 786 100
rect 979 53 1009 121
rect 1092 95 1122 121
rect 1204 53 1234 165
rect 1303 95 1333 121
rect 1402 95 1432 121
rect 1518 95 1548 121
rect 979 23 1234 53
<< polycont >>
rect 101 284 135 318
rect 215 286 249 320
rect 519 312 553 346
rect 757 286 791 320
rect 825 286 859 320
rect 959 287 993 321
rect 1391 301 1425 335
rect 1499 301 1533 335
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 17 580 71 596
rect 17 546 37 580
rect 17 499 71 546
rect 17 465 37 499
rect 17 418 71 465
rect 111 580 161 649
rect 111 546 127 580
rect 111 508 161 546
rect 111 474 127 508
rect 111 458 161 474
rect 195 581 531 615
rect 195 424 229 581
rect 465 576 531 581
rect 375 531 425 547
rect 465 542 481 576
rect 515 542 531 576
rect 679 592 745 649
rect 679 558 695 592
rect 729 558 745 592
rect 679 542 745 558
rect 898 581 1418 615
rect 898 576 964 581
rect 898 542 914 576
rect 948 542 964 576
rect 17 384 37 418
rect 17 368 71 384
rect 123 390 229 424
rect 263 462 333 500
rect 297 428 333 462
rect 263 390 333 428
rect 409 508 425 531
rect 1003 508 1053 515
rect 409 499 1053 508
rect 409 497 1019 499
rect 375 474 1019 497
rect 375 440 425 474
rect 409 406 425 440
rect 570 406 586 440
rect 620 406 637 440
rect 375 390 425 406
rect 17 234 51 368
rect 123 334 157 390
rect 85 318 157 334
rect 85 284 101 318
rect 135 284 157 318
rect 85 268 157 284
rect 199 320 265 356
rect 199 286 215 320
rect 249 286 265 320
rect 199 270 265 286
rect 299 350 333 390
rect 503 350 569 362
rect 299 346 569 350
rect 299 316 519 346
rect 17 218 89 234
rect 17 184 39 218
rect 73 184 89 218
rect 17 144 89 184
rect 17 110 39 144
rect 73 110 89 144
rect 123 166 157 268
rect 299 234 333 316
rect 503 312 519 316
rect 553 312 569 346
rect 503 296 569 312
rect 227 200 243 234
rect 277 200 333 234
rect 367 276 455 282
rect 367 242 415 276
rect 449 262 455 276
rect 603 262 637 406
rect 449 242 637 262
rect 367 228 637 242
rect 367 179 433 228
rect 671 194 705 474
rect 1003 465 1019 474
rect 784 406 800 440
rect 834 406 943 440
rect 784 390 943 406
rect 741 320 875 356
rect 741 286 757 320
rect 791 286 825 320
rect 859 286 875 320
rect 741 270 875 286
rect 909 337 943 390
rect 1003 421 1053 465
rect 1110 513 1318 547
rect 1110 471 1176 513
rect 1110 437 1126 471
rect 1160 437 1176 471
rect 1110 421 1176 437
rect 1216 456 1250 479
rect 1003 387 1019 421
rect 1216 387 1250 422
rect 1003 371 1053 387
rect 1087 353 1250 387
rect 909 321 1009 337
rect 909 287 959 321
rect 993 287 1009 321
rect 909 271 1009 287
rect 1087 282 1121 353
rect 1284 319 1318 513
rect 1352 539 1418 581
rect 1352 505 1360 539
rect 1394 505 1418 539
rect 1352 440 1418 505
rect 1452 569 1518 649
rect 1452 535 1468 569
rect 1502 535 1518 569
rect 1452 492 1518 535
rect 1452 458 1468 492
rect 1502 458 1518 492
rect 1558 570 1615 586
rect 1592 536 1615 570
rect 1558 488 1615 536
rect 1352 406 1360 440
rect 1394 424 1418 440
rect 1592 454 1615 488
rect 1558 438 1615 454
rect 1394 406 1524 424
rect 1352 390 1524 406
rect 1063 276 1121 282
rect 909 236 943 271
rect 1063 242 1087 276
rect 1063 237 1121 242
rect 781 202 797 236
rect 831 202 943 236
rect 1004 203 1033 237
rect 1067 236 1121 237
rect 1155 285 1318 319
rect 1369 335 1441 356
rect 1369 301 1391 335
rect 1425 301 1441 335
rect 1369 285 1441 301
rect 1483 351 1524 390
rect 1483 335 1533 351
rect 1483 301 1499 335
rect 1483 285 1533 301
rect 1155 276 1217 285
rect 1155 242 1183 276
rect 1483 251 1524 285
rect 1567 276 1615 438
rect 1155 237 1217 242
rect 1067 203 1097 236
rect 1189 203 1217 237
rect 123 132 333 166
rect 17 88 89 110
rect 125 82 191 98
rect 125 48 141 82
rect 175 48 191 82
rect 299 85 333 132
rect 367 145 383 179
rect 417 145 433 179
rect 367 119 433 145
rect 467 160 483 194
rect 517 160 533 194
rect 467 126 533 160
rect 467 92 483 126
rect 517 92 533 126
rect 467 85 533 92
rect 299 51 533 85
rect 567 188 705 194
rect 567 154 583 188
rect 617 168 705 188
rect 1155 187 1217 203
rect 1251 226 1307 242
rect 1251 192 1258 226
rect 1292 192 1307 226
rect 617 154 1036 168
rect 567 153 1036 154
rect 1251 153 1307 192
rect 567 134 1307 153
rect 567 120 633 134
rect 567 86 569 120
rect 603 86 633 120
rect 1002 119 1307 134
rect 1341 235 1524 251
rect 1341 201 1357 235
rect 1391 217 1524 235
rect 1559 242 1567 251
rect 1601 242 1615 276
rect 1559 235 1615 242
rect 1391 201 1407 217
rect 1341 167 1407 201
rect 1593 201 1615 235
rect 1341 133 1357 167
rect 1391 133 1407 167
rect 567 70 633 86
rect 679 84 745 100
rect 125 17 191 48
rect 679 50 695 84
rect 729 50 745 84
rect 893 66 913 100
rect 947 85 968 100
rect 1341 85 1407 133
rect 947 66 1407 85
rect 893 51 1407 66
rect 1441 167 1523 183
rect 1441 133 1465 167
rect 1499 133 1523 167
rect 679 17 745 50
rect 1441 17 1523 133
rect 1559 167 1615 201
rect 1593 133 1615 167
rect 1559 117 1615 133
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 415 242 449 276
rect 1087 242 1121 276
rect 1183 242 1217 276
rect 1567 242 1601 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 403 276 461 282
rect 403 242 415 276
rect 449 273 461 276
rect 1075 276 1133 282
rect 1075 273 1087 276
rect 449 245 1087 273
rect 449 242 461 245
rect 403 236 461 242
rect 1075 242 1087 245
rect 1121 242 1133 276
rect 1075 236 1133 242
rect 1171 276 1229 282
rect 1171 242 1183 276
rect 1217 273 1229 276
rect 1555 276 1613 282
rect 1555 273 1567 276
rect 1217 245 1567 273
rect 1217 242 1229 245
rect 1171 236 1229 242
rect 1555 242 1567 245
rect 1601 242 1613 276
rect 1555 236 1613 242
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xnor3_1
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 712606
string GDS_START 700458
<< end >>
