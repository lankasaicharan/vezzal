magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2770 1852
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 79 21 1417 203
rect 29 -17 63 17
<< scnmos >>
rect 168 47 198 177
rect 264 47 294 177
rect 360 47 390 177
rect 469 47 499 177
rect 566 47 596 177
rect 660 47 690 177
rect 777 47 807 177
rect 895 47 925 177
rect 1021 47 1051 177
rect 1107 47 1137 177
rect 1213 47 1243 177
rect 1299 47 1329 177
<< scpmoshvt >>
rect 81 297 117 497
rect 177 297 213 497
rect 273 297 309 497
rect 369 297 405 497
rect 577 297 613 497
rect 673 297 709 497
rect 769 297 805 497
rect 873 297 909 497
rect 991 297 1027 497
rect 1109 297 1145 497
rect 1205 297 1241 497
rect 1301 297 1337 497
<< ndiff >>
rect 105 93 168 177
rect 105 59 123 93
rect 157 59 168 93
rect 105 47 168 59
rect 198 101 264 177
rect 198 67 219 101
rect 253 67 264 101
rect 198 47 264 67
rect 294 89 360 177
rect 294 55 315 89
rect 349 55 360 89
rect 294 47 360 55
rect 390 101 469 177
rect 390 67 411 101
rect 445 67 469 101
rect 390 47 469 67
rect 499 89 566 177
rect 499 55 511 89
rect 545 55 566 89
rect 499 47 566 55
rect 596 114 660 177
rect 596 80 607 114
rect 641 80 660 114
rect 596 47 660 80
rect 690 89 777 177
rect 690 55 714 89
rect 748 55 777 89
rect 690 47 777 55
rect 807 161 895 177
rect 807 127 830 161
rect 864 127 895 161
rect 807 93 895 127
rect 807 59 830 93
rect 864 59 895 93
rect 807 47 895 59
rect 925 89 1021 177
rect 925 55 944 89
rect 978 55 1021 89
rect 925 47 1021 55
rect 1051 47 1107 177
rect 1137 157 1213 177
rect 1137 123 1158 157
rect 1192 123 1213 157
rect 1137 89 1213 123
rect 1137 55 1158 89
rect 1192 55 1213 89
rect 1137 47 1213 55
rect 1243 47 1299 177
rect 1329 161 1391 177
rect 1329 127 1349 161
rect 1383 127 1391 161
rect 1329 93 1391 127
rect 1329 59 1349 93
rect 1383 59 1391 93
rect 1329 47 1391 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 409 81 451
rect 27 375 35 409
rect 69 375 81 409
rect 27 297 81 375
rect 117 477 177 497
rect 117 443 130 477
rect 164 443 177 477
rect 117 388 177 443
rect 117 354 130 388
rect 164 354 177 388
rect 117 297 177 354
rect 213 485 273 497
rect 213 451 226 485
rect 260 451 273 485
rect 213 409 273 451
rect 213 375 226 409
rect 260 375 273 409
rect 213 297 273 375
rect 309 477 369 497
rect 309 443 322 477
rect 356 443 369 477
rect 309 388 369 443
rect 309 354 322 388
rect 356 354 369 388
rect 309 297 369 354
rect 405 485 459 497
rect 405 451 417 485
rect 451 451 459 485
rect 405 417 459 451
rect 405 383 417 417
rect 451 383 459 417
rect 405 297 459 383
rect 523 485 577 497
rect 523 451 531 485
rect 565 451 577 485
rect 523 297 577 451
rect 613 297 673 497
rect 709 408 769 497
rect 709 374 722 408
rect 756 374 769 408
rect 709 297 769 374
rect 805 297 873 497
rect 909 485 991 497
rect 909 451 930 485
rect 964 451 991 485
rect 909 417 991 451
rect 909 383 930 417
rect 964 383 991 417
rect 909 297 991 383
rect 1027 489 1109 497
rect 1027 455 1040 489
rect 1074 455 1109 489
rect 1027 297 1109 455
rect 1145 477 1205 497
rect 1145 443 1158 477
rect 1192 443 1205 477
rect 1145 297 1205 443
rect 1241 489 1301 497
rect 1241 455 1254 489
rect 1288 455 1301 489
rect 1241 297 1301 455
rect 1337 477 1391 497
rect 1337 443 1349 477
rect 1383 443 1391 477
rect 1337 343 1391 443
rect 1337 309 1349 343
rect 1383 309 1391 343
rect 1337 297 1391 309
<< ndiffc >>
rect 123 59 157 93
rect 219 67 253 101
rect 315 55 349 89
rect 411 67 445 101
rect 511 55 545 89
rect 607 80 641 114
rect 714 55 748 89
rect 830 127 864 161
rect 830 59 864 93
rect 944 55 978 89
rect 1158 123 1192 157
rect 1158 55 1192 89
rect 1349 127 1383 161
rect 1349 59 1383 93
<< pdiffc >>
rect 35 451 69 485
rect 35 375 69 409
rect 130 443 164 477
rect 130 354 164 388
rect 226 451 260 485
rect 226 375 260 409
rect 322 443 356 477
rect 322 354 356 388
rect 417 451 451 485
rect 417 383 451 417
rect 531 451 565 485
rect 722 374 756 408
rect 930 451 964 485
rect 930 383 964 417
rect 1040 455 1074 489
rect 1158 443 1192 477
rect 1254 455 1288 489
rect 1349 443 1383 477
rect 1349 309 1383 343
<< poly >>
rect 81 497 117 523
rect 177 497 213 523
rect 273 497 309 523
rect 369 497 405 523
rect 577 497 613 523
rect 673 497 709 523
rect 769 497 805 523
rect 873 497 909 523
rect 991 497 1027 523
rect 1109 497 1145 523
rect 1205 497 1241 523
rect 1301 497 1337 523
rect 81 282 117 297
rect 177 282 213 297
rect 273 282 309 297
rect 369 282 405 297
rect 577 282 613 297
rect 673 282 709 297
rect 769 282 805 297
rect 873 282 909 297
rect 991 282 1027 297
rect 1109 282 1145 297
rect 1205 282 1241 297
rect 1301 282 1337 297
rect 79 270 119 282
rect 175 270 215 282
rect 271 270 311 282
rect 367 270 407 282
rect 575 270 615 282
rect 671 271 711 282
rect 767 271 807 282
rect 79 249 499 270
rect 79 215 141 249
rect 175 215 219 249
rect 253 215 287 249
rect 321 215 365 249
rect 399 215 499 249
rect 79 204 499 215
rect 542 249 618 270
rect 542 215 558 249
rect 592 215 618 249
rect 542 204 618 215
rect 660 249 807 271
rect 871 270 911 282
rect 989 280 1029 282
rect 660 215 671 249
rect 705 215 749 249
rect 783 215 807 249
rect 168 177 198 204
rect 264 177 294 204
rect 360 177 390 204
rect 469 177 499 204
rect 566 177 596 204
rect 660 198 807 215
rect 660 177 690 198
rect 777 177 807 198
rect 849 249 925 270
rect 849 215 865 249
rect 899 215 925 249
rect 849 197 925 215
rect 989 249 1065 280
rect 989 215 1005 249
rect 1039 215 1065 249
rect 989 204 1065 215
rect 1107 270 1147 282
rect 1203 270 1243 282
rect 1107 249 1243 270
rect 1107 215 1123 249
rect 1157 215 1243 249
rect 1107 204 1243 215
rect 895 177 925 197
rect 1021 177 1051 204
rect 1107 177 1137 204
rect 1213 177 1243 204
rect 1299 270 1339 282
rect 1299 249 1375 270
rect 1299 215 1315 249
rect 1349 215 1375 249
rect 1299 202 1375 215
rect 1299 177 1329 202
rect 168 21 198 47
rect 264 21 294 47
rect 360 21 390 47
rect 469 21 499 47
rect 566 21 596 47
rect 660 21 690 47
rect 777 21 807 47
rect 895 21 925 47
rect 1021 21 1051 47
rect 1107 21 1137 47
rect 1213 21 1243 47
rect 1299 21 1329 47
<< polycont >>
rect 141 215 175 249
rect 219 215 253 249
rect 287 215 321 249
rect 365 215 399 249
rect 558 215 592 249
rect 671 215 705 249
rect 749 215 783 249
rect 865 215 899 249
rect 1005 215 1039 249
rect 1123 215 1157 249
rect 1315 215 1349 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 18 485 85 527
rect 18 451 35 485
rect 69 451 85 485
rect 18 409 85 451
rect 18 375 35 409
rect 69 375 85 409
rect 129 477 166 493
rect 129 443 130 477
rect 164 443 166 477
rect 129 388 166 443
rect 129 354 130 388
rect 164 354 166 388
rect 210 485 276 527
rect 210 451 226 485
rect 260 451 276 485
rect 210 409 276 451
rect 210 375 226 409
rect 260 375 276 409
rect 320 477 358 493
rect 320 443 322 477
rect 356 443 358 477
rect 320 388 358 443
rect 129 341 166 354
rect 320 354 322 388
rect 356 354 358 388
rect 402 485 452 527
rect 402 451 417 485
rect 451 451 452 485
rect 402 417 452 451
rect 514 485 980 493
rect 514 451 531 485
rect 565 451 930 485
rect 964 451 980 485
rect 1014 489 1090 527
rect 1014 455 1040 489
rect 1074 455 1090 489
rect 1132 477 1194 493
rect 514 442 980 451
rect 402 383 417 417
rect 451 383 452 417
rect 914 421 980 442
rect 1132 443 1158 477
rect 1192 443 1194 477
rect 1228 489 1304 527
rect 1228 455 1254 489
rect 1288 455 1304 489
rect 1348 477 1399 493
rect 1132 421 1194 443
rect 1348 443 1349 477
rect 1383 443 1399 477
rect 1348 421 1399 443
rect 914 417 1399 421
rect 402 367 452 383
rect 506 374 722 408
rect 756 374 772 408
rect 914 383 930 417
rect 964 383 1399 417
rect 914 376 1399 383
rect 320 341 358 354
rect 17 299 358 341
rect 506 335 541 374
rect 1323 343 1399 376
rect 477 301 541 335
rect 17 175 68 299
rect 477 265 524 301
rect 575 289 925 340
rect 575 265 621 289
rect 105 249 524 265
rect 105 215 141 249
rect 175 215 219 249
rect 253 215 287 249
rect 321 215 365 249
rect 399 215 524 249
rect 105 209 524 215
rect 17 127 445 175
rect 217 123 445 127
rect 479 161 524 209
rect 558 249 621 265
rect 592 215 621 249
rect 558 197 621 215
rect 655 249 809 255
rect 655 215 671 249
rect 705 215 749 249
rect 783 215 809 249
rect 655 197 809 215
rect 849 249 925 289
rect 849 215 865 249
rect 899 215 925 249
rect 849 197 925 215
rect 989 302 1289 340
rect 1323 309 1349 343
rect 1383 309 1399 343
rect 1323 307 1399 309
rect 989 249 1065 302
rect 989 215 1005 249
rect 1039 215 1065 249
rect 989 204 1065 215
rect 1107 249 1186 266
rect 1107 215 1123 249
rect 1157 215 1186 249
rect 1107 204 1186 215
rect 1225 264 1289 302
rect 1225 249 1375 264
rect 1225 215 1315 249
rect 1349 215 1375 249
rect 1225 204 1375 215
rect 479 127 830 161
rect 864 157 1208 161
rect 864 127 1158 157
rect 479 123 1158 127
rect 1192 123 1208 157
rect 217 101 255 123
rect 97 59 123 93
rect 157 59 173 93
rect 97 17 173 59
rect 217 67 219 101
rect 253 67 255 101
rect 409 101 445 123
rect 217 51 255 67
rect 289 55 315 89
rect 349 55 365 89
rect 289 17 365 55
rect 409 67 411 101
rect 605 114 654 123
rect 409 51 445 67
rect 484 55 511 89
rect 545 55 561 89
rect 484 17 561 55
rect 605 80 607 114
rect 641 80 654 114
rect 808 93 884 123
rect 605 51 654 80
rect 688 55 714 89
rect 748 55 764 89
rect 688 17 764 55
rect 808 59 830 93
rect 864 59 884 93
rect 1132 89 1208 123
rect 808 51 884 59
rect 928 55 944 89
rect 978 55 1002 89
rect 1132 55 1158 89
rect 1192 55 1208 89
rect 1323 127 1349 161
rect 1383 127 1399 161
rect 1323 93 1399 127
rect 1323 59 1349 93
rect 1383 59 1399 93
rect 928 17 1002 55
rect 1323 17 1399 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
flabel locali s 655 197 809 255 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 849 197 925 289 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 29 153 63 187 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 1225 264 1289 302 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1107 204 1186 266 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
rlabel comment s 0 0 0 0 4 a211o_4
rlabel locali s 1225 204 1375 264 1 A2
port 2 nsew signal input
rlabel locali s 989 302 1289 340 1 A2
port 2 nsew signal input
rlabel locali s 989 204 1065 302 1 A2
port 2 nsew signal input
rlabel locali s 575 289 925 340 1 B1
port 3 nsew signal input
rlabel locali s 575 265 621 289 1 B1
port 3 nsew signal input
rlabel locali s 558 197 621 265 1 B1
port 3 nsew signal input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1472 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 801778
string GDS_START 792110
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
