magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 43 49 575 251
rect 0 0 576 49
<< scnmos >>
rect 126 141 156 225
rect 204 141 234 225
rect 282 141 312 225
rect 390 141 420 225
rect 462 141 492 225
<< scpmoshvt >>
rect 100 416 150 616
rect 206 416 256 616
rect 312 416 362 616
rect 426 416 476 616
<< ndiff >>
rect 69 187 126 225
rect 69 153 81 187
rect 115 153 126 187
rect 69 141 126 153
rect 156 141 204 225
rect 234 141 282 225
rect 312 187 390 225
rect 312 153 323 187
rect 357 153 390 187
rect 312 141 390 153
rect 420 141 462 225
rect 492 208 549 225
rect 492 174 503 208
rect 537 174 549 208
rect 492 141 549 174
<< pdiff >>
rect 43 597 100 616
rect 43 563 55 597
rect 89 563 100 597
rect 43 467 100 563
rect 43 433 55 467
rect 89 433 100 467
rect 43 416 100 433
rect 150 572 206 616
rect 150 538 161 572
rect 195 538 206 572
rect 150 416 206 538
rect 256 597 312 616
rect 256 563 267 597
rect 301 563 312 597
rect 256 470 312 563
rect 256 436 267 470
rect 301 436 312 470
rect 256 416 312 436
rect 362 604 426 616
rect 362 570 373 604
rect 407 570 426 604
rect 362 533 426 570
rect 362 499 373 533
rect 407 499 426 533
rect 362 462 426 499
rect 362 428 373 462
rect 407 428 426 462
rect 362 416 426 428
rect 476 597 533 616
rect 476 563 487 597
rect 521 563 533 597
rect 476 462 533 563
rect 476 428 487 462
rect 521 428 533 462
rect 476 416 533 428
<< ndiffc >>
rect 81 153 115 187
rect 323 153 357 187
rect 503 174 537 208
<< pdiffc >>
rect 55 563 89 597
rect 55 433 89 467
rect 161 538 195 572
rect 267 563 301 597
rect 267 436 301 470
rect 373 570 407 604
rect 373 499 407 533
rect 373 428 407 462
rect 487 563 521 597
rect 487 428 521 462
<< poly >>
rect 100 616 150 642
rect 206 616 256 642
rect 312 616 362 642
rect 426 616 476 642
rect 100 381 150 416
rect 206 384 256 416
rect 90 365 156 381
rect 90 331 106 365
rect 140 331 156 365
rect 90 297 156 331
rect 198 368 264 384
rect 198 334 214 368
rect 248 334 264 368
rect 198 318 264 334
rect 312 376 362 416
rect 312 360 378 376
rect 312 326 328 360
rect 362 326 378 360
rect 90 263 106 297
rect 140 263 156 297
rect 90 247 156 263
rect 126 225 156 247
rect 204 225 234 318
rect 312 310 378 326
rect 426 329 476 416
rect 312 270 342 310
rect 426 299 492 329
rect 282 240 342 270
rect 282 225 312 240
rect 390 225 420 251
rect 462 225 492 299
rect 126 115 156 141
rect 204 115 234 141
rect 282 115 312 141
rect 390 119 420 141
rect 462 119 492 141
rect 390 103 492 119
rect 390 69 425 103
rect 459 69 492 103
rect 390 53 492 69
<< polycont >>
rect 106 331 140 365
rect 214 334 248 368
rect 328 326 362 360
rect 106 263 140 297
rect 425 69 459 103
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 20 597 105 613
rect 20 563 55 597
rect 89 563 105 597
rect 20 467 105 563
rect 145 572 211 649
rect 145 538 161 572
rect 195 538 211 572
rect 145 490 211 538
rect 251 597 317 613
rect 251 563 267 597
rect 301 563 317 597
rect 20 433 55 467
rect 89 454 105 467
rect 251 470 317 563
rect 251 454 267 470
rect 89 436 267 454
rect 301 436 317 470
rect 89 433 317 436
rect 20 420 317 433
rect 357 604 423 649
rect 357 570 373 604
rect 407 570 423 604
rect 357 533 423 570
rect 357 499 373 533
rect 407 499 423 533
rect 357 462 423 499
rect 357 428 373 462
rect 407 428 423 462
rect 20 417 105 420
rect 20 204 54 417
rect 357 412 423 428
rect 471 597 553 613
rect 471 563 487 597
rect 521 563 553 597
rect 471 462 553 563
rect 471 428 487 462
rect 521 428 553 462
rect 471 412 553 428
rect 90 365 156 381
rect 90 331 106 365
rect 140 331 156 365
rect 90 297 156 331
rect 198 368 264 384
rect 198 334 214 368
rect 248 334 264 368
rect 198 310 264 334
rect 312 360 455 376
rect 312 326 328 360
rect 362 326 455 360
rect 312 310 455 326
rect 90 263 106 297
rect 140 274 156 297
rect 519 274 553 412
rect 140 263 553 274
rect 90 240 553 263
rect 487 208 553 240
rect 20 187 263 204
rect 20 153 81 187
rect 115 153 263 187
rect 20 88 263 153
rect 307 187 373 204
rect 307 153 323 187
rect 357 153 373 187
rect 487 174 503 208
rect 537 174 553 208
rect 487 170 553 174
rect 307 17 373 153
rect 409 103 551 134
rect 409 69 425 103
rect 459 69 551 103
rect 409 53 551 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand3b_lp
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3636650
string GDS_START 3631014
<< end >>
