magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3986 1975
<< nwell >>
rect -38 331 2726 704
<< pwell >>
rect 2027 241 2348 267
rect 2027 229 2687 241
rect 775 223 1161 229
rect 1676 223 2687 229
rect 775 191 2687 223
rect 9 160 197 184
rect 376 160 2687 191
rect 9 49 2687 160
rect 0 0 2688 49
<< scnmos >>
rect 88 74 118 158
rect 278 50 308 134
rect 350 50 380 134
rect 482 81 512 165
rect 554 81 584 165
rect 649 81 679 165
rect 875 119 905 203
rect 961 119 991 203
rect 1055 119 1085 203
rect 1157 113 1187 197
rect 1290 69 1320 197
rect 1415 69 1445 197
rect 1569 113 1599 197
rect 1641 113 1671 197
rect 1788 119 1818 203
rect 1860 119 1890 203
rect 2110 73 2140 241
rect 2235 73 2265 241
rect 2476 47 2506 131
rect 2578 47 2608 215
<< scpmoshvt >>
rect 239 463 269 591
rect 325 463 355 591
rect 397 463 427 591
rect 483 463 513 591
rect 577 463 607 591
rect 674 463 704 591
rect 779 463 809 547
rect 865 463 895 547
rect 937 463 967 547
rect 1045 463 1075 547
rect 1338 379 1368 547
rect 1424 379 1454 547
rect 1548 533 1578 617
rect 1666 533 1696 617
rect 1833 533 1863 617
rect 1919 533 1949 617
rect 2118 367 2148 619
rect 2235 367 2265 619
rect 2461 367 2491 495
rect 2578 367 2608 619
<< ndiff >>
rect 35 133 88 158
rect 35 99 43 133
rect 77 99 88 133
rect 35 74 88 99
rect 118 122 171 158
rect 402 157 482 165
rect 402 134 414 157
rect 118 88 129 122
rect 163 88 171 122
rect 118 74 171 88
rect 225 103 278 134
rect 225 69 233 103
rect 267 69 278 103
rect 225 50 278 69
rect 308 50 350 134
rect 380 123 414 134
rect 448 123 482 157
rect 380 81 482 123
rect 512 81 554 165
rect 584 123 649 165
rect 584 89 595 123
rect 629 89 649 123
rect 584 81 649 89
rect 679 127 739 165
rect 679 93 697 127
rect 731 93 739 127
rect 679 81 739 93
rect 380 50 460 81
rect 801 181 875 203
rect 801 147 809 181
rect 843 147 875 181
rect 801 119 875 147
rect 905 195 961 203
rect 905 161 916 195
rect 950 161 961 195
rect 905 119 961 161
rect 991 119 1055 203
rect 1085 197 1135 203
rect 2053 233 2110 241
rect 1702 197 1788 203
rect 1085 119 1157 197
rect 1107 113 1157 119
rect 1187 120 1290 197
rect 1187 113 1245 120
rect 1237 86 1245 113
rect 1279 86 1290 120
rect 1237 69 1290 86
rect 1320 189 1415 197
rect 1320 155 1331 189
rect 1365 155 1415 189
rect 1320 111 1415 155
rect 1320 77 1370 111
rect 1404 77 1415 111
rect 1320 69 1415 77
rect 1445 183 1569 197
rect 1445 149 1456 183
rect 1490 149 1524 183
rect 1558 149 1569 183
rect 1445 115 1569 149
rect 1445 81 1456 115
rect 1490 113 1569 115
rect 1599 113 1641 197
rect 1671 177 1788 197
rect 1671 143 1714 177
rect 1748 143 1788 177
rect 1671 119 1788 143
rect 1818 119 1860 203
rect 1890 177 1943 203
rect 1890 143 1901 177
rect 1935 143 1943 177
rect 1890 119 1943 143
rect 2053 199 2065 233
rect 2099 199 2110 233
rect 1671 113 1752 119
rect 1490 81 1498 113
rect 1445 69 1498 81
rect 2053 73 2110 199
rect 2140 93 2235 241
rect 2140 73 2167 93
rect 2155 59 2167 73
rect 2201 73 2235 93
rect 2265 233 2322 241
rect 2265 199 2276 233
rect 2310 199 2322 233
rect 2265 73 2322 199
rect 2528 131 2578 215
rect 2423 105 2476 131
rect 2201 59 2213 73
rect 2155 51 2213 59
rect 2423 71 2431 105
rect 2465 71 2476 105
rect 2423 47 2476 71
rect 2506 91 2578 131
rect 2506 57 2533 91
rect 2567 57 2578 91
rect 2506 47 2578 57
rect 2608 203 2661 215
rect 2608 169 2619 203
rect 2653 169 2661 203
rect 2608 101 2661 169
rect 2608 67 2619 101
rect 2653 67 2661 101
rect 2608 47 2661 67
<< pdiff >>
rect 118 577 239 591
rect 118 475 126 577
rect 228 475 239 577
rect 118 463 239 475
rect 269 583 325 591
rect 269 549 280 583
rect 314 549 325 583
rect 269 509 325 549
rect 269 475 280 509
rect 314 475 325 509
rect 269 463 325 475
rect 355 463 397 591
rect 427 583 483 591
rect 427 549 438 583
rect 472 549 483 583
rect 427 509 483 549
rect 427 475 438 509
rect 472 475 483 509
rect 427 463 483 475
rect 513 463 577 591
rect 607 571 674 591
rect 607 537 624 571
rect 658 537 674 571
rect 607 463 674 537
rect 704 577 757 591
rect 704 543 715 577
rect 749 547 757 577
rect 1258 568 1316 576
rect 749 543 779 547
rect 704 509 779 543
rect 704 475 727 509
rect 761 475 779 509
rect 704 463 779 475
rect 809 522 865 547
rect 809 488 820 522
rect 854 488 865 522
rect 809 463 865 488
rect 895 463 937 547
rect 967 539 1045 547
rect 967 505 989 539
rect 1023 505 1045 539
rect 967 463 1045 505
rect 1075 522 1128 547
rect 1075 488 1086 522
rect 1120 488 1128 522
rect 1258 534 1270 568
rect 1304 547 1316 568
rect 1476 547 1548 617
rect 1304 534 1338 547
rect 1075 463 1128 488
rect 1258 379 1338 534
rect 1368 428 1424 547
rect 1368 394 1379 428
rect 1413 394 1424 428
rect 1368 379 1424 394
rect 1454 533 1548 547
rect 1578 533 1666 617
rect 1696 609 1833 617
rect 1696 575 1707 609
rect 1741 575 1788 609
rect 1822 575 1833 609
rect 1696 533 1833 575
rect 1863 599 1919 617
rect 1863 565 1874 599
rect 1908 565 1919 599
rect 1863 533 1919 565
rect 1949 592 2002 617
rect 1949 558 1960 592
rect 1994 558 2002 592
rect 1949 533 2002 558
rect 1454 531 1526 533
rect 1454 497 1465 531
rect 1499 497 1526 531
rect 1454 425 1526 497
rect 1454 391 1465 425
rect 1499 391 1526 425
rect 1454 379 1526 391
rect 2065 424 2118 619
rect 2065 390 2073 424
rect 2107 390 2118 424
rect 2065 367 2118 390
rect 2148 592 2235 619
rect 2148 558 2167 592
rect 2201 558 2235 592
rect 2148 367 2235 558
rect 2265 572 2318 619
rect 2265 538 2276 572
rect 2310 538 2318 572
rect 2265 367 2318 538
rect 2525 607 2578 619
rect 2525 573 2533 607
rect 2567 573 2578 607
rect 2525 518 2578 573
rect 2525 495 2533 518
rect 2408 483 2461 495
rect 2408 449 2416 483
rect 2450 449 2461 483
rect 2408 413 2461 449
rect 2408 379 2416 413
rect 2450 379 2461 413
rect 2408 367 2461 379
rect 2491 484 2533 495
rect 2567 484 2578 518
rect 2491 437 2578 484
rect 2491 403 2502 437
rect 2536 403 2578 437
rect 2491 367 2578 403
rect 2608 599 2661 619
rect 2608 565 2619 599
rect 2653 565 2661 599
rect 2608 506 2661 565
rect 2608 472 2619 506
rect 2653 472 2661 506
rect 2608 413 2661 472
rect 2608 379 2619 413
rect 2653 379 2661 413
rect 2608 367 2661 379
<< ndiffc >>
rect 43 99 77 133
rect 129 88 163 122
rect 233 69 267 103
rect 414 123 448 157
rect 595 89 629 123
rect 697 93 731 127
rect 809 147 843 181
rect 916 161 950 195
rect 1245 86 1279 120
rect 1331 155 1365 189
rect 1370 77 1404 111
rect 1456 149 1490 183
rect 1524 149 1558 183
rect 1456 81 1490 115
rect 1714 143 1748 177
rect 1901 143 1935 177
rect 2065 199 2099 233
rect 2167 59 2201 93
rect 2276 199 2310 233
rect 2431 71 2465 105
rect 2533 57 2567 91
rect 2619 169 2653 203
rect 2619 67 2653 101
<< pdiffc >>
rect 126 475 228 577
rect 280 549 314 583
rect 280 475 314 509
rect 438 549 472 583
rect 438 475 472 509
rect 624 537 658 571
rect 715 543 749 577
rect 727 475 761 509
rect 820 488 854 522
rect 989 505 1023 539
rect 1086 488 1120 522
rect 1270 534 1304 568
rect 1379 394 1413 428
rect 1707 575 1741 609
rect 1788 575 1822 609
rect 1874 565 1908 599
rect 1960 558 1994 592
rect 1465 497 1499 531
rect 1465 391 1499 425
rect 2073 390 2107 424
rect 2167 558 2201 592
rect 2276 538 2310 572
rect 2533 573 2567 607
rect 2416 449 2450 483
rect 2416 379 2450 413
rect 2533 484 2567 518
rect 2502 403 2536 437
rect 2619 565 2653 599
rect 2619 472 2653 506
rect 2619 379 2653 413
<< poly >>
rect 239 591 269 617
rect 325 591 355 617
rect 397 591 427 617
rect 483 591 513 617
rect 577 591 607 617
rect 674 591 704 617
rect 865 615 1454 645
rect 1548 617 1578 643
rect 1666 617 1696 643
rect 1833 617 1863 643
rect 1919 617 1949 643
rect 2118 619 2148 645
rect 2235 619 2265 645
rect 2578 619 2608 645
rect 779 547 809 573
rect 865 547 895 615
rect 937 547 967 573
rect 1045 547 1075 573
rect 1338 547 1368 573
rect 1424 547 1454 615
rect 1151 493 1226 509
rect 239 436 269 463
rect 325 436 355 463
rect 88 406 355 436
rect 88 276 183 406
rect 397 364 427 463
rect 483 429 513 463
rect 332 348 427 364
rect 469 413 535 429
rect 469 379 485 413
rect 519 379 535 413
rect 469 363 535 379
rect 577 369 607 463
rect 674 441 704 463
rect 674 411 715 441
rect 332 314 348 348
rect 382 334 427 348
rect 577 353 643 369
rect 382 314 398 334
rect 332 292 398 314
rect 577 319 593 353
rect 627 319 643 353
rect 88 242 133 276
rect 167 242 183 276
rect 88 226 183 242
rect 88 158 118 226
rect 236 206 302 222
rect 236 172 252 206
rect 286 186 302 206
rect 286 172 308 186
rect 236 156 308 172
rect 278 134 308 156
rect 350 134 380 292
rect 446 276 512 292
rect 446 242 462 276
rect 496 242 512 276
rect 577 285 643 319
rect 577 265 593 285
rect 446 226 512 242
rect 482 165 512 226
rect 554 251 593 265
rect 627 251 643 285
rect 554 235 643 251
rect 685 269 715 411
rect 779 383 809 463
rect 757 367 823 383
rect 757 333 773 367
rect 807 333 823 367
rect 757 317 823 333
rect 865 285 895 463
rect 937 399 967 463
rect 1045 441 1075 463
rect 1151 459 1176 493
rect 1210 459 1226 493
rect 1151 441 1226 459
rect 1045 425 1226 441
rect 1045 411 1176 425
rect 937 383 1003 399
rect 937 349 953 383
rect 987 369 1003 383
rect 1151 391 1176 411
rect 1210 391 1226 425
rect 1151 375 1226 391
rect 1548 477 1578 533
rect 1666 477 1696 533
rect 1833 501 1863 533
rect 1788 485 1863 501
rect 1548 461 1624 477
rect 1548 427 1574 461
rect 1608 427 1624 461
rect 1548 411 1624 427
rect 1666 461 1746 477
rect 1666 427 1696 461
rect 1730 427 1746 461
rect 1666 411 1746 427
rect 987 349 1091 369
rect 937 339 1091 349
rect 937 333 1003 339
rect 685 239 784 269
rect 865 255 905 285
rect 554 165 584 235
rect 649 165 679 191
rect 88 48 118 74
rect 482 55 512 81
rect 554 55 584 81
rect 649 51 679 81
rect 754 51 784 239
rect 875 203 905 255
rect 947 275 1013 291
rect 1061 285 1091 339
rect 947 241 963 275
rect 997 241 1013 275
rect 947 225 1013 241
rect 1055 255 1091 285
rect 961 203 991 225
rect 1055 203 1085 255
rect 1151 249 1181 375
rect 1338 327 1368 379
rect 1424 357 1454 379
rect 1563 357 1674 363
rect 1424 347 1674 357
rect 1424 327 1624 347
rect 1229 297 1368 327
rect 1569 313 1624 327
rect 1658 313 1674 347
rect 1569 297 1674 313
rect 1229 284 1320 297
rect 1229 250 1245 284
rect 1279 250 1320 284
rect 1151 219 1187 249
rect 1229 234 1320 250
rect 1455 269 1521 285
rect 1455 249 1471 269
rect 1157 197 1187 219
rect 1290 197 1320 234
rect 1415 235 1471 249
rect 1505 235 1521 269
rect 1415 219 1521 235
rect 1415 197 1445 219
rect 1569 197 1599 297
rect 1716 249 1746 411
rect 1641 219 1746 249
rect 1788 451 1804 485
rect 1838 451 1863 485
rect 1788 435 1863 451
rect 1641 197 1671 219
rect 1788 203 1818 435
rect 1919 291 1949 533
rect 2461 495 2491 521
rect 2118 335 2148 367
rect 2110 319 2193 335
rect 1896 275 1962 291
rect 1896 255 1912 275
rect 1860 241 1912 255
rect 1946 241 1962 275
rect 2110 285 2143 319
rect 2177 285 2193 319
rect 2110 269 2193 285
rect 2235 299 2265 367
rect 2310 319 2376 335
rect 2310 299 2326 319
rect 2235 285 2326 299
rect 2360 285 2376 319
rect 2461 317 2491 367
rect 2578 327 2608 367
rect 2235 269 2376 285
rect 2425 301 2491 317
rect 2110 241 2140 269
rect 2235 241 2265 269
rect 2425 267 2441 301
rect 2475 267 2491 301
rect 1860 225 1962 241
rect 1860 203 1890 225
rect 875 93 905 119
rect 961 93 991 119
rect 1055 93 1085 119
rect 1157 51 1187 113
rect 1569 87 1599 113
rect 278 24 308 50
rect 350 24 380 50
rect 649 21 1187 51
rect 1290 43 1320 69
rect 1415 43 1445 69
rect 1641 51 1671 113
rect 1788 93 1818 119
rect 1860 93 1890 119
rect 1965 87 2031 103
rect 1965 53 1981 87
rect 2015 53 2031 87
rect 1965 51 2031 53
rect 1641 21 2031 51
rect 2110 47 2140 73
rect 2425 233 2491 267
rect 2533 311 2608 327
rect 2533 277 2549 311
rect 2583 277 2608 311
rect 2533 261 2608 277
rect 2425 199 2441 233
rect 2475 213 2491 233
rect 2578 215 2608 261
rect 2475 199 2506 213
rect 2425 183 2506 199
rect 2476 131 2506 183
rect 2235 47 2265 73
rect 2476 21 2506 47
rect 2578 21 2608 47
<< polycont >>
rect 485 379 519 413
rect 348 314 382 348
rect 593 319 627 353
rect 133 242 167 276
rect 252 172 286 206
rect 462 242 496 276
rect 593 251 627 285
rect 773 333 807 367
rect 1176 459 1210 493
rect 953 349 987 383
rect 1176 391 1210 425
rect 1574 427 1608 461
rect 1696 427 1730 461
rect 963 241 997 275
rect 1624 313 1658 347
rect 1245 250 1279 284
rect 1471 235 1505 269
rect 1804 451 1838 485
rect 1912 241 1946 275
rect 2143 285 2177 319
rect 2326 285 2360 319
rect 2441 267 2475 301
rect 1981 53 2015 87
rect 2549 277 2583 311
rect 2441 199 2475 233
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 18 577 230 593
rect 18 475 126 577
rect 228 475 230 577
rect 18 429 230 475
rect 264 583 330 649
rect 264 549 280 583
rect 314 549 330 583
rect 264 509 330 549
rect 264 475 280 509
rect 314 475 330 509
rect 264 463 330 475
rect 422 583 488 599
rect 422 549 438 583
rect 472 549 488 583
rect 422 509 488 549
rect 608 571 674 649
rect 608 537 624 571
rect 658 537 674 571
rect 608 531 674 537
rect 708 577 765 593
rect 708 543 715 577
rect 749 543 765 577
rect 422 475 438 509
rect 472 497 488 509
rect 708 509 765 543
rect 973 539 1039 649
rect 708 497 727 509
rect 472 475 727 497
rect 761 475 765 509
rect 422 463 765 475
rect 696 459 765 463
rect 804 522 877 538
rect 804 488 820 522
rect 854 488 877 522
rect 973 505 989 539
rect 1023 505 1039 539
rect 1254 568 1320 649
rect 973 501 1039 505
rect 1073 522 1126 538
rect 1254 534 1270 568
rect 1304 534 1320 568
rect 1254 532 1320 534
rect 1354 581 1657 615
rect 804 467 877 488
rect 1073 488 1086 522
rect 1120 488 1126 522
rect 1073 467 1126 488
rect 18 413 535 429
rect 18 395 485 413
rect 18 206 74 395
rect 519 379 535 413
rect 485 363 535 379
rect 127 348 451 361
rect 127 314 348 348
rect 382 314 451 348
rect 127 313 451 314
rect 593 353 662 429
rect 627 319 662 353
rect 593 285 662 319
rect 108 276 559 279
rect 108 242 133 276
rect 167 242 462 276
rect 496 242 559 276
rect 108 240 559 242
rect 627 251 662 285
rect 593 235 662 251
rect 18 172 252 206
rect 286 172 302 206
rect 696 197 737 459
rect 804 433 1126 467
rect 1160 498 1226 509
rect 1354 498 1390 581
rect 1160 493 1390 498
rect 1160 459 1176 493
rect 1210 464 1390 493
rect 1463 531 1515 547
rect 1463 497 1465 531
rect 1499 497 1515 531
rect 1210 459 1226 464
rect 804 417 911 433
rect 771 367 843 383
rect 771 333 773 367
rect 807 333 843 367
rect 771 276 843 333
rect 771 242 799 276
rect 833 242 843 276
rect 771 231 843 242
rect 877 199 911 417
rect 1160 425 1226 459
rect 945 383 1003 399
rect 1160 391 1176 425
rect 1210 391 1226 425
rect 1160 388 1226 391
rect 1331 428 1429 430
rect 1331 394 1379 428
rect 1413 394 1429 428
rect 1331 392 1429 394
rect 1463 425 1515 497
rect 1607 529 1657 581
rect 1691 609 1838 649
rect 1691 575 1707 609
rect 1741 575 1788 609
rect 1822 575 1838 609
rect 1691 571 1838 575
rect 1872 599 1924 615
rect 1872 565 1874 599
rect 1908 565 1924 599
rect 1872 549 1924 565
rect 1607 514 1843 529
rect 1607 495 1854 514
rect 1788 485 1854 495
rect 945 349 953 383
rect 987 354 1003 383
rect 1331 354 1367 392
rect 1463 391 1465 425
rect 1499 391 1515 425
rect 1463 358 1515 391
rect 987 349 1367 354
rect 945 320 1367 349
rect 947 276 1025 286
rect 947 275 991 276
rect 947 241 963 275
rect 997 241 1025 242
rect 947 233 1025 241
rect 1229 284 1295 286
rect 1229 250 1245 284
rect 1279 250 1295 284
rect 1229 199 1295 250
rect 398 181 843 197
rect 18 133 86 172
rect 398 163 809 181
rect 398 157 464 163
rect 18 99 43 133
rect 77 99 86 133
rect 18 83 86 99
rect 120 122 179 138
rect 398 123 414 157
rect 448 123 464 157
rect 803 147 809 163
rect 877 195 1295 199
rect 877 161 916 195
rect 950 161 1295 195
rect 877 157 1295 161
rect 1329 189 1367 320
rect 803 131 843 147
rect 1329 155 1331 189
rect 1365 155 1367 189
rect 579 123 645 127
rect 120 88 129 122
rect 163 88 179 122
rect 120 17 179 88
rect 229 103 271 119
rect 229 69 233 103
rect 267 87 271 103
rect 579 89 595 123
rect 629 89 645 123
rect 579 87 645 89
rect 267 69 645 87
rect 229 53 645 69
rect 681 93 697 127
rect 731 93 747 127
rect 681 17 747 93
rect 1229 120 1295 123
rect 1229 86 1245 120
rect 1279 86 1295 120
rect 1229 17 1295 86
rect 1329 115 1367 155
rect 1401 324 1515 358
rect 1554 427 1574 461
rect 1608 427 1624 461
rect 1554 411 1624 427
rect 1680 427 1696 461
rect 1730 427 1746 461
rect 1788 451 1804 485
rect 1838 451 1854 485
rect 1680 415 1746 427
rect 1890 415 1924 549
rect 1958 592 2010 649
rect 1958 558 1960 592
rect 1994 558 2010 592
rect 1958 542 2010 558
rect 2143 592 2208 649
rect 2143 558 2167 592
rect 2201 558 2208 592
rect 2486 607 2583 649
rect 2143 542 2208 558
rect 2242 572 2326 588
rect 2242 538 2276 572
rect 2310 538 2326 572
rect 2242 534 2326 538
rect 2486 573 2533 607
rect 2567 573 2583 607
rect 2242 508 2276 534
rect 1680 411 1924 415
rect 1401 183 1435 324
rect 1554 285 1588 411
rect 1712 381 1924 411
rect 1960 474 2276 508
rect 2486 518 2583 573
rect 1622 347 1674 363
rect 1622 313 1624 347
rect 1658 345 1674 347
rect 1960 345 2009 474
rect 1658 313 2009 345
rect 1622 311 2009 313
rect 2043 424 2109 440
rect 2043 390 2073 424
rect 2107 390 2109 424
rect 1622 297 1674 311
rect 1469 276 1588 285
rect 1469 235 1471 276
rect 1505 235 1588 276
rect 1896 275 2009 277
rect 1896 261 1912 275
rect 1469 219 1588 235
rect 1622 241 1912 261
rect 1946 241 2009 275
rect 1622 227 2009 241
rect 1622 183 1664 227
rect 1401 149 1456 183
rect 1490 149 1524 183
rect 1558 149 1664 183
rect 1698 177 1764 193
rect 1454 115 1506 149
rect 1329 111 1420 115
rect 1329 77 1370 111
rect 1404 77 1420 111
rect 1329 71 1420 77
rect 1454 81 1456 115
rect 1490 81 1506 115
rect 1454 65 1506 81
rect 1698 143 1714 177
rect 1748 143 1764 177
rect 1698 17 1764 143
rect 1885 177 1941 193
rect 1885 143 1901 177
rect 1935 143 1941 177
rect 1885 95 1941 143
rect 1975 163 2009 227
rect 2043 276 2109 390
rect 2043 242 2047 276
rect 2081 242 2109 276
rect 2143 319 2276 474
rect 2177 285 2276 319
rect 2310 319 2376 500
rect 2410 483 2452 499
rect 2410 449 2416 483
rect 2450 449 2452 483
rect 2410 413 2452 449
rect 2410 379 2416 413
rect 2450 379 2452 413
rect 2486 484 2533 518
rect 2567 484 2583 518
rect 2486 437 2583 484
rect 2486 403 2502 437
rect 2536 403 2583 437
rect 2617 599 2671 615
rect 2617 565 2619 599
rect 2653 565 2671 599
rect 2617 506 2671 565
rect 2617 472 2619 506
rect 2653 472 2671 506
rect 2617 413 2671 472
rect 2410 369 2452 379
rect 2617 379 2619 413
rect 2653 379 2671 413
rect 2410 335 2583 369
rect 2310 285 2326 319
rect 2360 285 2376 319
rect 2533 311 2583 335
rect 2143 269 2276 285
rect 2043 233 2109 242
rect 2240 237 2276 269
rect 2425 267 2441 301
rect 2475 267 2491 301
rect 2240 233 2326 237
rect 2425 233 2491 267
rect 2043 199 2065 233
rect 2099 199 2115 233
rect 2043 197 2115 199
rect 2240 199 2276 233
rect 2310 199 2326 233
rect 2240 197 2326 199
rect 2362 199 2441 233
rect 2475 199 2491 233
rect 2362 197 2491 199
rect 2533 277 2549 311
rect 2362 163 2396 197
rect 2533 163 2583 277
rect 1975 129 2396 163
rect 2430 129 2583 163
rect 2617 203 2671 379
rect 2617 169 2619 203
rect 2653 169 2671 203
rect 2430 105 2481 129
rect 1885 87 2031 95
rect 1885 53 1981 87
rect 2015 53 2031 87
rect 1885 51 2031 53
rect 2151 93 2217 95
rect 2151 59 2167 93
rect 2201 59 2217 93
rect 2151 17 2217 59
rect 2430 71 2431 105
rect 2465 71 2481 105
rect 2617 101 2671 169
rect 2430 55 2481 71
rect 2515 91 2583 95
rect 2515 57 2533 91
rect 2567 57 2583 91
rect 2515 17 2583 57
rect 2617 67 2619 101
rect 2653 67 2671 101
rect 2617 51 2671 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 799 242 833 276
rect 991 275 1025 276
rect 991 242 997 275
rect 997 242 1025 275
rect 1471 269 1505 276
rect 1471 242 1505 269
rect 2047 242 2081 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 787 276 845 282
rect 787 242 799 276
rect 833 273 845 276
rect 979 276 1037 282
rect 979 273 991 276
rect 833 245 991 273
rect 833 242 845 245
rect 787 236 845 242
rect 979 242 991 245
rect 1025 273 1037 276
rect 1459 276 1517 282
rect 1459 273 1471 276
rect 1025 245 1471 273
rect 1025 242 1037 245
rect 979 236 1037 242
rect 1459 242 1471 245
rect 1505 273 1517 276
rect 2035 276 2093 282
rect 2035 273 2047 276
rect 1505 245 2047 273
rect 1505 242 1517 245
rect 1459 236 1517 242
rect 2035 242 2047 245
rect 2081 242 2093 276
rect 2035 236 2093 242
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
flabel pwell s 0 0 2688 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2688 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfrtp_1
flabel comment s 1729 347 1729 347 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 2688 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2688 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 1183 390 1217 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1183 464 1217 498 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 2335 316 2369 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2335 390 2369 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2335 464 2369 498 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2623 168 2657 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 242 2657 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 316 2657 350 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 390 2657 424 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 464 2657 498 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2623 538 2657 572 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2688 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3145054
string GDS_START 3124212
<< end >>
