magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3986 1975
<< nwell >>
rect -38 331 2726 704
rect 2065 303 2335 331
<< pwell >>
rect 684 219 1975 235
rect 263 167 1975 219
rect 1 157 1975 167
rect 2261 157 2687 184
rect 1 49 2687 157
rect 0 0 2688 49
<< scnmos >>
rect 80 57 110 141
rect 152 57 182 141
rect 343 109 373 193
rect 415 109 445 193
rect 501 109 531 193
rect 573 109 603 193
rect 763 125 793 209
rect 874 125 904 209
rect 946 125 976 209
rect 1226 125 1256 209
rect 1304 125 1334 209
rect 1418 125 1448 209
rect 1496 125 1526 209
rect 1653 125 1683 209
rect 1731 125 1761 209
rect 1862 125 1892 209
rect 2074 47 2104 131
rect 2146 47 2176 131
rect 2344 74 2374 158
rect 2416 74 2446 158
rect 2502 74 2532 158
rect 2574 74 2604 158
<< scpmoshvt >>
rect 85 409 135 609
rect 323 409 373 609
rect 429 409 479 609
rect 659 419 709 619
rect 831 419 881 619
rect 943 419 993 619
rect 1120 419 1170 619
rect 1229 419 1279 619
rect 1398 419 1448 619
rect 1496 419 1546 619
rect 1676 419 1726 619
rect 1784 419 1834 619
rect 1940 419 1990 619
rect 2158 339 2208 539
rect 2410 374 2460 574
rect 2516 374 2566 574
<< ndiff >>
rect 289 177 343 193
rect 289 143 298 177
rect 332 143 343 177
rect 27 116 80 141
rect 27 82 35 116
rect 69 82 80 116
rect 27 57 80 82
rect 110 57 152 141
rect 182 116 235 141
rect 182 82 193 116
rect 227 82 235 116
rect 289 109 343 143
rect 373 109 415 193
rect 445 161 501 193
rect 445 127 456 161
rect 490 127 501 161
rect 445 109 501 127
rect 531 109 573 193
rect 603 177 656 193
rect 603 143 614 177
rect 648 143 656 177
rect 603 109 656 143
rect 710 184 763 209
rect 710 150 718 184
rect 752 150 763 184
rect 710 125 763 150
rect 793 184 874 209
rect 793 150 817 184
rect 851 150 874 184
rect 793 125 874 150
rect 904 125 946 209
rect 976 125 1045 209
rect 1169 180 1226 209
rect 1169 146 1181 180
rect 1215 146 1226 180
rect 1169 125 1226 146
rect 1256 125 1304 209
rect 1334 179 1418 209
rect 1334 145 1353 179
rect 1387 145 1418 179
rect 1334 125 1418 145
rect 1448 125 1496 209
rect 1526 184 1653 209
rect 1526 150 1608 184
rect 1642 150 1653 184
rect 1526 125 1653 150
rect 1683 125 1731 209
rect 1761 125 1862 209
rect 1892 175 1949 209
rect 1892 141 1903 175
rect 1937 141 1949 175
rect 1892 125 1949 141
rect 2287 133 2344 158
rect 182 57 235 82
rect 991 123 1045 125
rect 991 89 999 123
rect 1033 89 1045 123
rect 991 77 1045 89
rect 2017 111 2074 131
rect 2017 77 2029 111
rect 2063 77 2074 111
rect 2017 47 2074 77
rect 2104 47 2146 131
rect 2176 103 2233 131
rect 2176 69 2187 103
rect 2221 69 2233 103
rect 2287 99 2299 133
rect 2333 99 2344 133
rect 2287 74 2344 99
rect 2374 74 2416 158
rect 2446 133 2502 158
rect 2446 99 2457 133
rect 2491 99 2502 133
rect 2446 74 2502 99
rect 2532 74 2574 158
rect 2604 133 2661 158
rect 2604 99 2615 133
rect 2649 99 2661 133
rect 2604 74 2661 99
rect 2176 47 2233 69
<< pdiff >>
rect 28 597 85 609
rect 28 563 40 597
rect 74 563 85 597
rect 28 526 85 563
rect 28 492 40 526
rect 74 492 85 526
rect 28 455 85 492
rect 28 421 40 455
rect 74 421 85 455
rect 28 409 85 421
rect 135 597 192 609
rect 135 563 146 597
rect 180 563 192 597
rect 135 526 192 563
rect 135 492 146 526
rect 180 492 192 526
rect 135 455 192 492
rect 135 421 146 455
rect 180 421 192 455
rect 135 409 192 421
rect 266 597 323 609
rect 266 563 278 597
rect 312 563 323 597
rect 266 526 323 563
rect 266 492 278 526
rect 312 492 323 526
rect 266 455 323 492
rect 266 421 278 455
rect 312 421 323 455
rect 266 409 323 421
rect 373 597 429 609
rect 373 563 384 597
rect 418 563 429 597
rect 373 512 429 563
rect 373 478 384 512
rect 418 478 429 512
rect 373 409 429 478
rect 479 597 536 609
rect 479 563 490 597
rect 524 563 536 597
rect 479 526 536 563
rect 479 492 490 526
rect 524 492 536 526
rect 479 455 536 492
rect 479 421 490 455
rect 524 421 536 455
rect 479 409 536 421
rect 602 496 659 619
rect 602 462 614 496
rect 648 462 659 496
rect 602 419 659 462
rect 709 496 831 619
rect 709 462 786 496
rect 820 462 831 496
rect 709 419 831 462
rect 881 419 943 619
rect 993 607 1120 619
rect 993 573 1004 607
rect 1038 573 1120 607
rect 993 419 1120 573
rect 1170 497 1229 619
rect 1170 463 1181 497
rect 1215 463 1229 497
rect 1170 419 1229 463
rect 1279 607 1398 619
rect 1279 573 1353 607
rect 1387 573 1398 607
rect 1279 532 1398 573
rect 1279 498 1353 532
rect 1387 498 1398 532
rect 1279 419 1398 498
rect 1448 419 1496 619
rect 1546 597 1676 619
rect 1546 563 1625 597
rect 1659 563 1676 597
rect 1546 465 1676 563
rect 1546 431 1625 465
rect 1659 431 1676 465
rect 1546 419 1676 431
rect 1726 419 1784 619
rect 1834 607 1940 619
rect 1834 573 1845 607
rect 1879 573 1940 607
rect 1834 524 1940 573
rect 1834 490 1845 524
rect 1879 490 1940 524
rect 1834 419 1940 490
rect 1990 597 2047 619
rect 1990 563 2001 597
rect 2035 563 2047 597
rect 1990 465 2047 563
rect 2353 562 2410 574
rect 1990 431 2001 465
rect 2035 431 2047 465
rect 1990 419 2047 431
rect 2101 527 2158 539
rect 2101 493 2113 527
rect 2147 493 2158 527
rect 2101 456 2158 493
rect 2101 422 2113 456
rect 2147 422 2158 456
rect 2101 385 2158 422
rect 2101 351 2113 385
rect 2147 351 2158 385
rect 2101 339 2158 351
rect 2208 527 2299 539
rect 2208 493 2253 527
rect 2287 493 2299 527
rect 2208 456 2299 493
rect 2208 422 2253 456
rect 2287 422 2299 456
rect 2208 385 2299 422
rect 2208 351 2253 385
rect 2287 351 2299 385
rect 2353 528 2365 562
rect 2399 528 2410 562
rect 2353 491 2410 528
rect 2353 457 2365 491
rect 2399 457 2410 491
rect 2353 420 2410 457
rect 2353 386 2365 420
rect 2399 386 2410 420
rect 2353 374 2410 386
rect 2460 562 2516 574
rect 2460 528 2471 562
rect 2505 528 2516 562
rect 2460 491 2516 528
rect 2460 457 2471 491
rect 2505 457 2516 491
rect 2460 420 2516 457
rect 2460 386 2471 420
rect 2505 386 2516 420
rect 2460 374 2516 386
rect 2566 562 2623 574
rect 2566 528 2577 562
rect 2611 528 2623 562
rect 2566 491 2623 528
rect 2566 457 2577 491
rect 2611 457 2623 491
rect 2566 420 2623 457
rect 2566 386 2577 420
rect 2611 386 2623 420
rect 2566 374 2623 386
rect 2208 339 2299 351
<< ndiffc >>
rect 298 143 332 177
rect 35 82 69 116
rect 193 82 227 116
rect 456 127 490 161
rect 614 143 648 177
rect 718 150 752 184
rect 817 150 851 184
rect 1181 146 1215 180
rect 1353 145 1387 179
rect 1608 150 1642 184
rect 1903 141 1937 175
rect 999 89 1033 123
rect 2029 77 2063 111
rect 2187 69 2221 103
rect 2299 99 2333 133
rect 2457 99 2491 133
rect 2615 99 2649 133
<< pdiffc >>
rect 40 563 74 597
rect 40 492 74 526
rect 40 421 74 455
rect 146 563 180 597
rect 146 492 180 526
rect 146 421 180 455
rect 278 563 312 597
rect 278 492 312 526
rect 278 421 312 455
rect 384 563 418 597
rect 384 478 418 512
rect 490 563 524 597
rect 490 492 524 526
rect 490 421 524 455
rect 614 462 648 496
rect 786 462 820 496
rect 1004 573 1038 607
rect 1181 463 1215 497
rect 1353 573 1387 607
rect 1353 498 1387 532
rect 1625 563 1659 597
rect 1625 431 1659 465
rect 1845 573 1879 607
rect 1845 490 1879 524
rect 2001 563 2035 597
rect 2001 431 2035 465
rect 2113 493 2147 527
rect 2113 422 2147 456
rect 2113 351 2147 385
rect 2253 493 2287 527
rect 2253 422 2287 456
rect 2253 351 2287 385
rect 2365 528 2399 562
rect 2365 457 2399 491
rect 2365 386 2399 420
rect 2471 528 2505 562
rect 2471 457 2505 491
rect 2471 386 2505 420
rect 2577 528 2611 562
rect 2577 457 2611 491
rect 2577 386 2611 420
<< poly >>
rect 85 609 135 635
rect 323 609 373 635
rect 429 609 479 635
rect 659 619 709 645
rect 831 619 881 645
rect 943 619 993 645
rect 1120 619 1170 645
rect 1229 619 1279 645
rect 1398 619 1448 645
rect 1496 619 1546 645
rect 1676 619 1726 645
rect 1784 619 1834 645
rect 1940 619 1990 645
rect 2410 574 2460 600
rect 2516 574 2566 600
rect 2158 539 2208 565
rect 85 356 135 409
rect 323 356 373 409
rect 44 340 135 356
rect 44 306 60 340
rect 94 306 135 340
rect 44 272 135 306
rect 302 340 373 356
rect 302 306 318 340
rect 352 306 373 340
rect 302 290 373 306
rect 429 369 479 409
rect 429 353 531 369
rect 659 368 709 419
rect 831 393 881 419
rect 429 319 445 353
rect 479 319 531 353
rect 429 303 531 319
rect 44 238 60 272
rect 94 238 135 272
rect 44 222 135 238
rect 80 186 135 222
rect 343 238 373 290
rect 501 254 531 303
rect 643 352 709 368
rect 643 318 659 352
rect 693 318 709 352
rect 643 302 709 318
rect 757 363 881 393
rect 943 387 993 419
rect 943 371 1073 387
rect 1120 381 1170 419
rect 757 254 787 363
rect 943 337 1023 371
rect 1057 337 1073 371
rect 943 321 1073 337
rect 1115 365 1181 381
rect 1115 331 1131 365
rect 1165 331 1181 365
rect 835 299 901 315
rect 835 265 851 299
rect 885 273 901 299
rect 885 265 904 273
rect 343 208 445 238
rect 343 193 373 208
rect 415 193 445 208
rect 501 224 793 254
rect 835 243 904 265
rect 501 193 531 224
rect 573 193 603 224
rect 763 209 793 224
rect 874 209 904 243
rect 946 209 976 321
rect 1115 315 1181 331
rect 1151 254 1181 315
rect 1229 376 1279 419
rect 1229 360 1340 376
rect 1398 374 1448 419
rect 1496 404 1546 419
rect 1496 374 1628 404
rect 1229 326 1290 360
rect 1324 326 1340 360
rect 1229 310 1340 326
rect 1382 358 1448 374
rect 1382 324 1398 358
rect 1432 324 1448 358
rect 1151 224 1256 254
rect 1226 209 1256 224
rect 1304 209 1334 310
rect 1382 290 1448 324
rect 1382 256 1398 290
rect 1432 256 1448 290
rect 1490 310 1556 326
rect 1490 276 1506 310
rect 1540 276 1556 310
rect 1490 260 1556 276
rect 1382 240 1448 256
rect 1418 209 1448 240
rect 1496 209 1526 260
rect 1598 254 1628 374
rect 1676 368 1726 419
rect 1784 368 1834 419
rect 1940 368 1990 419
rect 1670 352 1736 368
rect 1670 318 1686 352
rect 1720 318 1736 352
rect 1670 302 1736 318
rect 1784 352 1898 368
rect 1784 318 1848 352
rect 1882 318 1898 352
rect 1784 302 1898 318
rect 1940 352 2006 368
rect 1940 318 1956 352
rect 1990 318 2006 352
rect 1940 302 2006 318
rect 1784 254 1814 302
rect 1976 254 2006 302
rect 2158 299 2208 339
rect 2410 299 2460 374
rect 2516 332 2566 374
rect 1598 224 1683 254
rect 1653 209 1683 224
rect 1731 224 1814 254
rect 1862 224 2006 254
rect 2146 283 2460 299
rect 2146 249 2183 283
rect 2217 269 2460 283
rect 2502 316 2568 332
rect 2502 282 2518 316
rect 2552 282 2568 316
rect 2217 249 2233 269
rect 1731 209 1761 224
rect 1862 209 1892 224
rect 2146 215 2233 249
rect 80 156 182 186
rect 80 141 110 156
rect 152 141 182 156
rect 2146 181 2183 215
rect 2217 181 2233 215
rect 2146 176 2233 181
rect 2074 165 2233 176
rect 2074 146 2176 165
rect 2344 158 2374 269
rect 2416 158 2446 269
rect 2502 248 2568 282
rect 2502 214 2518 248
rect 2552 228 2568 248
rect 2552 214 2604 228
rect 2502 198 2604 214
rect 2502 158 2532 198
rect 2574 158 2604 198
rect 2074 131 2104 146
rect 2146 131 2176 146
rect 343 83 373 109
rect 415 83 445 109
rect 501 83 531 109
rect 573 83 603 109
rect 80 31 110 57
rect 152 31 182 57
rect 763 51 793 125
rect 874 99 904 125
rect 946 99 976 125
rect 1226 99 1256 125
rect 1304 99 1334 125
rect 1418 99 1448 125
rect 1496 99 1526 125
rect 1653 51 1683 125
rect 1731 99 1761 125
rect 1862 99 1892 125
rect 763 21 1683 51
rect 2344 48 2374 74
rect 2416 48 2446 74
rect 2502 48 2532 74
rect 2574 48 2604 74
rect 2074 21 2104 47
rect 2146 21 2176 47
<< polycont >>
rect 60 306 94 340
rect 318 306 352 340
rect 445 319 479 353
rect 60 238 94 272
rect 659 318 693 352
rect 1023 337 1057 371
rect 1131 331 1165 365
rect 851 265 885 299
rect 1290 326 1324 360
rect 1398 324 1432 358
rect 1398 256 1432 290
rect 1506 276 1540 310
rect 1686 318 1720 352
rect 1848 318 1882 352
rect 1956 318 1990 352
rect 2183 249 2217 283
rect 2518 282 2552 316
rect 2183 181 2217 215
rect 2518 214 2552 248
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 24 597 90 649
rect 24 563 40 597
rect 74 563 90 597
rect 24 526 90 563
rect 24 492 40 526
rect 74 492 90 526
rect 24 455 90 492
rect 24 421 40 455
rect 74 421 90 455
rect 24 405 90 421
rect 130 597 196 613
rect 130 563 146 597
rect 180 563 196 597
rect 130 526 196 563
rect 130 492 146 526
rect 180 492 196 526
rect 130 455 196 492
rect 130 421 146 455
rect 180 421 196 455
rect 130 405 196 421
rect 25 340 110 356
rect 25 306 60 340
rect 94 306 110 340
rect 25 272 110 306
rect 25 238 60 272
rect 94 238 110 272
rect 25 222 110 238
rect 162 145 196 405
rect 232 597 328 613
rect 232 563 278 597
rect 312 563 328 597
rect 232 526 328 563
rect 232 492 278 526
rect 312 492 328 526
rect 232 455 328 492
rect 368 597 434 649
rect 368 563 384 597
rect 418 563 434 597
rect 368 512 434 563
rect 368 478 384 512
rect 418 478 434 512
rect 368 462 434 478
rect 474 597 952 613
rect 474 563 490 597
rect 524 579 952 597
rect 474 526 524 563
rect 474 492 490 526
rect 232 421 278 455
rect 312 426 328 455
rect 474 455 524 492
rect 312 421 438 426
rect 232 392 438 421
rect 474 421 490 455
rect 474 405 524 421
rect 560 496 664 543
rect 560 462 614 496
rect 648 462 664 496
rect 560 415 664 462
rect 232 254 266 392
rect 404 369 438 392
rect 302 340 368 356
rect 302 306 318 340
rect 352 306 368 340
rect 302 290 368 306
rect 404 353 495 369
rect 404 319 445 353
rect 479 319 495 353
rect 404 303 495 319
rect 560 267 594 415
rect 700 368 734 579
rect 770 496 836 543
rect 770 462 786 496
rect 820 462 836 496
rect 918 521 952 579
rect 988 607 1054 649
rect 988 573 1004 607
rect 1038 573 1054 607
rect 988 557 1054 573
rect 1090 579 1301 613
rect 1090 521 1124 579
rect 918 487 1124 521
rect 1165 497 1231 543
rect 770 449 836 462
rect 1165 463 1181 497
rect 1215 463 1231 497
rect 1165 451 1231 463
rect 770 415 971 449
rect 420 254 594 267
rect 232 220 348 254
rect 282 177 348 220
rect 19 116 85 145
rect 19 82 35 116
rect 69 82 85 116
rect 19 17 85 82
rect 162 116 243 145
rect 282 143 298 177
rect 332 143 348 177
rect 282 123 348 143
rect 386 233 594 254
rect 630 352 734 368
rect 630 318 659 352
rect 693 318 734 352
rect 630 315 734 318
rect 630 299 901 315
rect 630 265 851 299
rect 885 265 901 299
rect 630 249 901 265
rect 386 220 560 233
rect 162 82 193 116
rect 227 87 243 116
rect 386 87 420 220
rect 227 82 420 87
rect 162 53 420 82
rect 456 161 490 184
rect 456 17 490 127
rect 526 87 560 220
rect 630 197 664 249
rect 937 213 971 415
rect 1007 417 1231 451
rect 1267 446 1301 579
rect 1337 607 1403 649
rect 1337 573 1353 607
rect 1387 573 1403 607
rect 1337 532 1403 573
rect 1337 498 1353 532
rect 1387 498 1403 532
rect 1337 482 1403 498
rect 1609 597 1675 613
rect 1609 563 1625 597
rect 1659 563 1675 597
rect 1609 465 1675 563
rect 1829 607 1895 649
rect 1829 573 1845 607
rect 1879 573 1895 607
rect 1829 524 1895 573
rect 1829 490 1845 524
rect 1879 490 1895 524
rect 1829 474 1895 490
rect 1985 597 2217 613
rect 1985 563 2001 597
rect 2035 579 2217 597
rect 2035 563 2051 579
rect 1007 371 1073 417
rect 1267 412 1556 446
rect 1007 337 1023 371
rect 1057 337 1073 371
rect 1007 279 1073 337
rect 1115 365 1181 381
rect 1115 331 1131 365
rect 1165 349 1181 365
rect 1279 360 1340 376
rect 1279 350 1290 360
rect 1165 331 1243 349
rect 1115 315 1243 331
rect 1007 245 1173 279
rect 598 177 664 197
rect 598 143 614 177
rect 648 143 664 177
rect 598 123 664 143
rect 702 184 768 213
rect 702 150 718 184
rect 752 150 768 184
rect 702 87 768 150
rect 817 209 971 213
rect 817 184 1103 209
rect 851 175 1103 184
rect 851 150 867 175
rect 817 121 867 150
rect 983 123 1033 139
rect 526 53 768 87
rect 983 89 999 123
rect 983 17 1033 89
rect 1069 87 1103 175
rect 1139 204 1173 245
rect 1209 274 1243 315
rect 1324 326 1340 360
rect 1313 316 1340 326
rect 1279 310 1340 316
rect 1382 358 1448 374
rect 1382 324 1398 358
rect 1432 324 1448 358
rect 1382 290 1448 324
rect 1382 274 1398 290
rect 1209 256 1398 274
rect 1432 256 1448 290
rect 1490 368 1556 412
rect 1609 431 1625 465
rect 1659 438 1675 465
rect 1985 465 2051 563
rect 1985 438 2001 465
rect 1659 431 2001 438
rect 2035 431 2051 465
rect 1609 404 2051 431
rect 2097 527 2147 543
rect 2097 493 2113 527
rect 2097 456 2147 493
rect 2097 422 2113 456
rect 1490 352 1731 368
rect 1490 318 1686 352
rect 1720 318 1731 352
rect 1490 310 1731 318
rect 1490 276 1506 310
rect 1540 302 1731 310
rect 1540 276 1556 302
rect 1490 260 1556 276
rect 1209 240 1448 256
rect 1139 180 1231 204
rect 1139 146 1181 180
rect 1215 146 1231 180
rect 1139 123 1231 146
rect 1267 87 1301 240
rect 1767 213 1801 404
rect 2097 385 2147 422
rect 1837 352 1898 368
rect 1837 318 1848 352
rect 1882 318 1898 352
rect 1837 266 1898 318
rect 1940 352 2006 368
rect 1940 350 1956 352
rect 1940 316 1951 350
rect 1990 318 2006 352
rect 1985 316 2006 318
rect 1940 302 2006 316
rect 2097 351 2113 385
rect 2097 335 2147 351
rect 2097 266 2131 335
rect 2183 299 2217 579
rect 2253 527 2303 649
rect 2287 493 2303 527
rect 2253 456 2303 493
rect 2287 422 2303 456
rect 2253 385 2303 422
rect 2287 351 2303 385
rect 2253 335 2303 351
rect 2339 562 2415 578
rect 2339 528 2365 562
rect 2399 528 2415 562
rect 2339 491 2415 528
rect 2339 457 2365 491
rect 2399 457 2415 491
rect 2339 420 2415 457
rect 2339 386 2365 420
rect 2399 386 2415 420
rect 2339 332 2415 386
rect 2455 562 2521 649
rect 2455 528 2471 562
rect 2505 528 2521 562
rect 2455 491 2521 528
rect 2455 457 2471 491
rect 2505 457 2521 491
rect 2455 420 2521 457
rect 2455 386 2471 420
rect 2505 386 2521 420
rect 2455 370 2521 386
rect 2561 562 2665 578
rect 2561 528 2577 562
rect 2611 528 2665 562
rect 2561 491 2665 528
rect 2561 457 2577 491
rect 2611 457 2665 491
rect 2561 420 2665 457
rect 2561 386 2577 420
rect 2611 386 2665 420
rect 2561 370 2665 386
rect 2339 316 2568 332
rect 1837 232 2131 266
rect 2167 283 2233 299
rect 2167 249 2183 283
rect 2217 249 2233 283
rect 1069 53 1301 87
rect 1337 179 1403 204
rect 1337 145 1353 179
rect 1387 145 1403 179
rect 1337 17 1403 145
rect 1592 184 1801 213
rect 1592 150 1608 184
rect 1642 179 1801 184
rect 1642 150 1658 179
rect 1592 121 1658 150
rect 1887 175 1953 196
rect 1887 141 1903 175
rect 1937 141 1953 175
rect 1887 17 1953 141
rect 2013 111 2079 232
rect 2167 215 2233 249
rect 2167 181 2183 215
rect 2217 181 2233 215
rect 2167 165 2233 181
rect 2339 298 2518 316
rect 2339 162 2373 298
rect 2502 282 2518 298
rect 2552 282 2568 316
rect 2502 248 2568 282
rect 2502 214 2518 248
rect 2552 214 2568 248
rect 2502 198 2568 214
rect 2617 162 2665 370
rect 2283 133 2373 162
rect 2013 77 2029 111
rect 2063 77 2079 111
rect 2013 53 2079 77
rect 2171 103 2237 129
rect 2171 69 2187 103
rect 2221 69 2237 103
rect 2283 99 2299 133
rect 2333 99 2373 133
rect 2283 70 2373 99
rect 2441 133 2507 162
rect 2441 99 2457 133
rect 2491 99 2507 133
rect 2171 17 2237 69
rect 2441 17 2507 99
rect 2599 133 2665 162
rect 2599 99 2615 133
rect 2649 99 2665 133
rect 2599 70 2665 99
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 1279 326 1290 350
rect 1290 326 1313 350
rect 1279 316 1313 326
rect 1951 318 1956 350
rect 1956 318 1985 350
rect 1951 316 1985 318
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 683 2688 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2688 683
rect 0 617 2688 649
rect 1267 350 1325 356
rect 1267 316 1279 350
rect 1313 347 1325 350
rect 1939 350 1997 356
rect 1939 347 1951 350
rect 1313 319 1951 347
rect 1313 316 1325 319
rect 1267 310 1325 316
rect 1939 316 1951 319
rect 1985 316 1997 350
rect 1939 310 1997 316
rect 0 17 2688 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -49 2688 -17
<< labels >>
flabel pwell s 0 0 2688 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2688 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfstp_lp
flabel metal1 s 1951 316 1985 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel metal1 s 0 617 2688 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2688 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2623 94 2657 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2623 168 2657 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2623 242 2657 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2623 316 2657 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2623 390 2657 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2623 464 2657 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2623 538 2657 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2688 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 73606
string GDS_START 55896
<< end >>
