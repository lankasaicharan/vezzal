magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
<< pwell >>
rect 21 241 639 243
rect 21 49 1535 241
rect 0 0 1536 49
<< scnmos >>
rect 100 49 130 217
rect 186 49 216 217
rect 272 49 302 217
rect 358 49 388 217
rect 444 49 474 217
rect 530 49 560 217
rect 720 47 750 215
rect 806 47 836 215
rect 892 47 922 215
rect 978 47 1008 215
rect 1168 47 1198 215
rect 1254 47 1284 215
rect 1340 47 1370 215
rect 1426 47 1456 215
<< scpmoshvt >>
rect 100 367 130 619
rect 186 367 216 619
rect 272 367 302 619
rect 358 367 388 619
rect 548 367 578 619
rect 634 367 664 619
rect 720 367 750 619
rect 806 367 836 619
rect 892 367 922 619
rect 987 367 1017 619
rect 1073 367 1103 619
rect 1159 367 1189 619
rect 1245 367 1275 619
rect 1331 367 1361 619
<< ndiff >>
rect 47 177 100 217
rect 47 143 55 177
rect 89 143 100 177
rect 47 95 100 143
rect 47 61 55 95
rect 89 61 100 95
rect 47 49 100 61
rect 130 205 186 217
rect 130 171 141 205
rect 175 171 186 205
rect 130 101 186 171
rect 130 67 141 101
rect 175 67 186 101
rect 130 49 186 67
rect 216 177 272 217
rect 216 143 227 177
rect 261 143 272 177
rect 216 91 272 143
rect 216 57 227 91
rect 261 57 272 91
rect 216 49 272 57
rect 302 205 358 217
rect 302 171 313 205
rect 347 171 358 205
rect 302 101 358 171
rect 302 67 313 101
rect 347 67 358 101
rect 302 49 358 67
rect 388 205 444 217
rect 388 171 399 205
rect 433 171 444 205
rect 388 95 444 171
rect 388 61 399 95
rect 433 61 444 95
rect 388 49 444 61
rect 474 209 530 217
rect 474 175 485 209
rect 519 175 530 209
rect 474 101 530 175
rect 474 67 485 101
rect 519 67 530 101
rect 474 49 530 67
rect 560 99 613 217
rect 560 65 571 99
rect 605 65 613 99
rect 560 49 613 65
rect 667 97 720 215
rect 667 63 675 97
rect 709 63 720 97
rect 667 47 720 63
rect 750 187 806 215
rect 750 153 761 187
rect 795 153 806 187
rect 750 47 806 153
rect 836 192 892 215
rect 836 158 847 192
rect 881 158 892 192
rect 836 101 892 158
rect 836 67 847 101
rect 881 67 892 101
rect 836 47 892 67
rect 922 103 978 215
rect 922 69 933 103
rect 967 69 978 103
rect 922 47 978 69
rect 1008 193 1061 215
rect 1008 159 1019 193
rect 1053 159 1061 193
rect 1008 47 1061 159
rect 1115 193 1168 215
rect 1115 159 1123 193
rect 1157 159 1168 193
rect 1115 47 1168 159
rect 1198 103 1254 215
rect 1198 69 1209 103
rect 1243 69 1254 103
rect 1198 47 1254 69
rect 1284 192 1340 215
rect 1284 158 1295 192
rect 1329 158 1340 192
rect 1284 101 1340 158
rect 1284 67 1295 101
rect 1329 67 1340 101
rect 1284 47 1340 67
rect 1370 124 1426 215
rect 1370 90 1381 124
rect 1415 90 1426 124
rect 1370 47 1426 90
rect 1456 192 1509 215
rect 1456 158 1467 192
rect 1501 158 1509 192
rect 1456 101 1509 158
rect 1456 67 1467 101
rect 1501 67 1509 101
rect 1456 47 1509 67
<< pdiff >>
rect 47 607 100 619
rect 47 573 55 607
rect 89 573 100 607
rect 47 529 100 573
rect 47 495 55 529
rect 89 495 100 529
rect 47 453 100 495
rect 47 419 55 453
rect 89 419 100 453
rect 47 367 100 419
rect 130 599 186 619
rect 130 565 141 599
rect 175 565 186 599
rect 130 508 186 565
rect 130 474 141 508
rect 175 474 186 508
rect 130 413 186 474
rect 130 379 141 413
rect 175 379 186 413
rect 130 367 186 379
rect 216 607 272 619
rect 216 573 227 607
rect 261 573 272 607
rect 216 529 272 573
rect 216 495 227 529
rect 261 495 272 529
rect 216 453 272 495
rect 216 419 227 453
rect 261 419 272 453
rect 216 367 272 419
rect 302 599 358 619
rect 302 565 313 599
rect 347 565 358 599
rect 302 508 358 565
rect 302 474 313 508
rect 347 474 358 508
rect 302 413 358 474
rect 302 379 313 413
rect 347 379 358 413
rect 302 367 358 379
rect 388 607 441 619
rect 388 573 399 607
rect 433 573 441 607
rect 388 508 441 573
rect 388 474 399 508
rect 433 474 441 508
rect 388 413 441 474
rect 388 379 399 413
rect 433 379 441 413
rect 388 367 441 379
rect 495 599 548 619
rect 495 565 503 599
rect 537 565 548 599
rect 495 529 548 565
rect 495 495 503 529
rect 537 495 548 529
rect 495 459 548 495
rect 495 425 503 459
rect 537 425 548 459
rect 495 367 548 425
rect 578 539 634 619
rect 578 505 589 539
rect 623 505 634 539
rect 578 413 634 505
rect 578 379 589 413
rect 623 379 634 413
rect 578 367 634 379
rect 664 599 720 619
rect 664 565 675 599
rect 709 565 720 599
rect 664 508 720 565
rect 664 474 675 508
rect 709 474 720 508
rect 664 413 720 474
rect 664 379 675 413
rect 709 379 720 413
rect 664 367 720 379
rect 750 607 806 619
rect 750 573 761 607
rect 795 573 806 607
rect 750 529 806 573
rect 750 495 761 529
rect 795 495 806 529
rect 750 453 806 495
rect 750 419 761 453
rect 795 419 806 453
rect 750 367 806 419
rect 836 599 892 619
rect 836 565 847 599
rect 881 565 892 599
rect 836 508 892 565
rect 836 474 847 508
rect 881 474 892 508
rect 836 413 892 474
rect 836 379 847 413
rect 881 379 892 413
rect 836 367 892 379
rect 922 607 987 619
rect 922 573 937 607
rect 971 573 987 607
rect 922 529 987 573
rect 922 495 937 529
rect 971 495 987 529
rect 922 453 987 495
rect 922 419 937 453
rect 971 419 987 453
rect 922 367 987 419
rect 1017 599 1073 619
rect 1017 565 1028 599
rect 1062 565 1073 599
rect 1017 508 1073 565
rect 1017 474 1028 508
rect 1062 474 1073 508
rect 1017 413 1073 474
rect 1017 379 1028 413
rect 1062 379 1073 413
rect 1017 367 1073 379
rect 1103 607 1159 619
rect 1103 573 1114 607
rect 1148 573 1159 607
rect 1103 529 1159 573
rect 1103 495 1114 529
rect 1148 495 1159 529
rect 1103 453 1159 495
rect 1103 419 1114 453
rect 1148 419 1159 453
rect 1103 367 1159 419
rect 1189 599 1245 619
rect 1189 565 1200 599
rect 1234 565 1245 599
rect 1189 508 1245 565
rect 1189 474 1200 508
rect 1234 474 1245 508
rect 1189 413 1245 474
rect 1189 379 1200 413
rect 1234 379 1245 413
rect 1189 367 1245 379
rect 1275 607 1331 619
rect 1275 573 1286 607
rect 1320 573 1331 607
rect 1275 529 1331 573
rect 1275 495 1286 529
rect 1320 495 1331 529
rect 1275 453 1331 495
rect 1275 419 1286 453
rect 1320 419 1331 453
rect 1275 367 1331 419
rect 1361 599 1414 619
rect 1361 565 1372 599
rect 1406 565 1414 599
rect 1361 508 1414 565
rect 1361 474 1372 508
rect 1406 474 1414 508
rect 1361 413 1414 474
rect 1361 379 1372 413
rect 1406 379 1414 413
rect 1361 367 1414 379
<< ndiffc >>
rect 55 143 89 177
rect 55 61 89 95
rect 141 171 175 205
rect 141 67 175 101
rect 227 143 261 177
rect 227 57 261 91
rect 313 171 347 205
rect 313 67 347 101
rect 399 171 433 205
rect 399 61 433 95
rect 485 175 519 209
rect 485 67 519 101
rect 571 65 605 99
rect 675 63 709 97
rect 761 153 795 187
rect 847 158 881 192
rect 847 67 881 101
rect 933 69 967 103
rect 1019 159 1053 193
rect 1123 159 1157 193
rect 1209 69 1243 103
rect 1295 158 1329 192
rect 1295 67 1329 101
rect 1381 90 1415 124
rect 1467 158 1501 192
rect 1467 67 1501 101
<< pdiffc >>
rect 55 573 89 607
rect 55 495 89 529
rect 55 419 89 453
rect 141 565 175 599
rect 141 474 175 508
rect 141 379 175 413
rect 227 573 261 607
rect 227 495 261 529
rect 227 419 261 453
rect 313 565 347 599
rect 313 474 347 508
rect 313 379 347 413
rect 399 573 433 607
rect 399 474 433 508
rect 399 379 433 413
rect 503 565 537 599
rect 503 495 537 529
rect 503 425 537 459
rect 589 505 623 539
rect 589 379 623 413
rect 675 565 709 599
rect 675 474 709 508
rect 675 379 709 413
rect 761 573 795 607
rect 761 495 795 529
rect 761 419 795 453
rect 847 565 881 599
rect 847 474 881 508
rect 847 379 881 413
rect 937 573 971 607
rect 937 495 971 529
rect 937 419 971 453
rect 1028 565 1062 599
rect 1028 474 1062 508
rect 1028 379 1062 413
rect 1114 573 1148 607
rect 1114 495 1148 529
rect 1114 419 1148 453
rect 1200 565 1234 599
rect 1200 474 1234 508
rect 1200 379 1234 413
rect 1286 573 1320 607
rect 1286 495 1320 529
rect 1286 419 1320 453
rect 1372 565 1406 599
rect 1372 474 1406 508
rect 1372 379 1406 413
<< poly >>
rect 100 619 130 645
rect 186 619 216 645
rect 272 619 302 645
rect 358 619 388 645
rect 548 619 578 645
rect 634 619 664 645
rect 720 619 750 645
rect 806 619 836 645
rect 892 619 922 645
rect 987 619 1017 645
rect 1073 619 1103 645
rect 1159 619 1189 645
rect 1245 619 1275 645
rect 1331 619 1361 645
rect 100 331 130 367
rect 186 331 216 367
rect 272 331 302 367
rect 358 331 388 367
rect 100 315 388 331
rect 100 281 134 315
rect 168 281 202 315
rect 236 281 270 315
rect 304 281 338 315
rect 372 281 388 315
rect 548 305 578 367
rect 634 305 664 367
rect 100 265 388 281
rect 100 217 130 265
rect 186 217 216 265
rect 272 217 302 265
rect 358 217 388 265
rect 444 289 664 305
rect 444 255 555 289
rect 589 255 664 289
rect 444 239 664 255
rect 444 217 474 239
rect 530 238 664 239
rect 720 303 750 367
rect 806 303 836 367
rect 892 303 922 367
rect 987 303 1017 367
rect 1073 303 1103 367
rect 1159 303 1189 367
rect 1245 339 1275 367
rect 1331 339 1361 367
rect 1245 315 1456 339
rect 1245 309 1406 315
rect 720 287 844 303
rect 720 253 794 287
rect 828 253 844 287
rect 530 217 560 238
rect 720 237 844 253
rect 892 287 1031 303
rect 892 253 981 287
rect 1015 253 1031 287
rect 892 237 1031 253
rect 1073 287 1189 303
rect 1073 253 1114 287
rect 1148 267 1189 287
rect 1340 281 1406 309
rect 1440 281 1456 315
rect 1148 253 1284 267
rect 1073 237 1284 253
rect 720 215 750 237
rect 806 215 836 237
rect 892 215 922 237
rect 978 215 1008 237
rect 1168 215 1198 237
rect 1254 215 1284 237
rect 1340 265 1456 281
rect 1340 215 1370 265
rect 1426 215 1456 265
rect 100 23 130 49
rect 186 23 216 49
rect 272 23 302 49
rect 358 23 388 49
rect 444 23 474 49
rect 530 23 560 49
rect 720 21 750 47
rect 806 21 836 47
rect 892 21 922 47
rect 978 21 1008 47
rect 1168 21 1198 47
rect 1254 21 1284 47
rect 1340 21 1370 47
rect 1426 21 1456 47
<< polycont >>
rect 134 281 168 315
rect 202 281 236 315
rect 270 281 304 315
rect 338 281 372 315
rect 555 255 589 289
rect 794 253 828 287
rect 981 253 1015 287
rect 1114 253 1148 287
rect 1406 281 1440 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 39 607 105 649
rect 39 573 55 607
rect 89 573 105 607
rect 39 529 105 573
rect 39 495 55 529
rect 89 495 105 529
rect 39 453 105 495
rect 39 419 55 453
rect 89 419 105 453
rect 139 599 177 615
rect 139 565 141 599
rect 175 565 177 599
rect 139 508 177 565
rect 139 474 141 508
rect 175 474 177 508
rect 139 413 177 474
rect 211 607 277 649
rect 211 573 227 607
rect 261 573 277 607
rect 211 529 277 573
rect 211 495 227 529
rect 261 495 277 529
rect 211 453 277 495
rect 211 419 227 453
rect 261 419 277 453
rect 311 599 356 615
rect 311 565 313 599
rect 347 565 356 599
rect 311 508 356 565
rect 311 474 313 508
rect 347 474 356 508
rect 139 385 141 413
rect 20 379 141 385
rect 175 385 177 413
rect 311 413 356 474
rect 311 385 313 413
rect 175 379 313 385
rect 347 379 356 413
rect 20 351 356 379
rect 390 607 447 649
rect 390 573 399 607
rect 433 573 447 607
rect 390 508 447 573
rect 390 474 399 508
rect 433 474 447 508
rect 390 413 447 474
rect 390 379 399 413
rect 433 379 447 413
rect 487 599 711 615
rect 487 565 503 599
rect 537 581 675 599
rect 537 565 539 581
rect 487 529 539 565
rect 673 565 675 581
rect 709 565 711 599
rect 487 495 503 529
rect 537 495 539 529
rect 487 459 539 495
rect 487 425 503 459
rect 537 425 539 459
rect 487 409 539 425
rect 573 539 639 547
rect 573 505 589 539
rect 623 505 639 539
rect 573 413 639 505
rect 390 363 447 379
rect 573 379 589 413
rect 623 379 639 413
rect 573 375 639 379
rect 20 245 84 351
rect 481 341 639 375
rect 673 508 711 565
rect 673 474 675 508
rect 709 474 711 508
rect 673 413 711 474
rect 745 607 811 649
rect 745 573 761 607
rect 795 573 811 607
rect 745 529 811 573
rect 745 495 761 529
rect 795 495 811 529
rect 745 453 811 495
rect 745 419 761 453
rect 795 419 811 453
rect 845 599 883 615
rect 845 565 847 599
rect 881 565 883 599
rect 845 508 883 565
rect 845 474 847 508
rect 881 474 883 508
rect 673 379 675 413
rect 709 385 711 413
rect 845 413 883 474
rect 921 607 987 649
rect 921 573 937 607
rect 971 573 987 607
rect 921 529 987 573
rect 921 495 937 529
rect 971 495 987 529
rect 921 453 987 495
rect 921 419 937 453
rect 971 419 987 453
rect 1022 599 1064 615
rect 1022 565 1028 599
rect 1062 565 1064 599
rect 1022 508 1064 565
rect 1022 474 1028 508
rect 1062 474 1064 508
rect 845 385 847 413
rect 709 379 847 385
rect 881 385 883 413
rect 1022 413 1064 474
rect 1098 607 1164 649
rect 1098 573 1114 607
rect 1148 573 1164 607
rect 1098 529 1164 573
rect 1098 495 1114 529
rect 1148 495 1164 529
rect 1098 453 1164 495
rect 1098 419 1114 453
rect 1148 419 1164 453
rect 1198 599 1236 615
rect 1198 565 1200 599
rect 1234 565 1236 599
rect 1198 508 1236 565
rect 1198 474 1200 508
rect 1234 474 1236 508
rect 1022 385 1028 413
rect 881 379 1028 385
rect 1062 385 1064 413
rect 1198 413 1236 474
rect 1270 607 1336 649
rect 1270 573 1286 607
rect 1320 573 1336 607
rect 1270 529 1336 573
rect 1270 495 1286 529
rect 1320 495 1336 529
rect 1270 453 1336 495
rect 1270 419 1286 453
rect 1320 419 1336 453
rect 1370 599 1422 615
rect 1370 565 1372 599
rect 1406 565 1422 599
rect 1370 508 1422 565
rect 1370 474 1372 508
rect 1406 474 1422 508
rect 1198 385 1200 413
rect 1062 379 1200 385
rect 1234 385 1236 413
rect 1370 413 1422 474
rect 1370 385 1372 413
rect 1234 379 1372 385
rect 1406 379 1422 413
rect 673 351 1422 379
rect 481 315 519 341
rect 118 281 134 315
rect 168 281 202 315
rect 236 281 270 315
rect 304 281 338 315
rect 372 281 519 315
rect 20 211 356 245
rect 139 205 177 211
rect 39 143 55 177
rect 89 143 105 177
rect 39 95 105 143
rect 39 61 55 95
rect 89 61 105 95
rect 39 17 105 61
rect 139 171 141 205
rect 175 171 177 205
rect 311 205 356 211
rect 139 101 177 171
rect 139 67 141 101
rect 175 67 177 101
rect 139 51 177 67
rect 211 143 227 177
rect 261 143 277 177
rect 211 91 277 143
rect 211 57 227 91
rect 261 57 277 91
rect 211 17 277 57
rect 311 171 313 205
rect 347 171 356 205
rect 311 101 356 171
rect 311 67 313 101
rect 347 67 356 101
rect 311 51 356 67
rect 390 205 442 221
rect 390 171 399 205
rect 433 171 442 205
rect 390 95 442 171
rect 390 61 399 95
rect 433 61 442 95
rect 390 17 442 61
rect 476 209 519 281
rect 553 289 744 307
rect 553 255 555 289
rect 589 255 744 289
rect 553 239 744 255
rect 778 287 940 317
rect 778 253 794 287
rect 828 253 940 287
rect 778 242 940 253
rect 974 287 1034 303
rect 974 253 981 287
rect 1015 253 1034 287
rect 974 237 1034 253
rect 1073 287 1217 304
rect 1073 253 1114 287
rect 1148 253 1217 287
rect 1073 242 1217 253
rect 1279 281 1406 315
rect 1440 281 1516 315
rect 1279 242 1516 281
rect 476 175 485 209
rect 519 187 797 203
rect 519 175 761 187
rect 476 153 761 175
rect 795 153 797 187
rect 476 137 797 153
rect 831 193 1069 203
rect 831 192 1019 193
rect 831 158 847 192
rect 881 159 1019 192
rect 1053 159 1069 193
rect 881 158 1069 159
rect 831 153 1069 158
rect 1107 193 1517 208
rect 1107 159 1123 193
rect 1157 192 1517 193
rect 1157 159 1295 192
rect 1107 158 1295 159
rect 1329 174 1467 192
rect 1329 158 1331 174
rect 1107 153 1331 158
rect 476 101 521 137
rect 476 67 485 101
rect 519 67 521 101
rect 476 51 521 67
rect 555 99 621 103
rect 831 101 885 153
rect 555 65 571 99
rect 605 65 621 99
rect 555 17 621 65
rect 659 97 847 101
rect 659 63 675 97
rect 709 67 847 97
rect 881 67 885 101
rect 709 63 885 67
rect 659 51 885 63
rect 919 103 1247 119
rect 919 69 933 103
rect 967 69 1209 103
rect 1243 69 1247 103
rect 919 53 1247 69
rect 1281 101 1331 153
rect 1465 158 1467 174
rect 1501 158 1517 192
rect 1281 67 1295 101
rect 1329 67 1331 101
rect 1281 51 1331 67
rect 1365 124 1431 140
rect 1365 90 1381 124
rect 1415 90 1431 124
rect 1365 17 1431 90
rect 1465 101 1517 158
rect 1465 67 1467 101
rect 1501 67 1517 101
rect 1465 51 1517 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a41o_4
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5499798
string GDS_START 5486578
<< end >>
