magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1586 1975
<< nwell >>
rect -38 331 326 704
<< pwell >>
rect 1 49 287 241
rect 0 0 288 49
<< scnmos >>
rect 80 47 110 215
rect 178 131 208 215
<< scpmoshvt >>
rect 80 367 110 619
rect 178 367 208 495
<< ndiff >>
rect 27 190 80 215
rect 27 156 35 190
rect 69 156 80 190
rect 27 101 80 156
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 131 178 215
rect 208 188 261 215
rect 208 154 219 188
rect 253 154 261 188
rect 208 131 261 154
rect 110 128 163 131
rect 110 94 121 128
rect 155 94 163 128
rect 110 47 163 94
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 507 80 565
rect 27 473 35 507
rect 69 473 80 507
rect 27 423 80 473
rect 27 389 35 423
rect 69 389 80 423
rect 27 367 80 389
rect 110 607 163 619
rect 110 573 121 607
rect 155 573 163 607
rect 110 516 163 573
rect 110 482 121 516
rect 155 495 163 516
rect 155 482 178 495
rect 110 428 178 482
rect 110 394 121 428
rect 155 394 178 428
rect 110 367 178 394
rect 208 481 261 495
rect 208 447 219 481
rect 253 447 261 481
rect 208 413 261 447
rect 208 379 219 413
rect 253 379 261 413
rect 208 367 261 379
<< ndiffc >>
rect 35 156 69 190
rect 35 67 69 101
rect 219 154 253 188
rect 121 94 155 128
<< pdiffc >>
rect 35 565 69 599
rect 35 473 69 507
rect 35 389 69 423
rect 121 573 155 607
rect 121 482 155 516
rect 121 394 155 428
rect 219 447 253 481
rect 219 379 253 413
<< poly >>
rect 80 619 110 645
rect 178 495 208 521
rect 80 303 110 367
rect 178 303 208 367
rect 70 287 136 303
rect 70 253 86 287
rect 120 253 136 287
rect 70 237 136 253
rect 178 287 267 303
rect 178 253 217 287
rect 251 253 267 287
rect 178 237 267 253
rect 80 215 110 237
rect 178 215 208 237
rect 178 105 208 131
rect 80 21 110 47
<< polycont >>
rect 86 253 120 287
rect 217 253 251 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 17 599 71 615
rect 17 565 35 599
rect 69 565 71 599
rect 17 507 71 565
rect 17 473 35 507
rect 69 473 71 507
rect 17 423 71 473
rect 17 389 35 423
rect 69 389 71 423
rect 105 607 171 649
rect 105 573 121 607
rect 155 573 171 607
rect 105 516 171 573
rect 105 482 121 516
rect 155 482 171 516
rect 105 428 171 482
rect 105 394 121 428
rect 155 394 171 428
rect 105 389 171 394
rect 205 481 269 497
rect 205 447 219 481
rect 253 447 269 481
rect 205 413 269 447
rect 17 373 71 389
rect 205 379 219 413
rect 253 379 269 413
rect 17 206 52 373
rect 205 355 269 379
rect 101 341 269 355
rect 86 321 269 341
rect 86 287 139 321
rect 120 253 139 287
rect 86 237 139 253
rect 201 253 217 287
rect 251 253 271 287
rect 201 238 271 253
rect 17 190 71 206
rect 17 156 35 190
rect 69 156 71 190
rect 105 204 139 237
rect 105 188 269 204
rect 105 170 219 188
rect 17 101 71 156
rect 205 154 219 170
rect 253 154 269 188
rect 205 138 269 154
rect 17 67 35 101
rect 69 67 71 101
rect 17 51 71 67
rect 105 128 171 136
rect 105 94 121 128
rect 155 94 171 128
rect 105 17 171 94
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
<< metal1 >>
rect 0 683 288 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 0 617 288 649
rect 0 17 288 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
rect 0 -49 288 -17
<< labels >>
flabel pwell s 0 0 288 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 288 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 busreceiver_1
flabel metal1 s 0 617 288 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 288 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 288 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y
string GDS_END 2662034
string GDS_START 2657914
<< end >>
