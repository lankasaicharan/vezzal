magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
rect 770 318 938 331
<< pwell >>
rect 781 241 891 263
rect 6 230 191 241
rect 6 191 194 230
rect 781 191 1625 241
rect 6 49 1625 191
rect 0 0 1632 49
<< scnmos >>
rect 85 47 115 215
rect 223 81 253 165
rect 295 81 325 165
rect 381 81 411 165
rect 475 81 505 165
rect 584 81 614 165
rect 887 131 917 215
rect 996 47 1026 215
rect 1068 47 1098 215
rect 1258 47 1288 215
rect 1344 47 1374 215
rect 1430 47 1460 215
rect 1516 47 1546 215
<< scpmoshvt >>
rect 80 367 110 619
rect 205 465 235 593
rect 277 465 307 593
rect 385 465 415 549
rect 457 465 487 549
rect 626 419 656 547
rect 924 367 954 495
rect 1048 367 1078 619
rect 1134 367 1164 619
rect 1228 367 1258 619
rect 1314 367 1344 619
rect 1400 367 1430 619
rect 1486 367 1516 619
<< ndiff >>
rect 32 203 85 215
rect 32 169 40 203
rect 74 169 85 203
rect 32 101 85 169
rect 32 67 40 101
rect 74 67 85 101
rect 32 47 85 67
rect 115 204 165 215
rect 115 165 168 204
rect 807 229 865 237
rect 807 195 819 229
rect 853 215 865 229
rect 853 195 887 215
rect 115 124 223 165
rect 115 90 126 124
rect 160 90 223 124
rect 115 81 223 90
rect 253 81 295 165
rect 325 157 381 165
rect 325 123 336 157
rect 370 123 381 157
rect 325 81 381 123
rect 411 81 475 165
rect 505 140 584 165
rect 505 106 539 140
rect 573 106 584 140
rect 505 81 584 106
rect 614 143 667 165
rect 614 109 625 143
rect 659 109 667 143
rect 807 131 887 195
rect 917 131 996 215
rect 614 81 667 109
rect 939 89 996 131
rect 115 47 168 81
rect 939 55 951 89
rect 985 55 996 89
rect 939 47 996 55
rect 1026 47 1068 215
rect 1098 203 1151 215
rect 1098 169 1109 203
rect 1143 169 1151 203
rect 1098 101 1151 169
rect 1098 67 1109 101
rect 1143 67 1151 101
rect 1098 47 1151 67
rect 1205 179 1258 215
rect 1205 145 1213 179
rect 1247 145 1258 179
rect 1205 93 1258 145
rect 1205 59 1213 93
rect 1247 59 1258 93
rect 1205 47 1258 59
rect 1288 203 1344 215
rect 1288 169 1299 203
rect 1333 169 1344 203
rect 1288 101 1344 169
rect 1288 67 1299 101
rect 1333 67 1344 101
rect 1288 47 1344 67
rect 1374 181 1430 215
rect 1374 147 1385 181
rect 1419 147 1430 181
rect 1374 93 1430 147
rect 1374 59 1385 93
rect 1419 59 1430 93
rect 1374 47 1430 59
rect 1460 203 1516 215
rect 1460 169 1471 203
rect 1505 169 1516 203
rect 1460 101 1516 169
rect 1460 67 1471 101
rect 1505 67 1516 101
rect 1460 47 1516 67
rect 1546 203 1599 215
rect 1546 169 1557 203
rect 1591 169 1599 203
rect 1546 93 1599 169
rect 1546 59 1557 93
rect 1591 59 1599 93
rect 1546 47 1599 59
<< pdiff >>
rect 125 630 183 638
rect 125 619 137 630
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 513 80 565
rect 27 479 35 513
rect 69 479 80 513
rect 27 420 80 479
rect 27 386 35 420
rect 69 386 80 420
rect 27 367 80 386
rect 110 596 137 619
rect 171 596 183 630
rect 110 593 183 596
rect 110 465 205 593
rect 235 465 277 593
rect 307 549 360 593
rect 509 566 611 584
rect 509 549 521 566
rect 307 531 385 549
rect 307 497 318 531
rect 352 497 385 531
rect 307 465 385 497
rect 415 465 457 549
rect 487 532 521 549
rect 555 547 611 566
rect 976 607 1048 619
rect 976 573 984 607
rect 1018 573 1048 607
rect 555 532 626 547
rect 487 465 626 532
rect 110 367 183 465
rect 509 419 626 465
rect 656 523 706 547
rect 656 491 731 523
rect 976 495 1048 573
rect 656 457 681 491
rect 715 457 731 491
rect 656 419 731 457
rect 844 396 924 495
rect 844 362 856 396
rect 890 367 924 396
rect 954 367 1048 495
rect 1078 452 1134 619
rect 1078 418 1089 452
rect 1123 418 1134 452
rect 1078 367 1134 418
rect 1164 607 1228 619
rect 1164 573 1175 607
rect 1209 573 1228 607
rect 1164 367 1228 573
rect 1258 599 1314 619
rect 1258 565 1269 599
rect 1303 565 1314 599
rect 1258 506 1314 565
rect 1258 472 1269 506
rect 1303 472 1314 506
rect 1258 413 1314 472
rect 1258 379 1269 413
rect 1303 379 1314 413
rect 1258 367 1314 379
rect 1344 607 1400 619
rect 1344 573 1355 607
rect 1389 573 1400 607
rect 1344 539 1400 573
rect 1344 505 1355 539
rect 1389 505 1400 539
rect 1344 471 1400 505
rect 1344 437 1355 471
rect 1389 437 1400 471
rect 1344 367 1400 437
rect 1430 599 1486 619
rect 1430 565 1441 599
rect 1475 565 1486 599
rect 1430 504 1486 565
rect 1430 470 1441 504
rect 1475 470 1486 504
rect 1430 413 1486 470
rect 1430 379 1441 413
rect 1475 379 1486 413
rect 1430 367 1486 379
rect 1516 607 1583 619
rect 1516 573 1541 607
rect 1575 573 1583 607
rect 1516 506 1583 573
rect 1516 472 1541 506
rect 1575 472 1583 506
rect 1516 413 1583 472
rect 1516 379 1541 413
rect 1575 379 1583 413
rect 1516 367 1583 379
rect 890 362 902 367
rect 844 354 902 362
<< ndiffc >>
rect 40 169 74 203
rect 40 67 74 101
rect 819 195 853 229
rect 126 90 160 124
rect 336 123 370 157
rect 539 106 573 140
rect 625 109 659 143
rect 951 55 985 89
rect 1109 169 1143 203
rect 1109 67 1143 101
rect 1213 145 1247 179
rect 1213 59 1247 93
rect 1299 169 1333 203
rect 1299 67 1333 101
rect 1385 147 1419 181
rect 1385 59 1419 93
rect 1471 169 1505 203
rect 1471 67 1505 101
rect 1557 169 1591 203
rect 1557 59 1591 93
<< pdiffc >>
rect 35 565 69 599
rect 35 479 69 513
rect 35 386 69 420
rect 137 596 171 630
rect 318 497 352 531
rect 521 532 555 566
rect 984 573 1018 607
rect 681 457 715 491
rect 856 362 890 396
rect 1089 418 1123 452
rect 1175 573 1209 607
rect 1269 565 1303 599
rect 1269 472 1303 506
rect 1269 379 1303 413
rect 1355 573 1389 607
rect 1355 505 1389 539
rect 1355 437 1389 471
rect 1441 565 1475 599
rect 1441 470 1475 504
rect 1441 379 1475 413
rect 1541 573 1575 607
rect 1541 472 1575 506
rect 1541 379 1575 413
<< poly >>
rect 80 619 110 645
rect 205 593 235 619
rect 277 593 307 619
rect 457 615 829 645
rect 1048 619 1078 645
rect 1134 619 1164 645
rect 1228 619 1258 645
rect 1314 619 1344 645
rect 1400 619 1430 645
rect 1486 619 1516 645
rect 385 549 415 575
rect 457 549 487 615
rect 763 605 829 615
rect 626 547 656 573
rect 763 571 779 605
rect 813 571 829 605
rect 763 555 829 571
rect 80 335 110 367
rect 73 319 139 335
rect 73 285 89 319
rect 123 285 139 319
rect 205 292 235 465
rect 277 433 307 465
rect 277 417 343 433
rect 277 383 293 417
rect 327 383 343 417
rect 277 367 343 383
rect 385 361 415 465
rect 457 439 487 465
rect 924 495 954 521
rect 385 345 535 361
rect 385 325 485 345
rect 295 311 485 325
rect 519 311 535 345
rect 626 329 656 419
rect 924 339 954 367
rect 1048 339 1078 367
rect 295 295 535 311
rect 584 313 656 329
rect 73 269 139 285
rect 187 276 253 292
rect 85 215 115 269
rect 187 242 203 276
rect 237 242 253 276
rect 187 226 253 242
rect 223 165 253 226
rect 295 165 325 295
rect 584 279 600 313
rect 634 279 656 313
rect 367 237 433 253
rect 367 203 383 237
rect 417 203 433 237
rect 367 187 433 203
rect 475 237 541 253
rect 475 203 491 237
rect 525 203 541 237
rect 475 187 541 203
rect 584 245 656 279
rect 704 323 1078 339
rect 1134 333 1164 367
rect 1228 333 1258 367
rect 1314 333 1344 367
rect 1400 333 1430 367
rect 1486 333 1516 367
rect 704 289 720 323
rect 754 309 1078 323
rect 1120 317 1186 333
rect 754 289 770 309
rect 704 273 770 289
rect 584 211 600 245
rect 634 211 656 245
rect 584 195 656 211
rect 887 215 917 309
rect 996 215 1026 309
rect 1120 283 1136 317
rect 1170 283 1186 317
rect 1120 267 1186 283
rect 1228 317 1516 333
rect 1228 283 1245 317
rect 1279 283 1313 317
rect 1347 283 1381 317
rect 1415 297 1516 317
rect 1415 283 1546 297
rect 1228 267 1546 283
rect 1068 237 1186 267
rect 1068 215 1098 237
rect 1258 215 1288 267
rect 1344 215 1374 267
rect 1430 215 1460 267
rect 1516 215 1546 267
rect 381 165 411 187
rect 475 165 505 187
rect 584 165 614 195
rect 887 105 917 131
rect 223 55 253 81
rect 295 55 325 81
rect 381 55 411 81
rect 475 55 505 81
rect 584 55 614 81
rect 85 21 115 47
rect 996 21 1026 47
rect 1068 21 1098 47
rect 1258 21 1288 47
rect 1344 21 1374 47
rect 1430 21 1460 47
rect 1516 21 1546 47
<< polycont >>
rect 779 571 813 605
rect 89 285 123 319
rect 293 383 327 417
rect 485 311 519 345
rect 203 242 237 276
rect 600 279 634 313
rect 383 203 417 237
rect 491 203 525 237
rect 720 289 754 323
rect 600 211 634 245
rect 1136 283 1170 317
rect 1245 283 1279 317
rect 1313 283 1347 317
rect 1381 283 1415 317
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 121 630 187 649
rect 19 599 87 615
rect 19 565 35 599
rect 69 565 87 599
rect 121 596 137 630
rect 171 596 187 630
rect 121 594 187 596
rect 19 560 87 565
rect 223 581 438 615
rect 223 560 257 581
rect 19 526 257 560
rect 302 531 368 547
rect 19 513 85 526
rect 19 479 35 513
rect 69 479 85 513
rect 302 497 318 531
rect 352 497 368 531
rect 302 490 368 497
rect 19 420 85 479
rect 19 386 35 420
rect 69 386 85 420
rect 19 380 85 386
rect 207 456 368 490
rect 404 490 438 581
rect 505 566 571 649
rect 505 532 521 566
rect 555 532 571 566
rect 505 524 571 532
rect 605 605 908 615
rect 605 571 779 605
rect 813 571 908 605
rect 605 553 908 571
rect 968 607 1034 649
rect 968 573 984 607
rect 1018 573 1034 607
rect 968 570 1034 573
rect 1159 607 1225 649
rect 1159 573 1175 607
rect 1209 573 1225 607
rect 1159 570 1225 573
rect 1259 599 1305 615
rect 605 490 639 553
rect 761 536 908 553
rect 1259 565 1269 599
rect 1303 565 1305 599
rect 404 456 639 490
rect 673 491 727 507
rect 761 502 1195 536
rect 673 457 681 491
rect 715 468 727 491
rect 715 457 1016 468
rect 19 219 53 380
rect 207 346 241 456
rect 673 432 1016 457
rect 673 422 739 432
rect 277 417 739 422
rect 277 383 293 417
rect 327 386 739 417
rect 840 396 906 398
rect 327 383 433 386
rect 277 380 433 383
rect 87 319 331 346
rect 87 285 89 319
rect 123 312 331 319
rect 123 285 137 312
rect 87 269 137 285
rect 171 276 263 278
rect 171 242 203 276
rect 237 242 263 276
rect 171 234 263 242
rect 19 203 90 219
rect 19 169 40 203
rect 74 200 90 203
rect 74 169 246 200
rect 19 166 246 169
rect 19 101 76 166
rect 19 67 40 101
rect 74 67 76 101
rect 19 51 76 67
rect 110 124 178 132
rect 110 90 126 124
rect 160 90 178 124
rect 110 17 178 90
rect 212 87 246 166
rect 297 169 331 312
rect 367 237 433 380
rect 840 362 856 396
rect 890 362 906 396
rect 469 345 646 352
rect 469 311 485 345
rect 519 313 646 345
rect 519 311 600 313
rect 469 295 600 311
rect 584 279 600 295
rect 634 279 646 313
rect 367 203 383 237
rect 417 203 433 237
rect 469 237 541 253
rect 469 203 491 237
rect 525 203 541 237
rect 584 245 646 279
rect 680 323 770 352
rect 680 289 720 323
rect 754 289 770 323
rect 680 273 770 289
rect 584 211 600 245
rect 634 239 646 245
rect 840 239 906 362
rect 634 229 906 239
rect 634 211 819 229
rect 297 157 386 169
rect 297 123 336 157
rect 370 123 386 157
rect 297 121 386 123
rect 469 87 503 203
rect 584 195 819 211
rect 853 195 906 229
rect 584 193 906 195
rect 940 159 1016 432
rect 1050 452 1125 468
rect 1050 418 1089 452
rect 1123 418 1125 452
rect 1050 402 1125 418
rect 1050 247 1084 402
rect 1159 333 1195 502
rect 1259 506 1305 565
rect 1259 472 1269 506
rect 1303 472 1305 506
rect 1259 413 1305 472
rect 1339 607 1405 649
rect 1339 573 1355 607
rect 1389 573 1405 607
rect 1339 539 1405 573
rect 1339 505 1355 539
rect 1389 505 1405 539
rect 1339 471 1405 505
rect 1339 437 1355 471
rect 1389 437 1405 471
rect 1339 433 1405 437
rect 1439 599 1507 615
rect 1439 565 1441 599
rect 1475 565 1507 599
rect 1439 504 1507 565
rect 1439 470 1441 504
rect 1475 470 1507 504
rect 1259 379 1269 413
rect 1303 397 1305 413
rect 1439 413 1507 470
rect 1439 397 1441 413
rect 1303 379 1441 397
rect 1475 379 1507 413
rect 1259 363 1507 379
rect 1541 607 1591 649
rect 1575 573 1591 607
rect 1541 506 1591 573
rect 1575 472 1591 506
rect 1541 413 1591 472
rect 1575 379 1591 413
rect 1541 363 1591 379
rect 1120 317 1195 333
rect 1120 283 1136 317
rect 1170 283 1195 317
rect 1120 281 1195 283
rect 1229 283 1245 317
rect 1279 283 1313 317
rect 1347 283 1381 317
rect 1415 283 1431 317
rect 1229 247 1263 283
rect 1471 249 1507 363
rect 1050 213 1263 247
rect 1297 215 1507 249
rect 212 53 503 87
rect 537 140 589 156
rect 537 106 539 140
rect 573 106 589 140
rect 537 17 589 106
rect 623 143 1016 159
rect 623 109 625 143
rect 659 125 1016 143
rect 1093 203 1159 213
rect 1093 169 1109 203
rect 1143 169 1159 203
rect 1297 203 1335 215
rect 659 109 675 125
rect 623 93 675 109
rect 1093 101 1159 169
rect 935 89 1001 91
rect 935 55 951 89
rect 985 55 1001 89
rect 935 17 1001 55
rect 1093 67 1109 101
rect 1143 67 1159 101
rect 1093 51 1159 67
rect 1197 145 1213 179
rect 1247 145 1263 179
rect 1197 93 1263 145
rect 1197 59 1213 93
rect 1247 59 1263 93
rect 1197 17 1263 59
rect 1297 169 1299 203
rect 1333 169 1335 203
rect 1469 203 1507 215
rect 1297 101 1335 169
rect 1297 67 1299 101
rect 1333 67 1335 101
rect 1297 51 1335 67
rect 1369 147 1385 181
rect 1419 147 1435 181
rect 1369 93 1435 147
rect 1369 59 1385 93
rect 1419 59 1435 93
rect 1369 17 1435 59
rect 1469 169 1471 203
rect 1505 169 1507 203
rect 1469 101 1507 169
rect 1469 67 1471 101
rect 1505 67 1507 101
rect 1469 51 1507 67
rect 1548 203 1607 219
rect 1548 169 1557 203
rect 1591 169 1607 203
rect 1548 93 1607 169
rect 1548 59 1557 93
rect 1591 59 1607 93
rect 1548 17 1607 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlclkp_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1471 94 1505 128 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1471 168 1505 202 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1471 390 1505 424 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1471 464 1505 498 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1471 538 1505 572 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3525824
string GDS_START 3513298
<< end >>
