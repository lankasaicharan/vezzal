magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 306 165 863 235
rect 28 49 863 165
rect 0 0 864 49
<< scnmos >>
rect 107 55 137 139
rect 193 55 223 139
rect 385 125 415 209
rect 457 125 487 209
rect 565 125 595 209
rect 637 125 667 209
rect 754 125 784 209
<< scpmoshvt >>
rect 357 535 387 619
rect 443 535 473 619
rect 529 535 559 619
rect 615 535 645 619
rect 709 535 739 619
rect 107 397 137 481
rect 193 397 223 481
<< ndiff >>
rect 332 179 385 209
rect 332 145 340 179
rect 374 145 385 179
rect 54 109 107 139
rect 54 75 62 109
rect 96 75 107 109
rect 54 55 107 75
rect 137 101 193 139
rect 137 67 148 101
rect 182 67 193 101
rect 137 55 193 67
rect 223 103 276 139
rect 332 125 385 145
rect 415 125 457 209
rect 487 125 565 209
rect 595 125 637 209
rect 667 171 754 209
rect 667 137 705 171
rect 739 137 754 171
rect 667 125 754 137
rect 784 171 837 209
rect 784 137 795 171
rect 829 137 837 171
rect 784 125 837 137
rect 223 69 234 103
rect 268 69 276 103
rect 223 55 276 69
<< pdiff >>
rect 304 607 357 619
rect 304 573 312 607
rect 346 573 357 607
rect 304 535 357 573
rect 387 581 443 619
rect 387 547 398 581
rect 432 547 443 581
rect 387 535 443 547
rect 473 607 529 619
rect 473 573 484 607
rect 518 573 529 607
rect 473 535 529 573
rect 559 581 615 619
rect 559 547 570 581
rect 604 547 615 581
rect 559 535 615 547
rect 645 607 709 619
rect 645 573 660 607
rect 694 573 709 607
rect 645 535 709 573
rect 739 581 792 619
rect 739 547 750 581
rect 784 547 792 581
rect 739 535 792 547
rect 54 443 107 481
rect 54 409 62 443
rect 96 409 107 443
rect 54 397 107 409
rect 137 469 193 481
rect 137 435 148 469
rect 182 435 193 469
rect 137 397 193 435
rect 223 451 276 481
rect 223 417 234 451
rect 268 417 276 451
rect 223 397 276 417
<< ndiffc >>
rect 340 145 374 179
rect 62 75 96 109
rect 148 67 182 101
rect 705 137 739 171
rect 795 137 829 171
rect 234 69 268 103
<< pdiffc >>
rect 312 573 346 607
rect 398 547 432 581
rect 484 573 518 607
rect 570 547 604 581
rect 660 573 694 607
rect 750 547 784 581
rect 62 409 96 443
rect 148 435 182 469
rect 234 417 268 451
<< poly >>
rect 357 619 387 645
rect 443 619 473 645
rect 529 619 559 645
rect 615 619 645 645
rect 709 619 739 645
rect 357 513 387 535
rect 107 481 137 507
rect 193 481 223 507
rect 343 483 387 513
rect 107 295 137 397
rect 193 295 223 397
rect 343 365 373 483
rect 443 441 473 535
rect 307 349 373 365
rect 307 315 323 349
rect 357 315 373 349
rect 79 279 145 295
rect 79 245 95 279
rect 129 245 145 279
rect 79 211 145 245
rect 79 177 95 211
rect 129 177 145 211
rect 79 161 145 177
rect 193 279 259 295
rect 193 245 209 279
rect 243 245 259 279
rect 193 211 259 245
rect 307 281 373 315
rect 421 425 487 441
rect 421 391 437 425
rect 471 391 487 425
rect 421 357 487 391
rect 421 323 437 357
rect 471 323 487 357
rect 421 307 487 323
rect 307 247 323 281
rect 357 261 373 281
rect 357 247 415 261
rect 307 231 415 247
rect 193 177 209 211
rect 243 177 259 211
rect 385 209 415 231
rect 457 209 487 307
rect 529 297 559 535
rect 615 440 645 535
rect 709 451 739 535
rect 601 424 667 440
rect 601 390 617 424
rect 651 390 667 424
rect 601 374 667 390
rect 529 281 595 297
rect 529 247 545 281
rect 579 247 595 281
rect 529 231 595 247
rect 565 209 595 231
rect 637 209 667 374
rect 709 435 784 451
rect 709 401 725 435
rect 759 401 784 435
rect 709 367 784 401
rect 709 333 725 367
rect 759 333 784 367
rect 709 317 784 333
rect 754 209 784 317
rect 193 161 259 177
rect 107 139 137 161
rect 193 139 223 161
rect 385 99 415 125
rect 457 103 487 125
rect 457 87 523 103
rect 565 99 595 125
rect 637 99 667 125
rect 754 99 784 125
rect 107 29 137 55
rect 193 29 223 55
rect 457 53 473 87
rect 507 53 523 87
rect 457 37 523 53
<< polycont >>
rect 323 315 357 349
rect 95 245 129 279
rect 95 177 129 211
rect 209 245 243 279
rect 437 391 471 425
rect 437 323 471 357
rect 323 247 357 281
rect 209 177 243 211
rect 617 390 651 424
rect 545 247 579 281
rect 725 401 759 435
rect 725 333 759 367
rect 473 53 507 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 144 469 186 649
rect 308 607 350 649
rect 308 573 312 607
rect 346 573 350 607
rect 480 607 522 649
rect 308 557 350 573
rect 394 581 436 597
rect 394 547 398 581
rect 432 547 436 581
rect 480 573 484 607
rect 518 573 522 607
rect 644 607 710 649
rect 480 557 522 573
rect 566 581 608 597
rect 394 521 436 547
rect 566 547 570 581
rect 604 547 608 581
rect 644 573 660 607
rect 694 573 710 607
rect 644 569 710 573
rect 746 581 833 597
rect 566 521 608 547
rect 746 547 750 581
rect 784 547 833 581
rect 746 531 833 547
rect 394 487 608 521
rect 25 443 100 459
rect 25 409 62 443
rect 96 409 100 443
rect 144 435 148 469
rect 182 435 186 469
rect 144 419 186 435
rect 230 451 272 467
rect 25 365 100 409
rect 230 417 234 451
rect 268 435 272 451
rect 268 425 487 435
rect 268 417 437 425
rect 230 401 437 417
rect 421 391 437 401
rect 471 391 487 425
rect 25 349 357 365
rect 25 331 323 349
rect 25 125 59 331
rect 421 357 487 391
rect 421 323 437 357
rect 471 323 487 357
rect 531 351 565 487
rect 725 435 759 451
rect 601 390 617 424
rect 651 390 667 424
rect 725 367 759 401
rect 531 333 725 351
rect 531 317 759 333
rect 95 279 161 295
rect 129 245 161 279
rect 95 211 161 245
rect 129 177 161 211
rect 95 161 161 177
rect 209 279 257 295
rect 243 245 257 279
rect 209 211 257 245
rect 323 281 357 315
rect 323 231 357 247
rect 415 247 545 281
rect 579 247 595 281
rect 415 242 595 247
rect 243 177 257 211
rect 631 195 665 317
rect 209 161 257 177
rect 336 179 665 195
rect 336 145 340 179
rect 374 145 665 179
rect 336 129 665 145
rect 701 171 743 187
rect 701 137 705 171
rect 739 137 743 171
rect 25 109 100 125
rect 25 75 62 109
rect 96 75 100 109
rect 25 59 100 75
rect 144 101 186 117
rect 144 67 148 101
rect 182 67 186 101
rect 144 17 186 67
rect 230 103 272 119
rect 230 69 234 103
rect 268 87 272 103
rect 268 69 473 87
rect 230 53 473 69
rect 507 53 523 87
rect 701 17 743 137
rect 795 171 833 531
rect 829 137 833 171
rect 795 94 833 137
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 and4bb_m
flabel comment s 473 226 473 226 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5141462
string GDS_START 5133278
<< end >>
