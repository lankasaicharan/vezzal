magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 22 259 486 263
rect 22 49 1147 259
rect 0 0 1152 49
<< scnmos >>
rect 105 69 135 237
rect 191 69 221 237
rect 277 69 307 237
rect 363 69 393 237
rect 608 65 638 233
rect 694 65 724 233
rect 780 65 810 233
rect 866 65 896 233
rect 952 65 982 233
rect 1038 65 1068 233
<< scpmoshvt >>
rect 105 367 135 619
rect 191 367 221 619
rect 277 367 307 619
rect 363 367 393 619
rect 496 367 526 619
rect 582 367 612 619
rect 780 367 810 619
rect 866 367 896 619
rect 952 367 982 619
rect 1038 367 1068 619
<< ndiff >>
rect 48 225 105 237
rect 48 191 60 225
rect 94 191 105 225
rect 48 115 105 191
rect 48 81 60 115
rect 94 81 105 115
rect 48 69 105 81
rect 135 181 191 237
rect 135 147 146 181
rect 180 147 191 181
rect 135 111 191 147
rect 135 77 146 111
rect 180 77 191 111
rect 135 69 191 77
rect 221 225 277 237
rect 221 191 232 225
rect 266 191 277 225
rect 221 115 277 191
rect 221 81 232 115
rect 266 81 277 115
rect 221 69 277 81
rect 307 181 363 237
rect 307 147 318 181
rect 352 147 363 181
rect 307 111 363 147
rect 307 77 318 111
rect 352 77 363 111
rect 307 69 363 77
rect 393 225 460 237
rect 393 191 418 225
rect 452 191 460 225
rect 393 153 460 191
rect 393 119 418 153
rect 452 119 460 153
rect 393 69 460 119
rect 535 225 608 233
rect 535 191 549 225
rect 583 191 608 225
rect 535 153 608 191
rect 535 119 549 153
rect 583 119 608 153
rect 535 65 608 119
rect 638 179 694 233
rect 638 145 649 179
rect 683 145 694 179
rect 638 107 694 145
rect 638 73 649 107
rect 683 73 694 107
rect 638 65 694 73
rect 724 221 780 233
rect 724 187 735 221
rect 769 187 780 221
rect 724 111 780 187
rect 724 77 735 111
rect 769 77 780 111
rect 724 65 780 77
rect 810 183 866 233
rect 810 149 821 183
rect 855 149 866 183
rect 810 107 866 149
rect 810 73 821 107
rect 855 73 866 107
rect 810 65 866 73
rect 896 221 952 233
rect 896 187 907 221
rect 941 187 952 221
rect 896 111 952 187
rect 896 77 907 111
rect 941 77 952 111
rect 896 65 952 77
rect 982 183 1038 233
rect 982 149 993 183
rect 1027 149 1038 183
rect 982 107 1038 149
rect 982 73 993 107
rect 1027 73 1038 107
rect 982 65 1038 73
rect 1068 221 1121 233
rect 1068 187 1079 221
rect 1113 187 1121 221
rect 1068 111 1121 187
rect 1068 77 1079 111
rect 1113 77 1121 111
rect 1068 65 1121 77
<< pdiff >>
rect 52 607 105 619
rect 52 573 60 607
rect 94 573 105 607
rect 52 510 105 573
rect 52 476 60 510
rect 94 476 105 510
rect 52 418 105 476
rect 52 384 60 418
rect 94 384 105 418
rect 52 367 105 384
rect 135 599 191 619
rect 135 565 146 599
rect 180 565 191 599
rect 135 504 191 565
rect 135 470 146 504
rect 180 470 191 504
rect 135 413 191 470
rect 135 379 146 413
rect 180 379 191 413
rect 135 367 191 379
rect 221 607 277 619
rect 221 573 232 607
rect 266 573 277 607
rect 221 534 277 573
rect 221 500 232 534
rect 266 500 277 534
rect 221 453 277 500
rect 221 419 232 453
rect 266 419 277 453
rect 221 367 277 419
rect 307 599 363 619
rect 307 565 318 599
rect 352 565 363 599
rect 307 506 363 565
rect 307 472 318 506
rect 352 472 363 506
rect 307 413 363 472
rect 307 379 318 413
rect 352 379 363 413
rect 307 367 363 379
rect 393 569 496 619
rect 393 535 428 569
rect 462 535 496 569
rect 393 367 496 535
rect 526 599 582 619
rect 526 565 537 599
rect 571 565 582 599
rect 526 492 582 565
rect 526 458 537 492
rect 571 458 582 492
rect 526 367 582 458
rect 612 569 665 619
rect 612 535 623 569
rect 657 535 665 569
rect 612 367 665 535
rect 727 600 780 619
rect 727 566 735 600
rect 769 566 780 600
rect 727 367 780 566
rect 810 508 866 619
rect 810 474 821 508
rect 855 474 866 508
rect 810 367 866 474
rect 896 599 952 619
rect 896 565 907 599
rect 941 565 952 599
rect 896 508 952 565
rect 896 474 907 508
rect 941 474 952 508
rect 896 367 952 474
rect 982 531 1038 619
rect 982 497 993 531
rect 1027 497 1038 531
rect 982 440 1038 497
rect 982 406 993 440
rect 1027 406 1038 440
rect 982 367 1038 406
rect 1068 599 1121 619
rect 1068 565 1079 599
rect 1113 565 1121 599
rect 1068 516 1121 565
rect 1068 482 1079 516
rect 1113 482 1121 516
rect 1068 434 1121 482
rect 1068 400 1079 434
rect 1113 400 1121 434
rect 1068 367 1121 400
<< ndiffc >>
rect 60 191 94 225
rect 60 81 94 115
rect 146 147 180 181
rect 146 77 180 111
rect 232 191 266 225
rect 232 81 266 115
rect 318 147 352 181
rect 318 77 352 111
rect 418 191 452 225
rect 418 119 452 153
rect 549 191 583 225
rect 549 119 583 153
rect 649 145 683 179
rect 649 73 683 107
rect 735 187 769 221
rect 735 77 769 111
rect 821 149 855 183
rect 821 73 855 107
rect 907 187 941 221
rect 907 77 941 111
rect 993 149 1027 183
rect 993 73 1027 107
rect 1079 187 1113 221
rect 1079 77 1113 111
<< pdiffc >>
rect 60 573 94 607
rect 60 476 94 510
rect 60 384 94 418
rect 146 565 180 599
rect 146 470 180 504
rect 146 379 180 413
rect 232 573 266 607
rect 232 500 266 534
rect 232 419 266 453
rect 318 565 352 599
rect 318 472 352 506
rect 318 379 352 413
rect 428 535 462 569
rect 537 565 571 599
rect 537 458 571 492
rect 623 535 657 569
rect 735 566 769 600
rect 821 474 855 508
rect 907 565 941 599
rect 907 474 941 508
rect 993 497 1027 531
rect 993 406 1027 440
rect 1079 565 1113 599
rect 1079 482 1113 516
rect 1079 400 1113 434
<< poly >>
rect 105 619 135 645
rect 191 619 221 645
rect 277 619 307 645
rect 363 619 393 645
rect 496 619 526 645
rect 582 619 612 645
rect 780 619 810 645
rect 866 619 896 645
rect 952 619 982 645
rect 1038 619 1068 645
rect 105 335 135 367
rect 191 335 221 367
rect 44 319 221 335
rect 44 285 60 319
rect 94 317 221 319
rect 94 285 171 317
rect 44 283 171 285
rect 205 283 221 317
rect 44 269 221 283
rect 105 267 221 269
rect 105 237 135 267
rect 191 237 221 267
rect 277 335 307 367
rect 363 335 393 367
rect 496 335 526 367
rect 582 335 612 367
rect 780 335 810 367
rect 866 335 896 367
rect 277 319 454 335
rect 277 317 404 319
rect 277 283 293 317
rect 327 285 404 317
rect 438 285 454 319
rect 496 319 724 335
rect 496 305 674 319
rect 327 283 454 285
rect 277 269 454 283
rect 608 285 674 305
rect 708 285 724 319
rect 608 269 724 285
rect 277 267 393 269
rect 277 237 307 267
rect 363 237 393 267
rect 608 233 638 269
rect 694 233 724 269
rect 780 319 896 335
rect 780 285 796 319
rect 830 285 896 319
rect 780 269 896 285
rect 780 233 810 269
rect 866 233 896 269
rect 952 335 982 367
rect 1038 335 1068 367
rect 952 319 1068 335
rect 952 285 1018 319
rect 1052 285 1068 319
rect 952 269 1068 285
rect 952 233 982 269
rect 1038 233 1068 269
rect 105 43 135 69
rect 191 43 221 69
rect 277 43 307 69
rect 363 43 393 69
rect 608 39 638 65
rect 694 39 724 65
rect 780 39 810 65
rect 866 39 896 65
rect 952 39 982 65
rect 1038 39 1068 65
<< polycont >>
rect 60 285 94 319
rect 171 283 205 317
rect 293 283 327 317
rect 404 285 438 319
rect 674 285 708 319
rect 796 285 830 319
rect 1018 285 1052 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 44 607 110 649
rect 44 573 60 607
rect 94 573 110 607
rect 44 510 110 573
rect 44 476 60 510
rect 94 476 110 510
rect 44 418 110 476
rect 44 384 60 418
rect 94 384 110 418
rect 144 599 180 615
rect 144 565 146 599
rect 144 504 180 565
rect 144 470 146 504
rect 144 413 180 470
rect 216 607 282 649
rect 216 573 232 607
rect 266 573 282 607
rect 216 534 282 573
rect 216 500 232 534
rect 266 500 282 534
rect 216 453 282 500
rect 216 419 232 453
rect 266 419 282 453
rect 316 599 368 615
rect 316 565 318 599
rect 352 565 368 599
rect 316 506 368 565
rect 412 569 478 649
rect 412 535 428 569
rect 462 535 478 569
rect 412 526 478 535
rect 521 599 573 615
rect 521 565 537 599
rect 571 565 573 599
rect 316 472 318 506
rect 352 492 368 506
rect 521 492 573 565
rect 607 569 673 649
rect 607 535 623 569
rect 657 535 673 569
rect 719 600 1129 615
rect 719 566 735 600
rect 769 599 1129 600
rect 769 566 907 599
rect 719 565 907 566
rect 941 581 1079 599
rect 941 565 950 581
rect 719 560 950 565
rect 607 526 673 535
rect 805 508 864 526
rect 805 492 821 508
rect 352 472 537 492
rect 316 458 537 472
rect 571 474 821 492
rect 855 474 864 508
rect 571 458 864 474
rect 898 508 950 560
rect 1073 565 1079 581
rect 1113 565 1129 599
rect 898 474 907 508
rect 941 474 950 508
rect 898 458 950 474
rect 984 531 1039 547
rect 984 497 993 531
rect 1027 497 1039 531
rect 144 379 146 413
rect 316 413 354 458
rect 984 440 1039 497
rect 984 424 993 440
rect 316 385 318 413
rect 180 379 318 385
rect 352 379 354 413
rect 395 406 993 424
rect 1027 406 1039 440
rect 395 384 1039 406
rect 1073 516 1129 565
rect 1073 482 1079 516
rect 1113 482 1129 516
rect 1073 434 1129 482
rect 1073 400 1079 434
rect 1113 400 1129 434
rect 1073 384 1129 400
rect 144 351 354 379
rect 31 319 110 350
rect 31 285 60 319
rect 94 317 110 319
rect 388 319 547 350
rect 388 317 404 319
rect 94 285 171 317
rect 31 283 171 285
rect 205 283 221 317
rect 277 283 293 317
rect 327 285 404 317
rect 438 285 547 319
rect 327 283 547 285
rect 581 251 615 384
rect 658 319 737 350
rect 658 285 674 319
rect 708 285 737 319
rect 780 319 846 350
rect 780 285 796 319
rect 830 285 846 319
rect 880 319 1135 350
rect 880 285 1018 319
rect 1052 285 1135 319
rect 581 249 1133 251
rect 44 225 470 249
rect 44 191 60 225
rect 94 215 232 225
rect 94 191 96 215
rect 44 115 96 191
rect 230 191 232 215
rect 266 215 418 225
rect 266 191 268 215
rect 44 81 60 115
rect 94 81 96 115
rect 44 65 96 81
rect 130 147 146 181
rect 180 147 196 181
rect 130 111 196 147
rect 130 77 146 111
rect 180 77 196 111
rect 130 17 196 77
rect 230 115 268 191
rect 402 191 418 215
rect 452 191 470 225
rect 230 81 232 115
rect 266 81 268 115
rect 230 65 268 81
rect 302 147 318 181
rect 352 147 368 181
rect 302 111 368 147
rect 402 153 470 191
rect 402 119 418 153
rect 452 119 470 153
rect 531 225 1133 249
rect 531 191 549 225
rect 583 221 1133 225
rect 583 217 735 221
rect 583 191 599 217
rect 531 153 599 191
rect 733 187 735 217
rect 769 217 907 221
rect 769 187 771 217
rect 531 119 549 153
rect 583 119 599 153
rect 633 145 649 179
rect 683 145 699 179
rect 302 77 318 111
rect 352 85 368 111
rect 633 107 699 145
rect 633 85 649 107
rect 352 77 649 85
rect 302 73 649 77
rect 683 73 699 107
rect 302 51 699 73
rect 733 111 771 187
rect 905 187 907 217
rect 941 217 1079 221
rect 941 187 943 217
rect 733 77 735 111
rect 769 77 771 111
rect 733 61 771 77
rect 805 149 821 183
rect 855 149 871 183
rect 805 107 871 149
rect 805 73 821 107
rect 855 73 871 107
rect 805 17 871 73
rect 905 111 943 187
rect 1077 187 1079 217
rect 1113 187 1133 221
rect 905 77 907 111
rect 941 77 943 111
rect 905 61 943 77
rect 977 149 993 183
rect 1027 149 1043 183
rect 977 107 1043 149
rect 977 73 993 107
rect 1027 73 1043 107
rect 977 17 1043 73
rect 1077 111 1133 187
rect 1077 77 1079 111
rect 1113 77 1133 111
rect 1077 61 1133 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a311oi_2
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3237326
string GDS_START 3226858
<< end >>
