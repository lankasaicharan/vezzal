magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 23 49 902 243
rect 0 0 960 49
<< scnmos >>
rect 102 49 132 217
rect 188 49 218 217
rect 397 49 427 217
rect 483 49 513 217
rect 588 49 618 217
rect 685 49 715 217
rect 793 49 823 217
<< scpmoshvt >>
rect 86 367 116 619
rect 172 367 202 619
rect 397 367 427 619
rect 469 367 499 619
rect 577 367 607 619
rect 685 367 715 619
rect 793 367 823 619
<< ndiff >>
rect 49 205 102 217
rect 49 171 57 205
rect 91 171 102 205
rect 49 95 102 171
rect 49 61 57 95
rect 91 61 102 95
rect 49 49 102 61
rect 132 205 188 217
rect 132 171 143 205
rect 177 171 188 205
rect 132 101 188 171
rect 132 67 143 101
rect 177 67 188 101
rect 132 49 188 67
rect 218 167 397 217
rect 218 133 229 167
rect 263 133 352 167
rect 386 133 397 167
rect 218 91 397 133
rect 218 57 229 91
rect 263 57 352 91
rect 386 57 397 91
rect 218 49 397 57
rect 427 205 483 217
rect 427 171 438 205
rect 472 171 483 205
rect 427 101 483 171
rect 427 67 438 101
rect 472 67 483 101
rect 427 49 483 67
rect 513 159 588 217
rect 513 125 534 159
rect 568 125 588 159
rect 513 91 588 125
rect 513 57 534 91
rect 568 57 588 91
rect 513 49 588 57
rect 618 205 685 217
rect 618 171 629 205
rect 663 171 685 205
rect 618 101 685 171
rect 618 67 629 101
rect 663 67 685 101
rect 618 49 685 67
rect 715 49 793 217
rect 823 205 876 217
rect 823 171 834 205
rect 868 171 876 205
rect 823 95 876 171
rect 823 61 834 95
rect 868 61 876 95
rect 823 49 876 61
<< pdiff >>
rect 33 607 86 619
rect 33 573 41 607
rect 75 573 86 607
rect 33 503 86 573
rect 33 469 41 503
rect 75 469 86 503
rect 33 413 86 469
rect 33 379 41 413
rect 75 379 86 413
rect 33 367 86 379
rect 116 549 172 619
rect 116 515 127 549
rect 161 515 172 549
rect 116 481 172 515
rect 116 447 127 481
rect 161 447 172 481
rect 116 413 172 447
rect 116 379 127 413
rect 161 379 172 413
rect 116 367 172 379
rect 202 607 255 619
rect 202 573 213 607
rect 247 573 255 607
rect 202 495 255 573
rect 202 461 213 495
rect 247 461 255 495
rect 202 367 255 461
rect 344 607 397 619
rect 344 573 352 607
rect 386 573 397 607
rect 344 512 397 573
rect 344 478 352 512
rect 386 478 397 512
rect 344 418 397 478
rect 344 384 352 418
rect 386 384 397 418
rect 344 367 397 384
rect 427 367 469 619
rect 499 367 577 619
rect 607 607 685 619
rect 607 573 630 607
rect 664 573 685 607
rect 607 512 685 573
rect 607 478 630 512
rect 664 478 685 512
rect 607 420 685 478
rect 607 386 630 420
rect 664 386 685 420
rect 607 367 685 386
rect 715 607 793 619
rect 715 573 737 607
rect 771 573 793 607
rect 715 495 793 573
rect 715 461 737 495
rect 771 461 793 495
rect 715 367 793 461
rect 823 599 876 619
rect 823 565 834 599
rect 868 565 876 599
rect 823 510 876 565
rect 823 476 834 510
rect 868 476 876 510
rect 823 420 876 476
rect 823 386 834 420
rect 868 386 876 420
rect 823 367 876 386
<< ndiffc >>
rect 57 171 91 205
rect 57 61 91 95
rect 143 171 177 205
rect 143 67 177 101
rect 229 133 263 167
rect 352 133 386 167
rect 229 57 263 91
rect 352 57 386 91
rect 438 171 472 205
rect 438 67 472 101
rect 534 125 568 159
rect 534 57 568 91
rect 629 171 663 205
rect 629 67 663 101
rect 834 171 868 205
rect 834 61 868 95
<< pdiffc >>
rect 41 573 75 607
rect 41 469 75 503
rect 41 379 75 413
rect 127 515 161 549
rect 127 447 161 481
rect 127 379 161 413
rect 213 573 247 607
rect 213 461 247 495
rect 352 573 386 607
rect 352 478 386 512
rect 352 384 386 418
rect 630 573 664 607
rect 630 478 664 512
rect 630 386 664 420
rect 737 573 771 607
rect 737 461 771 495
rect 834 565 868 599
rect 834 476 868 510
rect 834 386 868 420
<< poly >>
rect 86 619 116 645
rect 172 619 202 645
rect 397 619 427 645
rect 469 619 499 645
rect 577 619 607 645
rect 685 619 715 645
rect 793 619 823 645
rect 86 305 116 367
rect 172 305 202 367
rect 397 335 427 367
rect 361 319 427 335
rect 86 289 283 305
rect 86 275 233 289
rect 102 255 233 275
rect 267 255 283 289
rect 361 285 377 319
rect 411 285 427 319
rect 361 269 427 285
rect 469 335 499 367
rect 577 335 607 367
rect 469 319 535 335
rect 469 285 485 319
rect 519 285 535 319
rect 469 269 535 285
rect 577 319 643 335
rect 577 285 593 319
rect 627 285 643 319
rect 577 269 643 285
rect 685 305 715 367
rect 793 308 823 367
rect 685 289 751 305
rect 102 239 283 255
rect 102 217 132 239
rect 188 217 218 239
rect 397 217 427 269
rect 483 217 513 269
rect 588 217 618 269
rect 685 255 701 289
rect 735 255 751 289
rect 685 239 751 255
rect 793 292 859 308
rect 793 258 809 292
rect 843 258 859 292
rect 793 242 859 258
rect 685 217 715 239
rect 793 217 823 242
rect 102 23 132 49
rect 188 23 218 49
rect 397 23 427 49
rect 483 23 513 49
rect 588 23 618 49
rect 685 23 715 49
rect 793 23 823 49
<< polycont >>
rect 233 255 267 289
rect 377 285 411 319
rect 485 285 519 319
rect 593 285 627 319
rect 701 255 735 289
rect 809 258 843 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 25 607 91 649
rect 25 573 41 607
rect 75 573 91 607
rect 197 607 263 649
rect 25 503 91 573
rect 25 469 41 503
rect 75 469 91 503
rect 25 413 91 469
rect 25 379 41 413
rect 75 379 91 413
rect 25 363 91 379
rect 125 549 163 600
rect 125 515 127 549
rect 161 515 163 549
rect 125 481 163 515
rect 125 447 127 481
rect 161 447 163 481
rect 197 573 213 607
rect 247 573 263 607
rect 197 495 263 573
rect 197 461 213 495
rect 247 461 263 495
rect 197 454 263 461
rect 336 607 402 615
rect 336 573 352 607
rect 386 573 402 607
rect 614 607 680 615
rect 336 512 402 573
rect 336 478 352 512
rect 386 478 402 512
rect 125 420 163 447
rect 336 420 402 478
rect 125 413 179 420
rect 125 379 127 413
rect 161 379 179 413
rect 41 205 91 221
rect 41 171 57 205
rect 41 95 91 171
rect 41 61 57 95
rect 41 17 91 61
rect 125 205 179 379
rect 125 171 143 205
rect 177 171 179 205
rect 213 418 402 420
rect 213 384 352 418
rect 386 384 402 418
rect 213 289 283 384
rect 213 255 233 289
rect 267 255 283 289
rect 317 319 451 350
rect 317 285 377 319
rect 411 285 451 319
rect 317 269 451 285
rect 485 319 559 593
rect 614 573 630 607
rect 664 573 680 607
rect 614 512 680 573
rect 614 478 630 512
rect 664 478 680 512
rect 614 420 680 478
rect 721 607 787 649
rect 721 573 737 607
rect 771 573 787 607
rect 721 495 787 573
rect 721 461 737 495
rect 771 461 787 495
rect 721 454 787 461
rect 821 599 884 615
rect 821 565 834 599
rect 868 565 884 599
rect 821 510 884 565
rect 821 476 834 510
rect 868 476 884 510
rect 821 420 884 476
rect 614 386 630 420
rect 664 386 834 420
rect 868 386 884 420
rect 519 285 559 319
rect 485 269 559 285
rect 593 319 662 350
rect 627 285 662 319
rect 593 269 662 285
rect 701 289 755 350
rect 213 235 283 255
rect 735 255 755 289
rect 213 205 667 235
rect 213 201 438 205
rect 125 101 179 171
rect 436 171 438 201
rect 472 201 629 205
rect 472 171 484 201
rect 125 67 143 101
rect 177 67 179 101
rect 125 51 179 67
rect 213 133 229 167
rect 263 133 352 167
rect 386 133 402 167
rect 213 91 402 133
rect 213 57 229 91
rect 263 57 352 91
rect 386 57 402 91
rect 213 17 402 57
rect 436 101 484 171
rect 618 171 629 201
rect 663 171 667 205
rect 436 67 438 101
rect 472 67 484 101
rect 436 51 484 67
rect 518 159 584 163
rect 518 125 534 159
rect 568 125 584 159
rect 518 91 584 125
rect 518 57 534 91
rect 568 57 584 91
rect 518 17 584 57
rect 618 101 667 171
rect 618 67 629 101
rect 663 67 667 101
rect 618 51 667 67
rect 701 60 755 255
rect 789 292 943 350
rect 789 258 809 292
rect 843 258 943 292
rect 789 242 943 258
rect 818 205 884 208
rect 818 171 834 205
rect 868 171 884 205
rect 818 95 884 171
rect 818 61 834 95
rect 868 61 884 95
rect 818 17 884 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2111o_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1105266
string GDS_START 1095408
<< end >>
