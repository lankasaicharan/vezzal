magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1778 1975
<< nwell >>
rect -38 331 518 704
<< pwell >>
rect 20 49 433 164
rect 0 0 480 49
<< scnmos >>
rect 99 54 129 138
rect 252 54 282 138
rect 324 54 354 138
<< scpmoshvt >>
rect 144 532 174 616
rect 230 532 260 616
rect 316 532 346 616
<< ndiff >>
rect 46 126 99 138
rect 46 92 54 126
rect 88 92 99 126
rect 46 54 99 92
rect 129 100 252 138
rect 129 66 201 100
rect 235 66 252 100
rect 129 54 252 66
rect 282 54 324 138
rect 354 126 407 138
rect 354 92 365 126
rect 399 92 407 126
rect 354 54 407 92
<< pdiff >>
rect 91 578 144 616
rect 91 544 99 578
rect 133 544 144 578
rect 91 532 144 544
rect 174 604 230 616
rect 174 570 185 604
rect 219 570 230 604
rect 174 532 230 570
rect 260 578 316 616
rect 260 544 271 578
rect 305 544 316 578
rect 260 532 316 544
rect 346 604 399 616
rect 346 570 357 604
rect 391 570 399 604
rect 346 532 399 570
<< ndiffc >>
rect 54 92 88 126
rect 201 66 235 100
rect 365 92 399 126
<< pdiffc >>
rect 99 544 133 578
rect 185 570 219 604
rect 271 544 305 578
rect 357 570 391 604
<< poly >>
rect 144 616 174 642
rect 230 616 260 642
rect 316 616 346 642
rect 144 342 174 532
rect 99 326 174 342
rect 99 292 124 326
rect 158 292 174 326
rect 230 294 260 532
rect 316 476 346 532
rect 308 460 374 476
rect 308 426 324 460
rect 358 426 374 460
rect 308 392 374 426
rect 308 358 324 392
rect 358 358 374 392
rect 308 342 374 358
rect 99 258 174 292
rect 99 224 124 258
rect 158 224 174 258
rect 99 208 174 224
rect 216 278 282 294
rect 216 244 232 278
rect 266 244 282 278
rect 216 210 282 244
rect 99 138 129 208
rect 216 176 232 210
rect 266 176 282 210
rect 330 190 360 342
rect 216 160 282 176
rect 252 138 282 160
rect 324 160 360 190
rect 324 138 354 160
rect 99 28 129 54
rect 252 28 282 54
rect 324 28 354 54
<< polycont >>
rect 124 292 158 326
rect 324 426 358 460
rect 324 358 358 392
rect 124 224 158 258
rect 232 244 266 278
rect 232 176 266 210
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 181 604 223 649
rect 95 578 137 594
rect 95 544 99 578
rect 133 544 137 578
rect 181 570 185 604
rect 219 570 223 604
rect 341 604 407 649
rect 181 554 223 570
rect 267 578 305 594
rect 95 494 137 544
rect 267 544 271 578
rect 341 570 357 604
rect 391 570 407 604
rect 341 566 407 570
rect 267 530 305 544
rect 267 496 449 530
rect 50 460 231 494
rect 50 126 88 460
rect 197 426 324 460
rect 358 426 374 460
rect 50 92 54 126
rect 124 326 161 424
rect 308 392 374 426
rect 308 358 324 392
rect 358 358 374 392
rect 158 292 161 326
rect 124 258 161 292
rect 158 224 161 258
rect 124 94 161 224
rect 223 278 266 294
rect 223 244 232 278
rect 223 210 266 244
rect 223 176 232 210
rect 223 160 266 176
rect 415 130 449 496
rect 349 126 449 130
rect 197 100 239 116
rect 50 76 88 92
rect 197 66 201 100
rect 235 66 239 100
rect 349 92 365 126
rect 399 92 449 126
rect 349 88 449 92
rect 197 17 239 66
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
<< metal1 >>
rect 0 683 480 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 480 683
rect 0 617 480 649
rect 0 17 480 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 480 17
rect 0 -49 480 -17
<< labels >>
flabel pwell s 0 0 480 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 480 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2b_m
flabel metal1 s 0 617 480 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 480 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 480 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4471178
string GDS_START 4465596
<< end >>
