magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 4 228 465 248
rect 4 49 1150 228
rect 0 0 1152 49
<< scnmos >>
rect 87 74 117 222
rect 173 74 203 222
rect 273 74 303 222
rect 359 74 389 222
rect 459 74 489 202
rect 545 74 575 202
rect 743 74 773 202
rect 837 74 867 202
rect 923 74 953 202
rect 1027 74 1057 202
<< scpmoshvt >>
rect 86 368 116 592
rect 176 368 206 592
rect 286 368 316 592
rect 376 368 406 592
rect 486 424 516 592
rect 576 424 606 592
rect 736 424 766 592
rect 834 424 864 592
rect 936 424 966 592
rect 1026 424 1056 592
<< ndiff >>
rect 30 210 87 222
rect 30 176 42 210
rect 76 176 87 210
rect 30 120 87 176
rect 30 86 42 120
rect 76 86 87 120
rect 30 74 87 86
rect 117 210 173 222
rect 117 176 128 210
rect 162 176 173 210
rect 117 120 173 176
rect 117 86 128 120
rect 162 86 173 120
rect 117 74 173 86
rect 203 142 273 222
rect 203 108 214 142
rect 248 108 273 142
rect 203 74 273 108
rect 303 210 359 222
rect 303 176 314 210
rect 348 176 359 210
rect 303 120 359 176
rect 303 86 314 120
rect 348 86 359 120
rect 303 74 359 86
rect 389 202 439 222
rect 389 190 459 202
rect 389 156 400 190
rect 434 156 459 190
rect 389 120 459 156
rect 389 86 400 120
rect 434 86 459 120
rect 389 74 459 86
rect 489 190 545 202
rect 489 156 500 190
rect 534 156 545 190
rect 489 120 545 156
rect 489 86 500 120
rect 534 86 545 120
rect 489 74 545 86
rect 575 147 632 202
rect 575 113 586 147
rect 620 113 632 147
rect 575 74 632 113
rect 686 147 743 202
rect 686 113 698 147
rect 732 113 743 147
rect 686 74 743 113
rect 773 179 837 202
rect 773 145 784 179
rect 818 145 837 179
rect 773 74 837 145
rect 867 190 923 202
rect 867 156 878 190
rect 912 156 923 190
rect 867 120 923 156
rect 867 86 878 120
rect 912 86 923 120
rect 867 74 923 86
rect 953 169 1027 202
rect 953 135 978 169
rect 1012 135 1027 169
rect 953 74 1027 135
rect 1057 188 1124 202
rect 1057 154 1078 188
rect 1112 154 1124 188
rect 1057 120 1124 154
rect 1057 86 1078 120
rect 1112 86 1124 120
rect 1057 74 1124 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 497 86 546
rect 27 463 39 497
rect 73 463 86 497
rect 27 414 86 463
rect 27 380 39 414
rect 73 380 86 414
rect 27 368 86 380
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 497 176 546
rect 116 463 129 497
rect 163 463 176 497
rect 116 414 176 463
rect 116 380 129 414
rect 163 380 176 414
rect 116 368 176 380
rect 206 580 286 592
rect 206 546 229 580
rect 263 546 286 580
rect 206 478 286 546
rect 206 444 229 478
rect 263 444 286 478
rect 206 368 286 444
rect 316 580 376 592
rect 316 546 329 580
rect 363 546 376 580
rect 316 497 376 546
rect 316 463 329 497
rect 363 463 376 497
rect 316 414 376 463
rect 316 380 329 414
rect 363 380 376 414
rect 316 368 376 380
rect 406 580 486 592
rect 406 546 429 580
rect 463 546 486 580
rect 406 508 486 546
rect 406 474 429 508
rect 463 474 486 508
rect 406 424 486 474
rect 516 580 576 592
rect 516 546 529 580
rect 563 546 576 580
rect 516 470 576 546
rect 516 436 529 470
rect 563 436 576 470
rect 516 424 576 436
rect 606 580 736 592
rect 606 546 620 580
rect 654 546 688 580
rect 722 546 736 580
rect 606 508 736 546
rect 606 474 620 508
rect 654 474 688 508
rect 722 474 736 508
rect 606 424 736 474
rect 766 580 834 592
rect 766 546 779 580
rect 813 546 834 580
rect 766 470 834 546
rect 766 436 779 470
rect 813 436 834 470
rect 766 424 834 436
rect 864 580 936 592
rect 864 546 879 580
rect 913 546 936 580
rect 864 508 936 546
rect 864 474 879 508
rect 913 474 936 508
rect 864 424 936 474
rect 966 580 1026 592
rect 966 546 979 580
rect 1013 546 1026 580
rect 966 470 1026 546
rect 966 436 979 470
rect 1013 436 1026 470
rect 966 424 1026 436
rect 1056 580 1125 592
rect 1056 546 1079 580
rect 1113 546 1125 580
rect 1056 508 1125 546
rect 1056 474 1079 508
rect 1113 474 1125 508
rect 1056 424 1125 474
rect 406 368 459 424
<< ndiffc >>
rect 42 176 76 210
rect 42 86 76 120
rect 128 176 162 210
rect 128 86 162 120
rect 214 108 248 142
rect 314 176 348 210
rect 314 86 348 120
rect 400 156 434 190
rect 400 86 434 120
rect 500 156 534 190
rect 500 86 534 120
rect 586 113 620 147
rect 698 113 732 147
rect 784 145 818 179
rect 878 156 912 190
rect 878 86 912 120
rect 978 135 1012 169
rect 1078 154 1112 188
rect 1078 86 1112 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 129 546 163 580
rect 129 463 163 497
rect 129 380 163 414
rect 229 546 263 580
rect 229 444 263 478
rect 329 546 363 580
rect 329 463 363 497
rect 329 380 363 414
rect 429 546 463 580
rect 429 474 463 508
rect 529 546 563 580
rect 529 436 563 470
rect 620 546 654 580
rect 688 546 722 580
rect 620 474 654 508
rect 688 474 722 508
rect 779 546 813 580
rect 779 436 813 470
rect 879 546 913 580
rect 879 474 913 508
rect 979 546 1013 580
rect 979 436 1013 470
rect 1079 546 1113 580
rect 1079 474 1113 508
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 286 592 316 618
rect 376 592 406 618
rect 486 592 516 618
rect 576 592 606 618
rect 736 592 766 618
rect 834 592 864 618
rect 936 592 966 618
rect 1026 592 1056 618
rect 486 409 516 424
rect 576 409 606 424
rect 736 409 766 424
rect 834 409 864 424
rect 936 409 966 424
rect 1026 409 1056 424
rect 86 353 116 368
rect 176 353 206 368
rect 286 353 316 368
rect 376 353 406 368
rect 483 356 519 409
rect 573 356 609 409
rect 83 326 119 353
rect 173 326 209 353
rect 283 326 319 353
rect 373 326 409 353
rect 83 310 409 326
rect 483 340 639 356
rect 483 320 521 340
rect 83 276 223 310
rect 257 276 291 310
rect 325 276 359 310
rect 393 276 409 310
rect 83 260 409 276
rect 459 306 521 320
rect 555 306 589 340
rect 623 306 639 340
rect 459 290 639 306
rect 733 331 769 409
rect 831 331 867 409
rect 933 379 1059 409
rect 933 356 1057 379
rect 733 315 867 331
rect 87 222 117 260
rect 173 222 203 260
rect 273 222 303 260
rect 359 222 389 260
rect 459 202 489 290
rect 545 202 575 290
rect 733 281 749 315
rect 783 281 817 315
rect 851 281 867 315
rect 733 265 867 281
rect 743 202 773 265
rect 837 202 867 265
rect 923 340 1057 356
rect 923 306 939 340
rect 973 306 1007 340
rect 1041 306 1057 340
rect 923 290 1057 306
rect 923 202 953 290
rect 1027 202 1057 290
rect 87 48 117 74
rect 173 48 203 74
rect 273 48 303 74
rect 359 48 389 74
rect 459 48 489 74
rect 545 48 575 74
rect 743 48 773 74
rect 837 48 867 74
rect 923 48 953 74
rect 1027 48 1057 74
<< polycont >>
rect 223 276 257 310
rect 291 276 325 310
rect 359 276 393 310
rect 521 306 555 340
rect 589 306 623 340
rect 749 281 783 315
rect 817 281 851 315
rect 939 306 973 340
rect 1007 306 1041 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 580 73 649
rect 23 546 39 580
rect 23 497 73 546
rect 23 463 39 497
rect 23 414 73 463
rect 23 380 39 414
rect 23 364 73 380
rect 112 580 179 596
rect 112 546 129 580
rect 163 546 179 580
rect 112 497 179 546
rect 112 463 129 497
rect 163 463 179 497
rect 112 414 179 463
rect 213 580 279 649
rect 213 546 229 580
rect 263 546 279 580
rect 213 478 279 546
rect 213 444 229 478
rect 263 444 279 478
rect 213 428 279 444
rect 313 580 379 596
rect 313 546 329 580
rect 363 546 379 580
rect 313 497 379 546
rect 313 463 329 497
rect 363 463 379 497
rect 112 380 129 414
rect 163 394 179 414
rect 313 414 379 463
rect 413 580 479 649
rect 413 546 429 580
rect 463 546 479 580
rect 413 508 479 546
rect 413 474 429 508
rect 463 474 479 508
rect 413 458 479 474
rect 513 580 579 596
rect 513 546 529 580
rect 563 546 579 580
rect 513 470 579 546
rect 513 436 529 470
rect 563 436 579 470
rect 613 580 729 649
rect 613 546 620 580
rect 654 546 688 580
rect 722 546 729 580
rect 613 508 729 546
rect 613 474 620 508
rect 654 474 688 508
rect 722 474 729 508
rect 613 458 729 474
rect 763 580 829 596
rect 763 546 779 580
rect 813 546 829 580
rect 763 470 829 546
rect 513 424 579 436
rect 763 436 779 470
rect 813 436 829 470
rect 863 580 929 649
rect 863 546 879 580
rect 913 546 929 580
rect 863 508 929 546
rect 863 474 879 508
rect 913 474 929 508
rect 863 458 929 474
rect 963 580 1029 596
rect 963 546 979 580
rect 1013 546 1029 580
rect 963 470 1029 546
rect 763 424 829 436
rect 963 436 979 470
rect 1013 436 1029 470
rect 1063 580 1129 649
rect 1063 546 1079 580
rect 1113 546 1129 580
rect 1063 508 1129 546
rect 1063 474 1079 508
rect 1113 474 1129 508
rect 1063 458 1129 474
rect 963 424 1029 436
rect 313 394 329 414
rect 163 380 329 394
rect 363 380 379 414
rect 112 360 379 380
rect 413 390 1125 424
rect 112 226 167 360
rect 413 326 447 390
rect 207 310 447 326
rect 207 276 223 310
rect 257 276 291 310
rect 325 276 359 310
rect 393 276 447 310
rect 505 340 646 356
rect 505 306 521 340
rect 555 306 589 340
rect 623 306 646 340
rect 505 290 646 306
rect 697 315 867 356
rect 207 260 447 276
rect 697 281 749 315
rect 783 281 817 315
rect 851 281 867 315
rect 923 340 1057 356
rect 923 306 939 340
rect 973 306 1007 340
rect 1041 306 1057 340
rect 923 290 1057 306
rect 697 265 867 281
rect 1091 256 1125 390
rect 26 210 76 226
rect 26 176 42 210
rect 26 120 76 176
rect 26 86 42 120
rect 26 17 76 86
rect 112 210 348 226
rect 112 176 128 210
rect 162 192 314 210
rect 162 176 178 192
rect 112 120 178 176
rect 298 176 314 192
rect 112 86 128 120
rect 162 86 178 120
rect 112 70 178 86
rect 214 142 264 158
rect 248 108 264 142
rect 214 17 264 108
rect 298 120 348 176
rect 298 86 314 120
rect 298 70 348 86
rect 384 190 450 206
rect 384 156 400 190
rect 434 156 450 190
rect 384 120 450 156
rect 384 86 400 120
rect 434 86 450 120
rect 384 17 450 86
rect 484 197 818 231
rect 962 222 1125 256
rect 484 190 534 197
rect 484 156 500 190
rect 784 179 818 197
rect 484 120 534 156
rect 484 86 500 120
rect 484 70 534 86
rect 570 147 636 163
rect 570 113 586 147
rect 620 113 636 147
rect 570 17 636 113
rect 682 147 748 163
rect 682 113 698 147
rect 732 113 748 147
rect 784 119 818 145
rect 862 190 928 206
rect 862 156 878 190
rect 912 156 928 190
rect 862 120 928 156
rect 682 85 748 113
rect 862 86 878 120
rect 912 86 928 120
rect 962 169 1028 222
rect 962 135 978 169
rect 1012 135 1028 169
rect 962 119 1028 135
rect 1062 154 1078 188
rect 1112 154 1128 188
rect 1062 120 1128 154
rect 862 85 928 86
rect 1062 86 1078 120
rect 1112 86 1128 120
rect 1062 85 1128 86
rect 682 51 1128 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and3_4
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 2974598
string GDS_START 2964178
<< end >>
