magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3122 1975
<< nwell >>
rect -38 331 1862 704
<< pwell >>
rect 5 229 513 241
rect 1269 229 1823 247
rect 5 49 1823 229
rect 0 0 1824 49
<< scnmos >>
rect 84 47 114 215
rect 170 47 200 215
rect 279 131 309 215
rect 404 131 434 215
rect 594 119 624 203
rect 680 119 710 203
rect 752 119 782 203
rect 824 119 854 203
rect 910 119 940 203
rect 996 119 1026 203
rect 1157 119 1187 203
rect 1243 119 1273 203
rect 1368 53 1398 221
rect 1454 53 1484 221
rect 1623 137 1653 221
rect 1695 137 1725 221
<< scpmoshvt >>
rect 84 367 114 619
rect 170 367 200 619
rect 279 398 309 526
rect 365 398 395 526
rect 578 419 608 547
rect 680 419 710 547
rect 752 419 782 547
rect 824 419 854 547
rect 911 419 941 547
rect 1043 444 1073 572
rect 1137 444 1167 572
rect 1223 444 1253 572
rect 1382 367 1412 619
rect 1468 367 1498 619
rect 1623 367 1653 495
rect 1695 367 1725 495
<< ndiff >>
rect 31 95 84 215
rect 31 61 39 95
rect 73 61 84 95
rect 31 47 84 61
rect 114 175 170 215
rect 114 141 125 175
rect 159 141 170 175
rect 114 93 170 141
rect 114 59 125 93
rect 159 59 170 93
rect 114 47 170 59
rect 200 131 279 215
rect 309 140 404 215
rect 309 131 343 140
rect 200 126 257 131
rect 200 92 215 126
rect 249 92 257 126
rect 200 47 257 92
rect 331 106 343 131
rect 377 131 404 140
rect 434 192 487 215
rect 1295 203 1368 221
rect 434 158 445 192
rect 479 158 487 192
rect 434 131 487 158
rect 541 178 594 203
rect 541 144 549 178
rect 583 144 594 178
rect 377 106 389 131
rect 331 98 389 106
rect 541 119 594 144
rect 624 167 680 203
rect 624 133 635 167
rect 669 133 680 167
rect 624 119 680 133
rect 710 119 752 203
rect 782 119 824 203
rect 854 178 910 203
rect 854 144 865 178
rect 899 144 910 178
rect 854 119 910 144
rect 940 178 996 203
rect 940 144 951 178
rect 985 144 996 178
rect 940 119 996 144
rect 1026 165 1157 203
rect 1026 131 1037 165
rect 1071 131 1112 165
rect 1146 131 1157 165
rect 1026 119 1157 131
rect 1187 191 1243 203
rect 1187 157 1198 191
rect 1232 157 1243 191
rect 1187 119 1243 157
rect 1273 119 1368 203
rect 1295 69 1368 119
rect 1295 35 1307 69
rect 1341 53 1368 69
rect 1398 211 1454 221
rect 1398 177 1409 211
rect 1443 177 1454 211
rect 1398 53 1454 177
rect 1484 137 1623 221
rect 1653 137 1695 221
rect 1725 209 1797 221
rect 1725 175 1755 209
rect 1789 175 1797 209
rect 1725 137 1797 175
rect 1484 69 1557 137
rect 1484 53 1511 69
rect 1341 35 1353 53
rect 1295 27 1353 35
rect 1499 35 1511 53
rect 1545 35 1557 69
rect 1499 27 1557 35
<< pdiff >>
rect 31 582 84 619
rect 31 548 39 582
rect 73 548 84 582
rect 31 367 84 548
rect 114 599 170 619
rect 114 565 125 599
rect 159 565 170 599
rect 114 514 170 565
rect 114 480 125 514
rect 159 480 170 514
rect 114 367 170 480
rect 200 607 253 619
rect 200 573 211 607
rect 245 573 253 607
rect 200 526 253 573
rect 200 502 279 526
rect 200 468 220 502
rect 254 468 279 502
rect 200 398 279 468
rect 309 502 365 526
rect 309 468 320 502
rect 354 468 365 502
rect 309 398 365 468
rect 395 512 452 526
rect 395 478 406 512
rect 440 478 452 512
rect 395 444 452 478
rect 395 410 406 444
rect 440 410 452 444
rect 395 398 452 410
rect 200 367 253 398
rect 1275 583 1382 619
rect 1275 572 1337 583
rect 963 562 1043 572
rect 963 547 975 562
rect 525 535 578 547
rect 525 501 533 535
rect 567 501 578 535
rect 525 467 578 501
rect 525 433 533 467
rect 567 433 578 467
rect 525 419 578 433
rect 608 535 680 547
rect 608 501 635 535
rect 669 501 680 535
rect 608 467 680 501
rect 608 433 635 467
rect 669 433 680 467
rect 608 419 680 433
rect 710 419 752 547
rect 782 419 824 547
rect 854 533 911 547
rect 854 499 865 533
rect 899 499 911 533
rect 854 465 911 499
rect 854 431 865 465
rect 899 431 911 465
rect 854 419 911 431
rect 941 528 975 547
rect 1009 528 1043 562
rect 941 492 1043 528
rect 941 458 975 492
rect 1009 458 1043 492
rect 941 444 1043 458
rect 1073 564 1137 572
rect 1073 530 1087 564
rect 1121 530 1137 564
rect 1073 444 1137 530
rect 1167 558 1223 572
rect 1167 524 1178 558
rect 1212 524 1223 558
rect 1167 490 1223 524
rect 1167 456 1178 490
rect 1212 456 1223 490
rect 1167 444 1223 456
rect 1253 560 1337 572
rect 1253 526 1264 560
rect 1298 549 1337 560
rect 1371 549 1382 583
rect 1298 526 1382 549
rect 1253 488 1382 526
rect 1253 454 1264 488
rect 1298 454 1382 488
rect 1253 444 1382 454
rect 941 419 1021 444
rect 1275 419 1382 444
rect 1332 367 1382 419
rect 1412 413 1468 619
rect 1412 379 1423 413
rect 1457 379 1468 413
rect 1412 367 1468 379
rect 1498 575 1551 619
rect 1498 541 1509 575
rect 1543 541 1551 575
rect 1498 495 1551 541
rect 1498 367 1623 495
rect 1653 367 1695 495
rect 1725 483 1782 495
rect 1725 449 1740 483
rect 1774 449 1782 483
rect 1725 415 1782 449
rect 1725 381 1740 415
rect 1774 381 1782 415
rect 1725 367 1782 381
<< ndiffc >>
rect 39 61 73 95
rect 125 141 159 175
rect 125 59 159 93
rect 215 92 249 126
rect 343 106 377 140
rect 445 158 479 192
rect 549 144 583 178
rect 635 133 669 167
rect 865 144 899 178
rect 951 144 985 178
rect 1037 131 1071 165
rect 1112 131 1146 165
rect 1198 157 1232 191
rect 1307 35 1341 69
rect 1409 177 1443 211
rect 1755 175 1789 209
rect 1511 35 1545 69
<< pdiffc >>
rect 39 548 73 582
rect 125 565 159 599
rect 125 480 159 514
rect 211 573 245 607
rect 220 468 254 502
rect 320 468 354 502
rect 406 478 440 512
rect 406 410 440 444
rect 533 501 567 535
rect 533 433 567 467
rect 635 501 669 535
rect 635 433 669 467
rect 865 499 899 533
rect 865 431 899 465
rect 975 528 1009 562
rect 975 458 1009 492
rect 1087 530 1121 564
rect 1178 524 1212 558
rect 1178 456 1212 490
rect 1264 526 1298 560
rect 1337 549 1371 583
rect 1264 454 1298 488
rect 1423 379 1457 413
rect 1509 541 1543 575
rect 1740 449 1774 483
rect 1740 381 1774 415
<< poly >>
rect 84 619 114 645
rect 170 619 200 645
rect 467 615 1073 645
rect 1382 619 1412 645
rect 1468 619 1498 645
rect 279 526 309 552
rect 365 526 395 552
rect 84 299 114 367
rect 170 335 200 367
rect 170 319 237 335
rect 170 299 187 319
rect 84 285 187 299
rect 221 285 237 319
rect 84 269 237 285
rect 84 215 114 269
rect 170 215 200 269
rect 279 215 309 398
rect 365 366 395 398
rect 467 366 497 615
rect 578 547 608 573
rect 680 547 710 573
rect 752 547 782 573
rect 824 547 854 615
rect 911 547 941 573
rect 1043 572 1073 615
rect 1137 572 1167 598
rect 1223 572 1253 598
rect 365 350 497 366
rect 365 316 431 350
rect 465 316 497 350
rect 365 300 497 316
rect 578 337 608 419
rect 680 337 710 419
rect 578 321 710 337
rect 404 215 434 300
rect 578 287 660 321
rect 694 287 710 321
rect 578 271 710 287
rect 279 51 309 131
rect 594 203 624 271
rect 680 203 710 271
rect 752 203 782 419
rect 824 203 854 419
rect 911 387 941 419
rect 910 371 1001 387
rect 910 337 951 371
rect 985 337 1001 371
rect 910 321 1001 337
rect 910 203 940 321
rect 1043 273 1073 444
rect 1137 333 1167 444
rect 1223 387 1253 444
rect 1223 371 1289 387
rect 1223 337 1239 371
rect 1273 337 1289 371
rect 1623 495 1653 521
rect 1695 495 1725 521
rect 996 243 1073 273
rect 1115 317 1181 333
rect 1223 321 1289 337
rect 1115 283 1131 317
rect 1165 283 1181 317
rect 1115 267 1181 283
rect 1151 255 1181 267
rect 996 203 1026 243
rect 1151 225 1187 255
rect 1157 203 1187 225
rect 1243 203 1273 321
rect 1382 273 1412 367
rect 1468 309 1498 367
rect 1623 335 1653 367
rect 1587 319 1653 335
rect 1454 293 1545 309
rect 1454 273 1495 293
rect 1368 259 1495 273
rect 1529 259 1545 293
rect 1587 285 1603 319
rect 1637 285 1653 319
rect 1587 269 1653 285
rect 1368 243 1545 259
rect 1368 221 1398 243
rect 1454 221 1484 243
rect 1623 221 1653 269
rect 1695 273 1725 367
rect 1695 243 1731 273
rect 1695 221 1725 243
rect 404 105 434 131
rect 594 93 624 119
rect 680 93 710 119
rect 752 51 782 119
rect 824 93 854 119
rect 910 93 940 119
rect 996 93 1026 119
rect 1157 51 1187 119
rect 1243 93 1273 119
rect 84 21 114 47
rect 170 21 200 47
rect 279 21 1187 51
rect 1623 111 1653 137
rect 1695 115 1725 137
rect 1368 27 1398 53
rect 1454 27 1484 53
rect 1695 99 1766 115
rect 1695 65 1716 99
rect 1750 65 1766 99
rect 1695 49 1766 65
<< polycont >>
rect 187 285 221 319
rect 431 316 465 350
rect 660 287 694 321
rect 951 337 985 371
rect 1239 337 1273 371
rect 1131 283 1165 317
rect 1495 259 1529 293
rect 1603 285 1637 319
rect 1716 65 1750 99
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 23 582 89 649
rect 23 548 39 582
rect 73 548 89 582
rect 23 532 89 548
rect 123 599 161 615
rect 123 565 125 599
rect 159 565 161 599
rect 123 514 161 565
rect 123 498 125 514
rect 17 480 125 498
rect 159 480 161 514
rect 17 464 161 480
rect 195 607 270 649
rect 195 573 211 607
rect 245 573 270 607
rect 195 502 270 573
rect 195 468 220 502
rect 254 468 270 502
rect 195 464 270 468
rect 304 564 583 598
rect 304 502 370 564
rect 517 535 583 564
rect 304 468 320 502
rect 354 468 370 502
rect 304 464 370 468
rect 404 512 456 528
rect 404 478 406 512
rect 440 478 456 512
rect 17 181 67 464
rect 404 444 456 478
rect 404 430 406 444
rect 101 424 406 430
rect 101 390 127 424
rect 161 410 406 424
rect 440 410 456 444
rect 517 501 533 535
rect 567 501 583 535
rect 517 467 583 501
rect 517 433 533 467
rect 567 433 583 467
rect 517 429 583 433
rect 619 535 685 649
rect 959 562 1025 578
rect 619 501 635 535
rect 669 501 685 535
rect 619 467 685 501
rect 619 433 635 467
rect 669 433 685 467
rect 849 533 901 549
rect 849 499 865 533
rect 899 499 901 533
rect 849 465 901 499
rect 849 449 865 465
rect 619 429 685 433
rect 721 431 865 449
rect 899 431 901 465
rect 959 528 975 562
rect 1009 528 1025 562
rect 1071 564 1137 649
rect 1248 583 1387 649
rect 1071 530 1087 564
rect 1121 530 1137 564
rect 1071 528 1137 530
rect 1171 558 1214 574
rect 959 494 1025 528
rect 1171 524 1178 558
rect 1212 524 1214 558
rect 1171 494 1214 524
rect 959 492 1214 494
rect 959 458 975 492
rect 1009 490 1214 492
rect 1009 458 1178 490
rect 1162 456 1178 458
rect 1212 456 1214 490
rect 1162 440 1214 456
rect 1248 560 1337 583
rect 1248 526 1264 560
rect 1298 549 1337 560
rect 1371 549 1387 583
rect 1298 533 1387 549
rect 1493 575 1559 649
rect 1493 541 1509 575
rect 1543 541 1559 575
rect 1493 533 1559 541
rect 1298 526 1314 533
rect 1248 488 1314 526
rect 1248 454 1264 488
rect 1298 454 1314 488
rect 1353 465 1601 499
rect 161 390 456 410
rect 721 415 901 431
rect 721 391 755 415
rect 101 384 456 390
rect 101 249 137 384
rect 574 357 755 391
rect 935 390 991 424
rect 1353 420 1387 465
rect 1255 403 1387 420
rect 935 371 1025 390
rect 171 285 187 319
rect 221 285 332 319
rect 366 316 431 350
rect 465 316 514 350
rect 366 314 514 316
rect 298 280 332 285
rect 574 280 608 357
rect 935 337 951 371
rect 985 337 1025 371
rect 935 335 1025 337
rect 1061 386 1387 403
rect 1423 413 1461 429
rect 1061 371 1289 386
rect 1061 369 1239 371
rect 644 321 899 323
rect 644 287 660 321
rect 694 301 899 321
rect 1061 301 1095 369
rect 1223 337 1239 369
rect 1273 337 1289 371
rect 1457 379 1461 413
rect 1423 363 1461 379
rect 1423 350 1459 363
rect 1223 335 1289 337
rect 694 287 1095 301
rect 298 251 608 280
rect 865 267 1095 287
rect 1129 317 1181 333
rect 1129 283 1131 317
rect 1165 301 1181 317
rect 1165 283 1339 301
rect 1129 267 1339 283
rect 101 215 245 249
rect 298 246 743 251
rect 574 217 743 246
rect 211 210 245 215
rect 211 192 495 210
rect 17 175 175 181
rect 211 176 445 192
rect 17 145 125 175
rect 109 141 125 145
rect 159 141 175 175
rect 429 158 445 176
rect 479 158 495 192
rect 709 194 743 217
rect 941 199 1236 233
rect 429 142 495 158
rect 533 178 599 183
rect 533 144 549 178
rect 583 144 599 178
rect 23 95 75 111
rect 23 61 39 95
rect 73 61 75 95
rect 23 17 75 61
rect 109 93 175 141
rect 109 59 125 93
rect 159 59 175 93
rect 109 51 175 59
rect 209 126 265 142
rect 209 92 215 126
rect 249 92 265 126
rect 209 17 265 92
rect 327 140 393 142
rect 327 106 343 140
rect 377 108 393 140
rect 533 108 599 144
rect 377 106 599 108
rect 327 74 599 106
rect 633 167 675 183
rect 633 133 635 167
rect 669 133 675 167
rect 633 17 675 133
rect 709 178 907 194
rect 709 144 865 178
rect 899 144 907 178
rect 709 128 907 144
rect 941 178 987 199
rect 941 144 951 178
rect 985 144 987 178
rect 1196 191 1236 199
rect 941 128 987 144
rect 1021 131 1037 165
rect 1071 131 1112 165
rect 1146 131 1162 165
rect 1196 157 1198 191
rect 1232 157 1236 191
rect 1196 141 1236 157
rect 1021 17 1162 131
rect 1305 139 1339 267
rect 1373 211 1459 350
rect 1563 350 1601 465
rect 1736 483 1805 499
rect 1736 449 1740 483
rect 1774 449 1805 483
rect 1736 424 1805 449
rect 1736 415 1759 424
rect 1736 381 1740 415
rect 1793 390 1805 424
rect 1774 381 1805 390
rect 1563 319 1653 350
rect 1493 293 1529 309
rect 1493 259 1495 293
rect 1563 285 1603 319
rect 1637 285 1653 319
rect 1563 283 1653 285
rect 1493 249 1529 259
rect 1736 249 1805 381
rect 1493 215 1805 249
rect 1373 177 1409 211
rect 1443 177 1459 211
rect 1373 173 1459 177
rect 1736 209 1805 215
rect 1736 175 1755 209
rect 1789 175 1805 209
rect 1736 173 1805 175
rect 1305 105 1805 139
rect 1700 99 1805 105
rect 1291 69 1357 71
rect 1291 35 1307 69
rect 1341 35 1357 69
rect 1291 17 1357 35
rect 1495 69 1561 71
rect 1495 35 1511 69
rect 1545 35 1561 69
rect 1700 65 1716 99
rect 1750 65 1805 99
rect 1700 51 1805 65
rect 1495 17 1561 35
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 127 390 161 424
rect 991 390 1025 424
rect 1759 415 1793 424
rect 1759 390 1774 415
rect 1774 390 1793 415
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 115 424 173 430
rect 115 390 127 424
rect 161 421 173 424
rect 979 424 1037 430
rect 979 421 991 424
rect 161 393 991 421
rect 161 390 173 393
rect 115 384 173 390
rect 979 390 991 393
rect 1025 421 1037 424
rect 1747 424 1805 430
rect 1747 421 1759 424
rect 1025 393 1759 421
rect 1025 390 1037 393
rect 979 384 1037 390
rect 1747 390 1759 393
rect 1793 390 1805 424
rect 1747 384 1805 390
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fa_2
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1759 94 1793 128 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2433104
string GDS_START 2420058
<< end >>
