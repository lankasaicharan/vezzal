magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 332 1286 704
<< pwell >>
rect 106 49 1180 248
rect 0 0 1248 49
<< scpmos >>
rect 81 368 117 592
rect 171 368 207 592
rect 367 368 403 592
rect 457 368 493 592
rect 574 368 610 592
rect 664 368 700 592
rect 861 368 897 592
rect 951 368 987 592
rect 1041 368 1077 592
rect 1131 368 1167 592
<< nmoslvt >>
rect 189 74 219 222
rect 275 74 305 222
rect 375 74 405 222
rect 475 74 505 222
rect 574 74 604 222
rect 661 74 691 222
rect 753 74 783 222
rect 867 74 897 222
rect 953 74 983 222
rect 1053 74 1083 222
<< ndiff >>
rect 132 186 189 222
rect 132 152 144 186
rect 178 152 189 186
rect 132 118 189 152
rect 132 84 144 118
rect 178 84 189 118
rect 132 74 189 84
rect 219 179 275 222
rect 219 145 230 179
rect 264 145 275 179
rect 219 74 275 145
rect 305 210 375 222
rect 305 176 330 210
rect 364 176 375 210
rect 305 120 375 176
rect 305 86 330 120
rect 364 86 375 120
rect 305 74 375 86
rect 405 143 475 222
rect 405 109 430 143
rect 464 109 475 143
rect 405 74 475 109
rect 505 210 574 222
rect 505 176 516 210
rect 550 176 574 210
rect 505 120 574 176
rect 505 86 516 120
rect 550 86 574 120
rect 505 74 574 86
rect 604 143 661 222
rect 604 109 616 143
rect 650 109 661 143
rect 604 74 661 109
rect 691 210 753 222
rect 691 176 705 210
rect 739 176 753 210
rect 691 120 753 176
rect 691 86 705 120
rect 739 86 753 120
rect 691 74 753 86
rect 783 143 867 222
rect 783 109 808 143
rect 842 109 867 143
rect 783 74 867 109
rect 897 210 953 222
rect 897 176 908 210
rect 942 176 953 210
rect 897 120 953 176
rect 897 86 908 120
rect 942 86 953 120
rect 897 74 953 86
rect 983 143 1053 222
rect 983 109 1008 143
rect 1042 109 1053 143
rect 983 74 1053 109
rect 1083 210 1154 222
rect 1083 176 1108 210
rect 1142 176 1154 210
rect 1083 120 1154 176
rect 1083 86 1108 120
rect 1142 86 1154 120
rect 1083 74 1154 86
<< pdiff >>
rect 27 580 81 592
rect 27 546 37 580
rect 71 546 81 580
rect 27 497 81 546
rect 27 463 37 497
rect 71 463 81 497
rect 27 414 81 463
rect 27 380 37 414
rect 71 380 81 414
rect 27 368 81 380
rect 117 580 171 592
rect 117 546 127 580
rect 161 546 171 580
rect 117 497 171 546
rect 117 463 127 497
rect 161 463 171 497
rect 117 414 171 463
rect 117 380 127 414
rect 161 380 171 414
rect 117 368 171 380
rect 207 580 260 592
rect 207 546 217 580
rect 251 546 260 580
rect 207 462 260 546
rect 207 428 217 462
rect 251 428 260 462
rect 207 368 260 428
rect 314 580 367 592
rect 314 546 323 580
rect 357 546 367 580
rect 314 462 367 546
rect 314 428 323 462
rect 357 428 367 462
rect 314 368 367 428
rect 403 531 457 592
rect 403 497 413 531
rect 447 497 457 531
rect 403 414 457 497
rect 403 380 413 414
rect 447 380 457 414
rect 403 368 457 380
rect 493 580 574 592
rect 493 546 503 580
rect 537 546 574 580
rect 493 510 574 546
rect 493 476 503 510
rect 537 476 574 510
rect 493 440 574 476
rect 493 406 503 440
rect 537 406 574 440
rect 493 368 574 406
rect 610 580 664 592
rect 610 546 620 580
rect 654 546 664 580
rect 610 508 664 546
rect 610 474 620 508
rect 654 474 664 508
rect 610 368 664 474
rect 700 531 753 592
rect 700 497 710 531
rect 744 497 753 531
rect 700 440 753 497
rect 700 406 710 440
rect 744 406 753 440
rect 700 368 753 406
rect 807 531 861 592
rect 807 497 817 531
rect 851 497 861 531
rect 807 420 861 497
rect 807 386 817 420
rect 851 386 861 420
rect 807 368 861 386
rect 897 580 951 592
rect 897 546 907 580
rect 941 546 951 580
rect 897 508 951 546
rect 897 474 907 508
rect 941 474 951 508
rect 897 368 951 474
rect 987 580 1041 592
rect 987 546 997 580
rect 1031 546 1041 580
rect 987 510 1041 546
rect 987 476 997 510
rect 1031 476 1041 510
rect 987 440 1041 476
rect 987 406 997 440
rect 1031 406 1041 440
rect 987 368 1041 406
rect 1077 580 1131 592
rect 1077 546 1087 580
rect 1121 546 1131 580
rect 1077 508 1131 546
rect 1077 474 1087 508
rect 1121 474 1131 508
rect 1077 368 1131 474
rect 1167 580 1221 592
rect 1167 546 1177 580
rect 1211 546 1221 580
rect 1167 510 1221 546
rect 1167 476 1177 510
rect 1211 476 1221 510
rect 1167 440 1221 476
rect 1167 406 1177 440
rect 1211 406 1221 440
rect 1167 368 1221 406
<< ndiffc >>
rect 144 152 178 186
rect 144 84 178 118
rect 230 145 264 179
rect 330 176 364 210
rect 330 86 364 120
rect 430 109 464 143
rect 516 176 550 210
rect 516 86 550 120
rect 616 109 650 143
rect 705 176 739 210
rect 705 86 739 120
rect 808 109 842 143
rect 908 176 942 210
rect 908 86 942 120
rect 1008 109 1042 143
rect 1108 176 1142 210
rect 1108 86 1142 120
<< pdiffc >>
rect 37 546 71 580
rect 37 463 71 497
rect 37 380 71 414
rect 127 546 161 580
rect 127 463 161 497
rect 127 380 161 414
rect 217 546 251 580
rect 217 428 251 462
rect 323 546 357 580
rect 323 428 357 462
rect 413 497 447 531
rect 413 380 447 414
rect 503 546 537 580
rect 503 476 537 510
rect 503 406 537 440
rect 620 546 654 580
rect 620 474 654 508
rect 710 497 744 531
rect 710 406 744 440
rect 817 497 851 531
rect 817 386 851 420
rect 907 546 941 580
rect 907 474 941 508
rect 997 546 1031 580
rect 997 476 1031 510
rect 997 406 1031 440
rect 1087 546 1121 580
rect 1087 474 1121 508
rect 1177 546 1211 580
rect 1177 476 1211 510
rect 1177 406 1211 440
<< poly >>
rect 81 592 117 618
rect 171 592 207 618
rect 367 592 403 618
rect 457 592 493 618
rect 574 592 610 618
rect 664 592 700 618
rect 861 592 897 618
rect 951 592 987 618
rect 1041 592 1077 618
rect 1131 592 1167 618
rect 81 326 117 368
rect 25 310 117 326
rect 171 310 207 368
rect 25 276 41 310
rect 75 294 207 310
rect 75 276 130 294
rect 25 260 130 276
rect 164 274 207 294
rect 367 325 403 368
rect 457 336 493 368
rect 574 336 610 368
rect 664 336 700 368
rect 861 345 897 368
rect 951 345 987 368
rect 457 325 532 336
rect 367 320 532 325
rect 367 286 482 320
rect 516 286 532 320
rect 164 260 305 274
rect 367 270 532 286
rect 574 320 700 336
rect 574 286 641 320
rect 675 306 700 320
rect 753 320 987 345
rect 675 286 691 306
rect 574 270 691 286
rect 25 244 305 260
rect 25 242 117 244
rect 25 208 41 242
rect 75 208 117 242
rect 189 222 219 244
rect 275 222 305 244
rect 375 222 405 270
rect 475 222 505 270
rect 574 222 604 270
rect 661 222 691 270
rect 753 286 769 320
rect 803 286 837 320
rect 871 315 987 320
rect 1041 336 1077 368
rect 1131 336 1167 368
rect 1041 320 1204 336
rect 871 286 897 315
rect 753 270 897 286
rect 753 222 783 270
rect 867 222 897 270
rect 1041 286 1086 320
rect 1120 286 1154 320
rect 1188 286 1204 320
rect 1041 267 1204 286
rect 953 237 1204 267
rect 953 222 983 237
rect 1053 222 1083 237
rect 25 174 117 208
rect 25 140 41 174
rect 75 140 117 174
rect 25 106 117 140
rect 25 72 41 106
rect 75 72 117 106
rect 25 56 117 72
rect 189 48 219 74
rect 275 48 305 74
rect 375 48 405 74
rect 475 48 505 74
rect 574 48 604 74
rect 661 48 691 74
rect 753 48 783 74
rect 867 48 897 74
rect 953 48 983 74
rect 1053 48 1083 74
<< polycont >>
rect 41 276 75 310
rect 130 260 164 294
rect 482 286 516 320
rect 641 286 675 320
rect 41 208 75 242
rect 769 286 803 320
rect 837 286 871 320
rect 1086 286 1120 320
rect 1154 286 1188 320
rect 41 140 75 174
rect 41 72 75 106
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 21 580 87 649
rect 21 546 37 580
rect 71 546 87 580
rect 21 497 87 546
rect 21 463 37 497
rect 71 463 87 497
rect 21 414 87 463
rect 21 380 37 414
rect 71 380 87 414
rect 21 364 87 380
rect 127 580 161 596
rect 127 497 161 546
rect 127 414 161 463
rect 201 580 267 649
rect 201 546 217 580
rect 251 546 267 580
rect 201 462 267 546
rect 201 428 217 462
rect 251 428 267 462
rect 201 412 267 428
rect 307 581 553 615
rect 307 580 373 581
rect 307 546 323 580
rect 357 546 373 580
rect 487 580 553 581
rect 307 462 373 546
rect 307 428 323 462
rect 357 428 373 462
rect 307 412 373 428
rect 407 531 447 547
rect 407 497 413 531
rect 407 414 447 497
rect 127 378 161 380
rect 407 380 413 414
rect 487 546 503 580
rect 537 546 553 580
rect 487 510 553 546
rect 487 476 503 510
rect 537 476 553 510
rect 487 440 553 476
rect 604 581 941 615
rect 604 580 654 581
rect 604 546 620 580
rect 907 580 941 581
rect 604 508 654 546
rect 604 474 620 508
rect 604 458 654 474
rect 694 531 760 547
rect 694 497 710 531
rect 744 497 760 531
rect 487 406 503 440
rect 537 424 553 440
rect 694 440 760 497
rect 694 424 710 440
rect 537 406 710 424
rect 744 406 760 440
rect 487 390 760 406
rect 801 531 867 547
rect 801 497 817 531
rect 851 497 867 531
rect 801 424 867 497
rect 907 508 941 546
rect 907 458 941 474
rect 981 580 1047 596
rect 981 546 997 580
rect 1031 546 1047 580
rect 981 510 1047 546
rect 981 476 997 510
rect 1031 476 1047 510
rect 981 440 1047 476
rect 1087 580 1121 649
rect 1087 508 1121 546
rect 1087 458 1121 474
rect 1161 580 1227 596
rect 1161 546 1177 580
rect 1211 546 1227 580
rect 1161 510 1227 546
rect 1161 476 1177 510
rect 1211 476 1227 510
rect 981 424 997 440
rect 801 420 997 424
rect 407 378 447 380
rect 127 344 447 378
rect 801 386 817 420
rect 851 406 997 420
rect 1031 424 1047 440
rect 1161 440 1227 476
rect 1161 424 1177 440
rect 1031 406 1177 424
rect 1211 406 1227 440
rect 851 390 1227 406
rect 851 386 867 390
rect 801 370 867 386
rect 25 310 91 326
rect 214 310 447 344
rect 481 320 551 356
rect 25 276 41 310
rect 75 294 180 310
rect 75 276 130 294
rect 25 260 130 276
rect 164 260 180 294
rect 25 242 180 260
rect 25 208 41 242
rect 75 236 180 242
rect 75 208 91 236
rect 25 174 91 208
rect 25 140 41 174
rect 75 140 91 174
rect 25 106 91 140
rect 25 72 41 106
rect 75 72 91 106
rect 25 56 91 72
rect 128 186 178 202
rect 128 152 144 186
rect 128 118 178 152
rect 214 179 280 310
rect 481 286 482 320
rect 516 286 551 320
rect 481 270 551 286
rect 601 320 691 356
rect 985 336 1031 356
rect 601 286 641 320
rect 675 286 691 320
rect 601 270 691 286
rect 753 320 1031 336
rect 753 286 769 320
rect 803 286 837 320
rect 871 286 1031 320
rect 753 270 1031 286
rect 1070 320 1223 356
rect 1070 286 1086 320
rect 1120 286 1154 320
rect 1188 286 1223 320
rect 1070 270 1223 286
rect 214 145 230 179
rect 264 145 280 179
rect 214 129 280 145
rect 314 210 1158 236
rect 314 176 330 210
rect 364 202 516 210
rect 364 176 380 202
rect 128 84 144 118
rect 314 120 380 176
rect 550 202 705 210
rect 550 176 566 202
rect 314 86 330 120
rect 364 86 380 120
rect 314 85 380 86
rect 178 84 380 85
rect 128 51 380 84
rect 414 143 480 159
rect 414 109 430 143
rect 464 109 480 143
rect 414 17 480 109
rect 516 120 566 176
rect 702 176 705 202
rect 739 202 908 210
rect 739 176 758 202
rect 550 86 566 120
rect 516 70 566 86
rect 600 143 666 159
rect 600 109 616 143
rect 650 109 666 143
rect 600 17 666 109
rect 702 120 758 176
rect 892 176 908 202
rect 942 202 1108 210
rect 942 176 958 202
rect 702 86 705 120
rect 739 86 758 120
rect 702 70 758 86
rect 792 143 858 159
rect 792 109 808 143
rect 842 109 858 143
rect 792 17 858 109
rect 892 120 958 176
rect 1092 176 1108 202
rect 1142 176 1158 210
rect 892 86 908 120
rect 942 86 958 120
rect 892 70 958 86
rect 992 143 1058 159
rect 992 109 1008 143
rect 1042 109 1058 143
rect 992 17 1058 109
rect 1092 120 1158 176
rect 1092 86 1108 120
rect 1142 86 1158 120
rect 1092 70 1158 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o41ai_2
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 3563556
string GDS_START 3553160
<< end >>
