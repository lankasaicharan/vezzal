magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 369 1574 704
rect -38 331 146 369
rect 491 331 1574 369
<< pwell >>
rect 188 232 449 295
rect 1 157 449 232
rect 1103 157 1535 167
rect 1 49 1535 157
rect 0 0 1536 49
<< scnmos >>
rect 84 122 114 206
rect 162 122 192 206
rect 264 185 294 269
rect 336 185 366 269
rect 470 47 500 131
rect 542 47 572 131
rect 628 47 658 131
rect 706 47 736 131
rect 820 47 850 131
rect 898 47 928 131
rect 1186 57 1216 141
rect 1264 57 1294 141
rect 1350 57 1380 141
rect 1422 57 1452 141
<< scpmoshvt >>
rect 84 419 134 619
rect 206 405 256 605
rect 478 419 528 619
rect 690 419 740 619
rect 788 419 838 619
rect 894 419 944 619
rect 994 419 1044 619
rect 1135 419 1185 619
rect 1241 419 1291 619
rect 1356 419 1406 619
<< ndiff >>
rect 214 206 264 269
rect 27 177 84 206
rect 27 143 39 177
rect 73 143 84 177
rect 27 122 84 143
rect 114 122 162 206
rect 192 185 264 206
rect 294 185 336 269
rect 366 235 423 269
rect 366 201 377 235
rect 411 201 423 235
rect 366 185 423 201
rect 192 177 249 185
rect 192 143 203 177
rect 237 143 249 177
rect 192 122 249 143
rect 413 111 470 131
rect 413 77 425 111
rect 459 77 470 111
rect 413 47 470 77
rect 500 47 542 131
rect 572 93 628 131
rect 572 59 583 93
rect 617 59 628 93
rect 572 47 628 59
rect 658 47 706 131
rect 736 93 820 131
rect 736 59 775 93
rect 809 59 820 93
rect 736 47 820 59
rect 850 47 898 131
rect 928 106 1072 131
rect 928 72 1026 106
rect 1060 72 1072 106
rect 928 47 1072 72
rect 1129 116 1186 141
rect 1129 82 1141 116
rect 1175 82 1186 116
rect 1129 57 1186 82
rect 1216 57 1264 141
rect 1294 113 1350 141
rect 1294 79 1305 113
rect 1339 79 1350 113
rect 1294 57 1350 79
rect 1380 57 1422 141
rect 1452 116 1509 141
rect 1452 82 1463 116
rect 1497 82 1509 116
rect 1452 57 1509 82
<< pdiff >>
rect 27 597 84 619
rect 27 563 39 597
rect 73 563 84 597
rect 27 465 84 563
rect 27 431 39 465
rect 73 431 84 465
rect 27 419 84 431
rect 134 607 191 619
rect 134 573 145 607
rect 179 605 191 607
rect 179 573 206 605
rect 134 419 206 573
rect 156 405 206 419
rect 256 451 313 605
rect 256 417 267 451
rect 301 417 313 451
rect 421 597 478 619
rect 421 563 433 597
rect 467 563 478 597
rect 421 513 478 563
rect 421 479 433 513
rect 467 479 478 513
rect 421 419 478 479
rect 528 587 690 619
rect 528 553 539 587
rect 573 553 690 587
rect 528 419 690 553
rect 740 419 788 619
rect 838 597 894 619
rect 838 563 849 597
rect 883 563 894 597
rect 838 489 894 563
rect 838 455 849 489
rect 883 455 894 489
rect 838 419 894 455
rect 944 419 994 619
rect 1044 607 1135 619
rect 1044 573 1074 607
rect 1108 573 1135 607
rect 1044 536 1135 573
rect 1044 502 1074 536
rect 1108 502 1135 536
rect 1044 465 1135 502
rect 1044 431 1074 465
rect 1108 431 1135 465
rect 1044 419 1135 431
rect 1185 597 1241 619
rect 1185 563 1196 597
rect 1230 563 1241 597
rect 1185 465 1241 563
rect 1185 431 1196 465
rect 1230 431 1241 465
rect 1185 419 1241 431
rect 1291 607 1356 619
rect 1291 573 1302 607
rect 1336 573 1356 607
rect 1291 536 1356 573
rect 1291 502 1302 536
rect 1336 502 1356 536
rect 1291 465 1356 502
rect 1291 431 1302 465
rect 1336 431 1356 465
rect 1291 419 1356 431
rect 1406 597 1463 619
rect 1406 563 1417 597
rect 1451 563 1463 597
rect 1406 465 1463 563
rect 1406 431 1417 465
rect 1451 431 1463 465
rect 1406 419 1463 431
rect 256 405 313 417
<< ndiffc >>
rect 39 143 73 177
rect 377 201 411 235
rect 203 143 237 177
rect 425 77 459 111
rect 583 59 617 93
rect 775 59 809 93
rect 1026 72 1060 106
rect 1141 82 1175 116
rect 1305 79 1339 113
rect 1463 82 1497 116
<< pdiffc >>
rect 39 563 73 597
rect 39 431 73 465
rect 145 573 179 607
rect 267 417 301 451
rect 433 563 467 597
rect 433 479 467 513
rect 539 553 573 587
rect 849 563 883 597
rect 849 455 883 489
rect 1074 573 1108 607
rect 1074 502 1108 536
rect 1074 431 1108 465
rect 1196 563 1230 597
rect 1196 431 1230 465
rect 1302 573 1336 607
rect 1302 502 1336 536
rect 1302 431 1336 465
rect 1417 563 1451 597
rect 1417 431 1451 465
<< poly >>
rect 84 619 134 645
rect 206 605 256 631
rect 478 619 528 645
rect 690 619 740 645
rect 788 619 838 645
rect 894 619 944 645
rect 994 619 1044 645
rect 1135 619 1185 645
rect 1241 619 1291 645
rect 1356 619 1406 645
rect 84 373 134 419
rect 84 357 154 373
rect 206 365 256 405
rect 478 393 528 419
rect 84 323 104 357
rect 138 323 154 357
rect 84 289 154 323
rect 196 349 294 365
rect 478 357 508 393
rect 196 315 212 349
rect 246 329 294 349
rect 442 341 508 357
rect 690 381 740 419
rect 690 351 720 381
rect 246 315 366 329
rect 196 299 366 315
rect 84 255 104 289
rect 138 255 154 289
rect 264 269 294 299
rect 336 269 366 299
rect 442 307 458 341
rect 492 307 508 341
rect 442 291 508 307
rect 550 335 720 351
rect 550 301 566 335
rect 600 301 720 335
rect 788 345 838 419
rect 894 387 944 419
rect 886 371 952 387
rect 788 333 834 345
rect 84 251 154 255
rect 84 221 192 251
rect 84 206 114 221
rect 162 206 192 221
rect 264 159 294 185
rect 336 159 366 185
rect 470 176 500 291
rect 550 285 720 301
rect 768 317 834 333
rect 470 146 572 176
rect 470 131 500 146
rect 542 131 572 146
rect 628 131 658 285
rect 768 283 784 317
rect 818 297 834 317
rect 886 337 902 371
rect 936 337 952 371
rect 886 303 952 337
rect 818 283 844 297
rect 768 267 844 283
rect 706 203 772 219
rect 706 169 722 203
rect 756 169 772 203
rect 706 153 772 169
rect 814 176 844 267
rect 886 269 902 303
rect 936 269 952 303
rect 886 253 952 269
rect 994 285 1044 419
rect 1135 351 1185 419
rect 1241 379 1291 419
rect 1241 363 1308 379
rect 1086 335 1196 351
rect 1086 301 1102 335
rect 1136 301 1196 335
rect 1086 285 1196 301
rect 994 237 1024 285
rect 994 221 1124 237
rect 994 201 1074 221
rect 898 187 1074 201
rect 1108 187 1124 221
rect 706 131 736 153
rect 814 146 850 176
rect 820 131 850 146
rect 898 171 1124 187
rect 1166 197 1196 285
rect 1241 329 1258 363
rect 1292 329 1308 363
rect 1241 295 1308 329
rect 1356 309 1406 419
rect 1241 261 1258 295
rect 1292 261 1308 295
rect 1241 245 1308 261
rect 1350 293 1452 309
rect 1350 259 1371 293
rect 1405 259 1452 293
rect 898 131 928 171
rect 1166 167 1216 197
rect 1186 141 1216 167
rect 1264 141 1294 245
rect 1350 225 1452 259
rect 1350 191 1371 225
rect 1405 191 1452 225
rect 1350 175 1452 191
rect 1350 141 1380 175
rect 1422 141 1452 175
rect 84 96 114 122
rect 162 96 192 122
rect 470 21 500 47
rect 542 21 572 47
rect 628 21 658 47
rect 706 21 736 47
rect 820 21 850 47
rect 898 21 928 47
rect 1186 31 1216 57
rect 1264 31 1294 57
rect 1350 31 1380 57
rect 1422 31 1452 57
<< polycont >>
rect 104 323 138 357
rect 212 315 246 349
rect 104 255 138 289
rect 458 307 492 341
rect 566 301 600 335
rect 784 283 818 317
rect 902 337 936 371
rect 722 169 756 203
rect 902 269 936 303
rect 1102 301 1136 335
rect 1074 187 1108 221
rect 1258 329 1292 363
rect 1258 261 1292 295
rect 1371 259 1405 293
rect 1371 191 1405 225
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 18 597 89 613
rect 18 563 39 597
rect 73 563 89 597
rect 18 521 89 563
rect 129 607 195 649
rect 129 573 145 607
rect 179 573 195 607
rect 129 557 195 573
rect 433 597 483 613
rect 467 563 483 597
rect 18 487 397 521
rect 18 465 89 487
rect 18 431 39 465
rect 73 431 89 465
rect 18 415 89 431
rect 251 417 267 451
rect 301 417 327 451
rect 18 203 52 415
rect 251 401 327 417
rect 88 357 161 373
rect 88 323 104 357
rect 138 323 161 357
rect 88 289 161 323
rect 197 349 257 365
rect 197 315 212 349
rect 246 315 257 349
rect 197 299 257 315
rect 293 357 327 401
rect 363 427 397 487
rect 433 513 483 563
rect 523 587 589 649
rect 523 553 539 587
rect 573 553 589 587
rect 523 533 589 553
rect 833 597 899 613
rect 833 563 849 597
rect 883 563 899 597
rect 467 497 483 513
rect 467 479 797 497
rect 433 463 797 479
rect 363 393 608 427
rect 293 341 508 357
rect 293 307 458 341
rect 492 307 508 341
rect 293 291 508 307
rect 88 255 104 289
rect 138 255 161 289
rect 88 239 161 255
rect 361 235 427 291
rect 18 177 89 203
rect 18 143 39 177
rect 73 143 89 177
rect 18 118 89 143
rect 187 177 253 203
rect 361 201 377 235
rect 411 201 427 235
rect 474 249 508 291
rect 550 335 608 393
rect 763 403 797 463
rect 833 489 899 563
rect 833 455 849 489
rect 883 473 899 489
rect 1058 607 1124 649
rect 1058 573 1074 607
rect 1108 573 1124 607
rect 1058 536 1124 573
rect 1058 502 1074 536
rect 1108 502 1124 536
rect 883 455 1022 473
rect 833 439 1022 455
rect 763 371 952 403
rect 763 369 902 371
rect 550 301 566 335
rect 600 301 608 335
rect 870 337 902 369
rect 936 337 952 371
rect 550 285 608 301
rect 644 317 834 333
rect 644 283 784 317
rect 818 283 834 317
rect 644 267 834 283
rect 870 303 952 337
rect 870 269 902 303
rect 936 269 952 303
rect 644 249 678 267
rect 474 215 678 249
rect 870 253 952 269
rect 988 351 1022 439
rect 1058 465 1124 502
rect 1058 431 1074 465
rect 1108 431 1124 465
rect 1058 415 1124 431
rect 1180 597 1246 613
rect 1180 563 1196 597
rect 1230 563 1246 597
rect 1180 465 1246 563
rect 1180 431 1196 465
rect 1230 431 1246 465
rect 1180 415 1246 431
rect 1286 607 1352 649
rect 1286 573 1302 607
rect 1336 573 1352 607
rect 1286 536 1352 573
rect 1286 502 1302 536
rect 1336 502 1352 536
rect 1286 465 1352 502
rect 1286 431 1302 465
rect 1336 431 1352 465
rect 1286 415 1352 431
rect 1401 597 1513 613
rect 1401 563 1417 597
rect 1451 563 1513 597
rect 1401 465 1513 563
rect 1401 431 1417 465
rect 1451 431 1513 465
rect 1401 415 1513 431
rect 988 335 1144 351
rect 988 301 1102 335
rect 1136 301 1144 335
rect 988 285 1144 301
rect 870 219 904 253
rect 361 181 427 201
rect 714 203 904 219
rect 988 205 1022 285
rect 714 179 722 203
rect 187 143 203 177
rect 237 143 253 177
rect 187 17 253 143
rect 463 169 722 179
rect 756 185 904 203
rect 756 169 772 185
rect 463 145 772 169
rect 940 171 1022 205
rect 1058 221 1124 237
rect 1058 187 1074 221
rect 1108 205 1124 221
rect 1180 209 1214 415
rect 1250 363 1319 379
rect 1250 329 1258 363
rect 1292 329 1319 363
rect 1250 295 1319 329
rect 1250 261 1258 295
rect 1292 261 1319 295
rect 1250 245 1319 261
rect 1355 293 1421 309
rect 1355 259 1371 293
rect 1405 259 1421 293
rect 1355 225 1421 259
rect 1355 209 1371 225
rect 1180 205 1371 209
rect 1108 191 1371 205
rect 1405 191 1421 225
rect 1108 187 1421 191
rect 1058 175 1421 187
rect 1058 171 1214 175
rect 463 135 497 145
rect 409 111 497 135
rect 409 77 425 111
rect 459 77 497 111
rect 940 109 974 171
rect 409 53 497 77
rect 567 93 633 109
rect 567 59 583 93
rect 617 59 633 93
rect 759 93 974 109
rect 759 59 775 93
rect 809 59 974 93
rect 1010 106 1076 135
rect 1010 72 1026 106
rect 1060 72 1076 106
rect 567 17 633 59
rect 1010 17 1076 72
rect 1125 116 1214 171
rect 1125 82 1141 116
rect 1175 82 1214 116
rect 1125 53 1214 82
rect 1289 113 1355 139
rect 1289 79 1305 113
rect 1339 79 1355 113
rect 1289 17 1355 79
rect 1463 116 1513 415
rect 1497 82 1513 116
rect 1463 53 1513 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrtp_lp2
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1471 94 1505 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 168 1505 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 390 1505 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 464 1505 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1471 538 1505 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1883576
string GDS_START 1872132
<< end >>
