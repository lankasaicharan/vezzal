magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3598 1852
<< nwell >>
rect -38 261 2338 582
<< pwell >>
rect 973 157 1169 201
rect 1793 157 2275 203
rect 1 21 2275 157
rect 29 -17 63 21
<< scnmos >>
rect 89 47 119 131
rect 183 47 213 131
rect 438 47 468 131
rect 553 47 583 119
rect 659 47 689 119
rect 835 47 865 131
rect 907 47 937 131
rect 1059 47 1089 175
rect 1158 47 1188 119
rect 1287 47 1317 119
rect 1403 47 1433 131
rect 1582 47 1612 131
rect 1683 47 1713 131
rect 1881 47 1911 177
rect 1975 47 2005 177
rect 2069 47 2099 177
rect 2163 47 2193 177
<< scpmoshvt >>
rect 81 363 117 491
rect 175 363 211 491
rect 452 413 488 497
rect 554 413 590 497
rect 663 413 699 497
rect 813 413 849 497
rect 920 413 956 497
rect 1137 329 1173 497
rect 1246 413 1282 497
rect 1352 413 1388 497
rect 1456 413 1492 497
rect 1574 413 1610 497
rect 1668 413 1704 497
rect 1873 297 1909 497
rect 1967 297 2003 497
rect 2061 297 2097 497
rect 2155 297 2191 497
<< ndiff >>
rect 27 119 89 131
rect 27 85 35 119
rect 69 85 89 119
rect 27 47 89 85
rect 119 93 183 131
rect 119 59 129 93
rect 163 59 183 93
rect 119 47 183 59
rect 213 119 265 131
rect 213 85 223 119
rect 257 85 265 119
rect 213 47 265 85
rect 333 89 438 131
rect 333 55 345 89
rect 379 55 438 89
rect 333 47 438 55
rect 468 119 528 131
rect 999 131 1059 175
rect 707 119 835 131
rect 468 95 553 119
rect 468 61 488 95
rect 522 61 553 95
rect 468 47 553 61
rect 583 95 659 119
rect 583 61 605 95
rect 639 61 659 95
rect 583 47 659 61
rect 689 47 835 119
rect 865 47 907 131
rect 937 93 1059 131
rect 937 59 981 93
rect 1015 59 1059 93
rect 937 47 1059 59
rect 1089 119 1143 175
rect 1819 163 1881 177
rect 1343 119 1403 131
rect 1089 89 1158 119
rect 1089 55 1103 89
rect 1137 55 1158 89
rect 1089 47 1158 55
rect 1188 93 1287 119
rect 1188 59 1223 93
rect 1257 59 1287 93
rect 1188 47 1287 59
rect 1317 47 1403 119
rect 1433 89 1582 131
rect 1433 55 1475 89
rect 1509 55 1582 89
rect 1433 47 1582 55
rect 1612 47 1683 131
rect 1713 109 1765 131
rect 1713 75 1723 109
rect 1757 75 1765 109
rect 1713 47 1765 75
rect 1819 129 1827 163
rect 1861 129 1881 163
rect 1819 95 1881 129
rect 1819 61 1827 95
rect 1861 61 1881 95
rect 1819 47 1881 61
rect 1911 163 1975 177
rect 1911 129 1921 163
rect 1955 129 1975 163
rect 1911 95 1975 129
rect 1911 61 1921 95
rect 1955 61 1975 95
rect 1911 47 1975 61
rect 2005 95 2069 177
rect 2005 61 2015 95
rect 2049 61 2069 95
rect 2005 47 2069 61
rect 2099 163 2163 177
rect 2099 129 2109 163
rect 2143 129 2163 163
rect 2099 95 2163 129
rect 2099 61 2109 95
rect 2143 61 2163 95
rect 2099 47 2163 61
rect 2193 95 2249 177
rect 2193 61 2203 95
rect 2237 61 2249 95
rect 2193 47 2249 61
<< pdiff >>
rect 27 477 81 491
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 363 81 375
rect 117 461 175 491
rect 117 427 129 461
rect 163 427 175 461
rect 117 363 175 427
rect 211 477 265 491
rect 211 443 223 477
rect 257 443 265 477
rect 211 409 265 443
rect 398 485 452 497
rect 398 451 406 485
rect 440 451 452 485
rect 398 413 452 451
rect 488 477 554 497
rect 488 443 500 477
rect 534 443 554 477
rect 488 413 554 443
rect 590 483 663 497
rect 590 449 603 483
rect 637 449 663 483
rect 590 413 663 449
rect 699 459 813 497
rect 699 425 767 459
rect 801 425 813 459
rect 699 413 813 425
rect 849 475 920 497
rect 849 441 874 475
rect 908 441 920 475
rect 849 413 920 441
rect 956 459 1010 497
rect 956 425 968 459
rect 1002 425 1010 459
rect 956 413 1010 425
rect 1073 485 1137 497
rect 1073 451 1091 485
rect 1125 451 1137 485
rect 211 375 223 409
rect 257 375 265 409
rect 211 363 265 375
rect 1073 329 1137 451
rect 1173 477 1246 497
rect 1173 443 1189 477
rect 1223 443 1246 477
rect 1173 413 1246 443
rect 1282 484 1352 497
rect 1282 450 1296 484
rect 1330 450 1352 484
rect 1282 413 1352 450
rect 1388 413 1456 497
rect 1492 485 1574 497
rect 1492 451 1528 485
rect 1562 451 1574 485
rect 1492 413 1574 451
rect 1610 459 1668 497
rect 1610 425 1622 459
rect 1656 425 1668 459
rect 1610 413 1668 425
rect 1704 485 1760 497
rect 1704 451 1718 485
rect 1752 451 1760 485
rect 1704 413 1760 451
rect 1819 485 1873 497
rect 1819 451 1827 485
rect 1861 451 1873 485
rect 1819 417 1873 451
rect 1173 329 1229 413
rect 1819 383 1827 417
rect 1861 383 1873 417
rect 1819 297 1873 383
rect 1909 477 1967 497
rect 1909 443 1921 477
rect 1955 443 1967 477
rect 1909 409 1967 443
rect 1909 375 1921 409
rect 1955 375 1967 409
rect 1909 341 1967 375
rect 1909 307 1921 341
rect 1955 307 1967 341
rect 1909 297 1967 307
rect 2003 477 2061 497
rect 2003 443 2015 477
rect 2049 443 2061 477
rect 2003 409 2061 443
rect 2003 375 2015 409
rect 2049 375 2061 409
rect 2003 297 2061 375
rect 2097 477 2155 497
rect 2097 443 2109 477
rect 2143 443 2155 477
rect 2097 409 2155 443
rect 2097 375 2109 409
rect 2143 375 2155 409
rect 2097 341 2155 375
rect 2097 307 2109 341
rect 2143 307 2155 341
rect 2097 297 2155 307
rect 2191 477 2254 497
rect 2191 443 2203 477
rect 2237 443 2254 477
rect 2191 409 2254 443
rect 2191 375 2203 409
rect 2237 375 2254 409
rect 2191 297 2254 375
<< ndiffc >>
rect 35 85 69 119
rect 129 59 163 93
rect 223 85 257 119
rect 345 55 379 89
rect 488 61 522 95
rect 605 61 639 95
rect 981 59 1015 93
rect 1103 55 1137 89
rect 1223 59 1257 93
rect 1475 55 1509 89
rect 1723 75 1757 109
rect 1827 129 1861 163
rect 1827 61 1861 95
rect 1921 129 1955 163
rect 1921 61 1955 95
rect 2015 61 2049 95
rect 2109 129 2143 163
rect 2109 61 2143 95
rect 2203 61 2237 95
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 129 427 163 461
rect 223 443 257 477
rect 406 451 440 485
rect 500 443 534 477
rect 603 449 637 483
rect 767 425 801 459
rect 874 441 908 475
rect 968 425 1002 459
rect 1091 451 1125 485
rect 223 375 257 409
rect 1189 443 1223 477
rect 1296 450 1330 484
rect 1528 451 1562 485
rect 1622 425 1656 459
rect 1718 451 1752 485
rect 1827 451 1861 485
rect 1827 383 1861 417
rect 1921 443 1955 477
rect 1921 375 1955 409
rect 1921 307 1955 341
rect 2015 443 2049 477
rect 2015 375 2049 409
rect 2109 443 2143 477
rect 2109 375 2143 409
rect 2109 307 2143 341
rect 2203 443 2237 477
rect 2203 375 2237 409
<< poly >>
rect 81 491 117 517
rect 175 491 211 517
rect 452 497 488 523
rect 554 497 590 523
rect 663 497 699 523
rect 813 497 849 523
rect 920 497 956 523
rect 1137 497 1173 523
rect 1246 497 1282 523
rect 1352 497 1388 523
rect 1456 497 1492 523
rect 1574 497 1610 523
rect 1668 497 1704 523
rect 1873 497 1909 523
rect 1967 497 2003 523
rect 2061 497 2097 523
rect 2155 497 2191 523
rect 452 398 488 413
rect 554 398 590 413
rect 663 398 699 413
rect 813 398 849 413
rect 920 398 956 413
rect 81 348 117 363
rect 175 348 211 363
rect 46 318 119 348
rect 46 265 76 318
rect 173 274 213 348
rect 450 326 490 398
rect 552 375 592 398
rect 22 249 76 265
rect 22 215 32 249
rect 66 215 76 249
rect 128 264 213 274
rect 128 230 144 264
rect 178 230 213 264
rect 351 310 490 326
rect 536 365 612 375
rect 536 331 552 365
rect 586 331 612 365
rect 536 321 612 331
rect 351 276 361 310
rect 395 296 490 310
rect 395 276 468 296
rect 661 279 701 398
rect 811 355 851 398
rect 811 339 876 355
rect 811 305 821 339
rect 855 305 876 339
rect 811 289 876 305
rect 351 260 468 276
rect 128 220 213 230
rect 22 199 76 215
rect 46 176 76 199
rect 46 146 119 176
rect 89 131 119 146
rect 183 131 213 220
rect 438 131 468 260
rect 543 249 701 279
rect 543 219 584 249
rect 520 203 584 219
rect 520 169 530 203
rect 564 169 584 203
rect 520 153 584 169
rect 626 197 702 207
rect 626 163 642 197
rect 676 163 702 197
rect 626 153 702 163
rect 553 119 583 153
rect 659 119 689 153
rect 835 131 865 289
rect 918 219 958 398
rect 1246 398 1282 413
rect 1352 398 1388 413
rect 1456 398 1492 413
rect 1574 398 1610 413
rect 1668 398 1704 413
rect 1137 314 1173 329
rect 1049 284 1175 314
rect 1049 267 1089 284
rect 1013 251 1089 267
rect 907 203 971 219
rect 907 169 917 203
rect 951 169 971 203
rect 1013 217 1023 251
rect 1057 217 1089 251
rect 1244 279 1284 398
rect 1350 381 1390 398
rect 1336 365 1400 381
rect 1336 331 1346 365
rect 1380 331 1400 365
rect 1336 315 1400 331
rect 1244 267 1304 279
rect 1244 255 1327 267
rect 1244 249 1351 255
rect 1265 239 1351 249
rect 1265 237 1297 239
rect 1013 201 1089 217
rect 1059 175 1089 201
rect 1158 191 1235 207
rect 907 153 971 169
rect 907 131 937 153
rect 1158 157 1191 191
rect 1225 157 1235 191
rect 1158 141 1235 157
rect 1287 205 1297 237
rect 1331 205 1351 239
rect 1287 189 1351 205
rect 1454 229 1494 398
rect 1572 257 1612 398
rect 1666 365 1706 398
rect 1654 349 1718 365
rect 1654 315 1664 349
rect 1698 315 1718 349
rect 1654 299 1718 315
rect 1567 241 1631 257
rect 1454 213 1525 229
rect 1454 193 1471 213
rect 1158 119 1188 141
rect 1287 119 1317 189
rect 1403 179 1471 193
rect 1505 179 1525 213
rect 1567 207 1577 241
rect 1611 207 1631 241
rect 1567 191 1631 207
rect 1403 163 1525 179
rect 1403 131 1433 163
rect 1582 131 1612 191
rect 1683 131 1713 299
rect 1873 282 1909 297
rect 1967 282 2003 297
rect 2061 282 2097 297
rect 2155 282 2191 297
rect 1871 265 1911 282
rect 1965 265 2005 282
rect 2059 265 2099 282
rect 2153 265 2193 282
rect 1859 249 2193 265
rect 1859 215 1875 249
rect 1909 215 1953 249
rect 1987 215 2031 249
rect 2065 215 2109 249
rect 2143 215 2193 249
rect 1859 199 2193 215
rect 1881 177 1911 199
rect 1975 177 2005 199
rect 2069 177 2099 199
rect 2163 177 2193 199
rect 89 21 119 47
rect 183 21 213 47
rect 438 21 468 47
rect 553 21 583 47
rect 659 21 689 47
rect 835 21 865 47
rect 907 21 937 47
rect 1059 21 1089 47
rect 1158 21 1188 47
rect 1287 21 1317 47
rect 1403 21 1433 47
rect 1582 21 1612 47
rect 1683 21 1713 47
rect 1881 21 1911 47
rect 1975 21 2005 47
rect 2069 21 2099 47
rect 2163 21 2193 47
<< polycont >>
rect 32 215 66 249
rect 144 230 178 264
rect 552 331 586 365
rect 361 276 395 310
rect 821 305 855 339
rect 530 169 564 203
rect 642 163 676 197
rect 917 169 951 203
rect 1023 217 1057 251
rect 1346 331 1380 365
rect 1191 157 1225 191
rect 1297 205 1331 239
rect 1664 315 1698 349
rect 1471 179 1505 213
rect 1577 207 1611 241
rect 1875 215 1909 249
rect 1953 215 1987 249
rect 2031 215 2065 249
rect 2109 215 2143 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 18 477 69 493
rect 18 443 35 477
rect 18 409 69 443
rect 103 461 179 527
rect 103 427 129 461
rect 163 427 179 461
rect 223 477 257 493
rect 18 375 35 409
rect 223 409 257 443
rect 69 375 178 393
rect 18 359 178 375
rect 18 249 88 325
rect 18 215 32 249
rect 66 215 88 249
rect 18 195 88 215
rect 132 264 178 359
rect 132 255 144 264
rect 166 221 178 230
rect 132 161 178 221
rect 18 127 178 161
rect 18 119 69 127
rect 18 85 35 119
rect 223 119 257 357
rect 291 333 356 490
rect 390 485 440 527
rect 390 451 406 485
rect 390 435 440 451
rect 484 477 534 493
rect 484 443 500 477
rect 484 427 534 443
rect 587 483 733 493
rect 587 449 603 483
rect 637 449 733 483
rect 858 475 924 527
rect 1061 485 1145 527
rect 587 427 733 449
rect 484 401 518 427
rect 429 367 518 401
rect 552 391 655 393
rect 291 310 395 333
rect 291 276 361 310
rect 291 123 395 276
rect 18 69 69 85
rect 103 59 129 93
rect 163 59 179 93
rect 429 95 463 367
rect 552 365 621 391
rect 586 357 621 365
rect 586 331 655 357
rect 552 315 655 331
rect 507 255 587 277
rect 507 221 519 255
rect 553 221 587 255
rect 507 203 587 221
rect 507 169 530 203
rect 564 169 587 203
rect 507 153 587 169
rect 621 197 655 315
rect 699 271 733 427
rect 767 459 801 475
rect 858 441 874 475
rect 908 441 924 475
rect 968 459 1002 475
rect 767 407 801 425
rect 1061 451 1091 485
rect 1125 451 1145 485
rect 1061 435 1145 451
rect 1189 477 1223 493
rect 968 407 1002 425
rect 767 373 1002 407
rect 1189 401 1223 443
rect 1270 484 1494 493
rect 1270 450 1296 484
rect 1330 450 1494 484
rect 1270 425 1494 450
rect 1528 485 1578 527
rect 1562 451 1578 485
rect 1692 485 1768 527
rect 1528 435 1578 451
rect 1622 459 1656 475
rect 1101 367 1223 401
rect 1101 339 1135 367
rect 805 305 821 339
rect 855 305 1135 339
rect 1294 357 1305 391
rect 1339 365 1406 391
rect 1339 357 1346 365
rect 1294 333 1346 357
rect 699 251 1057 271
rect 699 237 1023 251
rect 621 163 642 197
rect 676 163 702 197
rect 621 153 702 163
rect 736 95 770 237
rect 835 187 917 203
rect 951 187 989 203
rect 1023 201 1057 217
rect 835 153 857 187
rect 891 169 917 187
rect 891 153 929 169
rect 963 153 989 187
rect 1101 167 1135 305
rect 223 69 257 85
rect 103 17 179 59
rect 329 55 345 89
rect 379 55 395 89
rect 429 61 488 95
rect 522 61 538 95
rect 589 61 605 95
rect 639 61 770 95
rect 965 93 1031 109
rect 329 17 395 55
rect 965 59 981 93
rect 1015 59 1031 93
rect 965 17 1031 59
rect 1073 89 1135 167
rect 1183 331 1346 333
rect 1380 331 1406 365
rect 1450 349 1494 425
rect 1692 451 1718 485
rect 1752 451 1768 485
rect 1827 485 1861 527
rect 1622 417 1656 425
rect 1827 417 1861 451
rect 1622 383 1792 417
rect 1183 299 1338 331
rect 1450 315 1664 349
rect 1698 315 1724 349
rect 1183 191 1225 299
rect 1450 297 1494 315
rect 1183 157 1191 191
rect 1183 141 1225 157
rect 1259 255 1349 265
rect 1259 239 1305 255
rect 1259 205 1297 239
rect 1339 221 1349 255
rect 1331 205 1349 221
rect 1259 141 1349 205
rect 1393 263 1494 297
rect 1393 107 1427 263
rect 1561 250 1679 281
rect 1758 259 1792 383
rect 1827 315 1861 383
rect 1913 477 1971 493
rect 1913 443 1921 477
rect 1955 443 1971 477
rect 1913 409 1971 443
rect 1913 375 1921 409
rect 1955 375 1971 409
rect 1913 341 1971 375
rect 2015 477 2049 527
rect 2015 409 2049 443
rect 2015 359 2049 375
rect 2101 477 2151 493
rect 2101 443 2109 477
rect 2143 443 2151 477
rect 2101 409 2151 443
rect 2101 375 2109 409
rect 2143 375 2151 409
rect 1913 307 1921 341
rect 1955 325 1971 341
rect 2101 341 2151 375
rect 2203 477 2237 527
rect 2203 409 2237 443
rect 2203 359 2237 375
rect 2101 325 2109 341
rect 1955 307 2109 325
rect 2143 325 2151 341
rect 2143 307 2281 325
rect 1913 291 2281 307
rect 1471 213 1525 229
rect 1505 179 1525 213
rect 1561 216 1574 250
rect 1608 241 1679 250
rect 1561 207 1577 216
rect 1611 207 1679 241
rect 1471 173 1525 179
rect 1631 187 1679 207
rect 1471 139 1587 173
rect 1207 93 1427 107
rect 1073 55 1103 89
rect 1137 55 1153 89
rect 1207 59 1223 93
rect 1257 59 1427 93
rect 1207 51 1427 59
rect 1471 89 1519 105
rect 1471 55 1475 89
rect 1509 55 1519 89
rect 1553 93 1587 139
rect 1631 153 1633 187
rect 1667 153 1679 187
rect 1631 127 1679 153
rect 1723 257 1792 259
rect 1723 249 2159 257
rect 1723 215 1875 249
rect 1909 215 1953 249
rect 1987 215 2031 249
rect 2065 215 2109 249
rect 2143 215 2159 249
rect 1723 164 1788 215
rect 2199 181 2281 291
rect 1723 109 1787 164
rect 1553 75 1723 93
rect 1757 75 1787 109
rect 1553 59 1787 75
rect 1827 163 1861 179
rect 1827 95 1861 129
rect 1471 17 1519 55
rect 1827 17 1861 61
rect 1895 163 2281 181
rect 1895 129 1921 163
rect 1955 147 2109 163
rect 1955 129 1971 147
rect 1895 95 1971 129
rect 2083 129 2109 147
rect 2143 147 2281 163
rect 2143 129 2159 147
rect 1895 61 1921 95
rect 1955 61 1971 95
rect 1895 51 1971 61
rect 2015 95 2049 111
rect 2015 17 2049 61
rect 2083 95 2159 129
rect 2083 61 2109 95
rect 2143 61 2159 95
rect 2083 51 2159 61
rect 2203 95 2237 111
rect 2203 17 2237 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 132 230 144 255
rect 144 230 166 255
rect 132 221 166 230
rect 223 375 257 391
rect 223 357 257 375
rect 621 357 655 391
rect 519 221 553 255
rect 1305 357 1339 391
rect 857 153 891 187
rect 929 169 951 187
rect 951 169 963 187
rect 929 153 963 169
rect 1305 239 1339 255
rect 1305 221 1331 239
rect 1331 221 1339 239
rect 1574 241 1608 250
rect 1574 216 1577 241
rect 1577 216 1608 241
rect 1633 153 1667 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
<< metal1 >>
rect 0 561 2300 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2300 561
rect 0 496 2300 527
rect 201 391 269 397
rect 201 357 223 391
rect 257 388 269 391
rect 609 391 667 397
rect 609 388 621 391
rect 257 360 621 388
rect 257 357 269 360
rect 201 351 269 357
rect 609 357 621 360
rect 655 388 667 391
rect 1293 391 1361 397
rect 1293 388 1305 391
rect 655 360 1305 388
rect 655 357 667 360
rect 609 351 667 357
rect 1293 357 1305 360
rect 1339 357 1361 391
rect 1293 351 1361 357
rect 120 255 178 261
rect 120 221 132 255
rect 166 252 178 255
rect 507 255 565 261
rect 507 252 519 255
rect 166 224 519 252
rect 166 221 178 224
rect 120 215 178 221
rect 507 221 519 224
rect 553 252 565 255
rect 1293 255 1361 261
rect 1293 252 1305 255
rect 553 224 1305 252
rect 553 221 565 224
rect 507 215 565 221
rect 1293 221 1305 224
rect 1339 221 1361 255
rect 1293 215 1361 221
rect 1562 250 1679 256
rect 1562 216 1574 250
rect 1608 216 1679 250
rect 835 187 985 193
rect 835 153 857 187
rect 891 153 929 187
rect 963 184 985 187
rect 1562 187 1679 216
rect 1562 184 1633 187
rect 963 156 1633 184
rect 963 153 985 156
rect 835 147 985 153
rect 1621 153 1633 156
rect 1667 153 1679 187
rect 1621 147 1679 153
rect 0 17 2300 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2300 17
rect 0 -48 2300 -17
<< labels >>
flabel locali s 2237 289 2271 323 0 FreeSans 400 0 0 0 Q
port 8 nsew signal output
flabel locali s 305 289 339 323 0 FreeSans 400 0 0 0 D
port 2 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 400 0 0 0 CLK
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew signal input
flabel locali s 2237 153 2271 187 0 FreeSans 400 0 0 0 Q
port 8 nsew signal output
flabel locali s 2237 221 2271 255 0 FreeSans 400 0 0 0 Q
port 8 nsew signal output
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 1593 221 1627 255 0 FreeSans 400 0 0 0 RESET_B
port 3 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 dfrtp_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2300 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 708282
string GDS_START 691504
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
