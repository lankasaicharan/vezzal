magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 8 49 761 243
rect 0 0 768 49
<< scnmos >>
rect 109 49 139 217
rect 195 49 225 217
rect 310 49 340 217
rect 382 49 412 217
rect 580 49 610 217
rect 652 49 682 217
<< scpmoshvt >>
rect 94 367 124 619
rect 180 367 210 619
rect 296 367 326 619
rect 382 367 412 619
rect 572 367 602 619
rect 658 367 688 619
<< ndiff >>
rect 34 205 109 217
rect 34 171 42 205
rect 76 171 109 205
rect 34 95 109 171
rect 34 61 42 95
rect 76 61 109 95
rect 34 49 109 61
rect 139 197 195 217
rect 139 163 150 197
rect 184 163 195 197
rect 139 101 195 163
rect 139 67 150 101
rect 184 67 195 101
rect 139 49 195 67
rect 225 165 310 217
rect 225 131 252 165
rect 286 131 310 165
rect 225 91 310 131
rect 225 57 252 91
rect 286 57 310 91
rect 225 49 310 57
rect 340 49 382 217
rect 412 205 465 217
rect 412 171 423 205
rect 457 171 465 205
rect 412 101 465 171
rect 412 67 423 101
rect 457 67 465 101
rect 412 49 465 67
rect 523 165 580 217
rect 523 131 535 165
rect 569 131 580 165
rect 523 91 580 131
rect 523 57 535 91
rect 569 57 580 91
rect 523 49 580 57
rect 610 49 652 217
rect 682 205 735 217
rect 682 171 693 205
rect 727 171 735 205
rect 682 101 735 171
rect 682 67 693 101
rect 727 67 735 101
rect 682 49 735 67
<< pdiff >>
rect 41 607 94 619
rect 41 573 49 607
rect 83 573 94 607
rect 41 529 94 573
rect 41 495 49 529
rect 83 495 94 529
rect 41 450 94 495
rect 41 416 49 450
rect 83 416 94 450
rect 41 367 94 416
rect 124 599 180 619
rect 124 565 135 599
rect 169 565 180 599
rect 124 507 180 565
rect 124 473 135 507
rect 169 473 180 507
rect 124 413 180 473
rect 124 379 135 413
rect 169 379 180 413
rect 124 367 180 379
rect 210 607 296 619
rect 210 573 236 607
rect 270 573 296 607
rect 210 514 296 573
rect 210 480 236 514
rect 270 480 296 514
rect 210 418 296 480
rect 210 384 236 418
rect 270 384 296 418
rect 210 367 296 384
rect 326 599 382 619
rect 326 565 337 599
rect 371 565 382 599
rect 326 517 382 565
rect 326 483 337 517
rect 371 483 382 517
rect 326 434 382 483
rect 326 400 337 434
rect 371 400 382 434
rect 326 367 382 400
rect 412 570 465 619
rect 412 536 423 570
rect 457 536 465 570
rect 412 367 465 536
rect 519 424 572 619
rect 519 390 527 424
rect 561 390 572 424
rect 519 367 572 390
rect 602 599 658 619
rect 602 565 613 599
rect 647 565 658 599
rect 602 514 658 565
rect 602 480 613 514
rect 647 480 658 514
rect 602 367 658 480
rect 688 599 741 619
rect 688 565 699 599
rect 733 565 741 599
rect 688 512 741 565
rect 688 478 699 512
rect 733 478 741 512
rect 688 420 741 478
rect 688 386 699 420
rect 733 386 741 420
rect 688 367 741 386
<< ndiffc >>
rect 42 171 76 205
rect 42 61 76 95
rect 150 163 184 197
rect 150 67 184 101
rect 252 131 286 165
rect 252 57 286 91
rect 423 171 457 205
rect 423 67 457 101
rect 535 131 569 165
rect 535 57 569 91
rect 693 171 727 205
rect 693 67 727 101
<< pdiffc >>
rect 49 573 83 607
rect 49 495 83 529
rect 49 416 83 450
rect 135 565 169 599
rect 135 473 169 507
rect 135 379 169 413
rect 236 573 270 607
rect 236 480 270 514
rect 236 384 270 418
rect 337 565 371 599
rect 337 483 371 517
rect 337 400 371 434
rect 423 536 457 570
rect 527 390 561 424
rect 613 565 647 599
rect 613 480 647 514
rect 699 565 733 599
rect 699 478 733 512
rect 699 386 733 420
<< poly >>
rect 94 619 124 645
rect 180 619 210 645
rect 296 619 326 645
rect 382 619 412 645
rect 572 619 602 645
rect 658 619 688 645
rect 94 279 124 367
rect 180 315 210 367
rect 296 335 326 367
rect 382 335 412 367
rect 572 335 602 367
rect 274 319 340 335
rect 166 299 232 315
rect 166 279 182 299
rect 94 265 182 279
rect 216 265 232 299
rect 274 285 290 319
rect 324 285 340 319
rect 274 269 340 285
rect 94 249 232 265
rect 109 217 139 249
rect 195 217 225 249
rect 310 217 340 269
rect 382 319 465 335
rect 382 285 415 319
rect 449 285 465 319
rect 382 269 465 285
rect 544 319 610 335
rect 544 285 560 319
rect 594 285 610 319
rect 658 325 688 367
rect 658 309 743 325
rect 658 289 693 309
rect 544 269 610 285
rect 382 217 412 269
rect 580 217 610 269
rect 652 275 693 289
rect 727 275 743 309
rect 652 259 743 275
rect 652 217 682 259
rect 109 23 139 49
rect 195 23 225 49
rect 310 23 340 49
rect 382 23 412 49
rect 580 23 610 49
rect 652 23 682 49
<< polycont >>
rect 182 265 216 299
rect 290 285 324 319
rect 415 285 449 319
rect 560 285 594 319
rect 693 275 727 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 33 607 83 649
rect 33 573 49 607
rect 33 529 83 573
rect 33 495 49 529
rect 33 450 83 495
rect 33 416 49 450
rect 33 400 83 416
rect 121 599 186 615
rect 121 565 135 599
rect 169 565 186 599
rect 121 507 186 565
rect 121 473 135 507
rect 169 473 186 507
rect 121 413 186 473
rect 121 385 135 413
rect 114 379 135 385
rect 169 379 186 413
rect 220 607 286 649
rect 220 573 236 607
rect 270 573 286 607
rect 220 514 286 573
rect 220 480 236 514
rect 270 480 286 514
rect 220 418 286 480
rect 220 384 236 418
rect 270 384 286 418
rect 321 599 373 615
rect 321 565 337 599
rect 371 565 373 599
rect 321 517 373 565
rect 407 570 473 649
rect 407 536 423 570
rect 457 536 473 570
rect 407 530 473 536
rect 597 599 663 615
rect 597 565 613 599
rect 647 565 663 599
rect 321 483 337 517
rect 371 496 373 517
rect 597 514 663 565
rect 597 496 613 514
rect 371 483 613 496
rect 321 480 613 483
rect 647 480 663 514
rect 321 462 663 480
rect 697 599 749 615
rect 697 565 699 599
rect 733 565 749 599
rect 697 512 749 565
rect 697 478 699 512
rect 733 478 749 512
rect 321 434 377 462
rect 321 400 337 434
rect 371 400 377 434
rect 697 428 749 478
rect 321 384 377 400
rect 114 351 186 379
rect 26 205 80 221
rect 26 171 42 205
rect 76 171 80 205
rect 26 95 80 171
rect 26 61 42 95
rect 76 61 80 95
rect 26 17 80 61
rect 114 213 148 351
rect 290 319 377 350
rect 182 299 256 317
rect 216 265 256 299
rect 324 285 377 319
rect 290 269 377 285
rect 411 319 449 428
rect 411 285 415 319
rect 411 269 449 285
rect 490 424 749 428
rect 490 390 527 424
rect 561 420 749 424
rect 561 390 699 420
rect 490 386 699 390
rect 733 386 749 420
rect 182 249 256 265
rect 222 233 256 249
rect 490 233 524 386
rect 558 319 641 350
rect 558 285 560 319
rect 594 285 641 319
rect 558 269 641 285
rect 677 309 749 350
rect 677 275 693 309
rect 727 275 749 309
rect 114 197 188 213
rect 222 205 743 233
rect 222 199 423 205
rect 114 163 150 197
rect 184 163 188 197
rect 407 171 423 199
rect 457 199 693 205
rect 457 171 473 199
rect 114 101 188 163
rect 114 67 150 101
rect 184 67 188 101
rect 114 51 188 67
rect 236 131 252 165
rect 286 131 302 165
rect 236 91 302 131
rect 236 57 252 91
rect 286 57 302 91
rect 236 17 302 57
rect 407 101 473 171
rect 677 171 693 199
rect 727 171 743 205
rect 407 67 423 101
rect 457 67 473 101
rect 407 51 473 67
rect 519 131 535 165
rect 569 131 585 165
rect 519 91 585 131
rect 519 57 535 91
rect 569 57 585 91
rect 519 17 585 57
rect 677 101 743 171
rect 677 67 693 101
rect 727 67 743 101
rect 677 51 743 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a22o_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1146464
string GDS_START 1139138
<< end >>
