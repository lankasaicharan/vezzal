magic
tech sky130A
magscale 1 2
timestamp 1627202617
<< checkpaint >>
rect -1298 -1308 3230 1852
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1931 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1191 47 1221 177
rect 1275 47 1305 177
rect 1359 47 1389 177
rect 1443 47 1473 177
rect 1571 47 1601 177
rect 1655 47 1685 177
rect 1739 47 1769 177
rect 1823 47 1853 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 751 297 781 497
rect 835 297 865 497
rect 919 297 949 497
rect 1003 297 1033 497
rect 1191 297 1221 497
rect 1275 297 1305 497
rect 1359 297 1389 497
rect 1443 297 1473 497
rect 1571 297 1601 497
rect 1655 297 1685 497
rect 1739 297 1769 497
rect 1823 297 1853 497
<< ndiff >>
rect 27 101 79 177
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 101 247 177
rect 193 67 203 101
rect 237 67 247 101
rect 193 47 247 67
rect 277 93 331 177
rect 277 59 287 93
rect 321 59 331 93
rect 277 47 331 59
rect 361 101 415 177
rect 361 67 371 101
rect 405 67 415 101
rect 361 47 415 67
rect 445 93 499 177
rect 445 59 455 93
rect 489 59 499 93
rect 445 47 499 59
rect 529 161 583 177
rect 529 127 539 161
rect 573 127 583 161
rect 529 47 583 127
rect 613 93 667 177
rect 613 59 623 93
rect 657 59 667 93
rect 613 47 667 59
rect 697 161 749 177
rect 697 127 707 161
rect 741 127 749 161
rect 697 47 749 127
rect 803 161 855 177
rect 803 127 811 161
rect 845 127 855 161
rect 803 47 855 127
rect 885 93 939 177
rect 885 59 895 93
rect 929 59 939 93
rect 885 47 939 59
rect 969 161 1023 177
rect 969 127 979 161
rect 1013 127 1023 161
rect 969 47 1023 127
rect 1053 93 1107 177
rect 1053 59 1063 93
rect 1097 59 1107 93
rect 1053 47 1107 59
rect 1137 161 1191 177
rect 1137 127 1147 161
rect 1181 127 1191 161
rect 1137 47 1191 127
rect 1221 93 1275 177
rect 1221 59 1231 93
rect 1265 59 1275 93
rect 1221 47 1275 59
rect 1305 101 1359 177
rect 1305 67 1315 101
rect 1349 67 1359 101
rect 1305 47 1359 67
rect 1389 93 1443 177
rect 1389 59 1399 93
rect 1433 59 1443 93
rect 1389 47 1443 59
rect 1473 101 1571 177
rect 1473 67 1483 101
rect 1517 67 1571 101
rect 1473 47 1571 67
rect 1601 93 1655 177
rect 1601 59 1611 93
rect 1645 59 1655 93
rect 1601 47 1655 59
rect 1685 101 1739 177
rect 1685 67 1695 101
rect 1729 67 1739 101
rect 1685 47 1739 67
rect 1769 93 1823 177
rect 1769 59 1779 93
rect 1813 59 1823 93
rect 1769 47 1823 59
rect 1853 101 1905 177
rect 1853 67 1863 101
rect 1897 67 1905 101
rect 1853 47 1905 67
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 477 331 497
rect 277 443 287 477
rect 321 443 331 477
rect 277 409 331 443
rect 277 375 287 409
rect 321 375 331 409
rect 277 297 331 375
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 417 415 451
rect 361 383 371 417
rect 405 383 415 417
rect 361 297 415 383
rect 445 477 499 497
rect 445 443 455 477
rect 489 443 499 477
rect 445 409 499 443
rect 445 375 455 409
rect 489 375 499 409
rect 445 297 499 375
rect 529 485 583 497
rect 529 451 539 485
rect 573 451 583 485
rect 529 417 583 451
rect 529 383 539 417
rect 573 383 583 417
rect 529 297 583 383
rect 613 477 667 497
rect 613 443 623 477
rect 657 443 667 477
rect 613 409 667 443
rect 613 375 623 409
rect 657 375 667 409
rect 613 297 667 375
rect 697 485 751 497
rect 697 451 707 485
rect 741 451 751 485
rect 697 417 751 451
rect 697 383 707 417
rect 741 383 751 417
rect 697 297 751 383
rect 781 477 835 497
rect 781 443 791 477
rect 825 443 835 477
rect 781 409 835 443
rect 781 375 791 409
rect 825 375 835 409
rect 781 297 835 375
rect 865 485 919 497
rect 865 451 875 485
rect 909 451 919 485
rect 865 417 919 451
rect 865 383 875 417
rect 909 383 919 417
rect 865 297 919 383
rect 949 477 1003 497
rect 949 443 959 477
rect 993 443 1003 477
rect 949 409 1003 443
rect 949 375 959 409
rect 993 375 1003 409
rect 949 297 1003 375
rect 1033 485 1085 497
rect 1033 451 1043 485
rect 1077 451 1085 485
rect 1033 297 1085 451
rect 1139 485 1191 497
rect 1139 451 1147 485
rect 1181 451 1191 485
rect 1139 297 1191 451
rect 1221 417 1275 497
rect 1221 383 1231 417
rect 1265 383 1275 417
rect 1221 297 1275 383
rect 1305 485 1359 497
rect 1305 451 1315 485
rect 1349 451 1359 485
rect 1305 297 1359 451
rect 1389 417 1443 497
rect 1389 383 1399 417
rect 1433 383 1443 417
rect 1389 297 1443 383
rect 1473 485 1571 497
rect 1473 451 1483 485
rect 1517 451 1571 485
rect 1473 297 1571 451
rect 1601 417 1655 497
rect 1601 383 1611 417
rect 1645 383 1655 417
rect 1601 343 1655 383
rect 1601 309 1611 343
rect 1645 309 1655 343
rect 1601 297 1655 309
rect 1685 485 1739 497
rect 1685 451 1695 485
rect 1729 451 1739 485
rect 1685 297 1739 451
rect 1769 417 1823 497
rect 1769 383 1779 417
rect 1813 383 1823 417
rect 1769 343 1823 383
rect 1769 309 1779 343
rect 1813 309 1823 343
rect 1769 297 1823 309
rect 1853 485 1905 497
rect 1853 451 1863 485
rect 1897 451 1905 485
rect 1853 417 1905 451
rect 1853 383 1863 417
rect 1897 383 1905 417
rect 1853 297 1905 383
<< ndiffc >>
rect 35 67 69 101
rect 119 59 153 93
rect 203 67 237 101
rect 287 59 321 93
rect 371 67 405 101
rect 455 59 489 93
rect 539 127 573 161
rect 623 59 657 93
rect 707 127 741 161
rect 811 127 845 161
rect 895 59 929 93
rect 979 127 1013 161
rect 1063 59 1097 93
rect 1147 127 1181 161
rect 1231 59 1265 93
rect 1315 67 1349 101
rect 1399 59 1433 93
rect 1483 67 1517 101
rect 1611 59 1645 93
rect 1695 67 1729 101
rect 1779 59 1813 93
rect 1863 67 1897 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 443 153 477
rect 119 375 153 409
rect 203 451 237 485
rect 203 383 237 417
rect 287 443 321 477
rect 287 375 321 409
rect 371 451 405 485
rect 371 383 405 417
rect 455 443 489 477
rect 455 375 489 409
rect 539 451 573 485
rect 539 383 573 417
rect 623 443 657 477
rect 623 375 657 409
rect 707 451 741 485
rect 707 383 741 417
rect 791 443 825 477
rect 791 375 825 409
rect 875 451 909 485
rect 875 383 909 417
rect 959 443 993 477
rect 959 375 993 409
rect 1043 451 1077 485
rect 1147 451 1181 485
rect 1231 383 1265 417
rect 1315 451 1349 485
rect 1399 383 1433 417
rect 1483 451 1517 485
rect 1611 383 1645 417
rect 1611 309 1645 343
rect 1695 451 1729 485
rect 1779 383 1813 417
rect 1779 309 1813 343
rect 1863 451 1897 485
rect 1863 383 1897 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 751 497 781 523
rect 835 497 865 523
rect 919 497 949 523
rect 1003 497 1033 523
rect 1191 497 1221 523
rect 1275 497 1305 523
rect 1359 497 1389 523
rect 1443 497 1473 523
rect 1571 497 1601 523
rect 1655 497 1685 523
rect 1739 497 1769 523
rect 1823 497 1853 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 22 249 361 265
rect 22 215 40 249
rect 74 215 114 249
rect 148 215 188 249
rect 222 215 262 249
rect 296 215 361 249
rect 22 199 361 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 265 445 297
rect 499 265 529 297
rect 583 265 613 297
rect 667 265 697 297
rect 415 249 697 265
rect 415 215 425 249
rect 459 215 499 249
rect 533 215 573 249
rect 607 215 647 249
rect 681 215 697 249
rect 415 199 697 215
rect 751 269 781 297
rect 835 269 865 297
rect 919 269 949 297
rect 1003 269 1033 297
rect 751 265 1033 269
rect 1191 265 1221 297
rect 1275 265 1305 297
rect 1359 265 1389 297
rect 1443 265 1473 297
rect 751 249 1137 265
rect 751 215 761 249
rect 795 215 835 249
rect 869 215 909 249
rect 943 215 983 249
rect 1017 215 1137 249
rect 751 199 1137 215
rect 1179 249 1473 265
rect 1179 215 1189 249
rect 1223 215 1263 249
rect 1297 215 1337 249
rect 1371 215 1473 249
rect 1179 199 1473 215
rect 415 177 445 199
rect 499 177 529 199
rect 583 177 613 199
rect 667 177 697 199
rect 855 177 885 199
rect 939 177 969 199
rect 1023 177 1053 199
rect 1107 177 1137 199
rect 1191 177 1221 199
rect 1275 177 1305 199
rect 1359 177 1389 199
rect 1443 177 1473 199
rect 1571 265 1601 297
rect 1655 265 1685 297
rect 1739 265 1769 297
rect 1823 265 1853 297
rect 1571 249 1910 265
rect 1571 215 1644 249
rect 1678 215 1718 249
rect 1752 215 1792 249
rect 1826 215 1866 249
rect 1900 215 1910 249
rect 1571 199 1910 215
rect 1571 177 1601 199
rect 1655 177 1685 199
rect 1739 177 1769 199
rect 1823 177 1853 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1191 21 1221 47
rect 1275 21 1305 47
rect 1359 21 1389 47
rect 1443 21 1473 47
rect 1571 21 1601 47
rect 1655 21 1685 47
rect 1739 21 1769 47
rect 1823 21 1853 47
<< polycont >>
rect 40 215 74 249
rect 114 215 148 249
rect 188 215 222 249
rect 262 215 296 249
rect 425 215 459 249
rect 499 215 533 249
rect 573 215 607 249
rect 647 215 681 249
rect 761 215 795 249
rect 835 215 869 249
rect 909 215 943 249
rect 983 215 1017 249
rect 1189 215 1223 249
rect 1263 215 1297 249
rect 1337 215 1371 249
rect 1644 215 1678 249
rect 1718 215 1752 249
rect 1792 215 1826 249
rect 1866 215 1900 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 19 485 85 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 19 349 85 383
rect 19 315 35 349
rect 69 315 85 349
rect 119 477 153 493
rect 119 409 153 443
rect 187 485 253 527
rect 187 451 203 485
rect 237 451 253 485
rect 187 417 253 451
rect 187 383 203 417
rect 237 383 253 417
rect 287 477 321 493
rect 287 409 321 443
rect 119 333 153 375
rect 355 485 421 527
rect 355 451 371 485
rect 405 451 421 485
rect 355 417 421 451
rect 355 383 371 417
rect 405 383 421 417
rect 455 477 489 493
rect 455 409 489 443
rect 287 333 321 375
rect 523 485 589 527
rect 523 451 539 485
rect 573 451 589 485
rect 523 417 589 451
rect 523 383 539 417
rect 573 383 589 417
rect 623 477 657 493
rect 623 409 657 443
rect 455 333 489 375
rect 691 485 757 527
rect 691 451 707 485
rect 741 451 757 485
rect 691 417 757 451
rect 691 383 707 417
rect 741 383 757 417
rect 791 477 825 493
rect 791 409 825 443
rect 623 333 657 375
rect 859 485 925 527
rect 859 451 875 485
rect 909 451 925 485
rect 859 417 925 451
rect 859 383 875 417
rect 909 383 925 417
rect 959 477 993 493
rect 1027 485 1093 527
rect 1027 451 1043 485
rect 1077 451 1093 485
rect 1131 451 1147 485
rect 1181 451 1315 485
rect 1349 451 1483 485
rect 1517 451 1695 485
rect 1729 451 1863 485
rect 1897 451 1913 485
rect 959 417 993 443
rect 1863 417 1913 451
rect 959 409 1231 417
rect 791 333 825 375
rect 993 383 1231 409
rect 1265 383 1399 417
rect 1433 383 1449 417
rect 959 333 993 375
rect 119 299 993 333
rect 1483 343 1547 395
rect 1595 383 1611 417
rect 1645 383 1661 417
rect 1595 343 1661 383
rect 1763 383 1779 417
rect 1813 383 1829 417
rect 1763 343 1829 383
rect 1897 383 1913 417
rect 1863 367 1913 383
rect 24 249 347 265
rect 24 215 40 249
rect 74 215 114 249
rect 148 215 188 249
rect 222 215 262 249
rect 296 215 347 249
rect 24 199 347 215
rect 387 249 710 265
rect 387 215 425 249
rect 459 215 499 249
rect 533 215 573 249
rect 607 215 647 249
rect 681 215 710 249
rect 387 199 710 215
rect 761 249 1084 265
rect 795 215 835 249
rect 869 215 909 249
rect 943 215 983 249
rect 1017 215 1084 249
rect 761 199 1084 215
rect 1134 249 1371 326
rect 1134 215 1189 249
rect 1223 215 1263 249
rect 1297 215 1337 249
rect 1134 199 1371 215
rect 1483 309 1611 343
rect 1645 309 1779 343
rect 1813 309 1829 343
rect 1483 161 1547 309
rect 1595 306 1661 309
rect 1587 249 1906 265
rect 1587 215 1644 249
rect 1678 215 1718 249
rect 1752 215 1792 249
rect 1826 215 1866 249
rect 1900 215 1906 249
rect 1587 199 1906 215
rect 35 127 539 161
rect 573 127 707 161
rect 741 127 757 161
rect 795 127 811 161
rect 845 127 979 161
rect 1013 127 1147 161
rect 1181 127 1897 161
rect 35 101 69 127
rect 203 101 237 127
rect 35 51 69 67
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 371 101 405 127
rect 203 51 237 67
rect 271 59 287 93
rect 321 59 337 93
rect 271 17 337 59
rect 1315 101 1349 127
rect 371 51 405 67
rect 439 59 455 93
rect 489 59 623 93
rect 657 59 895 93
rect 929 59 1063 93
rect 1097 59 1113 93
rect 1215 59 1231 93
rect 1265 59 1281 93
rect 1215 17 1281 59
rect 1483 101 1517 127
rect 1315 51 1349 67
rect 1383 59 1399 93
rect 1433 59 1449 93
rect 1383 17 1449 59
rect 1695 101 1729 127
rect 1483 51 1517 67
rect 1595 59 1611 93
rect 1645 59 1661 93
rect 1595 17 1661 59
rect 1863 101 1897 127
rect 1695 51 1729 67
rect 1763 59 1779 93
rect 1813 59 1829 93
rect 1763 17 1829 59
rect 1863 51 1897 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 1506 153 1540 187 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1138 289 1172 323 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 766 221 800 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1506 221 1540 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1506 357 1540 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1506 289 1540 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1592 221 1626 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 1684 221 1718 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 1776 221 1810 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 1868 221 1902 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 1138 221 1172 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1322 289 1356 323 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1230 289 1264 323 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1322 221 1356 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1230 221 1264 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1042 221 1076 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 950 221 984 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 858 221 892 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 a311oi_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 1679658
string GDS_START 1664112
string path 0.000 0.000 48.300 0.000 
<< end >>
