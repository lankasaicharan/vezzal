magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 195 241 671 243
rect 5 49 671 241
rect 0 0 672 49
<< scnmos >>
rect 84 47 114 215
rect 274 49 304 217
rect 382 49 412 217
rect 468 49 498 217
rect 562 49 592 217
<< scpmoshvt >>
rect 120 367 150 619
rect 274 367 304 619
rect 346 367 376 619
rect 490 367 520 619
rect 562 367 592 619
<< ndiff >>
rect 31 203 84 215
rect 31 169 39 203
rect 73 169 84 203
rect 31 101 84 169
rect 31 67 39 101
rect 73 67 84 101
rect 31 47 84 67
rect 114 161 167 215
rect 114 127 125 161
rect 159 127 167 161
rect 114 93 167 127
rect 114 59 125 93
rect 159 59 167 93
rect 114 47 167 59
rect 221 169 274 217
rect 221 135 229 169
rect 263 135 274 169
rect 221 49 274 135
rect 304 159 382 217
rect 304 125 326 159
rect 360 125 382 159
rect 304 91 382 125
rect 304 57 326 91
rect 360 57 382 91
rect 304 49 382 57
rect 412 205 468 217
rect 412 171 423 205
rect 457 171 468 205
rect 412 101 468 171
rect 412 67 423 101
rect 457 67 468 101
rect 412 49 468 67
rect 498 159 562 217
rect 498 125 515 159
rect 549 125 562 159
rect 498 91 562 125
rect 498 57 515 91
rect 549 57 562 91
rect 498 49 562 57
rect 592 205 645 217
rect 592 171 603 205
rect 637 171 645 205
rect 592 101 645 171
rect 592 67 603 101
rect 637 67 645 101
rect 592 49 645 67
<< pdiff >>
rect 67 599 120 619
rect 67 565 75 599
rect 109 565 120 599
rect 67 513 120 565
rect 67 479 75 513
rect 109 479 120 513
rect 67 420 120 479
rect 67 386 75 420
rect 109 386 120 420
rect 67 367 120 386
rect 150 607 274 619
rect 150 573 161 607
rect 195 573 229 607
rect 263 573 274 607
rect 150 497 274 573
rect 150 463 161 497
rect 195 463 229 497
rect 263 463 274 497
rect 150 367 274 463
rect 304 367 346 619
rect 376 599 490 619
rect 376 565 414 599
rect 448 565 490 599
rect 376 513 490 565
rect 376 479 414 513
rect 448 479 490 513
rect 376 424 490 479
rect 376 390 414 424
rect 448 390 490 424
rect 376 367 490 390
rect 520 367 562 619
rect 592 607 645 619
rect 592 573 603 607
rect 637 573 645 607
rect 592 512 645 573
rect 592 478 603 512
rect 637 478 645 512
rect 592 418 645 478
rect 592 384 603 418
rect 637 384 645 418
rect 592 367 645 384
<< ndiffc >>
rect 39 169 73 203
rect 39 67 73 101
rect 125 127 159 161
rect 125 59 159 93
rect 229 135 263 169
rect 326 125 360 159
rect 326 57 360 91
rect 423 171 457 205
rect 423 67 457 101
rect 515 125 549 159
rect 515 57 549 91
rect 603 171 637 205
rect 603 67 637 101
<< pdiffc >>
rect 75 565 109 599
rect 75 479 109 513
rect 75 386 109 420
rect 161 573 195 607
rect 229 573 263 607
rect 161 463 195 497
rect 229 463 263 497
rect 414 565 448 599
rect 414 479 448 513
rect 414 390 448 424
rect 603 573 637 607
rect 603 478 637 512
rect 603 384 637 418
<< poly >>
rect 120 619 150 645
rect 274 619 304 645
rect 346 619 376 645
rect 490 619 520 645
rect 562 619 592 645
rect 120 325 150 367
rect 274 335 304 367
rect 25 309 150 325
rect 25 275 41 309
rect 75 295 150 309
rect 217 319 304 335
rect 75 275 114 295
rect 25 259 114 275
rect 217 285 233 319
rect 267 285 304 319
rect 217 269 304 285
rect 346 335 376 367
rect 490 335 520 367
rect 346 319 412 335
rect 346 285 362 319
rect 396 285 412 319
rect 346 269 412 285
rect 454 319 520 335
rect 454 285 470 319
rect 504 285 520 319
rect 454 269 520 285
rect 562 325 592 367
rect 562 309 647 325
rect 562 275 597 309
rect 631 275 647 309
rect 84 215 114 259
rect 274 217 304 269
rect 382 217 412 269
rect 468 217 498 269
rect 562 259 647 275
rect 562 217 592 259
rect 84 21 114 47
rect 274 23 304 49
rect 382 23 412 49
rect 468 23 498 49
rect 562 23 592 49
<< polycont >>
rect 41 275 75 309
rect 233 285 267 319
rect 362 285 396 319
rect 470 285 504 319
rect 597 275 631 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 59 599 111 615
rect 59 565 75 599
rect 109 565 111 599
rect 59 513 111 565
rect 59 479 75 513
rect 109 479 111 513
rect 59 424 111 479
rect 145 607 279 649
rect 145 573 161 607
rect 195 573 229 607
rect 263 573 279 607
rect 145 497 279 573
rect 145 463 161 497
rect 195 463 229 497
rect 263 463 279 497
rect 145 458 279 463
rect 398 599 464 615
rect 398 565 414 599
rect 448 565 464 599
rect 587 607 653 649
rect 398 513 464 565
rect 398 479 414 513
rect 448 479 464 513
rect 398 424 464 479
rect 59 420 414 424
rect 59 386 75 420
rect 109 390 414 420
rect 448 390 464 424
rect 109 386 177 390
rect 25 309 91 352
rect 25 275 41 309
rect 75 275 91 309
rect 25 269 91 275
rect 125 235 177 386
rect 211 319 275 356
rect 211 285 233 319
rect 267 285 275 319
rect 211 269 275 285
rect 309 319 412 355
rect 498 335 547 592
rect 587 573 603 607
rect 637 573 653 607
rect 587 512 653 573
rect 587 478 603 512
rect 637 478 653 512
rect 587 418 653 478
rect 587 384 603 418
rect 637 384 653 418
rect 309 285 362 319
rect 396 285 412 319
rect 309 269 412 285
rect 454 319 547 335
rect 454 285 470 319
rect 504 285 547 319
rect 454 269 547 285
rect 581 309 655 350
rect 581 275 597 309
rect 631 275 655 309
rect 581 269 655 275
rect 23 203 177 235
rect 23 169 39 203
rect 73 201 177 203
rect 213 205 653 235
rect 73 169 75 201
rect 23 101 75 169
rect 213 199 423 205
rect 213 169 276 199
rect 23 67 39 101
rect 73 67 75 101
rect 23 51 75 67
rect 109 161 175 167
rect 109 127 125 161
rect 159 127 175 161
rect 109 93 175 127
rect 213 135 229 169
rect 263 135 276 169
rect 410 171 423 199
rect 457 201 603 205
rect 457 171 465 201
rect 213 119 276 135
rect 310 159 376 163
rect 310 125 326 159
rect 360 125 376 159
rect 109 59 125 93
rect 159 85 175 93
rect 310 91 376 125
rect 310 85 326 91
rect 159 59 326 85
rect 109 57 326 59
rect 360 57 376 91
rect 109 51 376 57
rect 410 101 465 171
rect 599 171 603 201
rect 637 171 653 205
rect 410 67 423 101
rect 457 67 465 101
rect 410 51 465 67
rect 499 159 565 167
rect 499 125 515 159
rect 549 125 565 159
rect 499 91 565 125
rect 499 57 515 91
rect 549 57 565 91
rect 499 17 565 57
rect 599 101 653 171
rect 599 67 603 101
rect 637 67 653 101
rect 599 51 653 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221ai_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5840662
string GDS_START 5833282
<< end >>
