magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 332 1958 704
<< pwell >>
rect 1 229 333 248
rect 1356 234 1914 248
rect 1 212 716 229
rect 955 212 1914 234
rect 1 49 1914 212
rect 0 0 1920 49
<< scnmos >>
rect 84 74 114 222
rect 209 74 239 222
rect 524 119 554 203
rect 610 119 640 203
rect 705 102 735 186
rect 777 102 807 186
rect 936 76 966 186
rect 1031 98 1061 208
rect 1148 124 1178 208
rect 1241 124 1271 208
rect 1439 74 1469 222
rect 1531 74 1561 222
rect 1625 74 1655 222
rect 1715 74 1745 222
rect 1801 74 1831 222
<< scpmoshvt >>
rect 86 368 116 592
rect 176 368 206 592
rect 407 503 437 587
rect 514 485 544 569
rect 621 503 651 587
rect 699 503 729 587
rect 868 424 898 592
rect 1004 424 1034 592
rect 1111 508 1141 592
rect 1236 508 1266 592
rect 1337 424 1367 592
rect 1427 424 1457 592
rect 1534 368 1564 592
rect 1624 368 1654 592
rect 1714 368 1744 592
rect 1804 368 1834 592
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 131 209 222
rect 114 97 125 131
rect 159 97 209 131
rect 114 74 209 97
rect 239 189 307 222
rect 239 155 261 189
rect 295 155 307 189
rect 239 74 307 155
rect 401 119 524 203
rect 554 180 610 203
rect 554 146 565 180
rect 599 146 610 180
rect 554 119 610 146
rect 640 186 690 203
rect 981 186 1031 208
rect 640 174 705 186
rect 640 140 654 174
rect 688 140 705 174
rect 640 119 705 140
rect 401 112 474 119
rect 401 78 413 112
rect 447 78 474 112
rect 655 102 705 119
rect 735 102 777 186
rect 807 102 936 186
rect 401 66 474 78
rect 822 88 936 102
rect 822 54 834 88
rect 868 76 936 88
rect 966 171 1031 186
rect 966 137 986 171
rect 1020 137 1031 171
rect 966 98 1031 137
rect 1061 178 1148 208
rect 1061 144 1094 178
rect 1128 144 1148 178
rect 1061 124 1148 144
rect 1178 124 1241 208
rect 1271 174 1328 208
rect 1271 140 1282 174
rect 1316 140 1328 174
rect 1271 124 1328 140
rect 1382 194 1439 222
rect 1382 160 1394 194
rect 1428 160 1439 194
rect 1061 98 1111 124
rect 966 76 1016 98
rect 868 54 880 76
rect 822 42 880 54
rect 1382 120 1439 160
rect 1382 86 1394 120
rect 1428 86 1439 120
rect 1382 74 1439 86
rect 1469 123 1531 222
rect 1469 89 1480 123
rect 1514 89 1531 123
rect 1469 74 1531 89
rect 1561 210 1625 222
rect 1561 176 1580 210
rect 1614 176 1625 210
rect 1561 120 1625 176
rect 1561 86 1580 120
rect 1614 86 1625 120
rect 1561 74 1625 86
rect 1655 131 1715 222
rect 1655 97 1666 131
rect 1700 97 1715 131
rect 1655 74 1715 97
rect 1745 210 1801 222
rect 1745 176 1756 210
rect 1790 176 1801 210
rect 1745 120 1801 176
rect 1745 86 1756 120
rect 1790 86 1801 120
rect 1745 74 1801 86
rect 1831 210 1888 222
rect 1831 176 1842 210
rect 1876 176 1888 210
rect 1831 120 1888 176
rect 1831 86 1842 120
rect 1876 86 1888 120
rect 1831 74 1888 86
<< pdiff >>
rect 319 623 377 635
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 510 86 546
rect 27 476 39 510
rect 73 476 86 510
rect 27 440 86 476
rect 27 406 39 440
rect 73 406 86 440
rect 27 368 86 406
rect 116 580 176 592
rect 116 546 129 580
rect 163 546 176 580
rect 116 508 176 546
rect 116 474 129 508
rect 163 474 176 508
rect 116 368 176 474
rect 206 580 265 592
rect 206 546 219 580
rect 253 546 265 580
rect 206 497 265 546
rect 319 589 331 623
rect 365 589 377 623
rect 747 620 815 632
rect 319 587 377 589
rect 319 503 407 587
rect 437 569 490 587
rect 747 587 759 620
rect 568 569 621 587
rect 437 531 514 569
rect 437 503 467 531
rect 206 463 219 497
rect 253 463 265 497
rect 455 497 467 503
rect 501 497 514 531
rect 455 485 514 497
rect 544 547 621 569
rect 544 513 557 547
rect 591 513 621 547
rect 544 503 621 513
rect 651 503 699 587
rect 729 586 759 587
rect 793 592 815 620
rect 793 586 868 592
rect 729 503 868 586
rect 544 485 603 503
rect 206 414 265 463
rect 206 380 219 414
rect 253 380 265 414
rect 206 368 265 380
rect 815 424 868 503
rect 898 509 1004 592
rect 898 475 911 509
rect 945 475 1004 509
rect 898 424 1004 475
rect 1034 509 1111 592
rect 1034 475 1047 509
rect 1081 508 1111 509
rect 1141 508 1236 592
rect 1266 550 1337 592
rect 1266 516 1280 550
rect 1314 516 1337 550
rect 1266 508 1337 516
rect 1081 475 1093 508
rect 1034 424 1093 475
rect 1284 424 1337 508
rect 1367 580 1427 592
rect 1367 546 1380 580
rect 1414 546 1427 580
rect 1367 470 1427 546
rect 1367 436 1380 470
rect 1414 436 1427 470
rect 1367 424 1427 436
rect 1457 580 1534 592
rect 1457 546 1487 580
rect 1521 546 1534 580
rect 1457 462 1534 546
rect 1457 428 1487 462
rect 1521 428 1534 462
rect 1457 424 1534 428
rect 1475 368 1534 424
rect 1564 580 1624 592
rect 1564 546 1577 580
rect 1611 546 1624 580
rect 1564 497 1624 546
rect 1564 463 1577 497
rect 1611 463 1624 497
rect 1564 414 1624 463
rect 1564 380 1577 414
rect 1611 380 1624 414
rect 1564 368 1624 380
rect 1654 580 1714 592
rect 1654 546 1667 580
rect 1701 546 1714 580
rect 1654 478 1714 546
rect 1654 444 1667 478
rect 1701 444 1714 478
rect 1654 368 1714 444
rect 1744 580 1804 592
rect 1744 546 1757 580
rect 1791 546 1804 580
rect 1744 497 1804 546
rect 1744 463 1757 497
rect 1791 463 1804 497
rect 1744 414 1804 463
rect 1744 380 1757 414
rect 1791 380 1804 414
rect 1744 368 1804 380
rect 1834 580 1893 592
rect 1834 546 1847 580
rect 1881 546 1893 580
rect 1834 497 1893 546
rect 1834 463 1847 497
rect 1881 463 1893 497
rect 1834 414 1893 463
rect 1834 380 1847 414
rect 1881 380 1893 414
rect 1834 368 1893 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 97 159 131
rect 261 155 295 189
rect 565 146 599 180
rect 654 140 688 174
rect 413 78 447 112
rect 834 54 868 88
rect 986 137 1020 171
rect 1094 144 1128 178
rect 1282 140 1316 174
rect 1394 160 1428 194
rect 1394 86 1428 120
rect 1480 89 1514 123
rect 1580 176 1614 210
rect 1580 86 1614 120
rect 1666 97 1700 131
rect 1756 176 1790 210
rect 1756 86 1790 120
rect 1842 176 1876 210
rect 1842 86 1876 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 129 546 163 580
rect 129 474 163 508
rect 219 546 253 580
rect 331 589 365 623
rect 219 463 253 497
rect 467 497 501 531
rect 557 513 591 547
rect 759 586 793 620
rect 219 380 253 414
rect 911 475 945 509
rect 1047 475 1081 509
rect 1280 516 1314 550
rect 1380 546 1414 580
rect 1380 436 1414 470
rect 1487 546 1521 580
rect 1487 428 1521 462
rect 1577 546 1611 580
rect 1577 463 1611 497
rect 1577 380 1611 414
rect 1667 546 1701 580
rect 1667 444 1701 478
rect 1757 546 1791 580
rect 1757 463 1791 497
rect 1757 380 1791 414
rect 1847 546 1881 580
rect 1847 463 1881 497
rect 1847 380 1881 414
<< poly >>
rect 86 592 116 618
rect 176 592 206 618
rect 407 587 437 613
rect 514 569 544 595
rect 621 587 651 613
rect 699 587 729 613
rect 407 488 437 503
rect 404 471 440 488
rect 868 592 898 618
rect 1004 592 1034 618
rect 1111 592 1141 618
rect 1236 592 1266 618
rect 1337 592 1367 618
rect 1427 592 1457 618
rect 1534 592 1564 618
rect 1624 592 1654 618
rect 1714 592 1744 618
rect 1804 592 1834 618
rect 621 488 651 503
rect 699 488 729 503
rect 357 455 440 471
rect 514 470 544 485
rect 357 421 373 455
rect 407 421 440 455
rect 357 405 440 421
rect 511 369 547 470
rect 86 353 116 368
rect 176 353 206 368
rect 488 363 547 369
rect 83 326 119 353
rect 35 310 119 326
rect 173 310 209 353
rect 323 339 547 363
rect 618 416 654 488
rect 696 458 769 488
rect 618 400 697 416
rect 618 366 647 400
rect 681 366 697 400
rect 618 350 697 366
rect 323 333 518 339
rect 323 310 353 333
rect 35 276 51 310
rect 85 276 119 310
rect 35 260 119 276
rect 161 294 239 310
rect 161 260 177 294
rect 211 260 239 294
rect 84 222 114 260
rect 161 244 239 260
rect 287 294 353 310
rect 287 260 303 294
rect 337 260 353 294
rect 287 244 353 260
rect 209 222 239 244
rect 84 48 114 74
rect 209 48 239 74
rect 323 51 353 244
rect 395 275 461 291
rect 395 241 411 275
rect 445 255 461 275
rect 445 241 554 255
rect 618 248 648 350
rect 739 284 769 458
rect 1111 493 1141 508
rect 1236 493 1266 508
rect 1108 476 1144 493
rect 1108 460 1191 476
rect 1108 426 1141 460
rect 1175 426 1191 460
rect 868 409 898 424
rect 1004 409 1034 424
rect 1108 410 1191 426
rect 865 392 901 409
rect 811 376 953 392
rect 811 342 827 376
rect 861 342 953 376
rect 1001 368 1037 409
rect 1001 344 1178 368
rect 1233 362 1269 493
rect 1337 409 1367 424
rect 1427 409 1457 424
rect 1334 379 1460 409
rect 811 326 953 342
rect 1007 338 1178 344
rect 923 290 953 326
rect 739 274 807 284
rect 739 258 875 274
rect 923 260 966 290
rect 739 254 825 258
rect 395 225 554 241
rect 524 203 554 225
rect 610 218 648 248
rect 777 224 825 254
rect 859 224 875 258
rect 610 203 640 218
rect 705 186 735 212
rect 777 208 875 224
rect 777 186 807 208
rect 936 186 966 260
rect 1031 280 1104 296
rect 1031 246 1054 280
rect 1088 246 1104 280
rect 1031 230 1104 246
rect 1031 208 1061 230
rect 1148 208 1178 338
rect 1226 346 1292 362
rect 1226 312 1242 346
rect 1276 312 1292 346
rect 1226 296 1292 312
rect 1360 310 1390 379
rect 1534 353 1564 368
rect 1624 353 1654 368
rect 1714 353 1744 368
rect 1804 353 1834 368
rect 1531 326 1567 353
rect 1621 326 1657 353
rect 1711 326 1747 353
rect 1531 320 1747 326
rect 1801 320 1837 353
rect 1531 310 1837 320
rect 1241 208 1271 296
rect 1360 294 1426 310
rect 1360 260 1376 294
rect 1410 274 1426 294
rect 1531 276 1547 310
rect 1581 276 1615 310
rect 1649 276 1683 310
rect 1717 290 1837 310
rect 1717 276 1831 290
rect 1410 260 1469 274
rect 1360 244 1469 260
rect 1439 222 1469 244
rect 1531 260 1831 276
rect 1531 222 1561 260
rect 1625 222 1655 260
rect 1715 222 1745 260
rect 1801 222 1831 260
rect 524 93 554 119
rect 610 93 640 119
rect 705 51 735 102
rect 777 76 807 102
rect 323 21 735 51
rect 1148 102 1178 124
rect 936 50 966 76
rect 1031 72 1061 98
rect 1133 86 1199 102
rect 1241 98 1271 124
rect 1133 52 1149 86
rect 1183 52 1199 86
rect 1133 36 1199 52
rect 1439 48 1469 74
rect 1531 48 1561 74
rect 1625 48 1655 74
rect 1715 48 1745 74
rect 1801 48 1831 74
<< polycont >>
rect 373 421 407 455
rect 647 366 681 400
rect 51 276 85 310
rect 177 260 211 294
rect 303 260 337 294
rect 411 241 445 275
rect 1141 426 1175 460
rect 827 342 861 376
rect 825 224 859 258
rect 1054 246 1088 280
rect 1242 312 1276 346
rect 1376 260 1410 294
rect 1547 276 1581 310
rect 1615 276 1649 310
rect 1683 276 1717 310
rect 1149 52 1183 86
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 129 580 163 649
rect 331 623 365 649
rect 129 508 163 546
rect 129 458 163 474
rect 203 580 295 596
rect 203 546 219 580
rect 253 546 295 580
rect 743 620 809 649
rect 331 573 365 589
rect 399 581 675 615
rect 743 586 759 620
rect 793 586 809 620
rect 203 539 295 546
rect 399 539 433 581
rect 641 552 675 581
rect 843 581 1191 615
rect 843 552 877 581
rect 203 505 433 539
rect 467 531 501 547
rect 203 497 295 505
rect 203 463 219 497
rect 253 463 295 497
rect 541 513 557 547
rect 591 513 607 547
rect 641 518 877 552
rect 541 497 607 513
rect 23 406 39 440
rect 73 424 89 440
rect 73 406 169 424
rect 23 390 169 406
rect 25 310 101 356
rect 25 276 51 310
rect 85 276 101 310
rect 25 260 101 276
rect 135 310 169 390
rect 203 414 295 463
rect 203 380 219 414
rect 253 380 295 414
rect 357 455 423 471
rect 357 421 373 455
rect 407 421 423 455
rect 357 405 423 421
rect 203 364 295 380
rect 261 310 295 364
rect 389 356 423 405
rect 467 424 501 497
rect 563 484 607 497
rect 911 509 945 547
rect 563 450 877 484
rect 467 390 529 424
rect 135 294 227 310
rect 135 260 177 294
rect 211 260 227 294
rect 135 226 227 260
rect 23 210 227 226
rect 23 176 39 210
rect 73 192 227 210
rect 73 176 89 192
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 125 131 159 158
rect 125 17 159 97
rect 193 85 227 192
rect 261 294 353 310
rect 261 260 303 294
rect 337 260 353 294
rect 261 244 353 260
rect 389 275 461 356
rect 261 189 295 244
rect 389 241 411 275
rect 445 241 461 275
rect 389 225 461 241
rect 495 248 529 390
rect 563 316 597 450
rect 631 400 775 416
rect 631 366 647 400
rect 681 366 775 400
rect 631 350 775 366
rect 563 282 669 316
rect 495 214 599 248
rect 565 180 599 214
rect 261 119 295 155
rect 329 146 531 180
rect 329 85 363 146
rect 193 51 363 85
rect 397 78 413 112
rect 447 78 463 112
rect 397 17 463 78
rect 497 85 531 146
rect 565 119 599 146
rect 635 190 669 282
rect 635 174 707 190
rect 635 140 654 174
rect 688 140 707 174
rect 635 124 707 140
rect 741 172 775 350
rect 811 376 877 450
rect 811 342 827 376
rect 861 342 877 376
rect 811 326 877 342
rect 911 274 945 475
rect 979 308 1013 581
rect 1047 509 1081 547
rect 1047 376 1081 475
rect 1125 460 1191 581
rect 1263 550 1330 649
rect 1263 516 1280 550
rect 1314 516 1330 550
rect 1263 490 1330 516
rect 1364 580 1430 596
rect 1364 546 1380 580
rect 1414 546 1430 580
rect 1125 426 1141 460
rect 1175 426 1191 460
rect 1125 410 1191 426
rect 1364 470 1430 546
rect 1364 436 1380 470
rect 1414 436 1430 470
rect 1364 378 1430 436
rect 1471 580 1521 649
rect 1471 546 1487 580
rect 1471 462 1521 546
rect 1471 428 1487 462
rect 1471 412 1521 428
rect 1561 580 1627 596
rect 1561 546 1577 580
rect 1611 546 1627 580
rect 1561 497 1627 546
rect 1561 463 1577 497
rect 1611 463 1627 497
rect 1561 414 1627 463
rect 1667 580 1701 649
rect 1667 478 1701 546
rect 1667 428 1701 444
rect 1741 580 1807 596
rect 1741 546 1757 580
rect 1791 546 1807 580
rect 1741 497 1807 546
rect 1741 463 1757 497
rect 1791 463 1807 497
rect 1561 380 1577 414
rect 1611 394 1627 414
rect 1741 414 1807 463
rect 1741 394 1757 414
rect 1611 380 1757 394
rect 1791 380 1807 414
rect 1047 342 1172 376
rect 1258 362 1494 378
rect 979 280 1104 308
rect 979 274 1054 280
rect 809 258 945 274
rect 809 224 825 258
rect 859 240 945 258
rect 1038 246 1054 274
rect 1088 246 1104 280
rect 859 224 1004 240
rect 1038 230 1104 246
rect 1138 262 1172 342
rect 1226 346 1494 362
rect 1561 360 1807 380
rect 1847 580 1897 649
rect 1881 546 1897 580
rect 1847 497 1897 546
rect 1881 463 1897 497
rect 1847 414 1897 463
rect 1881 380 1897 414
rect 1847 364 1897 380
rect 1226 312 1242 346
rect 1276 344 1494 346
rect 1276 312 1292 344
rect 1226 296 1292 312
rect 1460 326 1494 344
rect 1460 310 1733 326
rect 1360 294 1426 310
rect 1360 278 1376 294
rect 1326 262 1376 278
rect 1138 260 1376 262
rect 1410 260 1426 294
rect 1138 244 1426 260
rect 1460 276 1547 310
rect 1581 276 1615 310
rect 1649 276 1683 310
rect 1717 276 1733 310
rect 1460 260 1733 276
rect 809 206 1004 224
rect 970 190 1004 206
rect 1138 228 1360 244
rect 1138 194 1172 228
rect 1460 210 1494 260
rect 1773 226 1807 360
rect 1394 194 1494 210
rect 741 138 936 172
rect 741 85 775 138
rect 497 51 775 85
rect 818 88 868 104
rect 818 54 834 88
rect 818 17 868 54
rect 902 85 936 138
rect 970 171 1036 190
rect 970 137 986 171
rect 1020 137 1036 171
rect 1070 178 1172 194
rect 1070 144 1094 178
rect 1128 144 1172 178
rect 1282 174 1332 194
rect 970 119 1036 137
rect 1316 140 1332 174
rect 1133 86 1199 102
rect 1133 85 1149 86
rect 902 52 1149 85
rect 1183 52 1199 86
rect 902 51 1199 52
rect 1282 17 1332 140
rect 1378 160 1394 194
rect 1428 176 1494 194
rect 1564 210 1807 226
rect 1564 176 1580 210
rect 1614 192 1756 210
rect 1614 176 1630 192
rect 1378 120 1428 160
rect 1378 86 1394 120
rect 1378 70 1428 86
rect 1464 123 1530 142
rect 1464 89 1480 123
rect 1514 89 1530 123
rect 1464 17 1530 89
rect 1564 120 1630 176
rect 1740 176 1756 192
rect 1790 176 1807 210
rect 1564 86 1580 120
rect 1614 86 1630 120
rect 1564 70 1630 86
rect 1666 131 1700 158
rect 1666 17 1700 97
rect 1740 120 1807 176
rect 1740 86 1756 120
rect 1790 86 1807 120
rect 1740 70 1807 86
rect 1842 210 1892 226
rect 1876 176 1892 210
rect 1842 120 1892 176
rect 1876 86 1892 120
rect 1842 17 1892 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dfxtp_4
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 1759 390 1793 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1759 464 1793 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1759 538 1793 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 24720
string GDS_START 9868
<< end >>
