magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 500 228 956 248
rect 20 49 956 228
rect 0 0 960 49
<< scnmos >>
rect 103 74 133 202
rect 203 74 233 202
rect 303 74 333 202
rect 389 74 419 202
rect 479 74 509 202
rect 576 74 606 222
rect 664 74 694 222
rect 757 74 787 222
rect 843 74 873 222
<< scpmoshvt >>
rect 84 392 114 592
rect 188 424 218 592
rect 278 424 308 592
rect 382 424 412 592
rect 472 424 502 592
rect 576 368 606 592
rect 666 368 696 592
rect 756 368 786 592
rect 846 368 876 592
<< ndiff >>
rect 526 202 576 222
rect 46 190 103 202
rect 46 156 58 190
rect 92 156 103 190
rect 46 120 103 156
rect 46 86 58 120
rect 92 86 103 120
rect 46 74 103 86
rect 133 184 203 202
rect 133 150 158 184
rect 192 150 203 184
rect 133 116 203 150
rect 133 82 158 116
rect 192 82 203 116
rect 133 74 203 82
rect 233 146 303 202
rect 233 112 250 146
rect 284 112 303 146
rect 233 74 303 112
rect 333 185 389 202
rect 333 151 344 185
rect 378 151 389 185
rect 333 74 389 151
rect 419 117 479 202
rect 419 83 430 117
rect 464 83 479 117
rect 419 74 479 83
rect 509 117 576 202
rect 509 83 530 117
rect 564 83 576 117
rect 509 74 576 83
rect 606 210 664 222
rect 606 176 619 210
rect 653 176 664 210
rect 606 120 664 176
rect 606 86 619 120
rect 653 86 664 120
rect 606 74 664 86
rect 694 146 757 222
rect 694 112 705 146
rect 739 112 757 146
rect 694 74 757 112
rect 787 210 843 222
rect 787 176 798 210
rect 832 176 843 210
rect 787 120 843 176
rect 787 86 798 120
rect 832 86 843 120
rect 787 74 843 86
rect 873 146 930 222
rect 873 112 884 146
rect 918 112 930 146
rect 873 74 930 112
<< pdiff >>
rect 27 580 84 592
rect 27 546 37 580
rect 71 546 84 580
rect 27 510 84 546
rect 27 476 37 510
rect 71 476 84 510
rect 27 440 84 476
rect 27 406 37 440
rect 71 406 84 440
rect 27 392 84 406
rect 114 580 188 592
rect 114 546 127 580
rect 161 546 188 580
rect 114 470 188 546
rect 114 436 127 470
rect 161 436 188 470
rect 114 424 188 436
rect 218 580 278 592
rect 218 546 231 580
rect 265 546 278 580
rect 218 470 278 546
rect 218 436 231 470
rect 265 436 278 470
rect 218 424 278 436
rect 308 580 382 592
rect 308 546 321 580
rect 355 546 382 580
rect 308 510 382 546
rect 308 476 321 510
rect 355 476 382 510
rect 308 424 382 476
rect 412 580 472 592
rect 412 546 425 580
rect 459 546 472 580
rect 412 470 472 546
rect 412 436 425 470
rect 459 436 472 470
rect 412 424 472 436
rect 502 580 576 592
rect 502 546 529 580
rect 563 546 576 580
rect 502 510 576 546
rect 502 476 529 510
rect 563 476 576 510
rect 502 424 576 476
rect 114 392 170 424
rect 523 368 576 424
rect 606 580 666 592
rect 606 546 619 580
rect 653 546 666 580
rect 606 497 666 546
rect 606 463 619 497
rect 653 463 666 497
rect 606 414 666 463
rect 606 380 619 414
rect 653 380 666 414
rect 606 368 666 380
rect 696 580 756 592
rect 696 546 709 580
rect 743 546 756 580
rect 696 482 756 546
rect 696 448 709 482
rect 743 448 756 482
rect 696 368 756 448
rect 786 580 846 592
rect 786 546 799 580
rect 833 546 846 580
rect 786 497 846 546
rect 786 463 799 497
rect 833 463 846 497
rect 786 414 846 463
rect 786 380 799 414
rect 833 380 846 414
rect 786 368 846 380
rect 876 580 933 592
rect 876 546 889 580
rect 923 546 933 580
rect 876 497 933 546
rect 876 463 889 497
rect 923 463 933 497
rect 876 414 933 463
rect 876 380 889 414
rect 923 380 933 414
rect 876 368 933 380
<< ndiffc >>
rect 58 156 92 190
rect 58 86 92 120
rect 158 150 192 184
rect 158 82 192 116
rect 250 112 284 146
rect 344 151 378 185
rect 430 83 464 117
rect 530 83 564 117
rect 619 176 653 210
rect 619 86 653 120
rect 705 112 739 146
rect 798 176 832 210
rect 798 86 832 120
rect 884 112 918 146
<< pdiffc >>
rect 37 546 71 580
rect 37 476 71 510
rect 37 406 71 440
rect 127 546 161 580
rect 127 436 161 470
rect 231 546 265 580
rect 231 436 265 470
rect 321 546 355 580
rect 321 476 355 510
rect 425 546 459 580
rect 425 436 459 470
rect 529 546 563 580
rect 529 476 563 510
rect 619 546 653 580
rect 619 463 653 497
rect 619 380 653 414
rect 709 546 743 580
rect 709 448 743 482
rect 799 546 833 580
rect 799 463 833 497
rect 799 380 833 414
rect 889 546 923 580
rect 889 463 923 497
rect 889 380 923 414
<< poly >>
rect 84 592 114 618
rect 188 592 218 618
rect 278 592 308 618
rect 382 592 412 618
rect 472 592 502 618
rect 576 592 606 618
rect 666 592 696 618
rect 756 592 786 618
rect 846 592 876 618
rect 188 409 218 424
rect 278 409 308 424
rect 382 409 412 424
rect 472 409 502 424
rect 84 377 114 392
rect 185 379 333 409
rect 379 379 505 409
rect 81 356 117 377
rect 81 340 149 356
rect 81 306 99 340
rect 133 306 149 340
rect 81 290 149 306
rect 195 321 261 337
rect 103 202 133 290
rect 195 287 211 321
rect 245 287 261 321
rect 195 271 261 287
rect 303 290 333 379
rect 461 310 491 379
rect 576 353 606 368
rect 666 353 696 368
rect 756 353 786 368
rect 846 353 876 368
rect 573 330 609 353
rect 663 330 699 353
rect 753 330 789 353
rect 573 314 789 330
rect 461 294 527 310
rect 573 294 592 314
rect 303 274 369 290
rect 203 202 233 271
rect 303 240 319 274
rect 353 254 369 274
rect 461 260 477 294
rect 511 260 527 294
rect 353 240 419 254
rect 461 244 527 260
rect 576 280 592 294
rect 626 280 660 314
rect 694 280 728 314
rect 762 280 789 314
rect 576 267 789 280
rect 843 267 879 353
rect 576 264 873 267
rect 303 224 419 240
rect 303 202 333 224
rect 389 202 419 224
rect 479 202 509 244
rect 576 222 606 264
rect 664 222 694 264
rect 757 237 873 264
rect 757 222 787 237
rect 843 222 873 237
rect 103 48 133 74
rect 203 48 233 74
rect 303 48 333 74
rect 389 48 419 74
rect 479 48 509 74
rect 576 48 606 74
rect 664 48 694 74
rect 757 48 787 74
rect 843 48 873 74
<< polycont >>
rect 99 306 133 340
rect 211 287 245 321
rect 319 240 353 274
rect 477 260 511 294
rect 592 280 626 314
rect 660 280 694 314
rect 728 280 762 314
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 17 580 71 596
rect 17 546 37 580
rect 17 510 71 546
rect 17 476 37 510
rect 17 440 71 476
rect 17 406 37 440
rect 111 580 177 649
rect 111 546 127 580
rect 161 546 177 580
rect 111 470 177 546
rect 111 436 127 470
rect 161 436 177 470
rect 111 420 177 436
rect 215 580 281 596
rect 215 546 231 580
rect 265 546 281 580
rect 215 470 281 546
rect 215 436 231 470
rect 265 436 281 470
rect 321 580 371 649
rect 355 546 371 580
rect 321 510 371 546
rect 355 476 371 510
rect 321 460 371 476
rect 409 580 475 596
rect 409 546 425 580
rect 459 546 475 580
rect 409 470 475 546
rect 215 426 281 436
rect 409 436 425 470
rect 459 436 475 470
rect 513 580 579 649
rect 513 546 529 580
rect 563 546 579 580
rect 513 510 579 546
rect 513 476 529 510
rect 563 476 579 510
rect 513 460 579 476
rect 619 580 653 596
rect 619 497 653 546
rect 409 426 475 436
rect 17 390 71 406
rect 215 392 585 426
rect 17 253 51 390
rect 85 340 161 356
rect 85 306 99 340
rect 133 306 161 340
rect 85 290 161 306
rect 195 324 517 358
rect 195 321 261 324
rect 195 287 211 321
rect 245 287 261 321
rect 409 294 517 324
rect 303 274 369 290
rect 303 253 319 274
rect 17 240 319 253
rect 353 240 369 274
rect 17 219 369 240
rect 409 260 477 294
rect 511 260 517 294
rect 409 236 517 260
rect 551 330 585 392
rect 619 414 653 463
rect 693 580 759 649
rect 693 546 709 580
rect 743 546 759 580
rect 693 482 759 546
rect 693 448 709 482
rect 743 448 759 482
rect 693 432 759 448
rect 799 580 833 596
rect 799 497 833 546
rect 799 414 833 463
rect 653 380 799 398
rect 619 364 833 380
rect 873 580 939 649
rect 873 546 889 580
rect 923 546 939 580
rect 873 497 939 546
rect 873 463 889 497
rect 923 463 939 497
rect 873 414 939 463
rect 873 380 889 414
rect 923 380 939 414
rect 873 364 939 380
rect 799 330 833 364
rect 551 314 765 330
rect 551 280 592 314
rect 626 280 660 314
rect 694 280 728 314
rect 762 280 765 314
rect 799 296 935 330
rect 551 264 765 280
rect 17 190 108 219
rect 17 156 58 190
rect 92 156 108 190
rect 551 185 585 264
rect 889 230 935 296
rect 17 120 108 156
rect 17 86 58 120
rect 92 86 108 120
rect 17 70 108 86
rect 142 184 208 185
rect 142 150 158 184
rect 192 150 208 184
rect 142 116 208 150
rect 142 82 158 116
rect 192 82 208 116
rect 142 17 208 82
rect 242 146 294 185
rect 328 151 344 185
rect 378 151 585 185
rect 619 210 935 230
rect 653 196 798 210
rect 242 112 250 146
rect 284 117 294 146
rect 619 120 653 176
rect 782 176 798 196
rect 832 196 935 210
rect 284 112 430 117
rect 242 83 430 112
rect 464 83 480 117
rect 242 67 480 83
rect 514 83 530 117
rect 564 83 580 117
rect 514 17 580 83
rect 619 70 653 86
rect 689 146 739 162
rect 689 112 705 146
rect 689 17 739 112
rect 782 120 832 176
rect 782 86 798 120
rect 782 70 832 86
rect 868 146 934 162
rect 868 112 884 146
rect 918 112 934 146
rect 868 17 934 112
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 and2b_4
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 3071504
string GDS_START 3063080
<< end >>
