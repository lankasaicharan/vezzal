magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 6 241 281 246
rect 6 49 667 241
rect 0 0 672 49
<< scnmos >>
rect 85 52 115 220
rect 157 52 187 220
rect 366 47 396 215
rect 452 47 482 215
rect 558 47 588 215
<< scpmoshvt >>
rect 85 367 115 619
rect 171 367 201 619
rect 372 367 402 619
rect 474 367 504 619
rect 558 367 588 619
<< ndiff >>
rect 32 202 85 220
rect 32 168 40 202
rect 74 168 85 202
rect 32 98 85 168
rect 32 64 40 98
rect 74 64 85 98
rect 32 52 85 64
rect 115 52 157 220
rect 187 202 255 220
rect 187 168 213 202
rect 247 168 255 202
rect 187 98 255 168
rect 187 64 213 98
rect 247 64 255 98
rect 187 52 255 64
rect 313 203 366 215
rect 313 169 321 203
rect 355 169 366 203
rect 313 101 366 169
rect 313 67 321 101
rect 355 67 366 101
rect 313 47 366 67
rect 396 163 452 215
rect 396 129 407 163
rect 441 129 452 163
rect 396 95 452 129
rect 396 61 407 95
rect 441 61 452 95
rect 396 47 452 61
rect 482 103 558 215
rect 482 69 507 103
rect 541 69 558 103
rect 482 47 558 69
rect 588 203 641 215
rect 588 169 599 203
rect 633 169 641 203
rect 588 103 641 169
rect 588 69 599 103
rect 633 69 641 103
rect 588 47 641 69
<< pdiff >>
rect 32 607 85 619
rect 32 573 40 607
rect 74 573 85 607
rect 32 515 85 573
rect 32 481 40 515
rect 74 481 85 515
rect 32 418 85 481
rect 32 384 40 418
rect 74 384 85 418
rect 32 367 85 384
rect 115 599 171 619
rect 115 565 126 599
rect 160 565 171 599
rect 115 506 171 565
rect 115 472 126 506
rect 160 472 171 506
rect 115 413 171 472
rect 115 379 126 413
rect 160 379 171 413
rect 115 367 171 379
rect 201 607 372 619
rect 201 573 212 607
rect 246 573 327 607
rect 361 573 372 607
rect 201 539 372 573
rect 201 534 327 539
rect 201 500 212 534
rect 246 505 327 534
rect 361 505 372 539
rect 246 500 372 505
rect 201 469 372 500
rect 201 453 327 469
rect 201 419 212 453
rect 246 435 327 453
rect 361 435 372 469
rect 246 419 372 435
rect 201 367 372 419
rect 402 599 474 619
rect 402 565 417 599
rect 451 565 474 599
rect 402 504 474 565
rect 402 470 417 504
rect 451 470 474 504
rect 402 413 474 470
rect 402 379 417 413
rect 451 379 474 413
rect 402 367 474 379
rect 504 367 558 619
rect 588 607 641 619
rect 588 573 599 607
rect 633 573 641 607
rect 588 511 641 573
rect 588 477 599 511
rect 633 477 641 511
rect 588 418 641 477
rect 588 384 599 418
rect 633 384 641 418
rect 588 367 641 384
<< ndiffc >>
rect 40 168 74 202
rect 40 64 74 98
rect 213 168 247 202
rect 213 64 247 98
rect 321 169 355 203
rect 321 67 355 101
rect 407 129 441 163
rect 407 61 441 95
rect 507 69 541 103
rect 599 169 633 203
rect 599 69 633 103
<< pdiffc >>
rect 40 573 74 607
rect 40 481 74 515
rect 40 384 74 418
rect 126 565 160 599
rect 126 472 160 506
rect 126 379 160 413
rect 212 573 246 607
rect 327 573 361 607
rect 212 500 246 534
rect 327 505 361 539
rect 212 419 246 453
rect 327 435 361 469
rect 417 565 451 599
rect 417 470 451 504
rect 417 379 451 413
rect 599 573 633 607
rect 599 477 633 511
rect 599 384 633 418
<< poly >>
rect 85 619 115 645
rect 171 619 201 645
rect 372 619 402 645
rect 474 619 504 645
rect 558 619 588 645
rect 85 308 115 367
rect 171 308 201 367
rect 372 335 402 367
rect 286 319 402 335
rect 40 292 115 308
rect 40 258 56 292
rect 90 258 115 292
rect 40 242 115 258
rect 85 220 115 242
rect 157 292 229 308
rect 157 258 173 292
rect 207 258 229 292
rect 157 242 229 258
rect 286 285 302 319
rect 336 287 402 319
rect 474 308 504 367
rect 558 308 588 367
rect 444 292 516 308
rect 336 285 396 287
rect 286 257 396 285
rect 157 220 187 242
rect 366 215 396 257
rect 444 258 466 292
rect 500 258 516 292
rect 444 242 516 258
rect 558 292 631 308
rect 558 258 581 292
rect 615 258 631 292
rect 558 242 631 258
rect 452 215 482 242
rect 558 215 588 242
rect 85 26 115 52
rect 157 26 187 52
rect 366 21 396 47
rect 452 21 482 47
rect 558 21 588 47
<< polycont >>
rect 56 258 90 292
rect 173 258 207 292
rect 302 285 336 319
rect 466 258 500 292
rect 581 258 615 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 24 607 90 649
rect 24 573 40 607
rect 74 573 90 607
rect 24 515 90 573
rect 24 481 40 515
rect 74 481 90 515
rect 24 418 90 481
rect 24 384 40 418
rect 74 384 90 418
rect 124 599 162 615
rect 124 565 126 599
rect 160 565 162 599
rect 124 506 162 565
rect 124 472 126 506
rect 160 472 162 506
rect 124 413 162 472
rect 196 607 364 649
rect 196 573 212 607
rect 246 573 327 607
rect 361 573 364 607
rect 196 539 364 573
rect 196 534 327 539
rect 196 500 212 534
rect 246 505 327 534
rect 361 505 364 539
rect 246 500 364 505
rect 196 469 364 500
rect 196 453 327 469
rect 196 419 212 453
rect 246 435 327 453
rect 361 435 364 469
rect 246 419 364 435
rect 398 599 467 615
rect 583 607 649 649
rect 398 565 417 599
rect 451 565 467 599
rect 398 504 467 565
rect 398 470 417 504
rect 451 470 467 504
rect 124 379 126 413
rect 160 385 162 413
rect 398 413 467 470
rect 398 385 417 413
rect 160 379 283 385
rect 124 351 283 379
rect 17 292 90 350
rect 241 335 283 351
rect 386 379 417 385
rect 451 379 467 413
rect 386 351 467 379
rect 241 319 352 335
rect 17 258 56 292
rect 17 242 90 258
rect 125 292 207 308
rect 125 258 173 292
rect 125 242 207 258
rect 241 285 302 319
rect 336 285 352 319
rect 241 281 352 285
rect 241 208 275 281
rect 386 247 420 351
rect 501 317 547 599
rect 583 573 599 607
rect 633 573 649 607
rect 583 511 649 573
rect 583 477 599 511
rect 633 477 649 511
rect 583 418 649 477
rect 583 384 599 418
rect 633 384 649 418
rect 24 202 90 208
rect 24 168 40 202
rect 74 168 90 202
rect 24 98 90 168
rect 24 64 40 98
rect 74 64 90 98
rect 24 17 90 64
rect 197 202 275 208
rect 197 168 213 202
rect 247 168 275 202
rect 197 164 275 168
rect 309 213 420 247
rect 466 292 547 317
rect 500 258 547 292
rect 466 237 547 258
rect 581 292 655 350
rect 615 258 655 292
rect 581 237 655 258
rect 309 203 357 213
rect 309 169 321 203
rect 355 169 357 203
rect 454 179 599 203
rect 197 98 263 164
rect 309 130 357 169
rect 197 64 213 98
rect 247 64 263 98
rect 197 51 263 64
rect 305 101 357 130
rect 305 67 321 101
rect 355 67 357 101
rect 305 51 357 67
rect 391 169 599 179
rect 633 169 649 203
rect 391 163 649 169
rect 391 129 407 163
rect 441 145 649 163
rect 441 129 457 145
rect 391 95 457 129
rect 391 61 407 95
rect 441 61 457 95
rect 391 57 457 61
rect 491 103 557 111
rect 491 69 507 103
rect 541 69 557 103
rect 491 17 557 69
rect 595 103 649 145
rect 595 69 599 103
rect 633 69 649 103
rect 595 53 649 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2bb2ai_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4131462
string GDS_START 4123486
<< end >>
