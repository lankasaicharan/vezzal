magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 263 241 742 250
rect 1 49 742 241
rect 0 0 768 49
<< scnmos >>
rect 80 47 110 215
rect 152 47 182 215
rect 342 56 372 224
rect 428 56 458 224
rect 522 56 552 224
rect 608 56 638 224
<< scpmoshvt >>
rect 114 367 144 619
rect 208 367 238 619
rect 342 367 372 619
rect 414 367 444 619
rect 568 367 598 619
rect 654 367 684 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 93 80 169
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 47 152 215
rect 182 203 235 215
rect 182 169 193 203
rect 227 169 235 203
rect 182 104 235 169
rect 182 70 193 104
rect 227 70 235 104
rect 182 47 235 70
rect 289 132 342 224
rect 289 98 297 132
rect 331 98 342 132
rect 289 56 342 98
rect 372 208 428 224
rect 372 174 383 208
rect 417 174 428 208
rect 372 104 428 174
rect 372 70 383 104
rect 417 70 428 104
rect 372 56 428 70
rect 458 192 522 224
rect 458 158 473 192
rect 507 158 522 192
rect 458 102 522 158
rect 458 68 473 102
rect 507 68 522 102
rect 458 56 522 68
rect 552 209 608 224
rect 552 175 563 209
rect 597 175 608 209
rect 552 101 608 175
rect 552 67 563 101
rect 597 67 608 101
rect 552 56 608 67
rect 638 195 716 224
rect 638 161 674 195
rect 708 161 716 195
rect 638 102 716 161
rect 638 68 649 102
rect 683 68 716 102
rect 638 56 716 68
<< pdiff >>
rect 61 599 114 619
rect 61 565 69 599
rect 103 565 114 599
rect 61 503 114 565
rect 61 469 69 503
rect 103 469 114 503
rect 61 413 114 469
rect 61 379 69 413
rect 103 379 114 413
rect 61 367 114 379
rect 144 607 208 619
rect 144 573 159 607
rect 193 573 208 607
rect 144 528 208 573
rect 144 494 159 528
rect 193 494 208 528
rect 144 451 208 494
rect 144 417 159 451
rect 193 417 208 451
rect 144 367 208 417
rect 238 599 342 619
rect 238 565 273 599
rect 307 565 342 599
rect 238 503 342 565
rect 238 469 273 503
rect 307 469 342 503
rect 238 413 342 469
rect 238 379 249 413
rect 283 379 342 413
rect 238 367 342 379
rect 372 367 414 619
rect 444 568 568 619
rect 444 534 455 568
rect 489 534 523 568
rect 557 534 568 568
rect 444 367 568 534
rect 598 599 654 619
rect 598 565 609 599
rect 643 565 654 599
rect 598 503 654 565
rect 598 469 609 503
rect 643 469 654 503
rect 598 419 654 469
rect 598 385 609 419
rect 643 385 654 419
rect 598 367 654 385
rect 684 607 737 619
rect 684 573 695 607
rect 729 573 737 607
rect 684 496 737 573
rect 684 462 695 496
rect 729 462 737 496
rect 684 367 737 462
<< ndiffc >>
rect 35 169 69 203
rect 35 59 69 93
rect 193 169 227 203
rect 193 70 227 104
rect 297 98 331 132
rect 383 174 417 208
rect 383 70 417 104
rect 473 158 507 192
rect 473 68 507 102
rect 563 175 597 209
rect 563 67 597 101
rect 674 161 708 195
rect 649 68 683 102
<< pdiffc >>
rect 69 565 103 599
rect 69 469 103 503
rect 69 379 103 413
rect 159 573 193 607
rect 159 494 193 528
rect 159 417 193 451
rect 273 565 307 599
rect 273 469 307 503
rect 249 379 283 413
rect 455 534 489 568
rect 523 534 557 568
rect 609 565 643 599
rect 609 469 643 503
rect 609 385 643 419
rect 695 573 729 607
rect 695 462 729 496
<< poly >>
rect 114 619 144 645
rect 208 619 238 645
rect 342 619 372 645
rect 414 619 444 645
rect 568 619 598 645
rect 654 619 684 645
rect 114 345 144 367
rect 21 315 144 345
rect 21 299 110 315
rect 208 303 238 367
rect 342 328 372 367
rect 298 325 372 328
rect 21 265 37 299
rect 71 265 110 299
rect 186 287 252 303
rect 186 267 202 287
rect 21 249 110 265
rect 80 215 110 249
rect 152 253 202 267
rect 236 253 252 287
rect 152 237 252 253
rect 294 296 372 325
rect 294 262 319 296
rect 353 262 372 296
rect 294 246 372 262
rect 414 312 444 367
rect 568 326 598 367
rect 533 325 598 326
rect 654 325 684 367
rect 414 296 480 312
rect 414 262 430 296
rect 464 262 480 296
rect 414 246 480 262
rect 522 309 684 325
rect 522 275 538 309
rect 572 275 684 309
rect 522 259 684 275
rect 152 215 182 237
rect 342 224 372 246
rect 428 224 458 246
rect 522 224 552 259
rect 608 224 638 259
rect 80 21 110 47
rect 152 21 182 47
rect 342 30 372 56
rect 428 30 458 56
rect 522 30 552 56
rect 608 30 638 56
<< polycont >>
rect 37 265 71 299
rect 202 253 236 287
rect 319 262 353 296
rect 430 262 464 296
rect 538 275 572 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 53 599 109 615
rect 53 565 69 599
rect 103 565 109 599
rect 53 503 109 565
rect 53 469 69 503
rect 103 469 109 503
rect 53 413 109 469
rect 143 607 209 649
rect 143 573 159 607
rect 193 573 209 607
rect 143 528 209 573
rect 143 494 159 528
rect 193 494 209 528
rect 143 451 209 494
rect 143 417 159 451
rect 193 417 209 451
rect 243 599 323 615
rect 243 565 273 599
rect 307 565 323 599
rect 243 503 323 565
rect 439 568 573 649
rect 439 534 455 568
rect 489 534 523 568
rect 557 534 573 568
rect 439 526 573 534
rect 607 599 645 615
rect 607 565 609 599
rect 643 565 645 599
rect 243 469 273 503
rect 307 492 323 503
rect 607 503 645 565
rect 607 492 609 503
rect 307 469 532 492
rect 243 458 532 469
rect 53 379 69 413
rect 103 383 109 413
rect 243 413 285 458
rect 243 383 249 413
rect 103 379 249 383
rect 283 379 285 413
rect 53 349 285 379
rect 105 328 285 349
rect 31 299 71 315
rect 31 265 37 299
rect 31 242 71 265
rect 105 208 141 328
rect 319 296 363 424
rect 186 287 257 294
rect 186 253 202 287
rect 236 253 257 287
rect 186 242 257 253
rect 353 262 363 296
rect 319 242 363 262
rect 405 296 464 424
rect 405 262 430 296
rect 405 242 464 262
rect 498 325 532 458
rect 606 469 609 492
rect 643 469 645 503
rect 606 424 645 469
rect 679 607 745 649
rect 679 573 695 607
rect 729 573 745 607
rect 679 496 745 573
rect 679 462 695 496
rect 729 462 745 496
rect 679 458 745 462
rect 606 419 697 424
rect 606 385 609 419
rect 643 385 697 419
rect 498 309 572 325
rect 498 275 538 309
rect 498 259 572 275
rect 606 250 697 385
rect 606 238 644 250
rect 606 225 640 238
rect 547 209 640 225
rect 19 203 141 208
rect 19 169 35 203
rect 69 172 141 203
rect 177 203 383 208
rect 69 169 85 172
rect 19 93 85 169
rect 19 59 35 93
rect 69 59 85 93
rect 19 51 85 59
rect 177 169 193 203
rect 227 174 383 203
rect 417 174 433 208
rect 227 169 243 174
rect 177 104 243 169
rect 177 70 193 104
rect 227 70 243 104
rect 177 54 243 70
rect 281 132 347 140
rect 281 98 297 132
rect 331 98 347 132
rect 281 17 347 98
rect 381 104 433 174
rect 381 70 383 104
rect 417 70 433 104
rect 381 54 433 70
rect 467 192 513 208
rect 467 158 473 192
rect 507 158 513 192
rect 467 102 513 158
rect 467 68 473 102
rect 507 68 513 102
rect 467 17 513 68
rect 547 175 563 209
rect 597 191 640 209
rect 674 195 724 211
rect 597 175 613 191
rect 547 101 613 175
rect 708 161 724 195
rect 674 157 724 161
rect 547 67 563 101
rect 597 67 613 101
rect 547 51 613 67
rect 647 102 724 157
rect 647 68 649 102
rect 683 68 724 102
rect 647 17 724 68
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o211a_2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1686014
string GDS_START 1678326
<< end >>
