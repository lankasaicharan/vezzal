magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1682 1975
<< nwell >>
rect -38 331 422 704
<< pwell >>
rect 72 49 346 203
rect 0 0 384 49
<< scnmos >>
rect 155 67 185 177
rect 233 67 263 177
<< scpmoshvt >>
rect 141 396 191 596
rect 247 396 297 596
<< ndiff >>
rect 98 139 155 177
rect 98 105 110 139
rect 144 105 155 139
rect 98 67 155 105
rect 185 67 233 177
rect 263 126 320 177
rect 263 92 274 126
rect 308 92 320 126
rect 263 67 320 92
<< pdiff >>
rect 88 584 141 596
rect 88 550 96 584
rect 130 550 141 584
rect 88 513 141 550
rect 88 479 96 513
rect 130 479 141 513
rect 88 442 141 479
rect 88 408 96 442
rect 130 408 141 442
rect 88 396 141 408
rect 191 584 247 596
rect 191 550 202 584
rect 236 550 247 584
rect 191 513 247 550
rect 191 479 202 513
rect 236 479 247 513
rect 191 442 247 479
rect 191 408 202 442
rect 236 408 247 442
rect 191 396 247 408
rect 297 584 350 596
rect 297 550 308 584
rect 342 550 350 584
rect 297 513 350 550
rect 297 479 308 513
rect 342 479 350 513
rect 297 442 350 479
rect 297 408 308 442
rect 342 408 350 442
rect 297 396 350 408
<< ndiffc >>
rect 110 105 144 139
rect 274 92 308 126
<< pdiffc >>
rect 96 550 130 584
rect 96 479 130 513
rect 96 408 130 442
rect 202 550 236 584
rect 202 479 236 513
rect 202 408 236 442
rect 308 550 342 584
rect 308 479 342 513
rect 308 408 342 442
<< poly >>
rect 141 596 191 622
rect 247 596 297 622
rect 141 333 191 396
rect 247 333 297 396
rect 75 317 297 333
rect 75 283 121 317
rect 155 283 297 317
rect 75 269 297 283
rect 75 249 263 269
rect 75 215 121 249
rect 155 215 263 249
rect 75 199 263 215
rect 155 177 185 199
rect 233 177 263 199
rect 155 41 185 67
rect 233 41 263 67
<< polycont >>
rect 121 283 155 317
rect 121 215 155 249
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 80 584 146 649
rect 80 550 96 584
rect 130 550 146 584
rect 80 513 146 550
rect 80 479 96 513
rect 130 479 146 513
rect 80 442 146 479
rect 80 408 96 442
rect 130 408 146 442
rect 80 392 146 408
rect 186 584 264 600
rect 186 550 202 584
rect 236 550 264 584
rect 186 513 264 550
rect 186 479 202 513
rect 236 479 264 513
rect 186 442 264 479
rect 186 408 202 442
rect 236 408 264 442
rect 186 392 264 408
rect 298 584 358 649
rect 298 550 308 584
rect 342 550 358 584
rect 298 513 358 550
rect 298 479 308 513
rect 342 479 358 513
rect 298 442 358 479
rect 298 408 308 442
rect 342 408 358 442
rect 298 392 358 408
rect 20 317 171 356
rect 20 283 121 317
rect 155 283 171 317
rect 20 249 171 283
rect 20 215 121 249
rect 155 215 171 249
rect 20 199 171 215
rect 207 156 264 392
rect 94 139 160 155
rect 94 105 110 139
rect 144 105 160 139
rect 94 17 160 105
rect 207 126 324 156
rect 207 92 274 126
rect 308 92 324 126
rect 207 63 324 92
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 683 384 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 617 384 649
rect 0 17 384 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -49 384 -17
<< labels >>
flabel pwell s 0 0 384 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 384 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkinvlp_2
flabel metal1 s 0 617 384 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 384 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 384 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2205924
string GDS_START 2201400
<< end >>
