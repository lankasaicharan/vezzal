magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 164 49 1343 241
rect 0 0 1344 49
<< scnmos >>
rect 243 47 273 215
rect 329 47 359 215
rect 415 47 445 215
rect 501 47 531 215
rect 602 47 632 215
rect 688 47 718 215
rect 774 47 804 215
rect 860 47 890 215
rect 976 47 1006 215
rect 1062 47 1092 215
rect 1148 47 1178 215
rect 1234 47 1264 215
<< scpmoshvt >>
rect 153 367 183 619
rect 239 367 269 619
rect 325 367 355 619
rect 411 367 441 619
rect 602 367 632 619
rect 688 367 718 619
rect 774 367 804 619
rect 860 367 890 619
rect 960 367 990 619
rect 1062 367 1092 619
rect 1148 367 1178 619
rect 1234 367 1264 619
<< ndiff >>
rect 190 175 243 215
rect 190 141 198 175
rect 232 141 243 175
rect 190 93 243 141
rect 190 59 198 93
rect 232 59 243 93
rect 190 47 243 59
rect 273 203 329 215
rect 273 169 284 203
rect 318 169 329 203
rect 273 101 329 169
rect 273 67 284 101
rect 318 67 329 101
rect 273 47 329 67
rect 359 173 415 215
rect 359 139 370 173
rect 404 139 415 173
rect 359 89 415 139
rect 359 55 370 89
rect 404 55 415 89
rect 359 47 415 55
rect 445 203 501 215
rect 445 169 456 203
rect 490 169 501 203
rect 445 101 501 169
rect 445 67 456 101
rect 490 67 501 101
rect 445 47 501 67
rect 531 130 602 215
rect 531 96 542 130
rect 576 96 602 130
rect 531 47 602 96
rect 632 114 688 215
rect 632 80 643 114
rect 677 80 688 114
rect 632 47 688 80
rect 718 202 774 215
rect 718 168 729 202
rect 763 168 774 202
rect 718 47 774 168
rect 804 114 860 215
rect 804 80 815 114
rect 849 80 860 114
rect 804 47 860 80
rect 890 114 976 215
rect 890 80 905 114
rect 939 80 976 114
rect 890 47 976 80
rect 1006 114 1062 215
rect 1006 80 1017 114
rect 1051 80 1062 114
rect 1006 47 1062 80
rect 1092 190 1148 215
rect 1092 156 1103 190
rect 1137 156 1148 190
rect 1092 47 1148 156
rect 1178 190 1234 215
rect 1178 156 1189 190
rect 1223 156 1234 190
rect 1178 101 1234 156
rect 1178 67 1189 101
rect 1223 67 1234 101
rect 1178 47 1234 67
rect 1264 190 1317 215
rect 1264 156 1275 190
rect 1309 156 1317 190
rect 1264 93 1317 156
rect 1264 59 1275 93
rect 1309 59 1317 93
rect 1264 47 1317 59
<< pdiff >>
rect 100 607 153 619
rect 100 573 108 607
rect 142 573 153 607
rect 100 539 153 573
rect 100 505 108 539
rect 142 505 153 539
rect 100 453 153 505
rect 100 419 108 453
rect 142 419 153 453
rect 100 367 153 419
rect 183 599 239 619
rect 183 565 194 599
rect 228 565 239 599
rect 183 516 239 565
rect 183 482 194 516
rect 228 482 239 516
rect 183 413 239 482
rect 183 379 194 413
rect 228 379 239 413
rect 183 367 239 379
rect 269 607 325 619
rect 269 573 280 607
rect 314 573 325 607
rect 269 539 325 573
rect 269 505 280 539
rect 314 505 325 539
rect 269 453 325 505
rect 269 419 280 453
rect 314 419 325 453
rect 269 367 325 419
rect 355 599 411 619
rect 355 565 366 599
rect 400 565 411 599
rect 355 516 411 565
rect 355 482 366 516
rect 400 482 411 516
rect 355 413 411 482
rect 355 379 366 413
rect 400 379 411 413
rect 355 367 411 379
rect 441 607 494 619
rect 441 573 452 607
rect 486 573 494 607
rect 441 510 494 573
rect 441 476 452 510
rect 486 476 494 510
rect 441 413 494 476
rect 441 379 452 413
rect 486 379 494 413
rect 441 367 494 379
rect 549 599 602 619
rect 549 565 557 599
rect 591 565 602 599
rect 549 495 602 565
rect 549 461 557 495
rect 591 461 602 495
rect 549 367 602 461
rect 632 531 688 619
rect 632 497 643 531
rect 677 497 688 531
rect 632 441 688 497
rect 632 407 643 441
rect 677 407 688 441
rect 632 367 688 407
rect 718 599 774 619
rect 718 565 729 599
rect 763 565 774 599
rect 718 495 774 565
rect 718 461 729 495
rect 763 461 774 495
rect 718 367 774 461
rect 804 531 860 619
rect 804 497 815 531
rect 849 497 860 531
rect 804 443 860 497
rect 804 409 815 443
rect 849 409 860 443
rect 804 367 860 409
rect 890 599 960 619
rect 890 565 909 599
rect 943 565 960 599
rect 890 513 960 565
rect 890 479 909 513
rect 943 479 960 513
rect 890 425 960 479
rect 890 391 909 425
rect 943 391 960 425
rect 890 367 960 391
rect 990 607 1062 619
rect 990 573 1009 607
rect 1043 573 1062 607
rect 990 493 1062 573
rect 990 459 1009 493
rect 1043 459 1062 493
rect 990 367 1062 459
rect 1092 599 1148 619
rect 1092 565 1103 599
rect 1137 565 1148 599
rect 1092 513 1148 565
rect 1092 479 1103 513
rect 1137 479 1148 513
rect 1092 441 1148 479
rect 1092 407 1103 441
rect 1137 407 1148 441
rect 1092 367 1148 407
rect 1178 607 1234 619
rect 1178 573 1189 607
rect 1223 573 1234 607
rect 1178 493 1234 573
rect 1178 459 1189 493
rect 1223 459 1234 493
rect 1178 367 1234 459
rect 1264 599 1317 619
rect 1264 565 1275 599
rect 1309 565 1317 599
rect 1264 520 1317 565
rect 1264 486 1275 520
rect 1309 486 1317 520
rect 1264 441 1317 486
rect 1264 407 1275 441
rect 1309 407 1317 441
rect 1264 367 1317 407
<< ndiffc >>
rect 198 141 232 175
rect 198 59 232 93
rect 284 169 318 203
rect 284 67 318 101
rect 370 139 404 173
rect 370 55 404 89
rect 456 169 490 203
rect 456 67 490 101
rect 542 96 576 130
rect 643 80 677 114
rect 729 168 763 202
rect 815 80 849 114
rect 905 80 939 114
rect 1017 80 1051 114
rect 1103 156 1137 190
rect 1189 156 1223 190
rect 1189 67 1223 101
rect 1275 156 1309 190
rect 1275 59 1309 93
<< pdiffc >>
rect 108 573 142 607
rect 108 505 142 539
rect 108 419 142 453
rect 194 565 228 599
rect 194 482 228 516
rect 194 379 228 413
rect 280 573 314 607
rect 280 505 314 539
rect 280 419 314 453
rect 366 565 400 599
rect 366 482 400 516
rect 366 379 400 413
rect 452 573 486 607
rect 452 476 486 510
rect 452 379 486 413
rect 557 565 591 599
rect 557 461 591 495
rect 643 497 677 531
rect 643 407 677 441
rect 729 565 763 599
rect 729 461 763 495
rect 815 497 849 531
rect 815 409 849 443
rect 909 565 943 599
rect 909 479 943 513
rect 909 391 943 425
rect 1009 573 1043 607
rect 1009 459 1043 493
rect 1103 565 1137 599
rect 1103 479 1137 513
rect 1103 407 1137 441
rect 1189 573 1223 607
rect 1189 459 1223 493
rect 1275 565 1309 599
rect 1275 486 1309 520
rect 1275 407 1309 441
<< poly >>
rect 153 619 183 645
rect 239 619 269 645
rect 325 619 355 645
rect 411 619 441 645
rect 602 619 632 645
rect 688 619 718 645
rect 774 619 804 645
rect 860 619 890 645
rect 960 619 990 645
rect 1062 619 1092 645
rect 1148 619 1178 645
rect 1234 619 1264 645
rect 153 329 183 367
rect 239 329 269 367
rect 325 329 355 367
rect 411 329 441 367
rect 602 335 632 367
rect 103 313 531 329
rect 103 279 119 313
rect 153 279 187 313
rect 221 279 255 313
rect 289 279 323 313
rect 357 279 391 313
rect 425 279 459 313
rect 493 279 531 313
rect 103 263 531 279
rect 580 319 646 335
rect 580 285 596 319
rect 630 285 646 319
rect 580 269 646 285
rect 688 303 718 367
rect 774 303 804 367
rect 860 335 890 367
rect 960 335 990 367
rect 688 287 804 303
rect 243 215 273 263
rect 329 215 359 263
rect 415 215 445 263
rect 501 215 531 263
rect 602 215 632 269
rect 688 253 727 287
rect 761 253 804 287
rect 846 319 912 335
rect 846 285 862 319
rect 896 285 912 319
rect 846 269 912 285
rect 954 319 1020 335
rect 954 285 970 319
rect 1004 285 1020 319
rect 954 269 1020 285
rect 1062 303 1092 367
rect 1148 303 1178 367
rect 1062 287 1178 303
rect 688 237 804 253
rect 688 215 718 237
rect 774 215 804 237
rect 860 215 890 269
rect 976 215 1006 269
rect 1062 253 1102 287
rect 1136 253 1178 287
rect 1062 237 1178 253
rect 1062 215 1092 237
rect 1148 215 1178 237
rect 1234 308 1264 367
rect 1234 292 1323 308
rect 1234 258 1273 292
rect 1307 258 1323 292
rect 1234 242 1323 258
rect 1234 215 1264 242
rect 243 21 273 47
rect 329 21 359 47
rect 415 21 445 47
rect 501 21 531 47
rect 602 21 632 47
rect 688 21 718 47
rect 774 21 804 47
rect 860 21 890 47
rect 976 21 1006 47
rect 1062 21 1092 47
rect 1148 21 1178 47
rect 1234 21 1264 47
<< polycont >>
rect 119 279 153 313
rect 187 279 221 313
rect 255 279 289 313
rect 323 279 357 313
rect 391 279 425 313
rect 459 279 493 313
rect 596 285 630 319
rect 727 253 761 287
rect 862 285 896 319
rect 970 285 1004 319
rect 1102 253 1136 287
rect 1273 258 1307 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 92 607 158 649
rect 92 573 108 607
rect 142 573 158 607
rect 92 539 158 573
rect 92 505 108 539
rect 142 505 158 539
rect 92 453 158 505
rect 92 419 108 453
rect 142 419 158 453
rect 192 599 230 615
rect 192 565 194 599
rect 228 565 230 599
rect 192 516 230 565
rect 192 482 194 516
rect 228 482 230 516
rect 192 413 230 482
rect 264 607 330 649
rect 264 573 280 607
rect 314 573 330 607
rect 264 539 330 573
rect 264 505 280 539
rect 314 505 330 539
rect 264 453 330 505
rect 264 419 280 453
rect 314 419 330 453
rect 364 599 410 615
rect 364 565 366 599
rect 400 565 410 599
rect 364 516 410 565
rect 364 482 366 516
rect 400 482 410 516
rect 192 385 194 413
rect 20 379 194 385
rect 228 385 230 413
rect 364 413 410 482
rect 364 385 366 413
rect 228 379 366 385
rect 400 379 410 413
rect 20 351 410 379
rect 444 607 492 649
rect 444 573 452 607
rect 486 573 492 607
rect 444 510 492 573
rect 444 476 452 510
rect 486 476 492 510
rect 444 413 492 476
rect 541 599 959 615
rect 541 565 557 599
rect 591 581 729 599
rect 591 565 607 581
rect 541 495 607 565
rect 713 565 729 581
rect 763 581 909 599
rect 763 565 779 581
rect 541 461 557 495
rect 591 461 607 495
rect 641 531 679 547
rect 641 497 643 531
rect 677 497 679 531
rect 641 441 679 497
rect 713 495 779 565
rect 893 565 909 581
rect 943 565 959 599
rect 713 461 729 495
rect 763 461 779 495
rect 813 531 859 547
rect 813 497 815 531
rect 849 497 859 531
rect 641 427 643 441
rect 444 379 452 413
rect 486 379 492 413
rect 444 363 492 379
rect 526 407 643 427
rect 677 427 679 441
rect 813 443 859 497
rect 813 427 815 443
rect 677 409 815 427
rect 849 409 859 443
rect 677 407 859 409
rect 526 391 859 407
rect 893 513 959 565
rect 893 479 909 513
rect 943 479 959 513
rect 893 425 959 479
rect 993 607 1059 649
rect 993 573 1009 607
rect 1043 573 1059 607
rect 993 493 1059 573
rect 993 459 1009 493
rect 1043 459 1059 493
rect 1093 599 1139 615
rect 1093 565 1103 599
rect 1137 565 1139 599
rect 1093 513 1139 565
rect 1093 479 1103 513
rect 1137 479 1139 513
rect 1093 441 1139 479
rect 1173 607 1239 649
rect 1173 573 1189 607
rect 1223 573 1239 607
rect 1173 493 1239 573
rect 1173 459 1189 493
rect 1223 459 1239 493
rect 1273 599 1325 615
rect 1273 565 1275 599
rect 1309 565 1325 599
rect 1273 520 1325 565
rect 1273 486 1275 520
rect 1309 486 1325 520
rect 1093 425 1103 441
rect 893 391 909 425
rect 943 407 1103 425
rect 1137 425 1139 441
rect 1273 441 1325 486
rect 1273 425 1275 441
rect 1137 407 1275 425
rect 1309 407 1325 441
rect 943 391 1325 407
rect 20 243 69 351
rect 526 317 560 391
rect 103 313 560 317
rect 103 279 119 313
rect 153 279 187 313
rect 221 279 255 313
rect 289 279 323 313
rect 357 279 391 313
rect 425 279 459 313
rect 493 279 560 313
rect 103 277 560 279
rect 20 209 492 243
rect 20 65 85 209
rect 282 203 318 209
rect 182 141 198 175
rect 232 141 248 175
rect 182 93 248 141
rect 182 59 198 93
rect 232 59 248 93
rect 182 17 248 59
rect 282 169 284 203
rect 454 203 492 209
rect 282 101 318 169
rect 282 67 284 101
rect 282 51 318 67
rect 354 139 370 173
rect 404 139 420 173
rect 354 89 420 139
rect 354 55 370 89
rect 404 55 420 89
rect 354 17 420 55
rect 454 169 456 203
rect 490 169 492 203
rect 454 101 492 169
rect 526 206 560 277
rect 594 323 912 357
rect 594 319 646 323
rect 594 285 596 319
rect 630 285 646 319
rect 846 319 912 323
rect 594 269 646 285
rect 680 287 804 289
rect 680 253 727 287
rect 761 253 804 287
rect 846 285 862 319
rect 896 285 912 319
rect 846 269 912 285
rect 954 323 1323 357
rect 954 319 1020 323
rect 954 285 970 319
rect 1004 285 1020 319
rect 1257 292 1323 323
rect 954 269 1020 285
rect 1062 287 1223 289
rect 680 240 804 253
rect 1062 253 1102 287
rect 1136 253 1223 287
rect 1062 240 1223 253
rect 1257 258 1273 292
rect 1307 258 1323 292
rect 1257 242 1323 258
rect 526 202 1153 206
rect 526 168 729 202
rect 763 190 1153 202
rect 763 168 1103 190
rect 526 164 1103 168
rect 1097 156 1103 164
rect 1137 156 1153 190
rect 1097 140 1153 156
rect 1187 190 1233 206
rect 1187 156 1189 190
rect 1223 156 1233 190
rect 454 67 456 101
rect 490 67 492 101
rect 454 51 492 67
rect 526 96 542 130
rect 576 96 592 130
rect 526 17 592 96
rect 626 114 855 130
rect 626 80 643 114
rect 677 80 815 114
rect 849 80 855 114
rect 626 51 855 80
rect 889 114 955 130
rect 889 80 905 114
rect 939 80 955 114
rect 889 17 955 80
rect 1001 114 1063 130
rect 1001 80 1017 114
rect 1051 106 1063 114
rect 1187 106 1233 156
rect 1051 101 1233 106
rect 1051 80 1189 101
rect 1001 67 1189 80
rect 1223 67 1233 101
rect 1001 51 1233 67
rect 1267 190 1325 206
rect 1267 156 1275 190
rect 1309 156 1325 190
rect 1267 93 1325 156
rect 1267 59 1275 93
rect 1309 59 1325 93
rect 1267 17 1325 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a22o_4
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1131416
string GDS_START 1119984
<< end >>
