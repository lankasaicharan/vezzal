magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 332 1094 704
<< pwell >>
rect 288 49 1055 248
rect 0 0 1056 49
<< scpmos >>
rect 83 388 119 588
rect 173 388 209 588
rect 269 388 305 588
rect 359 388 395 588
rect 460 388 496 588
rect 560 388 596 588
rect 667 368 703 592
rect 757 368 793 592
rect 847 368 883 592
rect 937 368 973 592
<< nmoslvt >>
rect 371 74 401 222
rect 473 74 503 222
rect 571 74 601 222
rect 671 74 701 222
rect 758 74 788 222
rect 856 74 886 222
rect 942 74 972 222
<< ndiff >>
rect 314 188 371 222
rect 314 154 326 188
rect 360 154 371 188
rect 314 120 371 154
rect 314 86 326 120
rect 360 86 371 120
rect 314 74 371 86
rect 401 120 473 222
rect 401 86 426 120
rect 460 86 473 120
rect 401 74 473 86
rect 503 188 571 222
rect 503 154 526 188
rect 560 154 571 188
rect 503 120 571 154
rect 503 86 526 120
rect 560 86 571 120
rect 503 74 571 86
rect 601 120 671 222
rect 601 86 626 120
rect 660 86 671 120
rect 601 74 671 86
rect 701 210 758 222
rect 701 176 713 210
rect 747 176 758 210
rect 701 120 758 176
rect 701 86 713 120
rect 747 86 758 120
rect 701 74 758 86
rect 788 131 856 222
rect 788 97 799 131
rect 833 97 856 131
rect 788 74 856 97
rect 886 210 942 222
rect 886 176 897 210
rect 931 176 942 210
rect 886 120 942 176
rect 886 86 897 120
rect 931 86 942 120
rect 886 74 942 86
rect 972 139 1029 222
rect 972 105 983 139
rect 1017 105 1029 139
rect 972 74 1029 105
<< pdiff >>
rect 611 588 667 592
rect 27 576 83 588
rect 27 542 39 576
rect 73 542 83 576
rect 27 505 83 542
rect 27 471 39 505
rect 73 471 83 505
rect 27 434 83 471
rect 27 400 39 434
rect 73 400 83 434
rect 27 388 83 400
rect 119 576 173 588
rect 119 542 129 576
rect 163 542 173 576
rect 119 508 173 542
rect 119 474 129 508
rect 163 474 173 508
rect 119 440 173 474
rect 119 406 129 440
rect 163 406 173 440
rect 119 388 173 406
rect 209 576 269 588
rect 209 542 222 576
rect 256 542 269 576
rect 209 388 269 542
rect 305 437 359 588
rect 305 403 315 437
rect 349 403 359 437
rect 305 388 359 403
rect 395 576 460 588
rect 395 542 410 576
rect 444 542 460 576
rect 395 388 460 542
rect 496 576 560 588
rect 496 542 516 576
rect 550 542 560 576
rect 496 508 560 542
rect 496 474 516 508
rect 550 474 560 508
rect 496 388 560 474
rect 596 580 667 588
rect 596 546 623 580
rect 657 546 667 580
rect 596 508 667 546
rect 596 474 623 508
rect 657 474 667 508
rect 596 388 667 474
rect 617 368 667 388
rect 703 580 757 592
rect 703 546 713 580
rect 747 546 757 580
rect 703 497 757 546
rect 703 463 713 497
rect 747 463 757 497
rect 703 414 757 463
rect 703 380 713 414
rect 747 380 757 414
rect 703 368 757 380
rect 793 580 847 592
rect 793 546 803 580
rect 837 546 847 580
rect 793 478 847 546
rect 793 444 803 478
rect 837 444 847 478
rect 793 368 847 444
rect 883 580 937 592
rect 883 546 893 580
rect 927 546 937 580
rect 883 497 937 546
rect 883 463 893 497
rect 927 463 937 497
rect 883 414 937 463
rect 883 380 893 414
rect 927 380 937 414
rect 883 368 937 380
rect 973 580 1029 592
rect 973 546 983 580
rect 1017 546 1029 580
rect 973 478 1029 546
rect 973 444 983 478
rect 1017 444 1029 478
rect 973 368 1029 444
<< ndiffc >>
rect 326 154 360 188
rect 326 86 360 120
rect 426 86 460 120
rect 526 154 560 188
rect 526 86 560 120
rect 626 86 660 120
rect 713 176 747 210
rect 713 86 747 120
rect 799 97 833 131
rect 897 176 931 210
rect 897 86 931 120
rect 983 105 1017 139
<< pdiffc >>
rect 39 542 73 576
rect 39 471 73 505
rect 39 400 73 434
rect 129 542 163 576
rect 129 474 163 508
rect 129 406 163 440
rect 222 542 256 576
rect 315 403 349 437
rect 410 542 444 576
rect 516 542 550 576
rect 516 474 550 508
rect 623 546 657 580
rect 623 474 657 508
rect 713 546 747 580
rect 713 463 747 497
rect 713 380 747 414
rect 803 546 837 580
rect 803 444 837 478
rect 893 546 927 580
rect 893 463 927 497
rect 893 380 927 414
rect 983 546 1017 580
rect 983 444 1017 478
<< poly >>
rect 83 588 119 614
rect 173 588 209 614
rect 269 588 305 614
rect 359 588 395 614
rect 460 588 496 614
rect 560 588 596 614
rect 667 592 703 618
rect 757 592 793 618
rect 847 592 883 618
rect 937 592 973 618
rect 83 326 119 388
rect 173 356 209 388
rect 21 310 119 326
rect 21 276 37 310
rect 71 276 119 310
rect 161 340 227 356
rect 161 306 177 340
rect 211 306 227 340
rect 161 290 227 306
rect 269 301 305 388
rect 359 301 395 388
rect 460 356 496 388
rect 21 242 119 276
rect 269 267 395 301
rect 443 340 509 356
rect 443 306 459 340
rect 493 306 509 340
rect 560 310 596 388
rect 667 326 703 368
rect 757 326 793 368
rect 847 326 883 368
rect 937 326 973 368
rect 667 310 973 326
rect 443 290 509 306
rect 551 294 617 310
rect 269 248 401 267
rect 21 208 37 242
rect 71 208 119 242
rect 21 174 119 208
rect 21 140 37 174
rect 71 140 119 174
rect 21 106 119 140
rect 21 72 37 106
rect 71 72 119 106
rect 21 56 119 72
rect 210 237 401 248
rect 210 172 299 237
rect 371 222 401 237
rect 473 222 503 290
rect 551 260 567 294
rect 601 260 617 294
rect 667 276 683 310
rect 717 276 751 310
rect 785 276 819 310
rect 853 276 887 310
rect 921 276 973 310
rect 667 260 973 276
rect 551 244 617 260
rect 571 222 601 244
rect 671 222 701 260
rect 758 222 788 260
rect 856 222 886 260
rect 942 222 972 260
rect 210 138 226 172
rect 260 138 299 172
rect 210 104 299 138
rect 210 70 226 104
rect 260 70 299 104
rect 210 54 299 70
rect 371 48 401 74
rect 473 48 503 74
rect 571 48 601 74
rect 671 48 701 74
rect 758 48 788 74
rect 856 48 886 74
rect 942 48 972 74
<< polycont >>
rect 37 276 71 310
rect 177 306 211 340
rect 459 306 493 340
rect 37 208 71 242
rect 37 140 71 174
rect 37 72 71 106
rect 567 260 601 294
rect 683 276 717 310
rect 751 276 785 310
rect 819 276 853 310
rect 887 276 921 310
rect 226 138 260 172
rect 226 70 260 104
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 576 73 649
rect 23 542 39 576
rect 23 505 73 542
rect 23 471 39 505
rect 23 434 73 471
rect 23 400 39 434
rect 23 384 73 400
rect 113 576 163 592
rect 113 542 129 576
rect 203 576 466 592
rect 203 542 222 576
rect 256 542 410 576
rect 444 542 466 576
rect 500 576 566 592
rect 500 542 516 576
rect 550 542 566 576
rect 113 508 163 542
rect 500 508 566 542
rect 113 474 129 508
rect 163 474 516 508
rect 550 474 566 508
rect 113 440 163 474
rect 500 458 566 474
rect 607 580 673 649
rect 607 546 623 580
rect 657 546 673 580
rect 607 508 673 546
rect 607 474 623 508
rect 657 474 673 508
rect 607 458 673 474
rect 713 580 747 596
rect 713 497 747 546
rect 113 406 129 440
rect 113 390 163 406
rect 299 437 365 440
rect 299 403 315 437
rect 349 424 365 437
rect 349 403 679 424
rect 299 390 679 403
rect 121 340 509 356
rect 21 310 87 326
rect 21 276 37 310
rect 71 276 87 310
rect 121 306 177 340
rect 211 306 459 340
rect 493 306 509 340
rect 645 326 679 390
rect 713 414 747 463
rect 787 580 837 649
rect 787 546 803 580
rect 787 478 837 546
rect 787 444 803 478
rect 787 428 837 444
rect 877 580 943 596
rect 877 546 893 580
rect 927 546 943 580
rect 877 497 943 546
rect 877 463 893 497
rect 927 463 943 497
rect 877 414 943 463
rect 983 580 1033 649
rect 1017 546 1033 580
rect 983 478 1033 546
rect 1017 444 1033 478
rect 983 428 1033 444
rect 877 394 893 414
rect 747 380 893 394
rect 927 394 943 414
rect 927 380 1031 394
rect 713 360 1031 380
rect 645 310 937 326
rect 121 290 509 306
rect 551 294 611 310
rect 21 256 87 276
rect 551 260 567 294
rect 601 260 611 294
rect 551 256 611 260
rect 21 242 611 256
rect 21 208 37 242
rect 71 222 611 242
rect 645 276 683 310
rect 717 276 751 310
rect 785 276 819 310
rect 853 276 887 310
rect 921 276 937 310
rect 645 260 937 276
rect 71 208 87 222
rect 21 174 87 208
rect 645 188 679 260
rect 985 226 1031 360
rect 21 140 37 174
rect 71 140 87 174
rect 21 106 87 140
rect 21 72 37 106
rect 71 72 87 106
rect 21 56 87 72
rect 210 172 276 188
rect 210 138 226 172
rect 260 138 276 172
rect 210 104 276 138
rect 210 70 226 104
rect 260 70 276 104
rect 310 154 326 188
rect 360 154 526 188
rect 560 154 679 188
rect 713 210 1031 226
rect 747 192 897 210
rect 310 120 376 154
rect 510 120 576 154
rect 713 120 747 176
rect 881 176 897 192
rect 931 192 1031 210
rect 310 86 326 120
rect 360 86 376 120
rect 310 70 376 86
rect 410 86 426 120
rect 460 86 476 120
rect 210 54 276 70
rect 410 17 476 86
rect 510 86 526 120
rect 560 86 576 120
rect 510 70 576 86
rect 610 86 626 120
rect 660 86 676 120
rect 610 17 676 86
rect 713 70 747 86
rect 783 131 833 158
rect 783 97 799 131
rect 783 17 833 97
rect 881 120 931 176
rect 881 86 897 120
rect 881 70 931 86
rect 967 139 1033 158
rect 967 105 983 139
rect 1017 105 1033 139
rect 967 17 1033 105
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or3_4
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 2028882
string GDS_START 2019766
<< end >>
