magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 331 1478 704
<< pwell >>
rect 14 157 357 164
rect 934 157 1417 267
rect 14 49 1417 157
rect 0 0 1440 49
<< scnmos >>
rect 93 54 123 138
rect 244 54 274 138
rect 458 47 488 131
rect 544 47 574 131
rect 616 47 646 131
rect 724 47 754 131
rect 796 47 826 131
rect 1013 73 1043 241
rect 1085 73 1115 241
rect 1193 73 1223 241
rect 1302 73 1332 241
<< scpmoshvt >>
rect 93 475 123 603
rect 221 475 251 603
rect 436 479 466 607
rect 581 479 611 607
rect 653 479 683 607
rect 755 479 785 563
rect 833 479 863 563
rect 1013 367 1043 619
rect 1099 367 1129 619
rect 1238 367 1268 619
rect 1324 367 1354 619
<< ndiff >>
rect 40 113 93 138
rect 40 79 48 113
rect 82 79 93 113
rect 40 54 93 79
rect 123 113 244 138
rect 123 79 197 113
rect 231 79 244 113
rect 123 54 244 79
rect 274 116 331 138
rect 274 82 289 116
rect 323 82 331 116
rect 274 54 331 82
rect 401 101 458 131
rect 401 67 409 101
rect 443 67 458 101
rect 401 47 458 67
rect 488 91 544 131
rect 488 57 499 91
rect 533 57 544 91
rect 488 47 544 57
rect 574 47 616 131
rect 646 101 724 131
rect 646 67 679 101
rect 713 67 724 101
rect 646 47 724 67
rect 754 47 796 131
rect 826 95 900 131
rect 826 61 856 95
rect 890 61 900 95
rect 826 47 900 61
rect 960 217 1013 241
rect 960 183 968 217
rect 1002 183 1013 217
rect 960 119 1013 183
rect 960 85 968 119
rect 1002 85 1013 119
rect 960 73 1013 85
rect 1043 73 1085 241
rect 1115 208 1193 241
rect 1115 174 1137 208
rect 1171 174 1193 208
rect 1115 119 1193 174
rect 1115 85 1137 119
rect 1171 85 1193 119
rect 1115 73 1193 85
rect 1223 219 1302 241
rect 1223 185 1248 219
rect 1282 185 1302 219
rect 1223 119 1302 185
rect 1223 85 1248 119
rect 1282 85 1302 119
rect 1223 73 1302 85
rect 1332 229 1391 241
rect 1332 195 1347 229
rect 1381 195 1391 229
rect 1332 119 1391 195
rect 1332 85 1347 119
rect 1381 85 1391 119
rect 1332 73 1391 85
<< pdiff >>
rect 40 589 93 603
rect 40 555 48 589
rect 82 555 93 589
rect 40 521 93 555
rect 40 487 48 521
rect 82 487 93 521
rect 40 475 93 487
rect 123 591 221 603
rect 123 557 134 591
rect 168 557 221 591
rect 123 475 221 557
rect 251 527 316 603
rect 251 493 272 527
rect 306 493 316 527
rect 251 475 316 493
rect 383 527 436 607
rect 383 493 391 527
rect 425 493 436 527
rect 383 479 436 493
rect 466 599 581 607
rect 466 565 531 599
rect 565 565 581 599
rect 466 531 581 565
rect 466 497 531 531
rect 565 497 581 531
rect 466 479 581 497
rect 611 479 653 607
rect 683 563 733 607
rect 960 576 1013 619
rect 960 563 968 576
rect 683 525 755 563
rect 683 491 694 525
rect 728 491 755 525
rect 683 479 755 491
rect 785 479 833 563
rect 863 542 968 563
rect 1002 542 1013 576
rect 863 538 1013 542
rect 863 504 874 538
rect 908 504 1013 538
rect 863 479 1013 504
rect 960 367 1013 479
rect 1043 599 1099 619
rect 1043 565 1054 599
rect 1088 565 1099 599
rect 1043 506 1099 565
rect 1043 472 1054 506
rect 1088 472 1099 506
rect 1043 419 1099 472
rect 1043 385 1054 419
rect 1088 385 1099 419
rect 1043 367 1099 385
rect 1129 607 1238 619
rect 1129 573 1166 607
rect 1200 573 1238 607
rect 1129 493 1238 573
rect 1129 459 1166 493
rect 1200 459 1238 493
rect 1129 367 1238 459
rect 1268 599 1324 619
rect 1268 565 1279 599
rect 1313 565 1324 599
rect 1268 496 1324 565
rect 1268 462 1279 496
rect 1313 462 1324 496
rect 1268 413 1324 462
rect 1268 379 1279 413
rect 1313 379 1324 413
rect 1268 367 1324 379
rect 1354 607 1407 619
rect 1354 573 1365 607
rect 1399 573 1407 607
rect 1354 505 1407 573
rect 1354 471 1365 505
rect 1399 471 1407 505
rect 1354 413 1407 471
rect 1354 379 1365 413
rect 1399 379 1407 413
rect 1354 367 1407 379
<< ndiffc >>
rect 48 79 82 113
rect 197 79 231 113
rect 289 82 323 116
rect 409 67 443 101
rect 499 57 533 91
rect 679 67 713 101
rect 856 61 890 95
rect 968 183 1002 217
rect 968 85 1002 119
rect 1137 174 1171 208
rect 1137 85 1171 119
rect 1248 185 1282 219
rect 1248 85 1282 119
rect 1347 195 1381 229
rect 1347 85 1381 119
<< pdiffc >>
rect 48 555 82 589
rect 48 487 82 521
rect 134 557 168 591
rect 272 493 306 527
rect 391 493 425 527
rect 531 565 565 599
rect 531 497 565 531
rect 694 491 728 525
rect 968 542 1002 576
rect 874 504 908 538
rect 1054 565 1088 599
rect 1054 472 1088 506
rect 1054 385 1088 419
rect 1166 573 1200 607
rect 1166 459 1200 493
rect 1279 565 1313 599
rect 1279 462 1313 496
rect 1279 379 1313 413
rect 1365 573 1399 607
rect 1365 471 1399 505
rect 1365 379 1399 413
<< poly >>
rect 93 603 123 629
rect 221 603 251 629
rect 436 607 466 633
rect 581 607 611 633
rect 653 607 683 633
rect 1013 619 1043 645
rect 1099 619 1129 645
rect 1238 619 1268 645
rect 1324 619 1354 645
rect 755 563 785 589
rect 833 563 863 589
rect 93 294 123 475
rect 221 302 251 475
rect 436 443 466 479
rect 581 445 611 479
rect 293 427 466 443
rect 293 393 309 427
rect 343 413 466 427
rect 508 429 611 445
rect 343 393 359 413
rect 293 377 359 393
rect 508 395 524 429
rect 558 415 611 429
rect 558 395 574 415
rect 508 379 574 395
rect 93 278 168 294
rect 93 244 118 278
rect 152 244 168 278
rect 93 210 168 244
rect 93 176 118 210
rect 152 176 168 210
rect 93 160 168 176
rect 210 286 276 302
rect 210 252 226 286
rect 260 252 276 286
rect 210 218 276 252
rect 210 184 226 218
rect 260 184 276 218
rect 210 168 276 184
rect 329 287 359 377
rect 329 271 502 287
rect 329 237 452 271
rect 486 237 502 271
rect 329 203 502 237
rect 329 169 452 203
rect 486 169 502 203
rect 93 138 123 160
rect 244 138 274 168
rect 329 153 502 169
rect 458 131 488 153
rect 544 131 574 379
rect 653 333 683 479
rect 755 447 785 479
rect 833 447 863 479
rect 725 431 791 447
rect 725 397 741 431
rect 775 397 791 431
rect 725 381 791 397
rect 833 431 900 447
rect 833 397 850 431
rect 884 397 900 431
rect 833 381 900 397
rect 653 303 790 333
rect 724 275 790 303
rect 616 245 682 261
rect 616 211 632 245
rect 666 211 682 245
rect 616 195 682 211
rect 724 241 740 275
rect 774 241 790 275
rect 724 225 790 241
rect 616 131 646 195
rect 724 131 754 225
rect 833 183 863 381
rect 1013 339 1043 367
rect 941 333 1043 339
rect 905 317 1043 333
rect 1099 329 1129 367
rect 1238 335 1268 367
rect 905 283 921 317
rect 955 309 1043 317
rect 1085 313 1151 329
rect 955 283 971 309
rect 905 267 971 283
rect 1085 279 1101 313
rect 1135 279 1151 313
rect 796 153 863 183
rect 796 131 826 153
rect 93 28 123 54
rect 244 28 274 54
rect 915 51 945 267
rect 1013 241 1043 267
rect 1085 263 1151 279
rect 1193 319 1268 335
rect 1193 285 1209 319
rect 1243 299 1268 319
rect 1324 299 1354 367
rect 1243 285 1354 299
rect 1193 269 1354 285
rect 1085 241 1115 263
rect 1193 241 1223 269
rect 1302 241 1332 269
rect 1013 51 1043 73
rect 458 21 488 47
rect 544 21 574 47
rect 616 21 646 47
rect 724 21 754 47
rect 796 21 826 47
rect 915 21 1043 51
rect 1085 47 1115 73
rect 1193 47 1223 73
rect 1302 47 1332 73
<< polycont >>
rect 309 393 343 427
rect 524 395 558 429
rect 118 244 152 278
rect 118 176 152 210
rect 226 252 260 286
rect 226 184 260 218
rect 452 237 486 271
rect 452 169 486 203
rect 741 397 775 431
rect 850 397 884 431
rect 632 211 666 245
rect 740 241 774 275
rect 921 283 955 317
rect 1101 279 1135 313
rect 1209 285 1243 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 32 589 86 605
rect 32 555 48 589
rect 82 555 86 589
rect 32 521 86 555
rect 120 591 170 649
rect 120 557 134 591
rect 168 557 170 591
rect 120 539 170 557
rect 204 577 495 611
rect 32 487 48 521
rect 82 505 86 521
rect 204 505 238 577
rect 82 487 238 505
rect 32 471 238 487
rect 272 527 343 543
rect 306 493 343 527
rect 272 471 343 493
rect 32 113 82 471
rect 296 427 343 471
rect 32 79 48 113
rect 32 63 82 79
rect 116 278 176 424
rect 116 244 118 278
rect 152 244 176 278
rect 116 210 176 244
rect 116 176 118 210
rect 152 176 176 210
rect 116 163 176 176
rect 210 286 260 424
rect 210 252 226 286
rect 210 218 260 252
rect 210 184 226 218
rect 210 163 260 184
rect 296 393 309 427
rect 296 377 343 393
rect 377 527 427 543
rect 377 493 391 527
rect 425 493 427 527
rect 116 63 161 163
rect 296 132 330 377
rect 377 341 427 493
rect 461 445 495 577
rect 529 599 567 649
rect 529 565 531 599
rect 565 565 567 599
rect 529 531 567 565
rect 529 497 531 531
rect 565 497 567 531
rect 529 479 567 497
rect 601 565 814 599
rect 461 429 567 445
rect 461 395 524 429
rect 558 395 567 429
rect 461 379 567 395
rect 601 341 635 565
rect 195 113 235 129
rect 195 79 197 113
rect 231 79 235 113
rect 195 17 235 79
rect 285 116 330 132
rect 285 82 289 116
rect 323 82 330 116
rect 285 66 330 82
rect 364 307 635 341
rect 671 525 744 531
rect 671 491 694 525
rect 728 491 744 525
rect 671 481 744 491
rect 671 345 705 481
rect 780 447 814 565
rect 858 576 1010 649
rect 858 542 968 576
rect 1002 542 1010 576
rect 858 538 1010 542
rect 858 504 874 538
rect 908 526 1010 538
rect 1044 599 1094 615
rect 1044 565 1054 599
rect 1088 565 1094 599
rect 908 504 957 526
rect 858 488 957 504
rect 1044 506 1094 565
rect 1044 492 1054 506
rect 991 472 1054 492
rect 1088 472 1094 506
rect 991 447 1094 472
rect 1150 607 1216 649
rect 1150 573 1166 607
rect 1200 573 1216 607
rect 1150 493 1216 573
rect 1150 459 1166 493
rect 1200 459 1216 493
rect 1150 453 1216 459
rect 1277 599 1313 615
rect 1277 565 1279 599
rect 1277 496 1313 565
rect 1277 462 1279 496
rect 741 431 814 447
rect 775 397 814 431
rect 741 381 814 397
rect 848 431 1094 447
rect 848 397 850 431
rect 884 419 1094 431
rect 884 397 1054 419
rect 848 385 1054 397
rect 1088 385 1243 419
rect 848 381 1025 385
rect 671 317 955 345
rect 671 311 921 317
rect 364 107 402 307
rect 436 271 502 273
rect 436 237 452 271
rect 486 237 502 271
rect 436 203 502 237
rect 601 261 635 307
rect 894 283 921 311
rect 718 275 790 277
rect 601 245 682 261
rect 601 211 632 245
rect 666 211 682 245
rect 601 209 682 211
rect 718 241 740 275
rect 774 241 790 275
rect 718 225 790 241
rect 894 267 955 283
rect 436 169 452 203
rect 486 175 502 203
rect 718 175 752 225
rect 894 179 928 267
rect 991 233 1025 381
rect 1071 313 1135 351
rect 1071 279 1101 313
rect 1071 242 1135 279
rect 1193 319 1243 385
rect 1193 285 1209 319
rect 1193 269 1243 285
rect 1277 413 1313 462
rect 1277 379 1279 413
rect 1277 235 1313 379
rect 1347 607 1415 649
rect 1347 573 1365 607
rect 1399 573 1415 607
rect 1347 505 1415 573
rect 1347 471 1365 505
rect 1399 471 1415 505
rect 1347 413 1415 471
rect 1347 379 1365 413
rect 1399 379 1415 413
rect 1347 363 1415 379
rect 486 169 752 175
rect 436 141 752 169
rect 788 145 928 179
rect 962 217 1025 233
rect 962 183 968 217
rect 1002 183 1025 217
rect 1232 219 1313 235
rect 788 107 822 145
rect 962 119 1025 183
rect 364 101 459 107
rect 364 67 409 101
rect 443 67 459 101
rect 364 51 459 67
rect 493 91 549 107
rect 493 57 499 91
rect 533 57 549 91
rect 493 17 549 57
rect 663 101 822 107
rect 663 67 679 101
rect 713 67 822 101
rect 663 51 822 67
rect 856 95 896 111
rect 890 61 896 95
rect 962 85 968 119
rect 1002 85 1025 119
rect 962 69 1025 85
rect 1121 174 1137 208
rect 1171 174 1187 208
rect 1121 119 1187 174
rect 1121 85 1137 119
rect 1171 85 1187 119
rect 856 17 896 61
rect 1121 17 1187 85
rect 1232 185 1248 219
rect 1282 185 1313 219
rect 1232 119 1313 185
rect 1232 85 1248 119
rect 1282 85 1313 119
rect 1232 69 1313 85
rect 1347 229 1397 245
rect 1381 195 1397 229
rect 1347 119 1397 195
rect 1381 85 1397 119
rect 1347 17 1397 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrtp_2
flabel comment s 340 292 340 292 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1279 94 1313 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 168 1313 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 464 1313 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 538 1313 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1935352
string GDS_START 1922738
<< end >>
