magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 332 1382 704
<< pwell >>
rect 1 49 1338 228
rect 0 0 1344 49
<< scpmos >>
rect 83 392 119 592
rect 173 392 209 592
rect 269 392 305 592
rect 359 392 395 592
rect 571 392 607 592
rect 661 392 697 592
rect 751 392 787 592
rect 859 392 895 592
rect 949 392 985 592
rect 1045 392 1081 592
rect 1135 392 1171 592
rect 1225 392 1261 592
<< nmoslvt >>
rect 107 74 137 202
rect 193 74 223 202
rect 279 74 309 202
rect 365 74 395 202
rect 563 74 593 202
rect 649 74 679 202
rect 779 74 809 202
rect 865 74 895 202
rect 951 74 981 202
rect 1051 74 1081 202
rect 1139 74 1169 202
rect 1225 74 1255 202
<< ndiff >>
rect 27 115 107 202
rect 27 81 42 115
rect 76 81 107 115
rect 27 74 107 81
rect 137 121 193 202
rect 137 87 148 121
rect 182 87 193 121
rect 137 74 193 87
rect 223 190 279 202
rect 223 156 234 190
rect 268 156 279 190
rect 223 74 279 156
rect 309 156 365 202
rect 309 122 320 156
rect 354 122 365 156
rect 309 74 365 122
rect 395 188 452 202
rect 395 154 406 188
rect 440 154 452 188
rect 395 120 452 154
rect 395 86 406 120
rect 440 86 452 120
rect 395 74 452 86
rect 506 190 563 202
rect 506 156 518 190
rect 552 156 563 190
rect 506 120 563 156
rect 506 86 518 120
rect 552 86 563 120
rect 506 74 563 86
rect 593 127 649 202
rect 593 93 604 127
rect 638 93 649 127
rect 593 74 649 93
rect 679 82 779 202
rect 679 74 712 82
rect 27 69 92 74
rect 694 48 712 74
rect 746 74 779 82
rect 809 127 865 202
rect 809 93 820 127
rect 854 93 865 127
rect 809 74 865 93
rect 895 190 951 202
rect 895 156 906 190
rect 940 156 951 190
rect 895 120 951 156
rect 895 86 906 120
rect 940 86 951 120
rect 895 74 951 86
rect 981 184 1051 202
rect 981 150 993 184
rect 1027 150 1051 184
rect 981 116 1051 150
rect 981 82 993 116
rect 1027 82 1051 116
rect 981 74 1051 82
rect 1081 120 1139 202
rect 1081 86 1093 120
rect 1127 86 1139 120
rect 1081 74 1139 86
rect 1169 188 1225 202
rect 1169 154 1180 188
rect 1214 154 1225 188
rect 1169 116 1225 154
rect 1169 82 1180 116
rect 1214 82 1225 116
rect 1169 74 1225 82
rect 1255 190 1312 202
rect 1255 156 1266 190
rect 1300 156 1312 190
rect 1255 120 1312 156
rect 1255 86 1266 120
rect 1300 86 1312 120
rect 1255 74 1312 86
rect 746 48 764 74
rect 694 36 764 48
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 509 83 546
rect 27 475 39 509
rect 73 475 83 509
rect 27 438 83 475
rect 27 404 39 438
rect 73 404 83 438
rect 27 392 83 404
rect 119 584 173 592
rect 119 550 129 584
rect 163 550 173 584
rect 119 503 173 550
rect 119 469 129 503
rect 163 469 173 503
rect 119 392 173 469
rect 209 531 269 592
rect 209 497 222 531
rect 256 497 269 531
rect 209 435 269 497
rect 209 401 222 435
rect 256 401 269 435
rect 209 392 269 401
rect 305 584 359 592
rect 305 550 315 584
rect 349 550 359 584
rect 305 503 359 550
rect 305 469 315 503
rect 349 469 359 503
rect 305 392 359 469
rect 395 531 461 592
rect 395 497 415 531
rect 449 497 461 531
rect 395 451 461 497
rect 395 417 415 451
rect 449 417 461 451
rect 395 392 461 417
rect 515 531 571 592
rect 515 497 527 531
rect 561 497 571 531
rect 515 444 571 497
rect 515 410 527 444
rect 561 410 571 444
rect 515 392 571 410
rect 607 578 661 592
rect 607 544 617 578
rect 651 544 661 578
rect 607 392 661 544
rect 697 492 751 592
rect 697 458 707 492
rect 741 458 751 492
rect 697 392 751 458
rect 787 580 859 592
rect 787 546 806 580
rect 840 546 859 580
rect 787 392 859 546
rect 895 580 949 592
rect 895 546 905 580
rect 939 546 949 580
rect 895 510 949 546
rect 895 476 905 510
rect 939 476 949 510
rect 895 440 949 476
rect 895 406 905 440
rect 939 406 949 440
rect 895 392 949 406
rect 985 570 1045 592
rect 985 536 998 570
rect 1032 536 1045 570
rect 985 392 1045 536
rect 1081 580 1135 592
rect 1081 546 1091 580
rect 1125 546 1135 580
rect 1081 494 1135 546
rect 1081 460 1091 494
rect 1125 460 1135 494
rect 1081 392 1135 460
rect 1171 570 1225 592
rect 1171 536 1181 570
rect 1215 536 1225 570
rect 1171 392 1225 536
rect 1261 584 1317 592
rect 1261 550 1271 584
rect 1305 550 1317 584
rect 1261 508 1317 550
rect 1261 474 1271 508
rect 1305 474 1317 508
rect 1261 434 1317 474
rect 1261 400 1271 434
rect 1305 400 1317 434
rect 1261 392 1317 400
<< ndiffc >>
rect 42 81 76 115
rect 148 87 182 121
rect 234 156 268 190
rect 320 122 354 156
rect 406 154 440 188
rect 406 86 440 120
rect 518 156 552 190
rect 518 86 552 120
rect 604 93 638 127
rect 712 48 746 82
rect 820 93 854 127
rect 906 156 940 190
rect 906 86 940 120
rect 993 150 1027 184
rect 993 82 1027 116
rect 1093 86 1127 120
rect 1180 154 1214 188
rect 1180 82 1214 116
rect 1266 156 1300 190
rect 1266 86 1300 120
<< pdiffc >>
rect 39 546 73 580
rect 39 475 73 509
rect 39 404 73 438
rect 129 550 163 584
rect 129 469 163 503
rect 222 497 256 531
rect 222 401 256 435
rect 315 550 349 584
rect 315 469 349 503
rect 415 497 449 531
rect 415 417 449 451
rect 527 497 561 531
rect 527 410 561 444
rect 617 544 651 578
rect 707 458 741 492
rect 806 546 840 580
rect 905 546 939 580
rect 905 476 939 510
rect 905 406 939 440
rect 998 536 1032 570
rect 1091 546 1125 580
rect 1091 460 1125 494
rect 1181 536 1215 570
rect 1271 550 1305 584
rect 1271 474 1305 508
rect 1271 400 1305 434
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 269 592 305 618
rect 359 592 395 618
rect 571 592 607 618
rect 661 592 697 618
rect 751 592 787 618
rect 859 592 895 618
rect 949 592 985 618
rect 1045 592 1081 618
rect 1135 592 1171 618
rect 1225 592 1261 618
rect 83 299 119 392
rect 173 377 209 392
rect 173 347 223 377
rect 193 299 223 347
rect 269 299 305 392
rect 359 360 395 392
rect 571 360 607 392
rect 359 344 425 360
rect 359 310 375 344
rect 409 310 425 344
rect 83 283 151 299
rect 83 249 101 283
rect 135 249 151 283
rect 83 233 151 249
rect 193 283 309 299
rect 193 249 217 283
rect 251 249 309 283
rect 193 233 309 249
rect 107 202 137 233
rect 193 202 223 233
rect 279 202 309 233
rect 359 276 425 310
rect 535 344 607 360
rect 535 310 551 344
rect 585 310 607 344
rect 661 318 697 392
rect 751 318 787 392
rect 859 356 895 392
rect 949 356 985 392
rect 1045 356 1081 392
rect 1135 356 1171 392
rect 535 294 607 310
rect 649 302 787 318
rect 359 242 375 276
rect 409 242 425 276
rect 359 226 425 242
rect 365 202 395 226
rect 563 202 593 294
rect 649 268 697 302
rect 731 268 787 302
rect 829 340 895 356
rect 829 306 845 340
rect 879 306 895 340
rect 829 290 895 306
rect 937 340 1003 356
rect 937 306 953 340
rect 987 306 1003 340
rect 937 290 1003 306
rect 1045 340 1171 356
rect 1045 306 1077 340
rect 1111 306 1171 340
rect 1045 290 1171 306
rect 1225 356 1261 392
rect 1225 340 1291 356
rect 1225 306 1241 340
rect 1275 306 1291 340
rect 1225 290 1291 306
rect 649 252 787 268
rect 649 202 679 252
rect 757 248 787 252
rect 757 218 809 248
rect 779 202 809 218
rect 865 202 895 290
rect 951 202 981 290
rect 1051 202 1081 290
rect 1139 202 1169 290
rect 1225 202 1255 290
rect 107 48 137 74
rect 193 48 223 74
rect 279 48 309 74
rect 365 48 395 74
rect 563 48 593 74
rect 649 48 679 74
rect 779 48 809 74
rect 865 48 895 74
rect 951 48 981 74
rect 1051 48 1081 74
rect 1139 48 1169 74
rect 1225 48 1255 74
<< polycont >>
rect 375 310 409 344
rect 101 249 135 283
rect 217 249 251 283
rect 551 310 585 344
rect 375 242 409 276
rect 697 268 731 302
rect 845 306 879 340
rect 953 306 987 340
rect 1077 306 1111 340
rect 1241 306 1275 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 113 596 667 615
rect 17 580 73 596
rect 17 546 39 580
rect 17 509 73 546
rect 17 475 39 509
rect 17 438 73 475
rect 113 584 865 596
rect 113 550 129 584
rect 163 581 315 584
rect 163 550 179 581
rect 113 503 179 550
rect 299 550 315 581
rect 349 581 865 584
rect 349 550 365 581
rect 113 469 129 503
rect 163 469 179 503
rect 213 531 265 547
rect 213 497 222 531
rect 256 497 265 531
rect 17 404 39 438
rect 213 435 265 497
rect 299 503 365 550
rect 601 580 865 581
rect 601 578 806 580
rect 299 469 315 503
rect 349 469 365 503
rect 399 531 493 547
rect 399 497 415 531
rect 449 497 493 531
rect 399 451 493 497
rect 399 435 415 451
rect 73 404 222 435
rect 17 401 222 404
rect 256 417 415 435
rect 449 417 493 451
rect 256 401 493 417
rect 17 384 73 401
rect 17 199 51 384
rect 121 344 425 367
rect 121 333 375 344
rect 121 299 167 333
rect 359 310 375 333
rect 409 310 425 344
rect 85 283 167 299
rect 85 249 101 283
rect 135 249 167 283
rect 85 233 167 249
rect 201 283 267 299
rect 201 249 217 283
rect 251 249 267 283
rect 201 233 267 249
rect 359 276 425 310
rect 359 242 375 276
rect 409 242 425 276
rect 359 226 425 242
rect 459 260 493 401
rect 527 531 561 547
rect 601 544 617 578
rect 651 546 806 578
rect 840 546 865 580
rect 651 544 865 546
rect 601 530 865 544
rect 900 580 943 596
rect 900 546 905 580
rect 939 546 943 580
rect 601 526 667 530
rect 527 492 561 497
rect 900 510 943 546
rect 979 570 1051 649
rect 979 536 998 570
rect 1032 536 1051 570
rect 979 530 1051 536
rect 1085 580 1131 596
rect 1085 546 1091 580
rect 1125 546 1131 580
rect 900 492 905 510
rect 527 458 707 492
rect 741 476 905 492
rect 939 496 943 510
rect 1085 496 1131 546
rect 1165 570 1231 649
rect 1165 536 1181 570
rect 1215 536 1231 570
rect 1165 530 1231 536
rect 1267 584 1321 600
rect 1267 550 1271 584
rect 1305 550 1321 584
rect 1267 508 1321 550
rect 1267 496 1271 508
rect 939 494 1271 496
rect 939 476 1091 494
rect 741 460 1091 476
rect 1125 474 1271 494
rect 1305 474 1321 508
rect 1125 460 1321 474
rect 741 458 1321 460
rect 527 444 561 458
rect 889 440 955 458
rect 527 394 561 410
rect 613 390 855 424
rect 889 406 905 440
rect 939 406 955 440
rect 1255 434 1321 458
rect 889 390 955 406
rect 989 390 1211 424
rect 1255 400 1271 434
rect 1305 400 1321 434
rect 1255 390 1321 400
rect 613 360 647 390
rect 535 344 647 360
rect 821 356 855 390
rect 989 356 1023 390
rect 1177 356 1211 390
rect 535 310 551 344
rect 585 310 647 344
rect 535 294 647 310
rect 681 302 747 356
rect 681 268 697 302
rect 731 268 747 302
rect 821 340 895 356
rect 821 306 845 340
rect 879 306 895 340
rect 821 290 895 306
rect 937 340 1023 356
rect 937 306 953 340
rect 987 306 1023 340
rect 937 290 1023 306
rect 1061 340 1127 356
rect 1061 306 1077 340
rect 1111 306 1127 340
rect 1061 290 1127 306
rect 1177 340 1291 356
rect 1177 306 1241 340
rect 1275 306 1291 340
rect 1177 290 1291 306
rect 459 226 568 260
rect 681 252 747 268
rect 502 218 568 226
rect 890 222 1316 256
rect 890 218 943 222
rect 17 190 284 199
rect 17 165 234 190
rect 218 156 234 165
rect 268 156 284 190
rect 502 190 943 218
rect 318 156 356 177
rect 23 115 96 131
rect 318 122 320 156
rect 354 122 356 156
rect 23 81 42 115
rect 76 81 96 115
rect 23 17 96 81
rect 132 121 356 122
rect 132 87 148 121
rect 182 87 356 121
rect 132 70 356 87
rect 390 154 406 188
rect 440 154 456 188
rect 390 120 456 154
rect 390 86 406 120
rect 440 86 456 120
rect 390 17 456 86
rect 502 156 518 190
rect 552 184 906 190
rect 552 156 568 184
rect 502 120 568 156
rect 890 156 906 184
rect 940 156 943 190
rect 1264 190 1316 222
rect 502 86 518 120
rect 552 86 568 120
rect 502 70 568 86
rect 604 127 854 150
rect 638 116 820 127
rect 638 93 654 116
rect 604 70 654 93
rect 804 93 820 116
rect 690 48 712 82
rect 746 48 768 82
rect 804 70 854 93
rect 890 120 943 156
rect 890 86 906 120
rect 940 86 943 120
rect 890 70 943 86
rect 977 184 1180 188
rect 977 150 993 184
rect 1027 154 1180 184
rect 1214 154 1230 188
rect 1027 150 1043 154
rect 977 116 1043 150
rect 977 82 993 116
rect 1027 82 1043 116
rect 977 70 1043 82
rect 1077 86 1093 120
rect 1127 86 1143 120
rect 690 17 768 48
rect 1077 17 1143 86
rect 1180 116 1230 154
rect 1214 82 1230 116
rect 1180 66 1230 82
rect 1264 156 1266 190
rect 1300 156 1316 190
rect 1264 120 1316 156
rect 1264 86 1266 120
rect 1300 86 1316 120
rect 1264 70 1316 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a222oi_2
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 Y
port 11 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 Y
port 11 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 Y
port 11 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C2
port 6 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 1869024
string GDS_START 1857812
<< end >>
