magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3602 1975
<< nwell >>
rect -38 343 2342 704
rect -38 331 263 343
rect 1050 331 2342 343
<< pwell >>
rect 287 282 1037 301
rect 287 238 1394 282
rect 1770 241 2106 263
rect 1770 238 2303 241
rect 287 218 2303 238
rect 2 49 2303 218
rect 0 0 2304 49
<< scnmos >>
rect 81 108 111 192
rect 167 108 197 192
rect 393 191 423 275
rect 465 191 495 275
rect 573 191 603 275
rect 732 191 762 275
rect 818 191 848 275
rect 912 191 942 275
rect 1129 128 1159 256
rect 1215 128 1245 256
rect 1390 128 1420 212
rect 1462 128 1492 212
rect 1548 128 1578 212
rect 1620 128 1650 212
rect 1876 139 1906 223
rect 1993 69 2023 237
rect 2194 47 2224 215
<< scpmoshvt >>
rect 81 472 111 600
rect 167 472 197 600
rect 357 463 387 547
rect 471 463 501 547
rect 673 463 703 547
rect 759 463 789 547
rect 831 463 861 547
rect 941 463 971 547
rect 1131 379 1161 547
rect 1263 412 1293 580
rect 1368 472 1398 556
rect 1440 472 1470 556
rect 1596 472 1626 556
rect 1682 472 1712 556
rect 1876 487 1906 615
rect 2081 367 2111 619
rect 2178 367 2208 619
<< ndiff >>
rect 28 167 81 192
rect 28 133 36 167
rect 70 133 81 167
rect 28 108 81 133
rect 111 164 167 192
rect 111 130 122 164
rect 156 130 167 164
rect 111 108 167 130
rect 197 167 254 192
rect 197 133 212 167
rect 246 133 254 167
rect 197 108 254 133
rect 313 191 393 275
rect 423 191 465 275
rect 495 244 573 275
rect 495 210 518 244
rect 552 210 573 244
rect 495 191 573 210
rect 603 244 732 275
rect 603 210 687 244
rect 721 210 732 244
rect 603 191 732 210
rect 762 191 818 275
rect 848 191 912 275
rect 942 256 1011 275
rect 942 191 1129 256
rect 313 135 371 191
rect 313 101 325 135
rect 359 101 371 135
rect 313 86 371 101
rect 957 172 1129 191
rect 1049 128 1129 172
rect 1159 248 1215 256
rect 1159 214 1170 248
rect 1204 214 1215 248
rect 1159 128 1215 214
rect 1245 244 1368 256
rect 1245 210 1324 244
rect 1358 212 1368 244
rect 1796 229 1854 237
rect 1358 210 1390 212
rect 1245 176 1390 210
rect 1245 142 1324 176
rect 1358 142 1390 176
rect 1245 128 1390 142
rect 1420 128 1462 212
rect 1492 174 1548 212
rect 1492 140 1503 174
rect 1537 140 1548 174
rect 1492 128 1548 140
rect 1578 128 1620 212
rect 1650 187 1703 212
rect 1650 153 1661 187
rect 1695 153 1703 187
rect 1650 128 1703 153
rect 1796 195 1808 229
rect 1842 223 1854 229
rect 1928 223 1993 237
rect 1842 195 1876 223
rect 1796 139 1876 195
rect 1906 139 1993 223
rect 1049 108 1107 128
rect 1049 74 1061 108
rect 1095 74 1107 108
rect 1049 66 1107 74
rect 1928 89 1993 139
rect 1928 55 1936 89
rect 1970 69 1993 89
rect 2023 229 2080 237
rect 2023 195 2034 229
rect 2068 195 2080 229
rect 2023 69 2080 195
rect 2137 89 2194 215
rect 1970 55 1978 69
rect 1928 43 1978 55
rect 2137 55 2149 89
rect 2183 55 2194 89
rect 2137 47 2194 55
rect 2224 203 2277 215
rect 2224 169 2235 203
rect 2269 169 2277 203
rect 2224 101 2277 169
rect 2224 67 2235 101
rect 2269 67 2277 101
rect 2224 47 2277 67
<< pdiff >>
rect 28 588 81 600
rect 28 554 36 588
rect 70 554 81 588
rect 28 520 81 554
rect 28 486 36 520
rect 70 486 81 520
rect 28 472 81 486
rect 111 588 167 600
rect 111 554 122 588
rect 156 554 167 588
rect 111 520 167 554
rect 111 486 122 520
rect 156 486 167 520
rect 111 472 167 486
rect 197 588 250 600
rect 197 554 208 588
rect 242 554 250 588
rect 197 520 250 554
rect 402 567 456 583
rect 402 547 412 567
rect 197 486 208 520
rect 242 486 250 520
rect 197 472 250 486
rect 304 515 357 547
rect 304 481 312 515
rect 346 481 357 515
rect 304 463 357 481
rect 387 533 412 547
rect 446 547 456 567
rect 446 533 471 547
rect 387 463 471 533
rect 501 521 558 547
rect 501 487 512 521
rect 546 487 558 521
rect 501 463 558 487
rect 876 567 926 583
rect 1819 597 1876 615
rect 876 547 884 567
rect 618 521 673 547
rect 618 487 628 521
rect 662 487 673 521
rect 618 463 673 487
rect 703 524 759 547
rect 703 490 714 524
rect 748 490 759 524
rect 703 463 759 490
rect 789 463 831 547
rect 861 533 884 547
rect 918 547 926 567
rect 1183 566 1263 580
rect 1183 547 1191 566
rect 918 533 941 547
rect 861 463 941 533
rect 971 523 1024 547
rect 971 489 982 523
rect 1016 489 1024 523
rect 971 463 1024 489
rect 1078 498 1131 547
rect 1078 464 1086 498
rect 1120 464 1131 498
rect 1078 379 1131 464
rect 1161 532 1191 547
rect 1225 532 1263 566
rect 1161 498 1263 532
rect 1161 464 1191 498
rect 1225 464 1263 498
rect 1161 430 1263 464
rect 1161 396 1191 430
rect 1225 412 1263 430
rect 1293 567 1346 580
rect 1293 533 1304 567
rect 1338 556 1346 567
rect 1819 563 1831 597
rect 1865 563 1876 597
rect 1338 533 1368 556
rect 1293 472 1368 533
rect 1398 472 1440 556
rect 1470 531 1596 556
rect 1470 497 1481 531
rect 1515 497 1551 531
rect 1585 497 1596 531
rect 1470 472 1596 497
rect 1626 531 1682 556
rect 1626 497 1637 531
rect 1671 497 1682 531
rect 1626 472 1682 497
rect 1712 531 1765 556
rect 1712 497 1723 531
rect 1757 497 1765 531
rect 1712 472 1765 497
rect 1819 529 1876 563
rect 1819 495 1831 529
rect 1865 495 1876 529
rect 1819 487 1876 495
rect 1906 607 1963 615
rect 1906 573 1917 607
rect 1951 573 1963 607
rect 1906 535 1963 573
rect 1906 501 1917 535
rect 1951 501 1963 535
rect 1906 487 1963 501
rect 2028 599 2081 619
rect 2028 565 2036 599
rect 2070 565 2081 599
rect 2028 503 2081 565
rect 1293 458 1346 472
rect 1293 424 1304 458
rect 1338 424 1346 458
rect 1293 412 1346 424
rect 1225 396 1233 412
rect 1161 379 1233 396
rect 2028 469 2036 503
rect 2070 469 2081 503
rect 2028 421 2081 469
rect 2028 387 2036 421
rect 2070 387 2081 421
rect 2028 367 2081 387
rect 2111 607 2178 619
rect 2111 573 2129 607
rect 2163 573 2178 607
rect 2111 510 2178 573
rect 2111 476 2129 510
rect 2163 476 2178 510
rect 2111 414 2178 476
rect 2111 380 2129 414
rect 2163 380 2178 414
rect 2111 367 2178 380
rect 2208 599 2265 619
rect 2208 565 2223 599
rect 2257 565 2265 599
rect 2208 506 2265 565
rect 2208 472 2223 506
rect 2257 472 2265 506
rect 2208 414 2265 472
rect 2208 380 2223 414
rect 2257 380 2265 414
rect 2208 367 2265 380
<< ndiffc >>
rect 36 133 70 167
rect 122 130 156 164
rect 212 133 246 167
rect 518 210 552 244
rect 687 210 721 244
rect 325 101 359 135
rect 1170 214 1204 248
rect 1324 210 1358 244
rect 1324 142 1358 176
rect 1503 140 1537 174
rect 1661 153 1695 187
rect 1808 195 1842 229
rect 1061 74 1095 108
rect 1936 55 1970 89
rect 2034 195 2068 229
rect 2149 55 2183 89
rect 2235 169 2269 203
rect 2235 67 2269 101
<< pdiffc >>
rect 36 554 70 588
rect 36 486 70 520
rect 122 554 156 588
rect 122 486 156 520
rect 208 554 242 588
rect 208 486 242 520
rect 312 481 346 515
rect 412 533 446 567
rect 512 487 546 521
rect 628 487 662 521
rect 714 490 748 524
rect 884 533 918 567
rect 982 489 1016 523
rect 1086 464 1120 498
rect 1191 532 1225 566
rect 1191 464 1225 498
rect 1191 396 1225 430
rect 1304 533 1338 567
rect 1831 563 1865 597
rect 1481 497 1515 531
rect 1551 497 1585 531
rect 1637 497 1671 531
rect 1723 497 1757 531
rect 1831 495 1865 529
rect 1917 573 1951 607
rect 1917 501 1951 535
rect 2036 565 2070 599
rect 1304 424 1338 458
rect 2036 469 2070 503
rect 2036 387 2070 421
rect 2129 573 2163 607
rect 2129 476 2163 510
rect 2129 380 2163 414
rect 2223 565 2257 599
rect 2223 472 2257 506
rect 2223 380 2257 414
<< poly >>
rect 81 600 111 626
rect 167 615 1293 645
rect 1876 615 1906 641
rect 2081 619 2111 645
rect 2178 619 2208 645
rect 167 600 197 615
rect 357 547 387 573
rect 81 394 111 472
rect 167 457 197 472
rect 471 547 501 573
rect 167 436 228 457
rect 174 432 228 436
rect 178 430 228 432
rect 357 431 387 463
rect 471 431 501 463
rect 182 427 228 430
rect 186 424 228 427
rect 81 378 156 394
rect 81 344 106 378
rect 140 344 156 378
rect 81 328 156 344
rect 81 192 111 328
rect 198 280 228 424
rect 322 415 388 431
rect 322 381 338 415
rect 372 381 388 415
rect 322 347 388 381
rect 322 313 338 347
rect 372 327 388 347
rect 465 415 531 431
rect 465 381 481 415
rect 515 381 531 415
rect 465 347 531 381
rect 372 313 423 327
rect 322 297 423 313
rect 153 264 228 280
rect 393 275 423 297
rect 465 313 481 347
rect 515 313 531 347
rect 465 297 531 313
rect 465 275 495 297
rect 573 275 603 615
rect 673 547 703 573
rect 759 547 789 615
rect 831 547 861 573
rect 1263 580 1293 615
rect 941 547 971 573
rect 1131 547 1161 573
rect 673 389 703 463
rect 759 437 789 463
rect 831 394 861 463
rect 941 424 971 463
rect 912 408 994 424
rect 648 373 714 389
rect 648 339 664 373
rect 698 339 714 373
rect 648 323 714 339
rect 804 378 870 394
rect 804 344 820 378
rect 854 344 870 378
rect 804 328 870 344
rect 912 374 944 408
rect 978 374 994 408
rect 1368 556 1398 582
rect 1440 556 1470 582
rect 1596 556 1626 582
rect 1682 556 1712 582
rect 1263 386 1293 412
rect 912 358 994 374
rect 648 290 762 323
rect 732 275 762 290
rect 818 275 848 328
rect 912 275 942 358
rect 1131 344 1161 379
rect 1368 344 1398 472
rect 1068 328 1161 344
rect 1068 294 1084 328
rect 1118 294 1161 328
rect 1068 278 1161 294
rect 1215 328 1398 344
rect 1215 294 1256 328
rect 1290 314 1398 328
rect 1440 438 1470 472
rect 1596 440 1626 472
rect 1440 422 1506 438
rect 1440 388 1456 422
rect 1490 388 1506 422
rect 1440 354 1506 388
rect 1440 320 1456 354
rect 1490 320 1506 354
rect 1290 294 1306 314
rect 1440 304 1506 320
rect 1548 424 1626 440
rect 1548 390 1564 424
rect 1598 390 1626 424
rect 1548 374 1626 390
rect 1215 278 1306 294
rect 153 230 169 264
rect 203 230 228 264
rect 153 214 228 230
rect 167 192 197 214
rect 1129 256 1159 278
rect 1215 256 1245 278
rect 81 82 111 108
rect 167 51 197 108
rect 393 123 423 191
rect 465 165 495 191
rect 573 165 603 191
rect 732 165 762 191
rect 818 165 848 191
rect 912 123 942 191
rect 393 93 942 123
rect 1390 212 1420 238
rect 1462 212 1492 304
rect 1548 212 1578 374
rect 1682 300 1712 472
rect 1876 399 1906 487
rect 1620 284 1712 300
rect 1620 250 1636 284
rect 1670 250 1712 284
rect 1853 383 1919 399
rect 1853 349 1869 383
rect 1903 349 1919 383
rect 1853 315 1919 349
rect 2081 335 2111 367
rect 1853 281 1869 315
rect 1903 281 1919 315
rect 1853 265 1919 281
rect 1961 319 2111 335
rect 1961 285 1977 319
rect 2011 305 2111 319
rect 2011 285 2027 305
rect 2178 303 2208 367
rect 1961 269 2027 285
rect 2153 287 2224 303
rect 1620 234 1712 250
rect 1620 212 1650 234
rect 1876 223 1906 265
rect 1993 237 2023 269
rect 2153 253 2169 287
rect 2203 253 2224 287
rect 2153 237 2224 253
rect 1129 102 1159 128
rect 1215 102 1245 128
rect 1390 51 1420 128
rect 1462 102 1492 128
rect 1548 102 1578 128
rect 1620 102 1650 128
rect 1876 113 1906 139
rect 167 21 1420 51
rect 2194 215 2224 237
rect 1993 43 2023 69
rect 2194 21 2224 47
<< polycont >>
rect 106 344 140 378
rect 338 381 372 415
rect 338 313 372 347
rect 481 381 515 415
rect 481 313 515 347
rect 664 339 698 373
rect 820 344 854 378
rect 944 374 978 408
rect 1084 294 1118 328
rect 1256 294 1290 328
rect 1456 388 1490 422
rect 1456 320 1490 354
rect 1564 390 1598 424
rect 169 230 203 264
rect 1636 250 1670 284
rect 1869 349 1903 383
rect 1869 281 1903 315
rect 1977 285 2011 319
rect 2169 253 2203 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 20 588 72 604
rect 20 554 36 588
rect 70 554 72 588
rect 20 520 72 554
rect 20 486 36 520
rect 70 486 72 520
rect 20 280 72 486
rect 106 588 172 649
rect 106 554 122 588
rect 156 554 172 588
rect 106 520 172 554
rect 106 486 122 520
rect 156 486 172 520
rect 106 470 172 486
rect 206 588 270 604
rect 206 554 208 588
rect 242 554 270 588
rect 206 520 270 554
rect 394 567 464 649
rect 206 486 208 520
rect 242 486 270 520
rect 206 470 270 486
rect 106 378 183 436
rect 140 344 183 378
rect 106 316 183 344
rect 222 420 270 470
rect 304 515 346 547
rect 394 533 412 567
rect 446 533 464 567
rect 868 567 934 649
rect 304 481 312 515
rect 508 521 669 547
rect 508 499 512 521
rect 346 487 512 499
rect 546 487 628 521
rect 662 487 669 521
rect 346 481 669 487
rect 304 465 669 481
rect 703 524 793 547
rect 868 533 884 567
rect 918 533 934 567
rect 868 530 934 533
rect 703 490 714 524
rect 748 494 793 524
rect 970 523 1019 547
rect 970 494 982 523
rect 748 490 982 494
rect 703 489 982 490
rect 1016 489 1019 523
rect 703 474 1019 489
rect 551 460 669 465
rect 736 460 1019 474
rect 1070 498 1136 649
rect 1070 464 1086 498
rect 1120 464 1136 498
rect 319 424 372 431
rect 222 316 279 420
rect 20 264 207 280
rect 20 230 169 264
rect 203 230 207 264
rect 20 214 207 230
rect 20 167 86 214
rect 241 208 279 316
rect 353 415 372 424
rect 319 381 338 390
rect 319 347 372 381
rect 319 313 338 347
rect 319 290 372 313
rect 406 415 515 431
rect 406 381 481 415
rect 406 347 515 381
rect 406 313 481 347
rect 406 278 515 313
rect 551 423 630 460
rect 406 242 463 278
rect 551 244 585 423
rect 497 210 518 244
rect 552 210 585 244
rect 241 180 451 208
rect 497 196 585 210
rect 619 373 700 389
rect 619 339 664 373
rect 698 339 700 373
rect 619 323 700 339
rect 20 133 36 167
rect 70 133 86 167
rect 20 117 86 133
rect 120 164 162 180
rect 120 130 122 164
rect 156 130 162 164
rect 120 17 162 130
rect 196 174 451 180
rect 196 167 275 174
rect 196 133 212 167
rect 246 133 275 167
rect 409 160 451 174
rect 619 160 653 323
rect 736 260 772 460
rect 1070 448 1136 464
rect 1186 566 1229 582
rect 1186 532 1191 566
rect 1225 532 1229 566
rect 1186 498 1229 532
rect 1186 464 1191 498
rect 1225 464 1229 498
rect 1186 430 1229 464
rect 808 378 859 406
rect 808 344 820 378
rect 854 344 859 378
rect 929 408 980 424
rect 1186 414 1191 430
rect 929 390 944 408
rect 895 374 944 390
rect 978 374 980 408
rect 895 358 980 374
rect 1014 396 1191 414
rect 1225 396 1229 430
rect 1300 567 1364 583
rect 1300 533 1304 567
rect 1338 533 1364 567
rect 1300 458 1364 533
rect 1465 531 1599 649
rect 1465 497 1481 531
rect 1515 497 1551 531
rect 1585 497 1599 531
rect 1465 481 1599 497
rect 1633 531 1684 547
rect 1633 497 1637 531
rect 1671 497 1684 531
rect 1633 469 1684 497
rect 1718 531 1765 649
rect 1718 497 1723 531
rect 1757 497 1765 531
rect 1718 481 1765 497
rect 1799 597 1865 613
rect 1799 563 1831 597
rect 1799 529 1865 563
rect 1799 495 1831 529
rect 1901 607 1967 649
rect 1901 573 1917 607
rect 1951 573 1967 607
rect 1901 535 1967 573
rect 1901 501 1917 535
rect 1951 501 1967 535
rect 2034 599 2086 615
rect 2034 565 2036 599
rect 2070 565 2086 599
rect 2034 503 2086 565
rect 1300 424 1304 458
rect 1338 424 1364 458
rect 1300 408 1364 424
rect 1014 380 1229 396
rect 808 322 859 344
rect 1014 322 1048 380
rect 808 288 1048 322
rect 1082 328 1120 344
rect 1082 294 1084 328
rect 1118 294 1120 328
rect 687 252 772 260
rect 1082 252 1120 294
rect 1186 264 1220 380
rect 687 244 1120 252
rect 721 212 1120 244
rect 1154 248 1220 264
rect 1154 214 1170 248
rect 1204 214 1220 248
rect 1154 212 1220 214
rect 1254 328 1290 344
rect 1254 294 1256 328
rect 721 210 843 212
rect 687 194 843 210
rect 1254 178 1290 294
rect 908 160 1290 178
rect 409 144 1290 160
rect 1324 286 1364 408
rect 1440 422 1506 438
rect 1440 388 1456 422
rect 1490 388 1506 422
rect 1548 424 1614 440
rect 1548 390 1564 424
rect 1601 390 1614 424
rect 1548 388 1614 390
rect 1650 394 1684 469
rect 1799 467 1865 495
rect 2034 469 2036 503
rect 2070 469 2086 503
rect 1799 433 2000 467
rect 1440 354 1506 388
rect 1650 354 1758 394
rect 1440 320 1456 354
rect 1490 320 1758 354
rect 1324 284 1686 286
rect 1324 250 1636 284
rect 1670 250 1686 284
rect 1324 244 1364 250
rect 1358 210 1364 244
rect 1324 176 1364 210
rect 1575 238 1686 250
rect 196 117 275 133
rect 309 135 375 140
rect 309 101 325 135
rect 359 101 375 135
rect 409 126 951 144
rect 1358 142 1364 176
rect 1324 126 1364 142
rect 1499 174 1537 190
rect 1499 140 1503 174
rect 309 17 375 101
rect 1045 108 1111 110
rect 1045 74 1061 108
rect 1095 74 1111 108
rect 1045 17 1111 74
rect 1499 17 1537 140
rect 1575 103 1609 238
rect 1722 203 1758 320
rect 1799 250 1833 433
rect 1869 383 1928 399
rect 1903 349 1928 383
rect 1869 315 1928 349
rect 1903 281 1928 315
rect 1869 265 1928 281
rect 1966 335 2000 433
rect 2034 421 2086 469
rect 2034 387 2036 421
rect 2070 387 2086 421
rect 2034 369 2086 387
rect 1966 319 2011 335
rect 1966 285 1977 319
rect 1966 269 2011 285
rect 1645 187 1758 203
rect 1792 229 1833 250
rect 1792 195 1808 229
rect 1842 195 1858 229
rect 1792 193 1858 195
rect 1645 153 1661 187
rect 1695 153 1758 187
rect 1892 159 1928 265
rect 2045 233 2086 369
rect 2120 607 2173 649
rect 2120 573 2129 607
rect 2163 573 2173 607
rect 2120 510 2173 573
rect 2120 476 2129 510
rect 2163 476 2173 510
rect 2120 414 2173 476
rect 2120 380 2129 414
rect 2163 380 2173 414
rect 2120 364 2173 380
rect 2207 599 2287 615
rect 2207 565 2223 599
rect 2257 565 2287 599
rect 2207 506 2287 565
rect 2207 472 2223 506
rect 2257 472 2287 506
rect 2207 414 2287 472
rect 2207 380 2223 414
rect 2257 380 2287 414
rect 2207 364 2287 380
rect 2018 229 2086 233
rect 2018 195 2034 229
rect 2068 195 2086 229
rect 2018 193 2086 195
rect 2165 287 2203 303
rect 2165 253 2169 287
rect 2165 237 2203 253
rect 2165 159 2199 237
rect 2237 219 2287 364
rect 1645 137 1758 153
rect 1792 125 2199 159
rect 2233 203 2287 219
rect 2233 169 2235 203
rect 2269 169 2287 203
rect 1792 103 1826 125
rect 1575 69 1826 103
rect 2233 101 2287 169
rect 1920 89 1986 91
rect 1920 55 1936 89
rect 1970 55 1986 89
rect 1920 17 1986 55
rect 2133 89 2199 91
rect 2133 55 2149 89
rect 2183 55 2199 89
rect 2133 17 2199 55
rect 2233 67 2235 101
rect 2269 67 2287 101
rect 2233 51 2287 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 319 415 353 424
rect 319 390 338 415
rect 338 390 353 415
rect 895 390 929 424
rect 1567 390 1598 424
rect 1598 390 1601 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 683 2304 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2304 683
rect 0 617 2304 649
rect 307 424 365 430
rect 307 390 319 424
rect 353 421 365 424
rect 883 424 941 430
rect 883 421 895 424
rect 353 393 895 421
rect 353 390 365 393
rect 307 384 365 390
rect 883 390 895 393
rect 929 421 941 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 929 393 1567 421
rect 929 390 941 393
rect 883 384 941 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2304 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -49 2304 -17
<< labels >>
flabel pwell s 0 0 2304 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2304 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfrbp_1
flabel comment s 676 630 676 630 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 676 108 676 108 0 FreeSans 300 0 0 0 no_jumper_check
flabel comment s 676 36 676 36 0 FreeSans 300 0 0 0 no_jumper_check
flabel metal1 s 1567 390 1601 424 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 2304 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2304 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 464 2081 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 538 2081 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2239 94 2273 128 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2239 168 2273 202 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2239 242 2273 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2239 316 2273 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2239 390 2273 424 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2239 464 2273 498 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2239 538 2273 572 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2304 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry R90
string GDS_END 4505506
string GDS_START 4487018
<< end >>
