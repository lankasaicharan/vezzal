magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 459 243 1129 259
rect 11 49 1129 243
rect 0 0 1152 49
<< scnmos >>
rect 90 49 120 217
rect 176 49 206 217
rect 262 49 292 217
rect 348 49 378 217
rect 558 65 588 233
rect 644 65 674 233
rect 746 65 776 233
rect 848 65 878 233
rect 934 65 964 233
rect 1020 65 1050 233
<< scpmoshvt >>
rect 154 367 184 619
rect 240 367 270 619
rect 326 367 356 619
rect 412 367 442 619
rect 498 367 528 619
rect 584 367 614 619
rect 762 367 792 619
rect 848 367 878 619
rect 934 367 964 619
rect 1020 367 1050 619
<< ndiff >>
rect 37 177 90 217
rect 37 143 45 177
rect 79 143 90 177
rect 37 95 90 143
rect 37 61 45 95
rect 79 61 90 95
rect 37 49 90 61
rect 120 205 176 217
rect 120 171 131 205
rect 165 171 176 205
rect 120 101 176 171
rect 120 67 131 101
rect 165 67 176 101
rect 120 49 176 67
rect 206 177 262 217
rect 206 143 217 177
rect 251 143 262 177
rect 206 91 262 143
rect 206 57 217 91
rect 251 57 262 91
rect 206 49 262 57
rect 292 205 348 217
rect 292 171 303 205
rect 337 171 348 205
rect 292 101 348 171
rect 292 67 303 101
rect 337 67 348 101
rect 292 49 348 67
rect 378 181 431 217
rect 378 147 389 181
rect 423 147 431 181
rect 378 95 431 147
rect 378 61 389 95
rect 423 61 431 95
rect 485 179 558 233
rect 485 145 499 179
rect 533 145 558 179
rect 485 107 558 145
rect 485 73 499 107
rect 533 73 558 107
rect 485 65 558 73
rect 588 225 644 233
rect 588 191 599 225
rect 633 191 644 225
rect 588 153 644 191
rect 588 119 599 153
rect 633 119 644 153
rect 588 65 644 119
rect 674 181 746 233
rect 674 147 701 181
rect 735 147 746 181
rect 674 107 746 147
rect 674 73 701 107
rect 735 73 746 107
rect 674 65 746 73
rect 776 107 848 233
rect 776 73 801 107
rect 835 73 848 107
rect 776 65 848 73
rect 878 221 934 233
rect 878 187 889 221
rect 923 187 934 221
rect 878 111 934 187
rect 878 77 889 111
rect 923 77 934 111
rect 878 65 934 77
rect 964 183 1020 233
rect 964 149 975 183
rect 1009 149 1020 183
rect 964 107 1020 149
rect 964 73 975 107
rect 1009 73 1020 107
rect 964 65 1020 73
rect 1050 221 1103 233
rect 1050 187 1061 221
rect 1095 187 1103 221
rect 1050 111 1103 187
rect 1050 77 1061 111
rect 1095 77 1103 111
rect 1050 65 1103 77
rect 378 49 431 61
<< pdiff >>
rect 101 607 154 619
rect 101 573 109 607
rect 143 573 154 607
rect 101 530 154 573
rect 101 496 109 530
rect 143 496 154 530
rect 101 453 154 496
rect 101 419 109 453
rect 143 419 154 453
rect 101 367 154 419
rect 184 599 240 619
rect 184 565 195 599
rect 229 565 240 599
rect 184 507 240 565
rect 184 473 195 507
rect 229 473 240 507
rect 184 413 240 473
rect 184 379 195 413
rect 229 379 240 413
rect 184 367 240 379
rect 270 607 326 619
rect 270 573 281 607
rect 315 573 326 607
rect 270 530 326 573
rect 270 496 281 530
rect 315 496 326 530
rect 270 453 326 496
rect 270 419 281 453
rect 315 419 326 453
rect 270 367 326 419
rect 356 599 412 619
rect 356 565 367 599
rect 401 565 412 599
rect 356 507 412 565
rect 356 473 367 507
rect 401 473 412 507
rect 356 413 412 473
rect 356 379 367 413
rect 401 379 412 413
rect 356 367 412 379
rect 442 607 498 619
rect 442 573 453 607
rect 487 573 498 607
rect 442 493 498 573
rect 442 459 453 493
rect 487 459 498 493
rect 442 367 498 459
rect 528 599 584 619
rect 528 565 539 599
rect 573 565 584 599
rect 528 514 584 565
rect 528 480 539 514
rect 573 480 584 514
rect 528 436 584 480
rect 528 402 539 436
rect 573 402 584 436
rect 528 367 584 402
rect 614 611 762 619
rect 614 577 625 611
rect 659 577 717 611
rect 751 577 762 611
rect 614 521 762 577
rect 614 487 665 521
rect 699 487 762 521
rect 614 419 762 487
rect 614 385 665 419
rect 699 385 762 419
rect 614 367 762 385
rect 792 584 848 619
rect 792 550 803 584
rect 837 550 848 584
rect 792 367 848 550
rect 878 424 934 619
rect 878 390 889 424
rect 923 390 934 424
rect 878 367 934 390
rect 964 584 1020 619
rect 964 550 975 584
rect 1009 550 1020 584
rect 964 367 1020 550
rect 1050 607 1103 619
rect 1050 573 1061 607
rect 1095 573 1103 607
rect 1050 508 1103 573
rect 1050 474 1061 508
rect 1095 474 1103 508
rect 1050 413 1103 474
rect 1050 379 1061 413
rect 1095 379 1103 413
rect 1050 367 1103 379
<< ndiffc >>
rect 45 143 79 177
rect 45 61 79 95
rect 131 171 165 205
rect 131 67 165 101
rect 217 143 251 177
rect 217 57 251 91
rect 303 171 337 205
rect 303 67 337 101
rect 389 147 423 181
rect 389 61 423 95
rect 499 145 533 179
rect 499 73 533 107
rect 599 191 633 225
rect 599 119 633 153
rect 701 147 735 181
rect 701 73 735 107
rect 801 73 835 107
rect 889 187 923 221
rect 889 77 923 111
rect 975 149 1009 183
rect 975 73 1009 107
rect 1061 187 1095 221
rect 1061 77 1095 111
<< pdiffc >>
rect 109 573 143 607
rect 109 496 143 530
rect 109 419 143 453
rect 195 565 229 599
rect 195 473 229 507
rect 195 379 229 413
rect 281 573 315 607
rect 281 496 315 530
rect 281 419 315 453
rect 367 565 401 599
rect 367 473 401 507
rect 367 379 401 413
rect 453 573 487 607
rect 453 459 487 493
rect 539 565 573 599
rect 539 480 573 514
rect 539 402 573 436
rect 625 577 659 611
rect 717 577 751 611
rect 665 487 699 521
rect 665 385 699 419
rect 803 550 837 584
rect 889 390 923 424
rect 975 550 1009 584
rect 1061 573 1095 607
rect 1061 474 1095 508
rect 1061 379 1095 413
<< poly >>
rect 154 619 184 645
rect 240 619 270 645
rect 326 619 356 645
rect 412 619 442 645
rect 498 619 528 645
rect 584 619 614 645
rect 762 619 792 645
rect 848 619 878 645
rect 934 619 964 645
rect 1020 619 1050 645
rect 154 331 184 367
rect 240 331 270 367
rect 326 331 356 367
rect 412 331 442 367
rect 90 315 442 331
rect 90 281 120 315
rect 154 281 188 315
rect 222 281 256 315
rect 290 281 324 315
rect 358 281 392 315
rect 426 281 442 315
rect 90 265 442 281
rect 498 335 528 367
rect 584 335 614 367
rect 762 335 792 367
rect 498 319 674 335
rect 498 285 519 319
rect 553 285 587 319
rect 621 285 674 319
rect 498 269 674 285
rect 717 319 792 335
rect 717 285 733 319
rect 767 285 792 319
rect 717 269 792 285
rect 848 335 878 367
rect 934 335 964 367
rect 848 319 964 335
rect 848 285 905 319
rect 939 285 964 319
rect 848 269 964 285
rect 90 217 120 265
rect 176 217 206 265
rect 262 217 292 265
rect 348 217 378 265
rect 558 233 588 269
rect 644 233 674 269
rect 746 233 776 269
rect 848 233 878 269
rect 934 233 964 269
rect 1020 335 1050 367
rect 1020 319 1086 335
rect 1020 285 1036 319
rect 1070 285 1086 319
rect 1020 269 1086 285
rect 1020 233 1050 269
rect 90 23 120 49
rect 176 23 206 49
rect 262 23 292 49
rect 348 23 378 49
rect 558 39 588 65
rect 644 39 674 65
rect 746 39 776 65
rect 848 39 878 65
rect 934 39 964 65
rect 1020 39 1050 65
<< polycont >>
rect 120 281 154 315
rect 188 281 222 315
rect 256 281 290 315
rect 324 281 358 315
rect 392 281 426 315
rect 519 285 553 319
rect 587 285 621 319
rect 733 285 767 319
rect 905 285 939 319
rect 1036 285 1070 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 93 607 159 649
rect 93 573 109 607
rect 143 573 159 607
rect 93 530 159 573
rect 93 496 109 530
rect 143 496 159 530
rect 93 453 159 496
rect 93 419 109 453
rect 143 419 159 453
rect 193 599 231 615
rect 193 565 195 599
rect 229 565 231 599
rect 193 507 231 565
rect 193 473 195 507
rect 229 473 231 507
rect 193 413 231 473
rect 265 607 331 649
rect 265 573 281 607
rect 315 573 331 607
rect 265 530 331 573
rect 265 496 281 530
rect 315 496 331 530
rect 265 453 331 496
rect 265 419 281 453
rect 315 419 331 453
rect 365 599 401 615
rect 365 565 367 599
rect 365 507 401 565
rect 365 473 367 507
rect 193 385 195 413
rect 17 379 195 385
rect 229 385 231 413
rect 365 413 401 473
rect 437 607 503 649
rect 437 573 453 607
rect 487 573 503 607
rect 437 493 503 573
rect 437 459 453 493
rect 487 459 503 493
rect 437 454 503 459
rect 537 599 575 615
rect 537 565 539 599
rect 573 565 575 599
rect 537 514 575 565
rect 609 611 763 649
rect 609 577 625 611
rect 659 577 717 611
rect 751 577 763 611
rect 1059 607 1111 649
rect 609 561 763 577
rect 799 584 1013 600
rect 537 480 539 514
rect 573 480 575 514
rect 537 436 575 480
rect 537 420 539 436
rect 365 385 367 413
rect 229 379 367 385
rect 17 351 401 379
rect 435 402 539 420
rect 573 402 575 436
rect 435 386 575 402
rect 649 521 715 561
rect 799 550 803 584
rect 837 550 975 584
rect 1009 550 1013 584
rect 799 534 1013 550
rect 1059 573 1061 607
rect 1095 573 1111 607
rect 649 487 665 521
rect 699 487 715 521
rect 1059 508 1111 573
rect 649 419 715 487
rect 17 245 70 351
rect 435 317 469 386
rect 649 385 665 419
rect 699 385 715 419
rect 749 462 1025 500
rect 104 315 469 317
rect 104 281 120 315
rect 154 281 188 315
rect 222 281 256 315
rect 290 281 324 315
rect 358 281 392 315
rect 426 281 469 315
rect 503 319 637 352
rect 749 335 783 462
rect 503 285 519 319
rect 553 285 587 319
rect 621 285 637 319
rect 717 319 783 335
rect 717 285 733 319
rect 767 285 783 319
rect 817 424 939 428
rect 817 390 889 424
rect 923 390 939 424
rect 817 386 939 390
rect 104 279 469 281
rect 435 249 469 279
rect 817 249 853 386
rect 889 319 955 352
rect 889 285 905 319
rect 939 285 955 319
rect 991 329 1025 462
rect 1059 474 1061 508
rect 1095 474 1111 508
rect 1059 413 1111 474
rect 1059 379 1061 413
rect 1095 379 1111 413
rect 1059 363 1111 379
rect 991 319 1086 329
rect 991 285 1036 319
rect 1070 285 1086 319
rect 17 211 339 245
rect 435 225 853 249
rect 435 215 599 225
rect 129 205 167 211
rect 29 143 45 177
rect 79 143 95 177
rect 29 95 95 143
rect 29 61 45 95
rect 79 61 95 95
rect 29 17 95 61
rect 129 171 131 205
rect 165 171 167 205
rect 301 205 339 211
rect 129 101 167 171
rect 129 67 131 101
rect 165 67 167 101
rect 129 51 167 67
rect 201 143 217 177
rect 251 143 267 177
rect 201 91 267 143
rect 201 57 217 91
rect 251 57 267 91
rect 201 17 267 57
rect 301 171 303 205
rect 337 171 339 205
rect 583 191 599 215
rect 633 215 853 225
rect 887 221 1111 251
rect 633 191 649 215
rect 301 101 339 171
rect 301 67 303 101
rect 337 67 339 101
rect 301 51 339 67
rect 373 147 389 181
rect 423 147 439 181
rect 373 95 439 147
rect 373 61 389 95
rect 423 61 439 95
rect 373 17 439 61
rect 483 145 499 179
rect 533 145 549 179
rect 483 107 549 145
rect 583 153 649 191
rect 887 187 889 221
rect 923 217 1061 221
rect 923 187 925 217
rect 887 181 925 187
rect 1059 187 1061 217
rect 1095 187 1111 221
rect 583 119 599 153
rect 633 119 649 153
rect 685 147 701 181
rect 735 147 925 181
rect 483 73 499 107
rect 533 85 549 107
rect 685 107 751 147
rect 685 85 701 107
rect 533 73 701 85
rect 735 73 751 107
rect 483 51 751 73
rect 785 107 853 113
rect 785 73 801 107
rect 835 73 853 107
rect 785 17 853 73
rect 887 111 925 147
rect 887 77 889 111
rect 923 77 925 111
rect 887 61 925 77
rect 959 149 975 183
rect 1009 149 1025 183
rect 959 107 1025 149
rect 959 73 975 107
rect 1009 73 1025 107
rect 959 17 1025 73
rect 1059 111 1111 187
rect 1059 77 1061 111
rect 1095 77 1111 111
rect 1059 61 1111 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21a_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 464 929 498 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 464 1025 498 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 818702
string GDS_START 808832
<< end >>
