magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 437 165 863 185
rect 8 49 863 165
rect 0 0 864 49
<< scnmos >>
rect 91 55 121 139
rect 209 55 239 139
rect 317 55 347 139
rect 520 75 550 159
rect 592 75 622 159
rect 678 75 708 159
rect 750 75 780 159
<< scpmoshvt >>
rect 105 389 155 589
rect 203 389 253 589
rect 317 389 367 589
rect 455 389 505 589
rect 730 419 780 619
<< ndiff >>
rect 34 115 91 139
rect 34 81 46 115
rect 80 81 91 115
rect 34 55 91 81
rect 121 101 209 139
rect 121 67 148 101
rect 182 67 209 101
rect 121 55 209 67
rect 239 115 317 139
rect 239 81 250 115
rect 284 81 317 115
rect 239 55 317 81
rect 347 115 404 139
rect 347 81 358 115
rect 392 81 404 115
rect 347 55 404 81
rect 463 134 520 159
rect 463 100 475 134
rect 509 100 520 134
rect 463 75 520 100
rect 550 75 592 159
rect 622 134 678 159
rect 622 100 633 134
rect 667 100 678 134
rect 622 75 678 100
rect 708 75 750 159
rect 780 134 837 159
rect 780 100 791 134
rect 825 100 837 134
rect 780 75 837 100
<< pdiff >>
rect 382 607 440 619
rect 382 589 394 607
rect 48 577 105 589
rect 48 543 60 577
rect 94 543 105 577
rect 48 443 105 543
rect 48 409 60 443
rect 94 409 105 443
rect 48 389 105 409
rect 155 389 203 589
rect 253 577 317 589
rect 253 543 272 577
rect 306 543 317 577
rect 253 443 317 543
rect 253 409 272 443
rect 306 409 317 443
rect 253 389 317 409
rect 367 573 394 589
rect 428 589 440 607
rect 428 573 455 589
rect 367 389 455 573
rect 505 435 562 589
rect 505 401 516 435
rect 550 401 562 435
rect 505 389 562 401
rect 673 607 730 619
rect 673 573 685 607
rect 719 573 730 607
rect 673 419 730 573
rect 780 597 837 619
rect 780 563 791 597
rect 825 563 837 597
rect 780 465 837 563
rect 780 431 791 465
rect 825 431 837 465
rect 780 419 837 431
<< ndiffc >>
rect 46 81 80 115
rect 148 67 182 101
rect 250 81 284 115
rect 358 81 392 115
rect 475 100 509 134
rect 633 100 667 134
rect 791 100 825 134
<< pdiffc >>
rect 60 543 94 577
rect 60 409 94 443
rect 272 543 306 577
rect 272 409 306 443
rect 394 573 428 607
rect 516 401 550 435
rect 685 573 719 607
rect 791 563 825 597
rect 791 431 825 465
<< poly >>
rect 105 589 155 615
rect 203 589 253 615
rect 317 589 367 615
rect 455 604 630 634
rect 730 619 780 645
rect 455 589 505 604
rect 105 357 155 389
rect 44 341 155 357
rect 44 307 60 341
rect 94 307 155 341
rect 44 273 155 307
rect 44 239 60 273
rect 94 239 155 273
rect 44 223 155 239
rect 203 357 253 389
rect 203 341 269 357
rect 203 307 219 341
rect 253 307 269 341
rect 203 273 269 307
rect 317 315 367 389
rect 455 363 505 389
rect 600 349 630 604
rect 564 333 630 349
rect 730 333 780 419
rect 317 299 472 315
rect 317 285 422 299
rect 203 239 219 273
rect 253 239 269 273
rect 203 223 269 239
rect 406 265 422 285
rect 456 265 472 299
rect 406 231 472 265
rect 564 299 580 333
rect 614 299 630 333
rect 564 265 630 299
rect 564 245 580 265
rect 91 139 121 223
rect 209 139 239 223
rect 406 211 422 231
rect 317 197 422 211
rect 456 197 472 231
rect 317 181 472 197
rect 520 231 580 245
rect 614 231 630 265
rect 520 215 630 231
rect 678 317 780 333
rect 678 283 699 317
rect 733 283 780 317
rect 678 249 780 283
rect 678 215 699 249
rect 733 215 780 249
rect 317 139 347 181
rect 520 159 550 215
rect 592 159 622 215
rect 678 199 780 215
rect 678 159 708 199
rect 750 159 780 199
rect 91 29 121 55
rect 209 29 239 55
rect 317 29 347 55
rect 520 49 550 75
rect 592 49 622 75
rect 678 49 708 75
rect 750 49 780 75
<< polycont >>
rect 60 307 94 341
rect 60 239 94 273
rect 219 307 253 341
rect 219 239 253 273
rect 422 265 456 299
rect 580 299 614 333
rect 422 197 456 231
rect 580 231 614 265
rect 699 283 733 317
rect 699 215 733 249
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 44 577 110 649
rect 378 607 444 649
rect 44 543 60 577
rect 94 543 110 577
rect 44 443 110 543
rect 44 409 60 443
rect 94 409 110 443
rect 44 393 110 409
rect 256 577 336 593
rect 256 543 272 577
rect 306 543 336 577
rect 378 573 394 607
rect 428 573 444 607
rect 378 557 444 573
rect 669 607 735 649
rect 669 573 685 607
rect 719 573 735 607
rect 669 557 735 573
rect 775 597 841 613
rect 775 563 791 597
rect 825 563 841 597
rect 256 521 336 543
rect 256 487 717 521
rect 256 443 370 487
rect 256 409 272 443
rect 306 409 370 443
rect 256 393 370 409
rect 25 341 167 357
rect 25 307 60 341
rect 94 307 167 341
rect 25 273 167 307
rect 25 239 60 273
rect 94 239 167 273
rect 25 223 167 239
rect 203 341 269 357
rect 203 307 219 341
rect 253 307 269 341
rect 203 273 269 307
rect 203 239 219 273
rect 253 239 269 273
rect 203 223 269 239
rect 30 153 300 187
rect 30 115 96 153
rect 30 81 46 115
rect 80 81 96 115
rect 30 53 96 81
rect 132 101 198 117
rect 132 67 148 101
rect 182 67 198 101
rect 132 17 198 67
rect 234 115 300 153
rect 234 81 250 115
rect 284 81 300 115
rect 234 53 300 81
rect 336 143 370 393
rect 491 435 566 451
rect 491 401 516 435
rect 550 401 566 435
rect 491 385 566 401
rect 491 315 525 385
rect 406 299 525 315
rect 406 265 422 299
rect 456 265 525 299
rect 406 231 525 265
rect 406 197 422 231
rect 456 197 525 231
rect 564 333 647 349
rect 564 299 580 333
rect 614 299 647 333
rect 564 265 647 299
rect 564 231 580 265
rect 614 231 647 265
rect 564 215 647 231
rect 683 333 717 487
rect 775 465 841 563
rect 775 431 791 465
rect 825 431 841 465
rect 775 415 841 431
rect 683 317 749 333
rect 683 283 699 317
rect 733 283 749 317
rect 683 249 749 283
rect 683 215 699 249
rect 733 215 749 249
rect 683 199 749 215
rect 406 181 525 197
rect 336 115 408 143
rect 336 81 358 115
rect 392 81 408 115
rect 336 53 408 81
rect 459 134 525 181
rect 793 163 841 415
rect 459 100 475 134
rect 509 100 525 134
rect 459 71 525 100
rect 617 134 683 163
rect 617 100 633 134
rect 667 100 683 134
rect 617 17 683 100
rect 775 134 841 163
rect 775 100 791 134
rect 825 100 841 134
rect 775 71 841 100
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21ba_lp
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6534196
string GDS_START 6526524
<< end >>
