magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 383 1478 704
rect -38 364 1000 383
rect -38 331 348 364
rect 1296 331 1478 383
<< pwell >>
rect 450 235 560 313
rect 1042 235 1254 295
rect 450 157 1254 235
rect 3 49 1439 157
rect 0 0 1440 49
<< scnmos >>
rect 86 47 116 131
rect 158 47 188 131
rect 244 47 274 131
rect 316 47 346 131
rect 549 125 579 209
rect 635 125 665 209
rect 707 125 737 209
rect 793 125 823 209
rect 865 125 895 209
rect 951 125 981 209
rect 1023 125 1053 209
rect 1141 185 1171 269
rect 1254 47 1284 131
rect 1326 47 1356 131
<< scpmoshvt >>
rect 162 409 212 609
rect 268 409 318 609
rect 562 400 612 600
rect 654 400 704 600
rect 1026 419 1076 619
rect 1124 419 1174 619
rect 1234 419 1284 619
<< ndiff >>
rect 476 275 534 287
rect 476 241 488 275
rect 522 241 534 275
rect 476 209 534 241
rect 1068 257 1141 269
rect 1068 223 1080 257
rect 1114 223 1141 257
rect 1068 209 1141 223
rect 29 103 86 131
rect 29 69 41 103
rect 75 69 86 103
rect 29 47 86 69
rect 116 47 158 131
rect 188 98 244 131
rect 188 64 199 98
rect 233 64 244 98
rect 188 47 244 64
rect 274 47 316 131
rect 346 103 403 131
rect 476 125 549 209
rect 579 184 635 209
rect 579 150 590 184
rect 624 150 635 184
rect 579 125 635 150
rect 665 125 707 209
rect 737 171 793 209
rect 737 137 748 171
rect 782 137 793 171
rect 737 125 793 137
rect 823 125 865 209
rect 895 184 951 209
rect 895 150 906 184
rect 940 150 951 184
rect 895 125 951 150
rect 981 125 1023 209
rect 1053 185 1141 209
rect 1171 244 1228 269
rect 1171 210 1182 244
rect 1216 210 1228 244
rect 1171 185 1228 210
rect 1053 171 1126 185
rect 1053 137 1080 171
rect 1114 137 1126 171
rect 1053 125 1126 137
rect 346 69 357 103
rect 391 69 403 103
rect 346 47 403 69
rect 1197 106 1254 131
rect 1197 72 1209 106
rect 1243 72 1254 106
rect 1197 47 1254 72
rect 1284 47 1326 131
rect 1356 111 1413 131
rect 1356 77 1367 111
rect 1401 77 1413 111
rect 1356 47 1413 77
<< pdiff >>
rect 105 597 162 609
rect 105 563 117 597
rect 151 563 162 597
rect 105 515 162 563
rect 105 481 117 515
rect 151 481 162 515
rect 105 409 162 481
rect 212 597 268 609
rect 212 563 223 597
rect 257 563 268 597
rect 212 517 268 563
rect 212 483 223 517
rect 257 483 268 517
rect 212 409 268 483
rect 318 597 375 609
rect 318 563 329 597
rect 363 563 375 597
rect 318 526 375 563
rect 318 492 329 526
rect 363 492 375 526
rect 505 587 562 600
rect 505 553 517 587
rect 551 553 562 587
rect 318 455 375 492
rect 318 421 329 455
rect 363 421 375 455
rect 318 409 375 421
rect 505 400 562 553
rect 612 400 654 600
rect 704 446 761 600
rect 969 607 1026 619
rect 969 573 981 607
rect 1015 573 1026 607
rect 704 412 715 446
rect 749 412 761 446
rect 704 400 761 412
rect 969 419 1026 573
rect 1076 419 1124 619
rect 1174 604 1234 619
rect 1174 570 1185 604
rect 1219 570 1234 604
rect 1174 419 1234 570
rect 1284 597 1341 619
rect 1284 563 1295 597
rect 1329 563 1341 597
rect 1284 465 1341 563
rect 1284 431 1295 465
rect 1329 431 1341 465
rect 1284 419 1341 431
<< ndiffc >>
rect 488 241 522 275
rect 1080 223 1114 257
rect 41 69 75 103
rect 199 64 233 98
rect 590 150 624 184
rect 748 137 782 171
rect 906 150 940 184
rect 1182 210 1216 244
rect 1080 137 1114 171
rect 357 69 391 103
rect 1209 72 1243 106
rect 1367 77 1401 111
<< pdiffc >>
rect 117 563 151 597
rect 117 481 151 515
rect 223 563 257 597
rect 223 483 257 517
rect 329 563 363 597
rect 329 492 363 526
rect 517 553 551 587
rect 329 421 363 455
rect 981 573 1015 607
rect 715 412 749 446
rect 1185 570 1219 604
rect 1295 563 1329 597
rect 1295 431 1329 465
<< poly >>
rect 162 609 212 635
rect 268 609 318 635
rect 562 600 612 626
rect 654 615 901 645
rect 1026 619 1076 645
rect 1124 619 1174 645
rect 1234 619 1284 645
rect 654 600 704 615
rect 407 481 473 497
rect 407 447 423 481
rect 457 447 473 481
rect 407 413 473 447
rect 162 359 212 409
rect 268 361 318 409
rect 407 379 423 413
rect 457 385 473 413
rect 871 537 901 615
rect 871 521 937 537
rect 871 487 887 521
rect 921 487 937 521
rect 871 471 937 487
rect 871 413 937 429
rect 562 385 612 400
rect 457 379 612 385
rect 158 343 226 359
rect 158 309 176 343
rect 210 309 226 343
rect 158 275 226 309
rect 268 345 346 361
rect 407 355 612 379
rect 654 385 704 400
rect 654 355 823 385
rect 871 379 887 413
rect 921 393 937 413
rect 1026 393 1076 419
rect 921 379 1076 393
rect 871 363 1076 379
rect 1124 375 1174 419
rect 268 311 296 345
rect 330 311 346 345
rect 268 295 346 311
rect 158 255 176 275
rect 86 241 176 255
rect 210 241 226 275
rect 86 225 226 241
rect 86 131 116 225
rect 158 131 188 225
rect 316 176 346 295
rect 582 307 612 355
rect 244 146 346 176
rect 244 131 274 146
rect 316 131 346 146
rect 582 277 737 307
rect 549 209 579 235
rect 635 209 665 277
rect 707 209 737 277
rect 793 254 823 355
rect 951 254 981 363
rect 1118 359 1184 375
rect 1118 325 1134 359
rect 1168 325 1184 359
rect 1234 356 1284 419
rect 1118 309 1184 325
rect 1254 340 1356 356
rect 1141 269 1171 309
rect 1254 306 1295 340
rect 1329 306 1356 340
rect 1254 272 1356 306
rect 793 224 895 254
rect 793 209 823 224
rect 865 209 895 224
rect 951 224 1053 254
rect 951 209 981 224
rect 1023 209 1053 224
rect 1254 238 1295 272
rect 1329 238 1356 272
rect 1254 222 1356 238
rect 549 51 579 125
rect 635 99 665 125
rect 707 99 737 125
rect 793 99 823 125
rect 865 99 895 125
rect 951 99 981 125
rect 1023 99 1053 125
rect 1141 51 1171 185
rect 1254 131 1284 222
rect 1326 131 1356 222
rect 86 21 116 47
rect 158 21 188 47
rect 244 21 274 47
rect 316 21 346 47
rect 549 21 1171 51
rect 1254 21 1284 47
rect 1326 21 1356 47
<< polycont >>
rect 423 447 457 481
rect 423 379 457 413
rect 887 487 921 521
rect 176 309 210 343
rect 887 379 921 413
rect 296 311 330 345
rect 176 241 210 275
rect 1134 325 1168 359
rect 1295 306 1329 340
rect 1295 238 1329 272
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 25 597 167 613
rect 25 563 117 597
rect 151 563 167 597
rect 25 515 167 563
rect 25 481 117 515
rect 151 481 167 515
rect 25 465 167 481
rect 207 597 273 649
rect 207 563 223 597
rect 257 563 273 597
rect 207 517 273 563
rect 207 483 223 517
rect 257 483 273 517
rect 207 467 273 483
rect 313 597 379 613
rect 313 563 329 597
rect 363 563 379 597
rect 313 526 379 563
rect 501 587 981 607
rect 501 553 517 587
rect 551 573 981 587
rect 1015 573 1031 607
rect 1169 604 1235 649
rect 551 553 567 573
rect 501 552 567 553
rect 1169 570 1185 604
rect 1219 570 1235 604
rect 1169 551 1235 570
rect 1279 597 1345 613
rect 1279 563 1295 597
rect 1329 563 1345 597
rect 313 492 329 526
rect 363 497 379 526
rect 871 521 937 537
rect 363 492 473 497
rect 313 481 473 492
rect 25 119 65 465
rect 313 455 423 481
rect 313 431 329 455
rect 210 429 329 431
rect 101 421 329 429
rect 363 447 423 455
rect 457 447 473 481
rect 363 421 473 447
rect 101 413 473 421
rect 101 397 423 413
rect 101 395 244 397
rect 101 189 135 395
rect 407 379 423 397
rect 457 379 473 413
rect 407 363 473 379
rect 509 482 835 516
rect 171 343 226 359
rect 171 309 176 343
rect 210 309 226 343
rect 171 275 226 309
rect 280 345 359 361
rect 280 311 296 345
rect 330 311 359 345
rect 509 327 543 482
rect 280 295 359 311
rect 171 241 176 275
rect 210 259 226 275
rect 472 293 543 327
rect 699 412 715 446
rect 749 412 765 446
rect 472 275 538 293
rect 210 241 389 259
rect 171 225 389 241
rect 472 241 488 275
rect 522 241 538 275
rect 699 257 765 412
rect 801 327 835 482
rect 871 487 887 521
rect 921 515 937 521
rect 1279 515 1345 563
rect 921 487 1345 515
rect 871 481 1345 487
rect 871 471 937 481
rect 1279 465 1345 481
rect 871 413 937 430
rect 871 379 887 413
rect 921 379 937 413
rect 871 363 937 379
rect 973 411 1243 445
rect 1279 431 1295 465
rect 1329 449 1345 465
rect 1329 431 1417 449
rect 1279 415 1417 431
rect 973 327 1007 411
rect 801 293 1007 327
rect 1081 359 1173 375
rect 1081 325 1134 359
rect 1168 325 1173 359
rect 1081 309 1173 325
rect 1209 273 1243 411
rect 1064 257 1130 273
rect 472 225 538 241
rect 355 189 389 225
rect 574 223 868 257
rect 574 189 640 223
rect 101 155 319 189
rect 355 184 640 189
rect 834 213 868 223
rect 1064 223 1080 257
rect 1114 223 1130 257
rect 355 155 590 184
rect 285 119 319 155
rect 574 150 590 155
rect 624 150 640 184
rect 574 121 640 150
rect 732 171 798 187
rect 834 184 956 213
rect 834 179 906 184
rect 732 137 748 171
rect 782 137 798 171
rect 25 103 91 119
rect 25 69 41 103
rect 75 69 91 103
rect 25 53 91 69
rect 183 98 249 119
rect 183 64 199 98
rect 233 64 249 98
rect 183 17 249 64
rect 285 103 407 119
rect 285 69 357 103
rect 391 69 407 103
rect 285 53 407 69
rect 732 17 798 137
rect 890 150 906 179
rect 940 150 956 184
rect 890 121 956 150
rect 1064 171 1130 223
rect 1166 244 1243 273
rect 1166 210 1182 244
rect 1216 210 1243 244
rect 1279 340 1345 356
rect 1279 306 1295 340
rect 1329 306 1345 340
rect 1279 272 1345 306
rect 1279 238 1295 272
rect 1329 238 1345 272
rect 1279 222 1345 238
rect 1166 181 1243 210
rect 1064 137 1080 171
rect 1114 137 1130 171
rect 1064 17 1130 137
rect 1383 135 1417 415
rect 1193 106 1259 135
rect 1193 72 1209 106
rect 1243 72 1259 106
rect 1193 17 1259 72
rect 1351 111 1417 135
rect 1351 77 1367 111
rect 1401 77 1417 111
rect 1351 53 1417 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or4bb_lp
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6669272
string GDS_START 6658636
<< end >>
