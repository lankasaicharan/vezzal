magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 17 49 862 248
rect 0 0 864 49
<< scpmos >>
rect 90 368 126 592
rect 180 368 216 592
rect 283 392 319 592
rect 373 392 409 592
rect 567 392 603 592
rect 657 392 693 592
rect 747 392 783 592
<< nmoslvt >>
rect 96 74 126 222
rect 182 74 212 222
rect 307 74 337 222
rect 379 74 409 222
rect 573 74 603 222
rect 645 74 675 222
rect 753 74 783 222
<< ndiff >>
rect 43 142 96 222
rect 43 108 51 142
rect 85 108 96 142
rect 43 74 96 108
rect 126 210 182 222
rect 126 176 137 210
rect 171 176 182 210
rect 126 120 182 176
rect 126 86 137 120
rect 171 86 182 120
rect 126 74 182 86
rect 212 139 307 222
rect 212 105 242 139
rect 276 105 307 139
rect 212 74 307 105
rect 337 74 379 222
rect 409 210 573 222
rect 409 176 420 210
rect 454 176 528 210
rect 562 176 573 210
rect 409 120 573 176
rect 409 86 420 120
rect 454 86 528 120
rect 562 86 573 120
rect 409 74 573 86
rect 603 74 645 222
rect 675 127 753 222
rect 675 93 690 127
rect 724 93 753 127
rect 675 74 753 93
rect 783 202 836 222
rect 783 168 794 202
rect 828 168 836 202
rect 783 120 836 168
rect 783 86 794 120
rect 828 86 836 120
rect 783 74 836 86
<< pdiff >>
rect 38 580 90 592
rect 38 546 46 580
rect 80 546 90 580
rect 38 478 90 546
rect 38 444 46 478
rect 80 444 90 478
rect 38 368 90 444
rect 126 580 180 592
rect 126 546 136 580
rect 170 546 180 580
rect 126 497 180 546
rect 126 463 136 497
rect 170 463 180 497
rect 126 414 180 463
rect 126 380 136 414
rect 170 380 180 414
rect 126 368 180 380
rect 216 580 283 592
rect 216 546 226 580
rect 260 546 283 580
rect 216 510 283 546
rect 216 476 226 510
rect 260 476 283 510
rect 216 440 283 476
rect 216 406 226 440
rect 260 406 283 440
rect 216 392 283 406
rect 319 580 373 592
rect 319 546 329 580
rect 363 546 373 580
rect 319 510 373 546
rect 319 476 329 510
rect 363 476 373 510
rect 319 440 373 476
rect 319 406 329 440
rect 363 406 373 440
rect 319 392 373 406
rect 409 580 461 592
rect 409 546 419 580
rect 453 546 461 580
rect 409 492 461 546
rect 409 458 419 492
rect 453 458 461 492
rect 409 392 461 458
rect 515 530 567 592
rect 515 496 523 530
rect 557 496 567 530
rect 515 392 567 496
rect 603 547 657 592
rect 603 513 613 547
rect 647 513 657 547
rect 603 446 657 513
rect 603 412 613 446
rect 647 412 657 446
rect 603 392 657 412
rect 693 580 747 592
rect 693 546 703 580
rect 737 546 747 580
rect 693 462 747 546
rect 693 428 703 462
rect 737 428 747 462
rect 693 392 747 428
rect 783 580 835 592
rect 783 546 793 580
rect 827 546 835 580
rect 783 509 835 546
rect 783 475 793 509
rect 827 475 835 509
rect 783 438 835 475
rect 783 404 793 438
rect 827 404 835 438
rect 783 392 835 404
rect 216 368 268 392
<< ndiffc >>
rect 51 108 85 142
rect 137 176 171 210
rect 137 86 171 120
rect 242 105 276 139
rect 420 176 454 210
rect 528 176 562 210
rect 420 86 454 120
rect 528 86 562 120
rect 690 93 724 127
rect 794 168 828 202
rect 794 86 828 120
<< pdiffc >>
rect 46 546 80 580
rect 46 444 80 478
rect 136 546 170 580
rect 136 463 170 497
rect 136 380 170 414
rect 226 546 260 580
rect 226 476 260 510
rect 226 406 260 440
rect 329 546 363 580
rect 329 476 363 510
rect 329 406 363 440
rect 419 546 453 580
rect 419 458 453 492
rect 523 496 557 530
rect 613 513 647 547
rect 613 412 647 446
rect 703 546 737 580
rect 703 428 737 462
rect 793 546 827 580
rect 793 475 827 509
rect 793 404 827 438
<< poly >>
rect 90 592 126 618
rect 180 592 216 618
rect 283 592 319 618
rect 373 592 409 618
rect 567 592 603 618
rect 657 592 693 618
rect 747 592 783 618
rect 90 326 126 368
rect 180 326 216 368
rect 89 310 223 326
rect 283 318 319 392
rect 373 356 409 392
rect 567 356 603 392
rect 373 346 449 356
rect 379 340 449 346
rect 89 276 105 310
rect 139 276 173 310
rect 207 276 223 310
rect 89 260 223 276
rect 271 302 337 318
rect 271 268 287 302
rect 321 268 337 302
rect 96 222 126 260
rect 182 222 212 260
rect 271 252 337 268
rect 307 222 337 252
rect 379 306 399 340
rect 433 306 449 340
rect 379 290 449 306
rect 491 340 603 356
rect 491 306 507 340
rect 541 306 603 340
rect 657 310 693 392
rect 747 358 783 392
rect 753 310 783 358
rect 491 290 603 306
rect 379 222 409 290
rect 573 222 603 290
rect 645 294 711 310
rect 645 260 661 294
rect 695 260 711 294
rect 645 244 711 260
rect 753 294 839 310
rect 753 260 789 294
rect 823 260 839 294
rect 753 244 839 260
rect 645 222 675 244
rect 753 222 783 244
rect 96 48 126 74
rect 182 48 212 74
rect 307 48 337 74
rect 379 48 409 74
rect 573 48 603 74
rect 645 48 675 74
rect 753 48 783 74
<< polycont >>
rect 105 276 139 310
rect 173 276 207 310
rect 287 268 321 302
rect 399 306 433 340
rect 507 306 541 340
rect 661 260 695 294
rect 789 260 823 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 30 580 80 649
rect 30 546 46 580
rect 30 478 80 546
rect 30 444 46 478
rect 30 428 80 444
rect 120 580 186 596
rect 120 546 136 580
rect 170 546 186 580
rect 120 497 186 546
rect 120 463 136 497
rect 170 463 186 497
rect 120 414 186 463
rect 120 394 136 414
rect 20 380 136 394
rect 170 380 186 414
rect 226 580 276 649
rect 260 546 276 580
rect 226 510 276 546
rect 260 476 276 510
rect 226 440 276 476
rect 260 406 276 440
rect 226 390 276 406
rect 313 580 363 596
rect 313 546 329 580
rect 313 510 363 546
rect 313 476 329 510
rect 313 440 363 476
rect 403 580 469 649
rect 403 546 419 580
rect 453 546 469 580
rect 403 492 469 546
rect 403 458 419 492
rect 453 458 469 492
rect 507 581 737 615
rect 507 530 557 581
rect 703 580 737 581
rect 507 496 523 530
rect 507 480 557 496
rect 597 513 613 547
rect 647 513 663 547
rect 597 446 663 513
rect 313 406 329 440
rect 508 424 613 446
rect 363 412 613 424
rect 647 412 663 446
rect 703 462 737 546
rect 703 412 737 428
rect 777 580 843 596
rect 777 546 793 580
rect 827 546 843 580
rect 777 509 843 546
rect 777 475 793 509
rect 827 475 843 509
rect 777 438 843 475
rect 363 406 546 412
rect 313 390 546 406
rect 777 404 793 438
rect 827 404 843 438
rect 20 360 186 380
rect 777 378 843 404
rect 20 226 67 360
rect 105 310 239 326
rect 139 276 173 310
rect 207 276 239 310
rect 105 260 239 276
rect 20 210 171 226
rect 20 192 137 210
rect 121 176 137 192
rect 205 218 239 260
rect 273 302 353 356
rect 273 268 287 302
rect 321 268 353 302
rect 387 340 455 356
rect 387 306 399 340
rect 433 306 455 340
rect 387 290 455 306
rect 491 340 552 356
rect 491 306 507 340
rect 541 306 552 340
rect 491 290 552 306
rect 586 344 843 378
rect 273 252 353 268
rect 586 226 620 344
rect 654 294 739 310
rect 654 260 661 294
rect 695 260 739 294
rect 654 236 739 260
rect 773 294 839 310
rect 773 260 789 294
rect 823 260 839 294
rect 773 236 839 260
rect 404 218 620 226
rect 205 210 620 218
rect 205 184 420 210
rect 35 142 85 158
rect 35 108 51 142
rect 35 17 85 108
rect 121 120 171 176
rect 404 176 420 184
rect 454 176 528 210
rect 562 202 620 210
rect 562 176 794 202
rect 404 168 794 176
rect 828 168 844 202
rect 121 86 137 120
rect 121 70 171 86
rect 207 139 312 150
rect 207 105 242 139
rect 276 105 312 139
rect 207 17 312 105
rect 404 120 578 168
rect 404 86 420 120
rect 454 86 528 120
rect 562 86 578 120
rect 404 70 578 86
rect 670 127 744 134
rect 670 93 690 127
rect 724 93 744 127
rect 670 17 744 93
rect 778 120 844 168
rect 778 86 794 120
rect 828 86 844 120
rect 778 70 844 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a221o_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 3890770
string GDS_START 3882660
<< end >>
