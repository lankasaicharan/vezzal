magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 765 219
rect 0 0 768 49
<< scnmos >>
rect 84 109 114 193
rect 156 109 186 193
rect 242 109 272 193
rect 320 109 350 193
rect 422 109 452 193
rect 494 109 524 193
rect 580 109 610 193
rect 652 109 682 193
<< scpmoshvt >>
rect 136 409 186 609
rect 250 409 300 609
rect 348 409 398 609
rect 632 409 682 609
<< ndiff >>
rect 27 168 84 193
rect 27 134 39 168
rect 73 134 84 168
rect 27 109 84 134
rect 114 109 156 193
rect 186 168 242 193
rect 186 134 197 168
rect 231 134 242 168
rect 186 109 242 134
rect 272 109 320 193
rect 350 177 422 193
rect 350 143 361 177
rect 395 143 422 177
rect 350 109 422 143
rect 452 109 494 193
rect 524 168 580 193
rect 524 134 535 168
rect 569 134 580 168
rect 524 109 580 134
rect 610 109 652 193
rect 682 168 739 193
rect 682 134 693 168
rect 727 134 739 168
rect 682 109 739 134
<< pdiff >>
rect 79 597 136 609
rect 79 563 91 597
rect 125 563 136 597
rect 79 526 136 563
rect 79 492 91 526
rect 125 492 136 526
rect 79 455 136 492
rect 79 421 91 455
rect 125 421 136 455
rect 79 409 136 421
rect 186 597 250 609
rect 186 563 197 597
rect 231 563 250 597
rect 186 526 250 563
rect 186 492 197 526
rect 231 492 250 526
rect 186 455 250 492
rect 186 421 197 455
rect 231 421 250 455
rect 186 409 250 421
rect 300 409 348 609
rect 398 597 455 609
rect 398 563 409 597
rect 443 563 455 597
rect 398 526 455 563
rect 398 492 409 526
rect 443 492 455 526
rect 398 455 455 492
rect 398 421 409 455
rect 443 421 455 455
rect 398 409 455 421
rect 575 597 632 609
rect 575 563 587 597
rect 621 563 632 597
rect 575 526 632 563
rect 575 492 587 526
rect 621 492 632 526
rect 575 455 632 492
rect 575 421 587 455
rect 621 421 632 455
rect 575 409 632 421
rect 682 597 739 609
rect 682 563 693 597
rect 727 563 739 597
rect 682 526 739 563
rect 682 492 693 526
rect 727 492 739 526
rect 682 455 739 492
rect 682 421 693 455
rect 727 421 739 455
rect 682 409 739 421
<< ndiffc >>
rect 39 134 73 168
rect 197 134 231 168
rect 361 143 395 177
rect 535 134 569 168
rect 693 134 727 168
<< pdiffc >>
rect 91 563 125 597
rect 91 492 125 526
rect 91 421 125 455
rect 197 563 231 597
rect 197 492 231 526
rect 197 421 231 455
rect 409 563 443 597
rect 409 492 443 526
rect 409 421 443 455
rect 587 563 621 597
rect 587 492 621 526
rect 587 421 621 455
rect 693 563 727 597
rect 693 492 727 526
rect 693 421 727 455
<< poly >>
rect 136 609 186 635
rect 250 609 300 635
rect 348 609 398 635
rect 632 609 682 635
rect 136 369 186 409
rect 84 353 186 369
rect 250 367 300 409
rect 84 319 117 353
rect 151 319 186 353
rect 84 303 186 319
rect 234 351 300 367
rect 234 317 250 351
rect 284 317 300 351
rect 84 238 114 303
rect 234 283 300 317
rect 348 341 398 409
rect 632 369 682 409
rect 580 353 682 369
rect 348 311 452 341
rect 234 249 250 283
rect 284 263 300 283
rect 404 299 452 311
rect 580 319 603 353
rect 637 319 682 353
rect 404 283 538 299
rect 284 249 350 263
rect 84 208 186 238
rect 234 233 350 249
rect 404 249 420 283
rect 454 249 488 283
rect 522 249 538 283
rect 404 233 538 249
rect 580 285 682 319
rect 580 251 603 285
rect 637 251 682 285
rect 580 235 682 251
rect 84 193 114 208
rect 156 193 186 208
rect 242 193 272 233
rect 320 193 350 233
rect 422 193 452 233
rect 494 193 524 233
rect 580 193 610 235
rect 652 193 682 235
rect 84 83 114 109
rect 156 83 186 109
rect 242 83 272 109
rect 320 83 350 109
rect 422 83 452 109
rect 494 83 524 109
rect 580 83 610 109
rect 652 83 682 109
<< polycont >>
rect 117 319 151 353
rect 250 317 284 351
rect 250 249 284 283
rect 603 319 637 353
rect 420 249 454 283
rect 488 249 522 283
rect 603 251 637 285
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 23 597 125 613
rect 23 563 91 597
rect 23 526 125 563
rect 23 492 91 526
rect 23 455 125 492
rect 23 421 91 455
rect 23 405 125 421
rect 181 597 247 649
rect 181 563 197 597
rect 231 563 247 597
rect 181 526 247 563
rect 181 492 197 526
rect 231 492 247 526
rect 181 455 247 492
rect 181 421 197 455
rect 231 421 247 455
rect 181 405 247 421
rect 339 597 459 613
rect 339 563 409 597
rect 443 563 459 597
rect 339 526 459 563
rect 339 492 409 526
rect 443 492 459 526
rect 339 455 459 492
rect 339 421 409 455
rect 443 421 459 455
rect 23 267 57 405
rect 339 369 459 421
rect 571 597 637 649
rect 571 563 587 597
rect 621 563 637 597
rect 571 526 637 563
rect 571 492 587 526
rect 621 492 637 526
rect 571 455 637 492
rect 571 421 587 455
rect 621 421 637 455
rect 571 405 637 421
rect 677 597 743 613
rect 677 563 693 597
rect 727 563 743 597
rect 677 526 743 563
rect 677 492 693 526
rect 727 492 743 526
rect 677 455 743 492
rect 677 421 693 455
rect 727 421 743 455
rect 677 405 743 421
rect 101 353 167 369
rect 101 319 117 353
rect 151 319 167 353
rect 101 303 167 319
rect 234 351 300 367
rect 234 317 250 351
rect 284 317 300 351
rect 234 283 300 317
rect 234 267 250 283
rect 23 249 250 267
rect 284 249 300 283
rect 23 233 300 249
rect 339 353 653 369
rect 339 335 603 353
rect 23 168 89 233
rect 339 197 373 335
rect 587 319 603 335
rect 637 319 653 353
rect 409 283 551 299
rect 409 249 420 283
rect 454 249 488 283
rect 522 249 551 283
rect 409 233 551 249
rect 587 285 653 319
rect 587 251 603 285
rect 637 251 653 285
rect 587 235 653 251
rect 687 197 743 405
rect 23 134 39 168
rect 73 134 89 168
rect 23 105 89 134
rect 151 168 277 197
rect 151 134 197 168
rect 231 134 277 168
rect 151 128 277 134
rect 151 94 161 128
rect 195 94 233 128
rect 267 94 277 128
rect 339 177 411 197
rect 339 143 361 177
rect 395 143 411 177
rect 339 123 411 143
rect 489 168 615 197
rect 489 134 535 168
rect 569 134 615 168
rect 489 128 615 134
rect 151 87 277 94
rect 489 94 499 128
rect 533 94 571 128
rect 605 94 615 128
rect 677 168 743 197
rect 677 134 693 168
rect 727 134 743 168
rect 677 105 743 134
rect 489 87 615 94
rect 151 53 615 87
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 161 94 195 128
rect 233 94 267 128
rect 499 94 533 128
rect 571 94 605 128
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 14 128 754 134
rect 14 94 161 128
rect 195 94 233 128
rect 267 94 499 128
rect 533 94 571 128
rect 605 94 754 128
rect 14 88 754 94
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 iso1n_lp2
flabel metal1 s 14 88 754 134 0 FreeSans 340 0 0 0 KAGND
port 3 nsew ground input
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SLEEP_B
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2848660
string GDS_START 2841500
<< end >>
