magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 2 49 571 241
rect 0 0 576 49
<< scnmos >>
rect 81 47 111 215
rect 239 47 269 215
rect 348 47 378 215
rect 462 47 492 215
<< scpmoshvt >>
rect 80 367 110 619
rect 270 367 300 619
rect 356 367 386 619
rect 462 367 492 619
<< ndiff >>
rect 28 203 81 215
rect 28 169 36 203
rect 70 169 81 203
rect 28 101 81 169
rect 28 67 36 101
rect 70 67 81 101
rect 28 47 81 67
rect 111 163 239 215
rect 111 129 122 163
rect 156 129 194 163
rect 228 129 239 163
rect 111 89 239 129
rect 111 55 122 89
rect 156 55 194 89
rect 228 55 239 89
rect 111 47 239 55
rect 269 203 348 215
rect 269 169 294 203
rect 328 169 348 203
rect 269 101 348 169
rect 269 67 294 101
rect 328 67 348 101
rect 269 47 348 67
rect 378 47 462 215
rect 492 203 545 215
rect 492 169 503 203
rect 537 169 545 203
rect 492 93 545 169
rect 492 59 503 93
rect 537 59 545 93
rect 492 47 545 59
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 504 80 565
rect 27 470 35 504
rect 69 470 80 504
rect 27 413 80 470
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 607 163 619
rect 110 573 121 607
rect 155 573 163 607
rect 110 488 163 573
rect 110 454 121 488
rect 155 454 163 488
rect 110 367 163 454
rect 217 599 270 619
rect 217 565 225 599
rect 259 565 270 599
rect 217 518 270 565
rect 217 484 225 518
rect 259 484 270 518
rect 217 434 270 484
rect 217 400 225 434
rect 259 400 270 434
rect 217 367 270 400
rect 300 599 356 619
rect 300 565 311 599
rect 345 565 356 599
rect 300 508 356 565
rect 300 474 311 508
rect 345 474 356 508
rect 300 413 356 474
rect 300 379 311 413
rect 345 379 356 413
rect 300 367 356 379
rect 386 607 462 619
rect 386 573 408 607
rect 442 573 462 607
rect 386 525 462 573
rect 386 491 408 525
rect 442 491 462 525
rect 386 439 462 491
rect 386 405 408 439
rect 442 405 462 439
rect 386 367 462 405
rect 492 599 545 619
rect 492 565 503 599
rect 537 565 545 599
rect 492 508 545 565
rect 492 474 503 508
rect 537 474 545 508
rect 492 413 545 474
rect 492 379 503 413
rect 537 379 545 413
rect 492 367 545 379
<< ndiffc >>
rect 36 169 70 203
rect 36 67 70 101
rect 122 129 156 163
rect 194 129 228 163
rect 122 55 156 89
rect 194 55 228 89
rect 294 169 328 203
rect 294 67 328 101
rect 503 169 537 203
rect 503 59 537 93
<< pdiffc >>
rect 35 565 69 599
rect 35 470 69 504
rect 35 379 69 413
rect 121 573 155 607
rect 121 454 155 488
rect 225 565 259 599
rect 225 484 259 518
rect 225 400 259 434
rect 311 565 345 599
rect 311 474 345 508
rect 311 379 345 413
rect 408 573 442 607
rect 408 491 442 525
rect 408 405 442 439
rect 503 565 537 599
rect 503 474 537 508
rect 503 379 537 413
<< poly >>
rect 80 619 110 645
rect 270 619 300 645
rect 356 619 386 645
rect 462 619 492 645
rect 80 303 110 367
rect 270 335 300 367
rect 225 319 300 335
rect 80 287 177 303
rect 80 253 121 287
rect 155 253 177 287
rect 225 285 241 319
rect 275 285 300 319
rect 356 303 386 367
rect 462 303 492 367
rect 225 269 300 285
rect 348 287 414 303
rect 80 237 177 253
rect 81 215 111 237
rect 239 215 269 269
rect 348 253 364 287
rect 398 253 414 287
rect 348 237 414 253
rect 462 287 535 303
rect 462 253 485 287
rect 519 253 535 287
rect 462 237 535 253
rect 348 215 378 237
rect 462 215 492 237
rect 81 21 111 47
rect 239 21 269 47
rect 348 21 378 47
rect 462 21 492 47
<< polycont >>
rect 121 253 155 287
rect 241 285 275 319
rect 364 253 398 287
rect 485 253 519 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 19 599 71 615
rect 19 565 35 599
rect 69 565 71 599
rect 19 504 71 565
rect 19 470 35 504
rect 69 470 71 504
rect 19 413 71 470
rect 105 607 171 649
rect 105 573 121 607
rect 155 573 171 607
rect 105 488 171 573
rect 105 454 121 488
rect 155 454 171 488
rect 209 599 263 615
rect 209 565 225 599
rect 259 565 263 599
rect 209 518 263 565
rect 209 484 225 518
rect 259 484 263 518
rect 209 434 263 484
rect 209 420 225 434
rect 19 379 35 413
rect 69 379 71 413
rect 19 203 71 379
rect 143 400 225 420
rect 259 400 263 434
rect 143 384 263 400
rect 311 599 349 615
rect 345 565 349 599
rect 311 508 349 565
rect 345 474 349 508
rect 311 413 349 474
rect 143 303 177 384
rect 345 379 349 413
rect 392 607 458 649
rect 392 573 408 607
rect 442 573 458 607
rect 392 525 458 573
rect 392 491 408 525
rect 442 491 458 525
rect 392 439 458 491
rect 392 405 408 439
rect 442 405 458 439
rect 492 599 553 615
rect 492 565 503 599
rect 537 565 553 599
rect 492 508 553 565
rect 492 474 503 508
rect 537 474 553 508
rect 492 413 553 474
rect 311 371 349 379
rect 492 379 503 413
rect 537 379 553 413
rect 492 371 553 379
rect 105 287 177 303
rect 105 253 121 287
rect 155 253 177 287
rect 211 319 277 350
rect 311 337 553 371
rect 211 285 241 319
rect 275 285 277 319
rect 211 269 277 285
rect 348 287 451 303
rect 105 237 177 253
rect 348 253 364 287
rect 398 253 451 287
rect 348 237 451 253
rect 485 287 559 303
rect 519 253 559 287
rect 485 237 559 253
rect 19 169 36 203
rect 70 169 71 203
rect 143 231 177 237
rect 143 203 314 231
rect 143 197 294 203
rect 19 101 71 169
rect 278 169 294 197
rect 328 169 344 203
rect 19 67 36 101
rect 70 67 71 101
rect 19 51 71 67
rect 106 129 122 163
rect 156 129 194 163
rect 228 129 244 163
rect 106 89 244 129
rect 106 55 122 89
rect 156 55 194 89
rect 228 55 244 89
rect 106 17 244 55
rect 278 101 344 169
rect 278 67 294 101
rect 328 67 344 101
rect 388 68 451 237
rect 487 169 503 203
rect 537 169 553 203
rect 487 93 553 169
rect 278 51 344 67
rect 487 59 503 93
rect 537 59 553 93
rect 487 17 553 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a21o_1
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2568404
string GDS_START 2561472
<< end >>
