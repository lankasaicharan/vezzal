magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3506 1975
<< nwell >>
rect -38 331 2246 704
rect 1629 289 1837 331
<< pwell >>
rect 291 184 723 229
rect 3 157 723 184
rect 961 157 1609 201
rect 1927 157 2205 241
rect 3 49 1609 157
rect 1829 49 2205 157
rect 0 0 2208 49
<< scnmos >>
rect 86 74 116 158
rect 180 74 210 158
rect 370 119 400 203
rect 456 119 486 203
rect 542 119 572 203
rect 614 119 644 203
rect 827 47 857 131
rect 899 47 929 131
rect 1056 47 1086 175
rect 1128 47 1158 175
rect 1237 91 1267 175
rect 1309 91 1339 175
rect 1381 91 1411 175
rect 1496 91 1526 175
rect 1908 47 1938 131
rect 2010 47 2040 215
rect 2096 47 2126 215
<< scpmoshvt >>
rect 80 465 110 593
rect 166 465 196 593
rect 370 463 400 547
rect 456 463 486 547
rect 542 463 572 547
rect 614 463 644 547
rect 722 463 752 547
rect 808 463 838 547
rect 958 379 988 547
rect 1148 425 1178 509
rect 1257 425 1287 593
rect 1472 463 1502 547
rect 1558 463 1588 547
rect 1718 325 1748 409
rect 1908 397 1938 525
rect 2010 367 2040 619
rect 2096 367 2126 619
<< ndiff >>
rect 317 178 370 203
rect 29 132 86 158
rect 29 98 37 132
rect 71 98 86 132
rect 29 74 86 98
rect 116 126 180 158
rect 116 92 131 126
rect 165 92 180 126
rect 116 74 180 92
rect 210 133 263 158
rect 210 99 221 133
rect 255 99 263 133
rect 317 144 325 178
rect 359 144 370 178
rect 317 119 370 144
rect 400 178 456 203
rect 400 144 411 178
rect 445 144 456 178
rect 400 119 456 144
rect 486 164 542 203
rect 486 130 497 164
rect 531 130 542 164
rect 486 119 542 130
rect 572 119 614 203
rect 644 165 697 203
rect 644 131 655 165
rect 689 131 697 165
rect 987 163 1056 175
rect 987 131 995 163
rect 644 119 697 131
rect 210 74 263 99
rect 774 106 827 131
rect 774 72 782 106
rect 816 72 827 106
rect 774 47 827 72
rect 857 47 899 131
rect 929 129 995 131
rect 1029 129 1056 163
rect 929 93 1056 129
rect 929 59 995 93
rect 1029 59 1056 93
rect 929 47 1056 59
rect 1086 47 1128 175
rect 1158 163 1237 175
rect 1158 129 1173 163
rect 1207 129 1237 163
rect 1158 95 1237 129
rect 1158 61 1173 95
rect 1207 91 1237 95
rect 1267 91 1309 175
rect 1339 91 1381 175
rect 1411 133 1496 175
rect 1411 99 1422 133
rect 1456 99 1496 133
rect 1411 91 1496 99
rect 1526 137 1583 175
rect 1526 103 1541 137
rect 1575 103 1583 137
rect 1526 91 1583 103
rect 1207 61 1215 91
rect 1953 187 2010 215
rect 1953 153 1965 187
rect 1999 153 2010 187
rect 1953 131 2010 153
rect 1158 47 1215 61
rect 1855 101 1908 131
rect 1855 67 1863 101
rect 1897 67 1908 101
rect 1855 47 1908 67
rect 1938 93 2010 131
rect 1938 59 1953 93
rect 1987 59 2010 93
rect 1938 47 2010 59
rect 2040 203 2096 215
rect 2040 169 2051 203
rect 2085 169 2096 203
rect 2040 101 2096 169
rect 2040 67 2051 101
rect 2085 67 2096 101
rect 2040 47 2096 67
rect 2126 203 2179 215
rect 2126 169 2137 203
rect 2171 169 2179 203
rect 2126 93 2179 169
rect 2126 59 2137 93
rect 2171 59 2179 93
rect 2126 47 2179 59
<< pdiff >>
rect 27 579 80 593
rect 27 545 35 579
rect 69 545 80 579
rect 27 511 80 545
rect 27 477 35 511
rect 69 477 80 511
rect 27 465 80 477
rect 110 581 166 593
rect 110 547 121 581
rect 155 547 166 581
rect 110 513 166 547
rect 110 479 121 513
rect 155 479 166 513
rect 110 465 166 479
rect 196 581 251 593
rect 196 547 209 581
rect 243 547 251 581
rect 1309 607 1359 619
rect 1309 593 1317 607
rect 196 513 251 547
rect 196 479 209 513
rect 243 479 251 513
rect 196 465 251 479
rect 317 522 370 547
rect 317 488 325 522
rect 359 488 370 522
rect 317 463 370 488
rect 400 522 456 547
rect 400 488 411 522
rect 445 488 456 522
rect 400 463 456 488
rect 486 526 542 547
rect 486 492 497 526
rect 531 492 542 526
rect 486 463 542 492
rect 572 463 614 547
rect 644 522 722 547
rect 644 488 657 522
rect 691 488 722 522
rect 644 463 722 488
rect 752 522 808 547
rect 752 488 763 522
rect 797 488 808 522
rect 752 463 808 488
rect 838 525 958 547
rect 838 491 849 525
rect 883 491 958 525
rect 838 471 958 491
rect 838 463 913 471
rect 905 437 913 463
rect 947 437 958 471
rect 905 379 958 437
rect 988 535 1041 547
rect 988 501 999 535
rect 1033 501 1041 535
rect 1200 509 1257 593
rect 988 455 1041 501
rect 988 421 999 455
rect 1033 421 1041 455
rect 1095 484 1148 509
rect 1095 450 1103 484
rect 1137 450 1148 484
rect 1095 425 1148 450
rect 1178 467 1257 509
rect 1178 433 1201 467
rect 1235 433 1257 467
rect 1178 425 1257 433
rect 1287 573 1317 593
rect 1351 573 1359 607
rect 1287 476 1359 573
rect 1287 425 1337 476
rect 1419 525 1472 547
rect 1419 491 1427 525
rect 1461 491 1472 525
rect 1419 463 1472 491
rect 1502 537 1558 547
rect 1502 503 1513 537
rect 1547 503 1558 537
rect 1502 463 1558 503
rect 1588 522 1641 547
rect 1588 488 1599 522
rect 1633 488 1641 522
rect 1588 463 1641 488
rect 1960 525 2010 619
rect 1855 511 1908 525
rect 1855 477 1863 511
rect 1897 477 1908 511
rect 988 379 1041 421
rect 1855 443 1908 477
rect 1855 409 1863 443
rect 1897 409 1908 443
rect 1665 384 1718 409
rect 1665 350 1673 384
rect 1707 350 1718 384
rect 1665 325 1718 350
rect 1748 384 1801 409
rect 1855 397 1908 409
rect 1938 513 2010 525
rect 1938 479 1949 513
rect 1983 479 2010 513
rect 1938 445 2010 479
rect 1938 411 1949 445
rect 1983 411 2010 445
rect 1938 397 2010 411
rect 1748 350 1759 384
rect 1793 350 1801 384
rect 1748 325 1801 350
rect 1960 367 2010 397
rect 2040 599 2096 619
rect 2040 565 2051 599
rect 2085 565 2096 599
rect 2040 504 2096 565
rect 2040 470 2051 504
rect 2085 470 2096 504
rect 2040 420 2096 470
rect 2040 386 2051 420
rect 2085 386 2096 420
rect 2040 367 2096 386
rect 2126 607 2179 619
rect 2126 573 2137 607
rect 2171 573 2179 607
rect 2126 505 2179 573
rect 2126 471 2137 505
rect 2171 471 2179 505
rect 2126 413 2179 471
rect 2126 379 2137 413
rect 2171 379 2179 413
rect 2126 367 2179 379
<< ndiffc >>
rect 37 98 71 132
rect 131 92 165 126
rect 221 99 255 133
rect 325 144 359 178
rect 411 144 445 178
rect 497 130 531 164
rect 655 131 689 165
rect 782 72 816 106
rect 995 129 1029 163
rect 995 59 1029 93
rect 1173 129 1207 163
rect 1173 61 1207 95
rect 1422 99 1456 133
rect 1541 103 1575 137
rect 1965 153 1999 187
rect 1863 67 1897 101
rect 1953 59 1987 93
rect 2051 169 2085 203
rect 2051 67 2085 101
rect 2137 169 2171 203
rect 2137 59 2171 93
<< pdiffc >>
rect 35 545 69 579
rect 35 477 69 511
rect 121 547 155 581
rect 121 479 155 513
rect 209 547 243 581
rect 209 479 243 513
rect 325 488 359 522
rect 411 488 445 522
rect 497 492 531 526
rect 657 488 691 522
rect 763 488 797 522
rect 849 491 883 525
rect 913 437 947 471
rect 999 501 1033 535
rect 999 421 1033 455
rect 1103 450 1137 484
rect 1201 433 1235 467
rect 1317 573 1351 607
rect 1427 491 1461 525
rect 1513 503 1547 537
rect 1599 488 1633 522
rect 1863 477 1897 511
rect 1863 409 1897 443
rect 1673 350 1707 384
rect 1949 479 1983 513
rect 1949 411 1983 445
rect 1759 350 1793 384
rect 2051 565 2085 599
rect 2051 470 2085 504
rect 2051 386 2085 420
rect 2137 573 2171 607
rect 2137 471 2171 505
rect 2137 379 2171 413
<< poly >>
rect 80 593 110 619
rect 166 615 1287 645
rect 166 593 196 615
rect 370 547 400 573
rect 456 547 486 573
rect 542 547 572 615
rect 1257 593 1287 615
rect 614 547 644 573
rect 722 547 752 573
rect 808 547 838 573
rect 958 547 988 573
rect 80 443 110 465
rect 31 413 110 443
rect 31 251 61 413
rect 166 365 196 465
rect 370 441 400 463
rect 265 411 400 441
rect 265 377 281 411
rect 315 377 331 411
rect 103 349 210 365
rect 103 315 119 349
rect 153 315 210 349
rect 103 299 210 315
rect 31 235 138 251
rect 31 221 88 235
rect 72 201 88 221
rect 122 201 138 235
rect 72 185 138 201
rect 86 158 116 185
rect 180 158 210 299
rect 265 255 331 377
rect 456 369 486 463
rect 542 437 572 463
rect 373 353 486 369
rect 373 319 389 353
rect 423 333 486 353
rect 614 431 644 463
rect 614 415 680 431
rect 614 381 630 415
rect 664 381 680 415
rect 614 365 680 381
rect 423 319 564 333
rect 373 317 564 319
rect 373 303 572 317
rect 534 287 572 303
rect 265 225 400 255
rect 370 203 400 225
rect 456 203 486 229
rect 542 203 572 287
rect 614 291 644 365
rect 722 323 752 463
rect 808 431 838 463
rect 795 415 861 431
rect 795 381 811 415
rect 845 381 861 415
rect 795 365 861 381
rect 1148 509 1178 535
rect 1374 615 1813 645
rect 2010 619 2040 645
rect 2096 619 2126 645
rect 1374 461 1404 615
rect 1472 547 1502 615
rect 1747 605 1813 615
rect 1558 547 1588 573
rect 1747 571 1763 605
rect 1797 571 1813 605
rect 1747 537 1813 571
rect 1747 503 1763 537
rect 1797 503 1813 537
rect 1908 525 1938 551
rect 1747 487 1813 503
rect 1352 431 1404 461
rect 1472 437 1502 463
rect 958 323 988 379
rect 1148 335 1178 425
rect 1257 403 1287 425
rect 722 307 1037 323
rect 614 275 680 291
rect 614 241 630 275
rect 664 241 680 275
rect 722 273 739 307
rect 773 293 1037 307
rect 773 273 857 293
rect 722 257 857 273
rect 614 225 680 241
rect 614 203 644 225
rect 827 131 857 257
rect 899 231 965 247
rect 899 197 915 231
rect 949 197 965 231
rect 1007 227 1037 293
rect 1081 319 1178 335
rect 1081 285 1097 319
rect 1131 305 1178 319
rect 1237 373 1287 403
rect 1131 285 1158 305
rect 1081 269 1158 285
rect 1007 197 1086 227
rect 899 181 965 197
rect 899 131 929 181
rect 1056 175 1086 197
rect 1128 175 1158 269
rect 1237 175 1267 373
rect 1352 325 1382 431
rect 1558 383 1588 463
rect 1718 409 1748 435
rect 1309 295 1382 325
rect 1424 367 1588 383
rect 1424 333 1440 367
rect 1474 353 1588 367
rect 1474 333 1490 353
rect 1424 299 1490 333
rect 1908 375 1938 397
rect 1816 345 1938 375
rect 1309 175 1339 295
rect 1424 265 1440 299
rect 1474 265 1490 299
rect 1718 293 1748 325
rect 1816 293 1846 345
rect 2010 303 2040 367
rect 1424 249 1490 265
rect 1657 277 1846 293
rect 1424 227 1454 249
rect 1381 197 1454 227
rect 1657 243 1673 277
rect 1707 263 1846 277
rect 1707 243 1723 263
rect 1657 209 1723 243
rect 1381 175 1411 197
rect 1496 175 1526 201
rect 1657 175 1673 209
rect 1707 175 1723 209
rect 370 93 400 119
rect 86 48 116 74
rect 180 51 210 74
rect 456 51 486 119
rect 542 93 572 119
rect 614 93 644 119
rect 180 21 486 51
rect 1237 65 1267 91
rect 1309 65 1339 91
rect 1381 65 1411 91
rect 1496 69 1526 91
rect 1657 69 1723 175
rect 1816 189 1846 263
rect 1961 287 2040 303
rect 1961 253 1977 287
rect 2011 267 2040 287
rect 2096 267 2126 367
rect 2011 253 2126 267
rect 1961 237 2126 253
rect 2010 215 2040 237
rect 2096 215 2126 237
rect 1816 159 1938 189
rect 1908 131 1938 159
rect 827 21 857 47
rect 899 21 929 47
rect 1056 21 1086 47
rect 1128 21 1158 47
rect 1496 39 1723 69
rect 1908 21 1938 47
rect 2010 21 2040 47
rect 2096 21 2126 47
<< polycont >>
rect 281 377 315 411
rect 119 315 153 349
rect 88 201 122 235
rect 389 319 423 353
rect 630 381 664 415
rect 811 381 845 415
rect 1763 571 1797 605
rect 1763 503 1797 537
rect 630 241 664 275
rect 739 273 773 307
rect 915 197 949 231
rect 1097 285 1131 319
rect 1440 333 1474 367
rect 1440 265 1474 299
rect 1673 243 1707 277
rect 1673 175 1707 209
rect 1977 253 2011 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 18 579 73 595
rect 18 545 35 579
rect 69 545 73 579
rect 18 511 73 545
rect 18 477 35 511
rect 69 477 73 511
rect 18 365 73 477
rect 117 581 159 649
rect 117 547 121 581
rect 155 547 159 581
rect 117 513 159 547
rect 117 479 121 513
rect 155 479 159 513
rect 117 463 159 479
rect 205 581 247 597
rect 205 547 209 581
rect 243 547 247 581
rect 205 513 247 547
rect 205 479 209 513
rect 243 479 247 513
rect 205 463 247 479
rect 309 522 375 649
rect 309 488 325 522
rect 359 488 375 522
rect 309 472 375 488
rect 409 522 447 538
rect 409 488 411 522
rect 445 488 447 522
rect 18 349 169 365
rect 18 315 119 349
rect 153 315 169 349
rect 205 327 239 463
rect 409 453 447 488
rect 481 526 563 542
rect 481 492 497 526
rect 531 492 563 526
rect 481 487 563 492
rect 273 411 355 438
rect 409 419 493 453
rect 273 377 281 411
rect 315 377 355 411
rect 273 361 355 377
rect 389 353 425 369
rect 205 319 389 327
rect 423 319 425 353
rect 18 148 52 315
rect 205 291 425 319
rect 86 235 171 281
rect 86 201 88 235
rect 122 201 171 235
rect 86 185 171 201
rect 109 168 171 185
rect 205 276 271 291
rect 205 242 223 276
rect 257 242 271 276
rect 205 168 271 242
rect 459 235 493 419
rect 402 201 493 235
rect 529 345 563 487
rect 639 522 693 649
rect 639 488 657 522
rect 691 488 693 522
rect 639 472 693 488
rect 727 522 799 538
rect 727 488 763 522
rect 797 488 799 522
rect 727 472 799 488
rect 833 525 949 649
rect 833 491 849 525
rect 883 491 949 525
rect 833 472 949 491
rect 727 431 761 472
rect 897 471 949 472
rect 897 437 913 471
rect 947 437 949 471
rect 614 415 761 431
rect 614 381 630 415
rect 664 381 761 415
rect 614 379 761 381
rect 795 415 861 431
rect 897 421 949 437
rect 983 607 1367 611
rect 983 573 1317 607
rect 1351 573 1367 607
rect 983 571 1367 573
rect 983 535 1049 571
rect 1511 537 1557 649
rect 983 501 999 535
rect 1033 501 1049 535
rect 983 455 1049 501
rect 983 421 999 455
rect 1033 421 1049 455
rect 1087 525 1477 537
rect 1087 503 1427 525
rect 1087 484 1142 503
rect 1411 491 1427 503
rect 1461 491 1477 525
rect 1411 487 1477 491
rect 1511 503 1513 537
rect 1547 503 1557 537
rect 1511 487 1557 503
rect 1591 522 1639 538
rect 1591 488 1599 522
rect 1633 488 1639 522
rect 1087 450 1103 484
rect 1137 450 1142 484
rect 1087 434 1142 450
rect 1185 467 1270 469
rect 1185 433 1201 467
rect 1235 453 1270 467
rect 1591 453 1639 488
rect 1235 433 1639 453
rect 1185 421 1639 433
rect 1251 419 1639 421
rect 795 381 811 415
rect 845 387 861 415
rect 845 383 1217 387
rect 845 381 1527 383
rect 795 379 1527 381
rect 827 367 1527 379
rect 827 353 1440 367
rect 529 311 789 345
rect 18 132 81 148
rect 18 98 37 132
rect 71 98 81 132
rect 18 82 81 98
rect 115 126 181 134
rect 115 92 131 126
rect 165 92 181 126
rect 115 17 181 92
rect 215 133 271 168
rect 215 99 221 133
rect 255 99 271 133
rect 215 83 271 99
rect 309 178 368 194
rect 309 144 325 178
rect 359 144 368 178
rect 309 17 368 144
rect 402 178 447 201
rect 402 144 411 178
rect 445 144 447 178
rect 529 167 563 311
rect 723 307 789 311
rect 614 275 680 277
rect 614 241 630 275
rect 664 241 680 275
rect 723 273 739 307
rect 773 273 789 307
rect 723 271 789 273
rect 614 237 680 241
rect 827 247 861 353
rect 1181 333 1440 353
rect 1474 333 1527 367
rect 1081 285 1097 319
rect 1131 285 1147 319
rect 1081 276 1147 285
rect 614 203 791 237
rect 402 128 447 144
rect 481 164 563 167
rect 481 130 497 164
rect 531 130 563 164
rect 481 123 563 130
rect 639 165 705 169
rect 639 131 655 165
rect 689 131 705 165
rect 639 17 705 131
rect 757 122 791 203
rect 827 231 965 247
rect 1081 242 1087 276
rect 1121 242 1147 276
rect 1181 299 1527 333
rect 1181 265 1440 299
rect 1474 265 1527 299
rect 1181 249 1527 265
rect 1595 293 1639 419
rect 1673 384 1713 649
rect 1707 350 1713 384
rect 1673 334 1713 350
rect 1747 605 1813 615
rect 1747 571 1763 605
rect 1797 571 1813 605
rect 1747 537 1813 571
rect 1747 503 1763 537
rect 1797 503 1813 537
rect 1747 384 1813 503
rect 1747 350 1759 384
rect 1793 350 1813 384
rect 1595 277 1707 293
rect 1081 241 1147 242
rect 1595 243 1673 277
rect 827 197 915 231
rect 949 197 965 231
rect 1595 209 1707 243
rect 1595 207 1673 209
rect 1157 175 1673 207
rect 1157 173 1707 175
rect 1157 163 1223 173
rect 979 129 995 163
rect 1029 129 1045 163
rect 757 106 820 122
rect 757 72 782 106
rect 816 72 820 106
rect 757 56 820 72
rect 979 93 1045 129
rect 979 59 995 93
rect 1029 59 1045 93
rect 979 17 1045 59
rect 1157 129 1173 163
rect 1207 129 1223 163
rect 1657 159 1707 173
rect 1525 137 1591 139
rect 1157 95 1223 129
rect 1157 61 1173 95
rect 1207 61 1223 95
rect 1157 51 1223 61
rect 1406 99 1422 133
rect 1456 99 1472 133
rect 1406 17 1472 99
rect 1525 103 1541 137
rect 1575 123 1591 137
rect 1747 123 1813 350
rect 1575 103 1813 123
rect 1525 89 1813 103
rect 1847 511 1901 527
rect 1847 477 1863 511
rect 1897 477 1901 511
rect 1847 443 1901 477
rect 1847 409 1863 443
rect 1897 409 1901 443
rect 1847 303 1901 409
rect 1945 513 1987 649
rect 1945 479 1949 513
rect 1983 479 1987 513
rect 1945 445 1987 479
rect 1945 411 1949 445
rect 1983 411 1987 445
rect 1945 395 1987 411
rect 2045 599 2093 615
rect 2045 565 2051 599
rect 2085 565 2093 599
rect 2045 504 2093 565
rect 2045 470 2051 504
rect 2085 470 2093 504
rect 2045 420 2093 470
rect 2045 386 2051 420
rect 2085 386 2093 420
rect 1847 287 2011 303
rect 1847 253 1977 287
rect 1847 237 2011 253
rect 1847 101 1903 237
rect 2045 203 2093 386
rect 2127 607 2187 649
rect 2127 573 2137 607
rect 2171 573 2187 607
rect 2127 505 2187 573
rect 2127 471 2137 505
rect 2171 471 2187 505
rect 2127 413 2187 471
rect 2127 379 2137 413
rect 2171 379 2187 413
rect 2127 363 2187 379
rect 1949 187 2011 203
rect 1949 153 1965 187
rect 1999 153 2011 187
rect 1949 109 2011 153
rect 1847 67 1863 101
rect 1897 67 1903 101
rect 1847 51 1903 67
rect 1937 93 2011 109
rect 1937 59 1953 93
rect 1987 59 2011 93
rect 1937 17 2011 59
rect 2045 169 2051 203
rect 2085 169 2093 203
rect 2045 101 2093 169
rect 2045 67 2051 101
rect 2085 67 2093 101
rect 2045 51 2093 67
rect 2127 203 2187 219
rect 2127 169 2137 203
rect 2171 169 2187 203
rect 2127 93 2187 169
rect 2127 59 2137 93
rect 2171 59 2187 93
rect 2127 17 2187 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 223 242 257 276
rect 1087 242 1121 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 211 276 269 282
rect 211 242 223 276
rect 257 273 269 276
rect 1075 276 1133 282
rect 1075 273 1087 276
rect 257 245 1087 273
rect 257 242 269 245
rect 211 236 269 242
rect 1075 242 1087 245
rect 1121 242 1133 276
rect 1075 236 1133 242
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfstp_2
flabel comment s 624 332 624 332 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2047 94 2081 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 168 2081 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 464 2081 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2047 538 2081 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 344078
string GDS_START 327216
<< end >>
