magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 675 157 863 241
rect 12 49 863 157
rect 0 0 864 49
<< scnmos >>
rect 95 47 125 131
rect 181 47 211 131
rect 371 47 401 131
rect 457 47 487 131
rect 551 47 581 131
rect 637 47 667 131
rect 754 47 784 215
<< scpmoshvt >>
rect 80 535 110 619
rect 166 535 196 619
rect 385 391 415 475
rect 457 391 487 475
rect 565 391 595 475
rect 637 391 667 475
rect 742 367 772 619
<< ndiff >>
rect 701 189 754 215
rect 701 155 709 189
rect 743 155 754 189
rect 701 131 754 155
rect 38 106 95 131
rect 38 72 50 106
rect 84 72 95 106
rect 38 47 95 72
rect 125 103 181 131
rect 125 69 136 103
rect 170 69 181 103
rect 125 47 181 69
rect 211 106 264 131
rect 211 72 222 106
rect 256 72 264 106
rect 211 47 264 72
rect 318 105 371 131
rect 318 71 326 105
rect 360 71 371 105
rect 318 47 371 71
rect 401 106 457 131
rect 401 72 412 106
rect 446 72 457 106
rect 401 47 457 72
rect 487 106 551 131
rect 487 72 502 106
rect 536 72 551 106
rect 487 47 551 72
rect 581 106 637 131
rect 581 72 592 106
rect 626 72 637 106
rect 581 47 637 72
rect 667 93 754 131
rect 667 59 702 93
rect 736 59 754 93
rect 667 47 754 59
rect 784 203 837 215
rect 784 169 795 203
rect 829 169 837 203
rect 784 101 837 169
rect 784 67 795 101
rect 829 67 837 101
rect 784 47 837 67
<< pdiff >>
rect 27 594 80 619
rect 27 560 35 594
rect 69 560 80 594
rect 27 535 80 560
rect 110 594 166 619
rect 110 560 121 594
rect 155 560 166 594
rect 110 535 166 560
rect 196 594 249 619
rect 196 560 207 594
rect 241 560 249 594
rect 196 535 249 560
rect 689 607 742 619
rect 689 573 697 607
rect 731 573 742 607
rect 689 511 742 573
rect 689 477 697 511
rect 731 477 742 511
rect 689 475 742 477
rect 332 450 385 475
rect 332 416 340 450
rect 374 416 385 450
rect 332 391 385 416
rect 415 391 457 475
rect 487 391 565 475
rect 595 391 637 475
rect 667 413 742 475
rect 667 391 697 413
rect 689 379 697 391
rect 731 379 742 413
rect 689 367 742 379
rect 772 599 825 619
rect 772 565 783 599
rect 817 565 825 599
rect 772 511 825 565
rect 772 477 783 511
rect 817 477 825 511
rect 772 413 825 477
rect 772 379 783 413
rect 817 379 825 413
rect 772 367 825 379
<< ndiffc >>
rect 709 155 743 189
rect 50 72 84 106
rect 136 69 170 103
rect 222 72 256 106
rect 326 71 360 105
rect 412 72 446 106
rect 502 72 536 106
rect 592 72 626 106
rect 702 59 736 93
rect 795 169 829 203
rect 795 67 829 101
<< pdiffc >>
rect 35 560 69 594
rect 121 560 155 594
rect 207 560 241 594
rect 697 573 731 607
rect 697 477 731 511
rect 340 416 374 450
rect 697 379 731 413
rect 783 565 817 599
rect 783 477 817 511
rect 783 379 817 413
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 742 619 772 645
rect 268 601 357 617
rect 268 567 307 601
rect 341 567 357 601
rect 268 551 357 567
rect 575 599 667 615
rect 575 565 591 599
rect 625 565 667 599
rect 80 287 110 535
rect 166 477 196 535
rect 158 461 224 477
rect 158 427 174 461
rect 208 427 224 461
rect 158 411 224 427
rect 187 317 217 411
rect 181 287 217 317
rect 268 287 298 551
rect 575 549 667 565
rect 385 475 415 501
rect 457 475 487 501
rect 565 475 595 501
rect 637 475 667 549
rect 385 287 415 391
rect 73 271 139 287
rect 73 237 89 271
rect 123 237 139 271
rect 73 203 139 237
rect 73 169 89 203
rect 123 169 139 203
rect 73 153 139 169
rect 95 131 125 153
rect 181 131 211 287
rect 268 271 415 287
rect 268 257 322 271
rect 306 237 322 257
rect 356 257 415 271
rect 457 359 487 391
rect 457 343 523 359
rect 457 309 473 343
rect 507 309 523 343
rect 457 293 523 309
rect 356 237 401 257
rect 306 203 401 237
rect 306 169 322 203
rect 356 169 401 203
rect 457 183 487 293
rect 565 219 595 391
rect 306 153 401 169
rect 451 153 487 183
rect 529 203 595 219
rect 529 169 545 203
rect 579 169 595 203
rect 529 153 595 169
rect 371 131 401 153
rect 457 131 487 153
rect 551 131 581 153
rect 637 131 667 391
rect 742 305 772 367
rect 709 289 784 305
rect 709 255 725 289
rect 759 255 784 289
rect 709 239 784 255
rect 754 215 784 239
rect 95 21 125 47
rect 181 21 211 47
rect 371 21 401 47
rect 457 21 487 47
rect 551 21 581 47
rect 637 21 667 47
rect 754 21 784 47
<< polycont >>
rect 307 567 341 601
rect 591 565 625 599
rect 174 427 208 461
rect 89 237 123 271
rect 89 169 123 203
rect 322 237 356 271
rect 473 309 507 343
rect 322 169 356 203
rect 545 169 579 203
rect 725 255 759 289
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 17 594 78 610
rect 17 560 35 594
rect 69 560 78 594
rect 17 359 78 560
rect 112 594 164 649
rect 112 560 121 594
rect 155 560 164 594
rect 112 544 164 560
rect 198 601 357 610
rect 198 594 307 601
rect 198 560 207 594
rect 241 567 307 594
rect 341 567 357 601
rect 675 607 735 649
rect 241 560 357 567
rect 198 544 357 560
rect 412 565 591 599
rect 625 565 641 599
rect 112 461 267 510
rect 112 427 174 461
rect 208 427 267 461
rect 112 409 267 427
rect 324 450 378 466
rect 412 461 641 565
rect 675 573 697 607
rect 731 573 735 607
rect 675 511 735 573
rect 675 477 697 511
rect 731 477 735 511
rect 324 416 340 450
rect 374 427 378 450
rect 374 416 593 427
rect 324 393 593 416
rect 17 343 523 359
rect 17 323 473 343
rect 17 119 53 323
rect 457 309 473 323
rect 507 309 523 343
rect 457 307 523 309
rect 559 305 593 393
rect 675 413 735 477
rect 675 379 697 413
rect 731 379 735 413
rect 675 363 735 379
rect 779 599 847 615
rect 779 565 783 599
rect 817 565 847 599
rect 779 511 847 565
rect 779 477 783 511
rect 817 477 847 511
rect 779 413 847 477
rect 779 379 783 413
rect 817 379 847 413
rect 779 363 847 379
rect 559 289 759 305
rect 87 271 184 287
rect 87 237 89 271
rect 123 237 184 271
rect 87 203 184 237
rect 87 169 89 203
rect 123 169 184 203
rect 306 271 372 287
rect 559 273 725 289
rect 306 237 322 271
rect 356 237 372 271
rect 306 203 372 237
rect 306 189 322 203
rect 87 153 184 169
rect 218 169 322 189
rect 356 169 372 203
rect 218 155 372 169
rect 406 255 725 273
rect 406 239 759 255
rect 17 106 100 119
rect 17 72 50 106
rect 84 72 100 106
rect 17 56 100 72
rect 134 103 184 119
rect 134 69 136 103
rect 170 69 184 103
rect 134 17 184 69
rect 218 106 272 155
rect 218 72 222 106
rect 256 72 272 106
rect 218 56 272 72
rect 310 105 372 121
rect 310 71 326 105
rect 360 71 372 105
rect 310 17 372 71
rect 406 106 452 239
rect 495 203 595 205
rect 495 169 545 203
rect 579 169 595 203
rect 495 156 595 169
rect 631 122 665 239
rect 406 72 412 106
rect 446 72 452 106
rect 406 56 452 72
rect 486 106 552 122
rect 486 72 502 106
rect 536 72 552 106
rect 486 17 552 72
rect 588 106 665 122
rect 588 72 592 106
rect 626 72 665 106
rect 588 56 665 72
rect 699 189 759 205
rect 699 155 709 189
rect 743 155 759 189
rect 699 93 759 155
rect 699 59 702 93
rect 736 59 759 93
rect 699 17 759 59
rect 793 203 847 363
rect 793 169 795 203
rect 829 169 847 203
rect 793 101 847 169
rect 793 67 795 101
rect 829 67 847 101
rect 793 51 847 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or4bb_1
flabel comment s 279 413 279 413 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6650124
string GDS_START 6641052
<< end >>
