magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 58 49 554 157
rect 0 0 576 49
<< scnmos >>
rect 141 47 171 131
rect 219 47 249 131
rect 327 47 357 131
rect 441 47 471 131
<< scpmoshvt >>
rect 121 409 171 609
rect 227 409 277 609
rect 333 409 383 609
rect 441 409 491 609
<< ndiff >>
rect 84 93 141 131
rect 84 59 96 93
rect 130 59 141 93
rect 84 47 141 59
rect 171 47 219 131
rect 249 111 327 131
rect 249 77 260 111
rect 294 77 327 111
rect 249 47 327 77
rect 357 47 441 131
rect 471 106 528 131
rect 471 72 482 106
rect 516 72 528 106
rect 471 47 528 72
<< pdiff >>
rect 64 597 121 609
rect 64 563 76 597
rect 110 563 121 597
rect 64 505 121 563
rect 64 471 76 505
rect 110 471 121 505
rect 64 409 121 471
rect 171 527 227 609
rect 171 493 182 527
rect 216 493 227 527
rect 171 455 227 493
rect 171 421 182 455
rect 216 421 227 455
rect 171 409 227 421
rect 277 597 333 609
rect 277 563 288 597
rect 322 563 333 597
rect 277 526 333 563
rect 277 492 288 526
rect 322 492 333 526
rect 277 455 333 492
rect 277 421 288 455
rect 322 421 333 455
rect 277 409 333 421
rect 383 597 441 609
rect 383 563 394 597
rect 428 563 441 597
rect 383 505 441 563
rect 383 471 394 505
rect 428 471 441 505
rect 383 409 441 471
rect 491 597 548 609
rect 491 563 502 597
rect 536 563 548 597
rect 491 526 548 563
rect 491 492 502 526
rect 536 492 548 526
rect 491 455 548 492
rect 491 421 502 455
rect 536 421 548 455
rect 491 409 548 421
<< ndiffc >>
rect 96 59 130 93
rect 260 77 294 111
rect 482 72 516 106
<< pdiffc >>
rect 76 563 110 597
rect 76 471 110 505
rect 182 493 216 527
rect 182 421 216 455
rect 288 563 322 597
rect 288 492 322 526
rect 288 421 322 455
rect 394 563 428 597
rect 394 471 428 505
rect 502 563 536 597
rect 502 492 536 526
rect 502 421 536 455
<< poly >>
rect 121 609 171 635
rect 227 609 277 635
rect 333 609 383 635
rect 441 609 491 635
rect 121 349 171 409
rect 227 349 277 409
rect 333 349 383 409
rect 105 333 171 349
rect 105 299 121 333
rect 155 299 171 333
rect 105 265 171 299
rect 105 231 121 265
rect 155 231 171 265
rect 105 215 171 231
rect 213 333 279 349
rect 213 299 229 333
rect 263 299 279 333
rect 213 265 279 299
rect 213 231 229 265
rect 263 231 279 265
rect 213 215 279 231
rect 327 333 393 349
rect 327 299 343 333
rect 377 299 393 333
rect 327 265 393 299
rect 327 231 343 265
rect 377 231 393 265
rect 327 215 393 231
rect 441 305 491 409
rect 441 289 532 305
rect 441 255 482 289
rect 516 255 532 289
rect 441 221 532 255
rect 141 131 171 215
rect 219 131 249 215
rect 327 131 357 215
rect 441 187 482 221
rect 516 187 532 221
rect 441 171 532 187
rect 441 131 471 171
rect 141 21 171 47
rect 219 21 249 47
rect 327 21 357 47
rect 441 21 471 47
<< polycont >>
rect 121 299 155 333
rect 121 231 155 265
rect 229 299 263 333
rect 229 231 263 265
rect 343 299 377 333
rect 343 231 377 265
rect 482 255 516 289
rect 482 187 516 221
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 60 597 338 613
rect 60 563 76 597
rect 110 579 288 597
rect 110 563 126 579
rect 60 505 126 563
rect 272 563 288 579
rect 322 563 338 597
rect 60 471 76 505
rect 110 471 126 505
rect 60 455 126 471
rect 166 527 232 543
rect 166 493 182 527
rect 216 493 232 527
rect 166 455 232 493
rect 166 421 182 455
rect 216 421 232 455
rect 166 419 232 421
rect 25 385 232 419
rect 272 526 338 563
rect 272 492 288 526
rect 322 492 338 526
rect 272 455 338 492
rect 378 597 444 649
rect 378 563 394 597
rect 428 563 444 597
rect 378 505 444 563
rect 378 471 394 505
rect 428 471 444 505
rect 378 455 444 471
rect 486 597 552 613
rect 486 563 502 597
rect 536 563 552 597
rect 486 526 552 563
rect 486 492 502 526
rect 536 492 552 526
rect 486 455 552 492
rect 272 421 288 455
rect 322 421 338 455
rect 272 419 338 421
rect 486 421 502 455
rect 536 421 552 455
rect 486 419 552 421
rect 272 385 552 419
rect 25 179 69 385
rect 105 333 171 349
rect 105 299 121 333
rect 155 299 171 333
rect 105 265 171 299
rect 105 231 121 265
rect 155 231 171 265
rect 105 215 171 231
rect 213 333 279 349
rect 213 299 229 333
rect 263 299 279 333
rect 213 265 279 299
rect 213 231 229 265
rect 263 231 279 265
rect 213 215 279 231
rect 315 333 393 349
rect 315 299 343 333
rect 377 299 393 333
rect 315 265 393 299
rect 315 231 343 265
rect 377 231 393 265
rect 315 215 393 231
rect 466 289 551 305
rect 466 255 482 289
rect 516 255 551 289
rect 466 221 551 255
rect 466 187 482 221
rect 516 187 551 221
rect 25 145 310 179
rect 466 171 551 187
rect 244 111 310 145
rect 80 93 146 109
rect 80 59 96 93
rect 130 59 146 93
rect 80 17 146 59
rect 244 77 260 111
rect 294 77 310 111
rect 244 53 310 77
rect 466 106 532 135
rect 466 72 482 106
rect 516 72 532 106
rect 466 17 532 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a22oi_lp
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 368492
string GDS_START 362764
<< end >>
