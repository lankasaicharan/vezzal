magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1261 3122 1975
<< nwell >>
rect -38 331 1862 704
<< scpmoshvt >>
rect 211 536 1611 566
<< pdiff >>
rect 211 611 1611 619
rect 211 577 248 611
rect 282 577 316 611
rect 350 577 384 611
rect 418 577 452 611
rect 486 577 520 611
rect 554 577 588 611
rect 622 577 656 611
rect 690 577 724 611
rect 758 577 792 611
rect 826 577 860 611
rect 894 577 928 611
rect 962 577 996 611
rect 1030 577 1064 611
rect 1098 577 1132 611
rect 1166 577 1200 611
rect 1234 577 1268 611
rect 1302 577 1336 611
rect 1370 577 1404 611
rect 1438 577 1472 611
rect 1506 577 1540 611
rect 1574 577 1611 611
rect 211 566 1611 577
rect 211 525 1611 536
rect 211 491 248 525
rect 282 491 316 525
rect 350 491 384 525
rect 418 491 452 525
rect 486 491 520 525
rect 554 491 588 525
rect 622 491 656 525
rect 690 491 724 525
rect 758 491 792 525
rect 826 491 860 525
rect 894 491 928 525
rect 962 491 996 525
rect 1030 491 1064 525
rect 1098 491 1132 525
rect 1166 491 1200 525
rect 1234 491 1268 525
rect 1302 491 1336 525
rect 1370 491 1404 525
rect 1438 491 1472 525
rect 1506 491 1540 525
rect 1574 491 1611 525
rect 211 483 1611 491
<< pdiffc >>
rect 248 577 282 611
rect 316 577 350 611
rect 384 577 418 611
rect 452 577 486 611
rect 520 577 554 611
rect 588 577 622 611
rect 656 577 690 611
rect 724 577 758 611
rect 792 577 826 611
rect 860 577 894 611
rect 928 577 962 611
rect 996 577 1030 611
rect 1064 577 1098 611
rect 1132 577 1166 611
rect 1200 577 1234 611
rect 1268 577 1302 611
rect 1336 577 1370 611
rect 1404 577 1438 611
rect 1472 577 1506 611
rect 1540 577 1574 611
rect 248 491 282 525
rect 316 491 350 525
rect 384 491 418 525
rect 452 491 486 525
rect 520 491 554 525
rect 588 491 622 525
rect 656 491 690 525
rect 724 491 758 525
rect 792 491 826 525
rect 860 491 894 525
rect 928 491 962 525
rect 996 491 1030 525
rect 1064 491 1098 525
rect 1132 491 1166 525
rect 1200 491 1234 525
rect 1268 491 1302 525
rect 1336 491 1370 525
rect 1404 491 1438 525
rect 1472 491 1506 525
rect 1540 491 1574 525
<< poly >>
rect 185 536 211 566
rect 1611 550 1717 566
rect 1611 536 1667 550
rect 1634 516 1667 536
rect 1701 516 1717 550
rect 1634 482 1717 516
rect 1634 448 1667 482
rect 1701 448 1717 482
rect 1634 414 1717 448
rect 1634 380 1667 414
rect 1701 380 1717 414
rect 1634 364 1717 380
<< polycont >>
rect 1667 516 1701 550
rect 1667 448 1701 482
rect 1667 380 1701 414
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 211 611 1611 649
rect 211 577 248 611
rect 282 577 316 611
rect 350 577 379 611
rect 418 577 451 611
rect 486 577 520 611
rect 554 577 588 611
rect 622 577 656 611
rect 758 577 762 611
rect 826 577 860 611
rect 894 577 928 611
rect 962 577 996 611
rect 1035 577 1064 611
rect 1107 577 1132 611
rect 1166 577 1200 611
rect 1234 577 1268 611
rect 1302 577 1312 611
rect 1370 577 1384 611
rect 1438 577 1472 611
rect 1506 577 1540 611
rect 1574 577 1611 611
rect 211 568 1611 577
rect 1651 550 1757 566
rect 211 525 1590 534
rect 211 491 223 525
rect 282 491 295 525
rect 350 491 384 525
rect 418 491 452 525
rect 486 491 520 525
rect 568 491 588 525
rect 640 491 656 525
rect 690 491 724 525
rect 758 491 792 525
rect 826 491 845 525
rect 894 491 917 525
rect 962 491 996 525
rect 1030 491 1064 525
rect 1098 491 1132 525
rect 1190 491 1200 525
rect 1262 491 1268 525
rect 1302 491 1336 525
rect 1370 491 1404 525
rect 1438 491 1471 525
rect 1506 491 1540 525
rect 1577 491 1590 525
rect 211 482 1590 491
rect 1651 516 1667 550
rect 1701 516 1757 550
rect 1651 482 1757 516
rect 1651 448 1667 482
rect 1701 448 1757 482
rect 1651 414 1757 448
rect 1651 380 1667 414
rect 1701 380 1757 414
rect 1651 160 1757 380
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 379 577 384 611
rect 384 577 413 611
rect 451 577 452 611
rect 452 577 485 611
rect 690 577 724 611
rect 762 577 792 611
rect 792 577 796 611
rect 1001 577 1030 611
rect 1030 577 1035 611
rect 1073 577 1098 611
rect 1098 577 1107 611
rect 1312 577 1336 611
rect 1336 577 1346 611
rect 1384 577 1404 611
rect 1404 577 1418 611
rect 223 491 248 525
rect 248 491 257 525
rect 295 491 316 525
rect 316 491 329 525
rect 534 491 554 525
rect 554 491 568 525
rect 606 491 622 525
rect 622 491 640 525
rect 845 491 860 525
rect 860 491 879 525
rect 917 491 928 525
rect 928 491 951 525
rect 1156 491 1166 525
rect 1166 491 1190 525
rect 1228 491 1234 525
rect 1234 491 1262 525
rect 1471 491 1472 525
rect 1472 491 1505 525
rect 1543 491 1574 525
rect 1574 491 1577 525
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 369 611 494 617
rect 369 577 379 611
rect 413 577 451 611
rect 485 577 494 611
rect 369 565 494 577
rect 680 611 805 617
rect 680 577 690 611
rect 724 577 762 611
rect 796 577 805 611
rect 680 565 805 577
rect 991 611 1116 617
rect 991 577 1001 611
rect 1035 577 1073 611
rect 1107 577 1116 611
rect 991 565 1116 577
rect 1302 611 1431 617
rect 1302 577 1312 611
rect 1346 577 1384 611
rect 1418 577 1431 611
rect 1302 565 1431 577
rect 211 482 219 534
rect 271 482 283 534
rect 335 482 341 534
rect 522 482 528 534
rect 580 482 592 534
rect 644 482 652 534
rect 833 482 839 534
rect 891 482 903 534
rect 955 482 963 534
rect 1144 482 1150 534
rect 1202 482 1214 534
rect 1266 482 1274 534
rect 1459 482 1465 534
rect 1517 482 1529 534
rect 1581 482 1589 534
<< via1 >>
rect 219 525 271 534
rect 219 491 223 525
rect 223 491 257 525
rect 257 491 271 525
rect 219 482 271 491
rect 283 525 335 534
rect 283 491 295 525
rect 295 491 329 525
rect 329 491 335 525
rect 283 482 335 491
rect 528 525 580 534
rect 528 491 534 525
rect 534 491 568 525
rect 568 491 580 525
rect 528 482 580 491
rect 592 525 644 534
rect 592 491 606 525
rect 606 491 640 525
rect 640 491 644 525
rect 592 482 644 491
rect 839 525 891 534
rect 839 491 845 525
rect 845 491 879 525
rect 879 491 891 525
rect 839 482 891 491
rect 903 525 955 534
rect 903 491 917 525
rect 917 491 951 525
rect 951 491 955 525
rect 903 482 955 491
rect 1150 525 1202 534
rect 1150 491 1156 525
rect 1156 491 1190 525
rect 1190 491 1202 525
rect 1150 482 1202 491
rect 1214 525 1266 534
rect 1214 491 1228 525
rect 1228 491 1262 525
rect 1262 491 1266 525
rect 1214 482 1266 491
rect 1465 525 1517 534
rect 1465 491 1471 525
rect 1471 491 1505 525
rect 1505 491 1517 525
rect 1465 482 1517 491
rect 1529 525 1581 534
rect 1529 491 1543 525
rect 1543 491 1577 525
rect 1577 491 1581 525
rect 1529 482 1581 491
<< metal2 >>
rect 56 534 1768 666
rect 56 482 219 534
rect 271 482 283 534
rect 335 482 528 534
rect 580 482 592 534
rect 644 482 839 534
rect 891 482 903 534
rect 955 482 1150 534
rect 1202 482 1214 534
rect 1266 482 1465 534
rect 1517 482 1529 534
rect 1581 482 1768 534
rect 56 0 1768 482
<< labels >>
flabel metal1 s 0 617 1824 666 0 FreeSans 200 0 0 0 VIRTPWR
port 1 nsew
flabel metal2 s 56 0 1768 34 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power default
flabel locali s 1663 168 1697 202 0 FreeSans 200 0 0 0 SLEEP
port 3 nsew
flabel locali s 1663 242 1697 276 0 FreeSans 200 0 0 0 SLEEP
port 3 nsew
flabel locali s 1663 316 1697 350 0 FreeSans 200 0 0 0 SLEEP
port 3 nsew
flabel locali s 1663 390 1697 424 0 FreeSans 200 0 0 0 SLEEP
port 3 nsew
flabel locali s 1663 464 1697 498 0 FreeSans 200 0 0 0 SLEEP
port 3 nsew
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew
rlabel comment s 0 -1 0 -1 4 sleep_pargate_plv_7
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 1824 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string GDS_END 5008830
string GDS_START 4999318
<< end >>
