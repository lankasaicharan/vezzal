magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -300 17731 15300 35331
<< metal4 >>
tri 1934 33739 2266 34071 se
rect 2266 34047 12734 34071
tri 12734 34047 12758 34071 sw
rect 2266 33811 2269 34047
rect 2505 33811 2589 34047
rect 2825 33811 2909 34047
rect 3145 33811 3229 34047
rect 3465 33811 3549 34047
rect 3785 33811 3869 34047
rect 4105 33811 4189 34047
rect 4425 33811 4509 34047
rect 4745 33811 4829 34047
rect 5065 33811 5149 34047
rect 5385 33811 5469 34047
rect 5705 33811 5789 34047
rect 6025 33811 6109 34047
rect 6345 33811 6429 34047
rect 6665 33811 6749 34047
rect 6985 33811 7069 34047
rect 7305 33811 7389 34047
rect 7625 33811 7709 34047
rect 7945 33811 8029 34047
rect 8265 33811 8349 34047
rect 8585 33811 8669 34047
rect 8905 33811 8989 34047
rect 9225 33811 9309 34047
rect 9545 33811 9629 34047
rect 9865 33811 9949 34047
rect 10185 33811 10269 34047
rect 10505 33811 10589 34047
rect 10825 33811 10909 34047
rect 11145 33811 11229 34047
rect 11465 33811 11549 34047
rect 11785 33811 11869 34047
rect 12105 33811 12189 34047
rect 12425 33811 12509 34047
rect 12745 33811 12758 34047
rect 2266 33739 12758 33811
tri 1726 33531 1934 33739 se
rect 1934 33531 1947 33739
tri 1614 33419 1726 33531 se
rect 1726 33503 1947 33531
rect 2183 33685 12758 33739
tri 12758 33685 13120 34047 sw
rect 2183 33531 12871 33685
rect 2183 33503 2462 33531
tri 2462 33503 2490 33531 nw
rect 1726 33419 2378 33503
tri 2378 33419 2462 33503 nw
tri 1500 33305 1614 33419 se
rect 1614 33305 1627 33419
tri 1294 33099 1500 33305 se
rect 1500 33183 1627 33305
rect 1863 33183 2142 33419
tri 2142 33183 2378 33419 nw
tri 12510 33305 12736 33531 ne
rect 12736 33449 12871 33531
rect 13107 33531 13120 33685
tri 13120 33531 13274 33685 sw
rect 13107 33449 13274 33531
rect 12736 33365 13274 33449
tri 13274 33365 13440 33531 sw
rect 12736 33305 13191 33365
rect 1500 33099 1726 33183
tri 971 32776 1294 33099 se
rect 1294 32863 1307 33099
rect 1543 32863 1726 33099
rect 1294 32776 1726 32863
tri 962 32767 971 32776 se
rect 971 32767 984 32776
tri 960 32765 962 32767 se
rect 962 32765 984 32767
rect 960 32540 984 32765
rect 1220 32767 1726 32776
tri 1726 32767 2142 33183 nw
tri 12736 33129 12912 33305 ne
rect 12912 33129 13191 33305
rect 13427 33305 13440 33365
tri 13440 33305 13500 33365 sw
rect 13427 33129 13500 33305
tri 12912 32767 13274 33129 ne
rect 13274 33045 13500 33129
tri 13500 33045 13760 33305 sw
rect 13274 32809 13511 33045
rect 13747 32809 13760 33045
rect 13274 32767 13760 32809
rect 1220 32540 1500 32767
tri 1500 32541 1726 32767 nw
tri 13274 32541 13500 32767 ne
rect 13500 32765 13760 32767
tri 13760 32765 14040 33045 sw
rect 13500 32682 14040 32765
rect 960 32456 1500 32540
rect 960 32220 984 32456
rect 1220 32220 1500 32456
rect 960 32136 1500 32220
rect 960 31900 984 32136
rect 1220 31900 1500 32136
rect 960 31816 1500 31900
rect 960 31580 984 31816
rect 1220 31580 1500 31816
rect 960 31496 1500 31580
rect 960 31260 984 31496
rect 1220 31260 1500 31496
rect 960 31176 1500 31260
rect 960 30940 984 31176
rect 1220 30940 1500 31176
rect 960 30856 1500 30940
rect 960 30620 984 30856
rect 1220 30620 1500 30856
rect 960 30536 1500 30620
rect 960 30300 984 30536
rect 1220 30300 1500 30536
rect 960 30216 1500 30300
rect 960 29980 984 30216
rect 1220 29980 1500 30216
rect 960 29896 1500 29980
rect 960 29660 984 29896
rect 1220 29660 1500 29896
rect 960 29576 1500 29660
rect 960 29340 984 29576
rect 1220 29340 1500 29576
rect 960 29256 1500 29340
rect 960 29020 984 29256
rect 1220 29020 1500 29256
rect 960 28936 1500 29020
rect 960 28700 984 28936
rect 1220 28700 1500 28936
rect 960 28616 1500 28700
rect 960 28380 984 28616
rect 1220 28380 1500 28616
rect 960 28296 1500 28380
rect 960 28060 984 28296
rect 1220 28060 1500 28296
rect 960 27976 1500 28060
rect 960 27740 984 27976
rect 1220 27740 1500 27976
rect 960 27656 1500 27740
rect 960 27420 984 27656
rect 1220 27420 1500 27656
rect 960 27336 1500 27420
rect 960 27100 984 27336
rect 1220 27100 1500 27336
rect 960 27016 1500 27100
rect 960 26780 984 27016
rect 1220 26780 1500 27016
rect 960 26696 1500 26780
rect 960 26460 984 26696
rect 1220 26460 1500 26696
rect 960 26376 1500 26460
rect 960 26140 984 26376
rect 1220 26140 1500 26376
rect 960 26056 1500 26140
rect 960 25820 984 26056
rect 1220 25820 1500 26056
rect 960 25736 1500 25820
rect 960 25500 984 25736
rect 1220 25500 1500 25736
rect 960 25416 1500 25500
rect 960 25180 984 25416
rect 1220 25180 1500 25416
rect 960 25096 1500 25180
rect 960 24860 984 25096
rect 1220 24860 1500 25096
rect 960 24776 1500 24860
rect 960 24540 984 24776
rect 1220 24540 1500 24776
rect 960 24456 1500 24540
rect 960 24220 984 24456
rect 1220 24220 1500 24456
rect 960 24136 1500 24220
rect 960 23900 984 24136
rect 1220 23900 1500 24136
rect 960 23816 1500 23900
rect 960 23580 984 23816
rect 1220 23580 1500 23816
rect 960 23496 1500 23580
rect 960 23260 984 23496
rect 1220 23260 1500 23496
rect 960 23176 1500 23260
rect 960 22940 984 23176
rect 1220 22940 1500 23176
rect 960 22856 1500 22940
rect 960 22620 984 22856
rect 1220 22620 1500 22856
rect 960 22536 1500 22620
rect 960 22300 984 22536
rect 1220 22300 1500 22536
rect 960 22216 1500 22300
rect 960 21980 984 22216
rect 1220 21980 1500 22216
rect 960 21896 1500 21980
rect 960 21660 984 21896
rect 1220 21660 1500 21896
rect 960 21576 1500 21660
rect 960 21340 984 21576
rect 1220 21340 1500 21576
rect 960 21256 1500 21340
rect 960 21020 984 21256
rect 1220 21020 1500 21256
rect 960 20936 1500 21020
rect 960 20700 984 20936
rect 1220 20700 1500 20936
rect 960 20616 1500 20700
rect 960 20380 984 20616
rect 1220 20380 1500 20616
rect 13500 32446 13780 32682
rect 14016 32446 14040 32682
rect 13500 32362 14040 32446
rect 13500 32126 13780 32362
rect 14016 32126 14040 32362
rect 13500 32042 14040 32126
rect 13500 31806 13780 32042
rect 14016 31806 14040 32042
rect 13500 31722 14040 31806
rect 13500 31486 13780 31722
rect 14016 31486 14040 31722
rect 13500 31402 14040 31486
rect 13500 31166 13780 31402
rect 14016 31166 14040 31402
rect 13500 31082 14040 31166
rect 13500 30846 13780 31082
rect 14016 30846 14040 31082
rect 13500 30762 14040 30846
rect 13500 30526 13780 30762
rect 14016 30526 14040 30762
rect 13500 30442 14040 30526
rect 13500 30206 13780 30442
rect 14016 30206 14040 30442
rect 13500 30122 14040 30206
rect 13500 29886 13780 30122
rect 14016 29886 14040 30122
rect 13500 29802 14040 29886
rect 13500 29566 13780 29802
rect 14016 29566 14040 29802
rect 13500 29482 14040 29566
rect 13500 29246 13780 29482
rect 14016 29246 14040 29482
rect 13500 29162 14040 29246
rect 13500 28926 13780 29162
rect 14016 28926 14040 29162
rect 13500 28842 14040 28926
rect 13500 28606 13780 28842
rect 14016 28606 14040 28842
rect 13500 28522 14040 28606
rect 13500 28286 13780 28522
rect 14016 28286 14040 28522
rect 13500 28202 14040 28286
rect 13500 27966 13780 28202
rect 14016 27966 14040 28202
rect 13500 27882 14040 27966
rect 13500 27646 13780 27882
rect 14016 27646 14040 27882
rect 13500 27562 14040 27646
rect 13500 27326 13780 27562
rect 14016 27326 14040 27562
rect 13500 27242 14040 27326
rect 13500 27006 13780 27242
rect 14016 27006 14040 27242
rect 13500 26922 14040 27006
rect 13500 26686 13780 26922
rect 14016 26686 14040 26922
rect 13500 26602 14040 26686
rect 13500 26366 13780 26602
rect 14016 26366 14040 26602
rect 13500 26282 14040 26366
rect 13500 26046 13780 26282
rect 14016 26046 14040 26282
rect 13500 25962 14040 26046
rect 13500 25726 13780 25962
rect 14016 25726 14040 25962
rect 13500 25642 14040 25726
rect 13500 25406 13780 25642
rect 14016 25406 14040 25642
rect 13500 25322 14040 25406
rect 13500 25086 13780 25322
rect 14016 25086 14040 25322
rect 13500 25002 14040 25086
rect 13500 24766 13780 25002
rect 14016 24766 14040 25002
rect 13500 24682 14040 24766
rect 13500 24446 13780 24682
rect 14016 24446 14040 24682
rect 13500 24362 14040 24446
rect 13500 24126 13780 24362
rect 14016 24126 14040 24362
rect 13500 24042 14040 24126
rect 13500 23806 13780 24042
rect 14016 23806 14040 24042
rect 13500 23722 14040 23806
rect 13500 23486 13780 23722
rect 14016 23486 14040 23722
rect 13500 23402 14040 23486
rect 13500 23166 13780 23402
rect 14016 23166 14040 23402
rect 13500 23082 14040 23166
rect 13500 22846 13780 23082
rect 14016 22846 14040 23082
rect 13500 22762 14040 22846
rect 13500 22526 13780 22762
rect 14016 22526 14040 22762
rect 13500 22442 14040 22526
rect 13500 22206 13780 22442
rect 14016 22206 14040 22442
rect 13500 22122 14040 22206
rect 13500 21886 13780 22122
rect 14016 21886 14040 22122
rect 13500 21802 14040 21886
rect 13500 21566 13780 21802
rect 14016 21566 14040 21802
rect 13500 21482 14040 21566
rect 13500 21246 13780 21482
rect 14016 21246 14040 21482
rect 13500 21162 14040 21246
rect 13500 20926 13780 21162
rect 14016 20926 14040 21162
rect 13500 20842 14040 20926
rect 13500 20606 13780 20842
rect 14016 20606 14040 20842
rect 13500 20522 14040 20606
rect 960 20297 1500 20380
tri 1500 20297 1724 20521 sw
tri 13276 20297 13500 20521 se
rect 13500 20297 13780 20522
tri 960 20253 1004 20297 ne
rect 1004 20295 1724 20297
tri 1724 20295 1726 20297 sw
tri 13274 20295 13276 20297 se
rect 13276 20295 13780 20297
rect 1004 20253 1726 20295
tri 1004 20017 1240 20253 ne
rect 1240 20017 1253 20253
rect 1489 20017 1726 20253
tri 1240 19757 1500 20017 ne
rect 1500 19933 1726 20017
tri 1726 19933 2088 20295 sw
rect 1500 19757 1573 19933
tri 1500 19697 1560 19757 ne
rect 1560 19697 1573 19757
rect 1809 19757 2088 19933
tri 2088 19757 2264 19933 sw
tri 12858 19879 13274 20295 se
rect 13274 20286 13780 20295
rect 14016 20297 14040 20522
rect 14016 20295 14038 20297
tri 14038 20295 14040 20297 nw
rect 14016 20286 14029 20295
tri 14029 20286 14038 20295 nw
rect 13274 20199 13942 20286
tri 13942 20199 14029 20286 nw
rect 13274 19963 13457 20199
rect 13693 19963 13706 20199
tri 13706 19963 13942 20199 nw
rect 13274 19879 13500 19963
tri 12736 19757 12858 19879 se
rect 12858 19757 13137 19879
rect 1809 19697 2264 19757
tri 1560 19531 1726 19697 ne
rect 1726 19613 2264 19697
rect 1726 19531 1893 19613
tri 1726 19377 1880 19531 ne
rect 1880 19377 1893 19531
rect 2129 19531 2264 19613
tri 2264 19531 2490 19757 sw
tri 12510 19531 12736 19757 se
rect 12736 19643 13137 19757
rect 13373 19757 13500 19879
tri 13500 19757 13706 19963 nw
rect 13373 19643 13386 19757
tri 13386 19643 13500 19757 nw
rect 12736 19559 13274 19643
rect 12736 19531 12817 19559
rect 2129 19377 12817 19531
tri 1880 19251 2006 19377 ne
rect 2006 19323 12817 19377
rect 13053 19531 13274 19559
tri 13274 19531 13386 19643 nw
rect 13053 19323 13066 19531
tri 13066 19323 13274 19531 nw
rect 2006 19251 12734 19323
tri 2006 19015 2242 19251 ne
rect 2242 19015 2255 19251
rect 2491 19015 2575 19251
rect 2811 19015 2895 19251
rect 3131 19015 3215 19251
rect 3451 19015 3535 19251
rect 3771 19015 3855 19251
rect 4091 19015 4175 19251
rect 4411 19015 4495 19251
rect 4731 19015 4815 19251
rect 5051 19015 5135 19251
rect 5371 19015 5455 19251
rect 5691 19015 5775 19251
rect 6011 19015 6095 19251
rect 6331 19015 6415 19251
rect 6651 19015 6735 19251
rect 6971 19015 7055 19251
rect 7291 19015 7375 19251
rect 7611 19015 7695 19251
rect 7931 19015 8015 19251
rect 8251 19015 8335 19251
rect 8571 19015 8655 19251
rect 8891 19015 8975 19251
rect 9211 19015 9295 19251
rect 9531 19015 9615 19251
rect 9851 19015 9935 19251
rect 10171 19015 10255 19251
rect 10491 19015 10575 19251
rect 10811 19015 10895 19251
rect 11131 19015 11215 19251
rect 11451 19015 11535 19251
rect 11771 19015 11855 19251
rect 12091 19015 12175 19251
rect 12411 19015 12495 19251
rect 12731 19015 12734 19251
tri 2242 18991 2266 19015 ne
rect 2266 18991 12734 19015
tri 12734 18991 13066 19323 nw
<< via4 >>
rect 2269 33811 2505 34047
rect 2589 33811 2825 34047
rect 2909 33811 3145 34047
rect 3229 33811 3465 34047
rect 3549 33811 3785 34047
rect 3869 33811 4105 34047
rect 4189 33811 4425 34047
rect 4509 33811 4745 34047
rect 4829 33811 5065 34047
rect 5149 33811 5385 34047
rect 5469 33811 5705 34047
rect 5789 33811 6025 34047
rect 6109 33811 6345 34047
rect 6429 33811 6665 34047
rect 6749 33811 6985 34047
rect 7069 33811 7305 34047
rect 7389 33811 7625 34047
rect 7709 33811 7945 34047
rect 8029 33811 8265 34047
rect 8349 33811 8585 34047
rect 8669 33811 8905 34047
rect 8989 33811 9225 34047
rect 9309 33811 9545 34047
rect 9629 33811 9865 34047
rect 9949 33811 10185 34047
rect 10269 33811 10505 34047
rect 10589 33811 10825 34047
rect 10909 33811 11145 34047
rect 11229 33811 11465 34047
rect 11549 33811 11785 34047
rect 11869 33811 12105 34047
rect 12189 33811 12425 34047
rect 12509 33811 12745 34047
rect 1947 33503 2183 33739
rect 1627 33183 1863 33419
rect 12871 33449 13107 33685
rect 1307 32863 1543 33099
rect 984 32540 1220 32776
rect 13191 33129 13427 33365
rect 13511 32809 13747 33045
rect 984 32220 1220 32456
rect 984 31900 1220 32136
rect 984 31580 1220 31816
rect 984 31260 1220 31496
rect 984 30940 1220 31176
rect 984 30620 1220 30856
rect 984 30300 1220 30536
rect 984 29980 1220 30216
rect 984 29660 1220 29896
rect 984 29340 1220 29576
rect 984 29020 1220 29256
rect 984 28700 1220 28936
rect 984 28380 1220 28616
rect 984 28060 1220 28296
rect 984 27740 1220 27976
rect 984 27420 1220 27656
rect 984 27100 1220 27336
rect 984 26780 1220 27016
rect 984 26460 1220 26696
rect 984 26140 1220 26376
rect 984 25820 1220 26056
rect 984 25500 1220 25736
rect 984 25180 1220 25416
rect 984 24860 1220 25096
rect 984 24540 1220 24776
rect 984 24220 1220 24456
rect 984 23900 1220 24136
rect 984 23580 1220 23816
rect 984 23260 1220 23496
rect 984 22940 1220 23176
rect 984 22620 1220 22856
rect 984 22300 1220 22536
rect 984 21980 1220 22216
rect 984 21660 1220 21896
rect 984 21340 1220 21576
rect 984 21020 1220 21256
rect 984 20700 1220 20936
rect 984 20380 1220 20616
rect 13780 32446 14016 32682
rect 13780 32126 14016 32362
rect 13780 31806 14016 32042
rect 13780 31486 14016 31722
rect 13780 31166 14016 31402
rect 13780 30846 14016 31082
rect 13780 30526 14016 30762
rect 13780 30206 14016 30442
rect 13780 29886 14016 30122
rect 13780 29566 14016 29802
rect 13780 29246 14016 29482
rect 13780 28926 14016 29162
rect 13780 28606 14016 28842
rect 13780 28286 14016 28522
rect 13780 27966 14016 28202
rect 13780 27646 14016 27882
rect 13780 27326 14016 27562
rect 13780 27006 14016 27242
rect 13780 26686 14016 26922
rect 13780 26366 14016 26602
rect 13780 26046 14016 26282
rect 13780 25726 14016 25962
rect 13780 25406 14016 25642
rect 13780 25086 14016 25322
rect 13780 24766 14016 25002
rect 13780 24446 14016 24682
rect 13780 24126 14016 24362
rect 13780 23806 14016 24042
rect 13780 23486 14016 23722
rect 13780 23166 14016 23402
rect 13780 22846 14016 23082
rect 13780 22526 14016 22762
rect 13780 22206 14016 22442
rect 13780 21886 14016 22122
rect 13780 21566 14016 21802
rect 13780 21246 14016 21482
rect 13780 20926 14016 21162
rect 13780 20606 14016 20842
rect 1253 20017 1489 20253
rect 1573 19697 1809 19933
rect 13780 20286 14016 20522
rect 13457 19963 13693 20199
rect 1893 19377 2129 19613
rect 13137 19643 13373 19879
rect 12817 19323 13053 19559
rect 2255 19015 2491 19251
rect 2575 19015 2811 19251
rect 2895 19015 3131 19251
rect 3215 19015 3451 19251
rect 3535 19015 3771 19251
rect 3855 19015 4091 19251
rect 4175 19015 4411 19251
rect 4495 19015 4731 19251
rect 4815 19015 5051 19251
rect 5135 19015 5371 19251
rect 5455 19015 5691 19251
rect 5775 19015 6011 19251
rect 6095 19015 6331 19251
rect 6415 19015 6651 19251
rect 6735 19015 6971 19251
rect 7055 19015 7291 19251
rect 7375 19015 7611 19251
rect 7695 19015 7931 19251
rect 8015 19015 8251 19251
rect 8335 19015 8571 19251
rect 8655 19015 8891 19251
rect 8975 19015 9211 19251
rect 9295 19015 9531 19251
rect 9615 19015 9851 19251
rect 9935 19015 10171 19251
rect 10255 19015 10491 19251
rect 10575 19015 10811 19251
rect 10895 19015 11131 19251
rect 11215 19015 11451 19251
rect 11535 19015 11771 19251
rect 11855 19015 12091 19251
rect 12175 19015 12411 19251
rect 12495 19015 12731 19251
<< metal5 >>
tri 1934 33739 2266 34071 se
rect 2266 34047 12734 34071
tri 12734 34047 12758 34071 sw
rect 2266 33811 2269 34047
rect 2505 33811 2589 34047
rect 2825 33811 2909 34047
rect 3145 33811 3229 34047
rect 3465 33811 3549 34047
rect 3785 33811 3869 34047
rect 4105 33811 4189 34047
rect 4425 33811 4509 34047
rect 4745 33811 4829 34047
rect 5065 33811 5149 34047
rect 5385 33811 5469 34047
rect 5705 33811 5789 34047
rect 6025 33811 6109 34047
rect 6345 33811 6429 34047
rect 6665 33811 6749 34047
rect 6985 33811 7069 34047
rect 7305 33811 7389 34047
rect 7625 33811 7709 34047
rect 7945 33811 8029 34047
rect 8265 33811 8349 34047
rect 8585 33811 8669 34047
rect 8905 33811 8989 34047
rect 9225 33811 9309 34047
rect 9545 33811 9629 34047
rect 9865 33811 9949 34047
rect 10185 33811 10269 34047
rect 10505 33811 10589 34047
rect 10825 33811 10909 34047
rect 11145 33811 11229 34047
rect 11465 33811 11549 34047
rect 11785 33811 11869 34047
rect 12105 33811 12189 34047
rect 12425 33811 12509 34047
rect 12745 33811 12758 34047
rect 2266 33739 12758 33811
tri 1614 33419 1934 33739 se
rect 1934 33503 1947 33739
rect 2183 33685 12758 33739
tri 12758 33685 13120 34047 sw
rect 2183 33503 12871 33685
rect 1934 33449 12871 33503
rect 13107 33449 13120 33685
rect 1934 33419 13120 33449
tri 1294 33099 1614 33419 se
rect 1614 33183 1627 33419
rect 1863 33365 13120 33419
tri 13120 33365 13440 33685 sw
rect 1863 33183 13191 33365
rect 1614 33129 13191 33183
rect 13427 33129 13440 33365
rect 1614 33099 13440 33129
tri 971 32776 1294 33099 se
rect 1294 32863 1307 33099
rect 1543 33045 13440 33099
tri 13440 33045 13760 33365 sw
rect 1543 32863 13511 33045
rect 1294 32809 13511 32863
rect 13747 32809 13760 33045
rect 1294 32776 13760 32809
tri 960 32765 971 32776 se
rect 971 32765 984 32776
rect 960 32540 984 32765
rect 1220 32765 13760 32776
tri 13760 32765 14040 33045 sw
rect 1220 32682 14040 32765
rect 1220 32540 13780 32682
rect 960 32456 13780 32540
rect 960 32220 984 32456
rect 1220 32446 13780 32456
rect 14016 32446 14040 32682
rect 1220 32362 14040 32446
rect 1220 32220 13780 32362
rect 960 32136 13780 32220
rect 960 31900 984 32136
rect 1220 32126 13780 32136
rect 14016 32126 14040 32362
rect 1220 32042 14040 32126
rect 1220 31900 13780 32042
rect 960 31816 13780 31900
rect 960 31580 984 31816
rect 1220 31806 13780 31816
rect 14016 31806 14040 32042
rect 1220 31722 14040 31806
rect 1220 31580 13780 31722
rect 960 31496 13780 31580
rect 960 31260 984 31496
rect 1220 31486 13780 31496
rect 14016 31486 14040 31722
rect 1220 31402 14040 31486
rect 1220 31260 13780 31402
rect 960 31176 13780 31260
rect 960 30940 984 31176
rect 1220 31166 13780 31176
rect 14016 31166 14040 31402
rect 1220 31082 14040 31166
rect 1220 30940 13780 31082
rect 960 30856 13780 30940
rect 960 30620 984 30856
rect 1220 30846 13780 30856
rect 14016 30846 14040 31082
rect 1220 30762 14040 30846
rect 1220 30620 13780 30762
rect 960 30536 13780 30620
rect 960 30300 984 30536
rect 1220 30526 13780 30536
rect 14016 30526 14040 30762
rect 1220 30442 14040 30526
rect 1220 30300 13780 30442
rect 960 30216 13780 30300
rect 960 29980 984 30216
rect 1220 30206 13780 30216
rect 14016 30206 14040 30442
rect 1220 30122 14040 30206
rect 1220 29980 13780 30122
rect 960 29896 13780 29980
rect 960 29660 984 29896
rect 1220 29886 13780 29896
rect 14016 29886 14040 30122
rect 1220 29802 14040 29886
rect 1220 29660 13780 29802
rect 960 29576 13780 29660
rect 960 29340 984 29576
rect 1220 29566 13780 29576
rect 14016 29566 14040 29802
rect 1220 29482 14040 29566
rect 1220 29340 13780 29482
rect 960 29256 13780 29340
rect 960 29020 984 29256
rect 1220 29246 13780 29256
rect 14016 29246 14040 29482
rect 1220 29162 14040 29246
rect 1220 29020 13780 29162
rect 960 28936 13780 29020
rect 960 28700 984 28936
rect 1220 28926 13780 28936
rect 14016 28926 14040 29162
rect 1220 28842 14040 28926
rect 1220 28700 13780 28842
rect 960 28616 13780 28700
rect 960 28380 984 28616
rect 1220 28606 13780 28616
rect 14016 28606 14040 28842
rect 1220 28522 14040 28606
rect 1220 28380 13780 28522
rect 960 28296 13780 28380
rect 960 28060 984 28296
rect 1220 28286 13780 28296
rect 14016 28286 14040 28522
rect 1220 28202 14040 28286
rect 1220 28060 13780 28202
rect 960 27976 13780 28060
rect 960 27740 984 27976
rect 1220 27966 13780 27976
rect 14016 27966 14040 28202
rect 1220 27882 14040 27966
rect 1220 27740 13780 27882
rect 960 27656 13780 27740
rect 960 27420 984 27656
rect 1220 27646 13780 27656
rect 14016 27646 14040 27882
rect 1220 27562 14040 27646
rect 1220 27420 13780 27562
rect 960 27336 13780 27420
rect 960 27100 984 27336
rect 1220 27326 13780 27336
rect 14016 27326 14040 27562
rect 1220 27242 14040 27326
rect 1220 27100 13780 27242
rect 960 27016 13780 27100
rect 960 26780 984 27016
rect 1220 27006 13780 27016
rect 14016 27006 14040 27242
rect 1220 26922 14040 27006
rect 1220 26780 13780 26922
rect 960 26696 13780 26780
rect 960 26460 984 26696
rect 1220 26686 13780 26696
rect 14016 26686 14040 26922
rect 1220 26602 14040 26686
rect 1220 26460 13780 26602
rect 960 26376 13780 26460
rect 960 26140 984 26376
rect 1220 26366 13780 26376
rect 14016 26366 14040 26602
rect 1220 26282 14040 26366
rect 1220 26140 13780 26282
rect 960 26056 13780 26140
rect 960 25820 984 26056
rect 1220 26046 13780 26056
rect 14016 26046 14040 26282
rect 1220 25962 14040 26046
rect 1220 25820 13780 25962
rect 960 25736 13780 25820
rect 960 25500 984 25736
rect 1220 25726 13780 25736
rect 14016 25726 14040 25962
rect 1220 25642 14040 25726
rect 1220 25500 13780 25642
rect 960 25416 13780 25500
rect 960 25180 984 25416
rect 1220 25406 13780 25416
rect 14016 25406 14040 25642
rect 1220 25322 14040 25406
rect 1220 25180 13780 25322
rect 960 25096 13780 25180
rect 960 24860 984 25096
rect 1220 25086 13780 25096
rect 14016 25086 14040 25322
rect 1220 25002 14040 25086
rect 1220 24860 13780 25002
rect 960 24776 13780 24860
rect 960 24540 984 24776
rect 1220 24766 13780 24776
rect 14016 24766 14040 25002
rect 1220 24682 14040 24766
rect 1220 24540 13780 24682
rect 960 24456 13780 24540
rect 960 24220 984 24456
rect 1220 24446 13780 24456
rect 14016 24446 14040 24682
rect 1220 24362 14040 24446
rect 1220 24220 13780 24362
rect 960 24136 13780 24220
rect 960 23900 984 24136
rect 1220 24126 13780 24136
rect 14016 24126 14040 24362
rect 1220 24042 14040 24126
rect 1220 23900 13780 24042
rect 960 23816 13780 23900
rect 960 23580 984 23816
rect 1220 23806 13780 23816
rect 14016 23806 14040 24042
rect 1220 23722 14040 23806
rect 1220 23580 13780 23722
rect 960 23496 13780 23580
rect 960 23260 984 23496
rect 1220 23486 13780 23496
rect 14016 23486 14040 23722
rect 1220 23402 14040 23486
rect 1220 23260 13780 23402
rect 960 23176 13780 23260
rect 960 22940 984 23176
rect 1220 23166 13780 23176
rect 14016 23166 14040 23402
rect 1220 23082 14040 23166
rect 1220 22940 13780 23082
rect 960 22856 13780 22940
rect 960 22620 984 22856
rect 1220 22846 13780 22856
rect 14016 22846 14040 23082
rect 1220 22762 14040 22846
rect 1220 22620 13780 22762
rect 960 22536 13780 22620
rect 960 22300 984 22536
rect 1220 22526 13780 22536
rect 14016 22526 14040 22762
rect 1220 22442 14040 22526
rect 1220 22300 13780 22442
rect 960 22216 13780 22300
rect 960 21980 984 22216
rect 1220 22206 13780 22216
rect 14016 22206 14040 22442
rect 1220 22122 14040 22206
rect 1220 21980 13780 22122
rect 960 21896 13780 21980
rect 960 21660 984 21896
rect 1220 21886 13780 21896
rect 14016 21886 14040 22122
rect 1220 21802 14040 21886
rect 1220 21660 13780 21802
rect 960 21576 13780 21660
rect 960 21340 984 21576
rect 1220 21566 13780 21576
rect 14016 21566 14040 21802
rect 1220 21482 14040 21566
rect 1220 21340 13780 21482
rect 960 21256 13780 21340
rect 960 21020 984 21256
rect 1220 21246 13780 21256
rect 14016 21246 14040 21482
rect 1220 21162 14040 21246
rect 1220 21020 13780 21162
rect 960 20936 13780 21020
rect 960 20700 984 20936
rect 1220 20926 13780 20936
rect 14016 20926 14040 21162
rect 1220 20842 14040 20926
rect 1220 20700 13780 20842
rect 960 20616 13780 20700
rect 960 20380 984 20616
rect 1220 20606 13780 20616
rect 14016 20606 14040 20842
rect 1220 20522 14040 20606
rect 1220 20380 13780 20522
rect 960 20297 13780 20380
tri 960 20253 1004 20297 ne
rect 1004 20286 13780 20297
rect 14016 20297 14040 20522
rect 14016 20286 14029 20297
tri 14029 20286 14040 20297 nw
rect 1004 20253 13942 20286
tri 1004 20017 1240 20253 ne
rect 1240 20017 1253 20253
rect 1489 20199 13942 20253
tri 13942 20199 14029 20286 nw
rect 1489 20017 13457 20199
tri 1240 19933 1324 20017 ne
rect 1324 19963 13457 20017
rect 13693 19963 13706 20199
tri 13706 19963 13942 20199 nw
rect 1324 19933 13622 19963
tri 1324 19697 1560 19933 ne
rect 1560 19697 1573 19933
rect 1809 19879 13622 19933
tri 13622 19879 13706 19963 nw
rect 1809 19697 13137 19879
tri 1560 19613 1644 19697 ne
rect 1644 19643 13137 19697
rect 13373 19643 13386 19879
tri 13386 19643 13622 19879 nw
rect 1644 19613 13302 19643
tri 1644 19377 1880 19613 ne
rect 1880 19377 1893 19613
rect 2129 19559 13302 19613
tri 13302 19559 13386 19643 nw
rect 2129 19377 12817 19559
tri 1880 19251 2006 19377 ne
rect 2006 19323 12817 19377
rect 13053 19323 13066 19559
tri 13066 19323 13302 19559 nw
rect 2006 19251 12734 19323
tri 2006 19015 2242 19251 ne
rect 2242 19015 2255 19251
rect 2491 19015 2575 19251
rect 2811 19015 2895 19251
rect 3131 19015 3215 19251
rect 3451 19015 3535 19251
rect 3771 19015 3855 19251
rect 4091 19015 4175 19251
rect 4411 19015 4495 19251
rect 4731 19015 4815 19251
rect 5051 19015 5135 19251
rect 5371 19015 5455 19251
rect 5691 19015 5775 19251
rect 6011 19015 6095 19251
rect 6331 19015 6415 19251
rect 6651 19015 6735 19251
rect 6971 19015 7055 19251
rect 7291 19015 7375 19251
rect 7611 19015 7695 19251
rect 7931 19015 8015 19251
rect 8251 19015 8335 19251
rect 8571 19015 8655 19251
rect 8891 19015 8975 19251
rect 9211 19015 9295 19251
rect 9531 19015 9615 19251
rect 9851 19015 9935 19251
rect 10171 19015 10255 19251
rect 10491 19015 10575 19251
rect 10811 19015 10895 19251
rect 11131 19015 11215 19251
rect 11451 19015 11535 19251
rect 11771 19015 11855 19251
rect 12091 19015 12175 19251
rect 12411 19015 12495 19251
rect 12731 19015 12734 19251
tri 2242 18991 2266 19015 ne
rect 2266 18991 12734 19015
tri 12734 18991 13066 19323 nw
<< glass >>
tri 1500 32541 2490 33531 se
rect 2490 32541 12510 33531
tri 12510 32541 13500 33531 sw
rect 1500 20521 13500 32541
tri 1500 19531 2490 20521 ne
rect 2490 19531 12510 20521
tri 12510 19531 13500 20521 nw
use sky130_fd_pr__padplhp__example_559591418080  sky130_fd_pr__padplhp__example_559591418080_0
timestamp 1627201311
transform 1 0 1500 0 1 19531
box -478 -478 6000 7000
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 12450
string GDS_START 12378
<< end >>
