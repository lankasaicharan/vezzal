magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 240 241 732 243
rect 13 49 732 241
rect 0 0 768 49
<< scnmos >>
rect 92 47 122 215
rect 319 49 349 217
rect 443 49 473 217
rect 551 49 581 217
rect 623 49 653 217
<< scpmoshvt >>
rect 181 367 211 619
rect 335 367 365 619
rect 407 367 437 619
rect 515 367 545 619
rect 623 367 653 619
<< ndiff >>
rect 39 184 92 215
rect 39 150 47 184
rect 81 150 92 184
rect 39 101 92 150
rect 39 67 47 101
rect 81 67 92 101
rect 39 47 92 67
rect 122 203 175 215
rect 122 169 133 203
rect 167 169 175 203
rect 122 93 175 169
rect 122 59 133 93
rect 167 59 175 93
rect 122 47 175 59
rect 266 171 319 217
rect 266 137 274 171
rect 308 137 319 171
rect 266 97 319 137
rect 266 63 274 97
rect 308 63 319 97
rect 266 49 319 63
rect 349 99 443 217
rect 349 65 379 99
rect 413 65 443 99
rect 349 49 443 65
rect 473 171 551 217
rect 473 137 495 171
rect 529 137 551 171
rect 473 97 551 137
rect 473 63 495 97
rect 529 63 551 97
rect 473 49 551 63
rect 581 49 623 217
rect 653 205 706 217
rect 653 171 664 205
rect 698 171 706 205
rect 653 101 706 171
rect 653 67 664 101
rect 698 67 706 101
rect 653 49 706 67
<< pdiff >>
rect 128 599 181 619
rect 128 565 136 599
rect 170 565 181 599
rect 128 506 181 565
rect 128 472 136 506
rect 170 472 181 506
rect 128 413 181 472
rect 128 379 136 413
rect 170 379 181 413
rect 128 367 181 379
rect 211 607 335 619
rect 211 573 222 607
rect 256 573 290 607
rect 324 573 335 607
rect 211 490 335 573
rect 211 456 222 490
rect 256 456 290 490
rect 324 456 335 490
rect 211 367 335 456
rect 365 367 407 619
rect 437 607 515 619
rect 437 573 459 607
rect 493 573 515 607
rect 437 512 515 573
rect 437 478 459 512
rect 493 478 515 512
rect 437 418 515 478
rect 437 384 459 418
rect 493 384 515 418
rect 437 367 515 384
rect 545 607 623 619
rect 545 573 566 607
rect 600 573 623 607
rect 545 490 623 573
rect 545 456 566 490
rect 600 456 623 490
rect 545 367 623 456
rect 653 599 706 619
rect 653 565 664 599
rect 698 565 706 599
rect 653 509 706 565
rect 653 475 664 509
rect 698 475 706 509
rect 653 418 706 475
rect 653 384 664 418
rect 698 384 706 418
rect 653 367 706 384
<< ndiffc >>
rect 47 150 81 184
rect 47 67 81 101
rect 133 169 167 203
rect 133 59 167 93
rect 274 137 308 171
rect 274 63 308 97
rect 379 65 413 99
rect 495 137 529 171
rect 495 63 529 97
rect 664 171 698 205
rect 664 67 698 101
<< pdiffc >>
rect 136 565 170 599
rect 136 472 170 506
rect 136 379 170 413
rect 222 573 256 607
rect 290 573 324 607
rect 222 456 256 490
rect 290 456 324 490
rect 459 573 493 607
rect 459 478 493 512
rect 459 384 493 418
rect 566 573 600 607
rect 566 456 600 490
rect 664 565 698 599
rect 664 475 698 509
rect 664 384 698 418
<< poly >>
rect 181 619 211 645
rect 335 619 365 645
rect 407 619 437 645
rect 515 619 545 645
rect 623 619 653 645
rect 181 304 211 367
rect 335 335 365 367
rect 299 319 365 335
rect 181 303 218 304
rect 80 287 218 303
rect 80 253 100 287
rect 134 253 168 287
rect 202 253 218 287
rect 299 285 315 319
rect 349 285 365 319
rect 299 269 365 285
rect 407 335 437 367
rect 515 335 545 367
rect 407 319 473 335
rect 407 285 423 319
rect 457 285 473 319
rect 407 269 473 285
rect 515 319 581 335
rect 515 285 531 319
rect 565 285 581 319
rect 515 269 581 285
rect 80 237 218 253
rect 92 215 122 237
rect 319 217 349 269
rect 443 217 473 269
rect 551 217 581 269
rect 623 325 653 367
rect 623 309 743 325
rect 623 275 693 309
rect 727 275 743 309
rect 623 259 743 275
rect 623 217 653 259
rect 92 21 122 47
rect 319 23 349 49
rect 443 23 473 49
rect 551 23 581 49
rect 623 23 653 49
<< polycont >>
rect 100 253 134 287
rect 168 253 202 287
rect 315 285 349 319
rect 423 285 457 319
rect 531 285 565 319
rect 693 275 727 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 599 172 615
rect 17 565 136 599
rect 170 565 172 599
rect 17 506 172 565
rect 17 472 136 506
rect 170 472 172 506
rect 17 413 172 472
rect 206 607 340 649
rect 206 573 222 607
rect 256 573 290 607
rect 324 573 340 607
rect 206 490 340 573
rect 206 456 222 490
rect 256 456 290 490
rect 324 456 340 490
rect 206 452 340 456
rect 443 607 509 615
rect 443 573 459 607
rect 493 573 509 607
rect 443 512 509 573
rect 443 478 459 512
rect 493 478 509 512
rect 443 418 509 478
rect 550 607 616 649
rect 550 573 566 607
rect 600 573 616 607
rect 550 490 616 573
rect 550 456 566 490
rect 600 456 616 490
rect 550 452 616 456
rect 650 599 714 615
rect 650 565 664 599
rect 698 565 714 599
rect 650 509 714 565
rect 650 475 664 509
rect 698 475 714 509
rect 650 418 714 475
rect 17 379 136 413
rect 170 379 172 413
rect 17 363 172 379
rect 217 384 459 418
rect 493 384 664 418
rect 698 384 714 418
rect 17 200 66 363
rect 217 303 265 384
rect 100 287 265 303
rect 134 253 168 287
rect 202 253 265 287
rect 299 319 365 350
rect 299 285 315 319
rect 349 285 365 319
rect 299 273 365 285
rect 407 319 473 350
rect 407 285 423 319
rect 457 285 473 319
rect 407 273 473 285
rect 507 319 641 350
rect 507 285 531 319
rect 565 285 641 319
rect 507 273 641 285
rect 677 309 751 350
rect 677 275 693 309
rect 727 275 751 309
rect 677 273 751 275
rect 100 239 265 253
rect 100 237 714 239
rect 217 205 714 237
rect 17 184 83 200
rect 17 150 47 184
rect 81 150 83 184
rect 17 101 83 150
rect 17 67 47 101
rect 81 67 83 101
rect 17 51 83 67
rect 117 169 133 203
rect 167 169 183 203
rect 648 171 664 205
rect 698 171 714 205
rect 117 93 183 169
rect 117 59 133 93
rect 167 59 183 93
rect 117 17 183 59
rect 258 137 274 171
rect 308 137 495 171
rect 529 137 545 171
rect 258 97 324 137
rect 258 63 274 97
rect 308 63 324 97
rect 258 51 324 63
rect 363 99 429 103
rect 363 65 379 99
rect 413 65 429 99
rect 363 17 429 65
rect 479 97 545 137
rect 479 63 495 97
rect 529 63 545 97
rect 479 51 545 63
rect 648 101 714 171
rect 648 67 664 101
rect 698 67 714 101
rect 648 51 714 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o211a_1
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1655968
string GDS_START 1648442
<< end >>
