magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 34 49 667 241
rect 0 0 672 49
<< scnmos >>
rect 113 47 143 215
rect 270 47 300 215
rect 342 47 372 215
rect 450 47 480 215
rect 558 47 588 215
<< scpmoshvt >>
rect 80 367 110 619
rect 270 367 300 619
rect 360 367 390 619
rect 456 367 486 619
rect 558 367 588 619
<< ndiff >>
rect 60 192 113 215
rect 60 158 68 192
rect 102 158 113 192
rect 60 103 113 158
rect 60 69 68 103
rect 102 69 113 103
rect 60 47 113 69
rect 143 127 270 215
rect 143 93 154 127
rect 188 93 225 127
rect 259 93 270 127
rect 143 47 270 93
rect 300 47 342 215
rect 372 192 450 215
rect 372 158 394 192
rect 428 158 450 192
rect 372 93 450 158
rect 372 59 394 93
rect 428 59 450 93
rect 372 47 450 59
rect 480 47 558 215
rect 588 200 641 215
rect 588 166 599 200
rect 633 166 641 200
rect 588 93 641 166
rect 588 59 599 93
rect 633 59 641 93
rect 588 47 641 59
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 503 80 565
rect 27 469 35 503
rect 69 469 80 503
rect 27 413 80 469
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 599 163 619
rect 110 565 121 599
rect 155 565 163 599
rect 110 518 163 565
rect 110 484 121 518
rect 155 484 163 518
rect 110 434 163 484
rect 110 400 121 434
rect 155 400 163 434
rect 110 367 163 400
rect 217 547 270 619
rect 217 513 225 547
rect 259 513 270 547
rect 217 413 270 513
rect 217 379 225 413
rect 259 379 270 413
rect 217 367 270 379
rect 300 597 360 619
rect 300 563 311 597
rect 345 563 360 597
rect 300 529 360 563
rect 300 495 311 529
rect 345 495 360 529
rect 300 459 360 495
rect 300 425 311 459
rect 345 425 360 459
rect 300 367 360 425
rect 390 599 456 619
rect 390 565 401 599
rect 435 565 456 599
rect 390 505 456 565
rect 390 471 401 505
rect 435 471 456 505
rect 390 413 456 471
rect 390 379 401 413
rect 435 379 456 413
rect 390 367 456 379
rect 486 607 558 619
rect 486 573 504 607
rect 538 573 558 607
rect 486 525 558 573
rect 486 491 504 525
rect 538 491 558 525
rect 486 443 558 491
rect 486 409 504 443
rect 538 409 558 443
rect 486 367 558 409
rect 588 599 641 619
rect 588 565 599 599
rect 633 565 641 599
rect 588 507 641 565
rect 588 473 599 507
rect 633 473 641 507
rect 588 413 641 473
rect 588 379 599 413
rect 633 379 641 413
rect 588 367 641 379
<< ndiffc >>
rect 68 158 102 192
rect 68 69 102 103
rect 154 93 188 127
rect 225 93 259 127
rect 394 158 428 192
rect 394 59 428 93
rect 599 166 633 200
rect 599 59 633 93
<< pdiffc >>
rect 35 565 69 599
rect 35 469 69 503
rect 35 379 69 413
rect 121 565 155 599
rect 121 484 155 518
rect 121 400 155 434
rect 225 513 259 547
rect 225 379 259 413
rect 311 563 345 597
rect 311 495 345 529
rect 311 425 345 459
rect 401 565 435 599
rect 401 471 435 505
rect 401 379 435 413
rect 504 573 538 607
rect 504 491 538 525
rect 504 409 538 443
rect 599 565 633 599
rect 599 473 633 507
rect 599 379 633 413
<< poly >>
rect 80 619 110 645
rect 270 619 300 645
rect 360 619 390 645
rect 456 619 486 645
rect 558 619 588 645
rect 80 308 110 367
rect 80 292 175 308
rect 270 303 300 367
rect 360 303 390 367
rect 456 303 486 367
rect 558 303 588 367
rect 80 258 125 292
rect 159 258 175 292
rect 80 242 175 258
rect 228 287 300 303
rect 228 253 244 287
rect 278 253 300 287
rect 113 215 143 242
rect 228 237 300 253
rect 270 215 300 237
rect 342 287 408 303
rect 342 253 358 287
rect 392 253 408 287
rect 342 237 408 253
rect 450 287 516 303
rect 450 253 466 287
rect 500 253 516 287
rect 450 237 516 253
rect 558 287 631 303
rect 558 253 581 287
rect 615 253 631 287
rect 558 237 631 253
rect 342 215 372 237
rect 450 215 480 237
rect 558 215 588 237
rect 113 21 143 47
rect 270 21 300 47
rect 342 21 372 47
rect 450 21 480 47
rect 558 21 588 47
<< polycont >>
rect 125 258 159 292
rect 244 253 278 287
rect 358 253 392 287
rect 466 253 500 287
rect 581 253 615 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 18 599 75 615
rect 18 565 35 599
rect 69 565 75 599
rect 18 503 75 565
rect 18 469 35 503
rect 69 469 75 503
rect 18 413 75 469
rect 18 379 35 413
rect 69 379 75 413
rect 109 599 356 615
rect 109 565 121 599
rect 155 597 356 599
rect 155 581 311 597
rect 155 565 171 581
rect 109 518 171 565
rect 309 563 311 581
rect 345 563 356 597
rect 109 484 121 518
rect 155 484 171 518
rect 109 434 171 484
rect 109 400 121 434
rect 155 400 171 434
rect 109 384 171 400
rect 209 513 225 547
rect 259 513 275 547
rect 209 413 275 513
rect 18 203 75 379
rect 209 379 225 413
rect 259 379 275 413
rect 309 529 356 563
rect 309 495 311 529
rect 345 495 356 529
rect 309 459 356 495
rect 309 425 311 459
rect 345 425 356 459
rect 309 409 356 425
rect 390 599 454 615
rect 390 565 401 599
rect 435 565 454 599
rect 390 505 454 565
rect 390 471 401 505
rect 435 471 454 505
rect 390 413 454 471
rect 209 375 275 379
rect 390 379 401 413
rect 435 379 454 413
rect 488 607 554 649
rect 488 573 504 607
rect 538 573 554 607
rect 488 525 554 573
rect 488 491 504 525
rect 538 491 554 525
rect 488 443 554 491
rect 488 409 504 443
rect 538 409 554 443
rect 595 599 649 615
rect 595 565 599 599
rect 633 565 649 599
rect 595 507 649 565
rect 595 473 599 507
rect 633 473 649 507
rect 595 413 649 473
rect 390 375 454 379
rect 595 379 599 413
rect 633 379 649 413
rect 595 375 649 379
rect 109 292 172 350
rect 209 341 649 375
rect 109 258 125 292
rect 159 258 172 292
rect 109 242 172 258
rect 206 287 278 303
rect 206 253 244 287
rect 206 237 278 253
rect 312 287 408 303
rect 312 253 358 287
rect 392 253 408 287
rect 312 242 408 253
rect 462 287 547 303
rect 462 253 466 287
rect 500 253 547 287
rect 462 237 547 253
rect 581 287 655 303
rect 615 253 655 287
rect 581 237 655 253
rect 18 192 444 203
rect 18 158 68 192
rect 102 169 394 192
rect 102 158 104 169
rect 18 103 104 158
rect 378 158 394 169
rect 428 158 444 192
rect 18 69 68 103
rect 102 69 104 103
rect 18 53 104 69
rect 138 127 275 135
rect 138 93 154 127
rect 188 93 225 127
rect 259 93 275 127
rect 138 17 275 93
rect 378 93 444 158
rect 378 59 394 93
rect 428 59 444 93
rect 490 65 547 237
rect 583 200 649 203
rect 583 166 599 200
rect 633 166 649 200
rect 583 93 649 166
rect 378 51 444 59
rect 583 59 599 93
rect 633 59 649 93
rect 583 17 649 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a221oi_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5032070
string GDS_START 5024358
<< end >>
