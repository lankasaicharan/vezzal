magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3122 1975
<< nwell >>
rect -38 331 1862 704
rect 1025 299 1498 331
<< pwell >>
rect 1 157 197 289
rect 1627 165 1823 249
rect 1518 157 1823 165
rect 1 49 1823 157
rect 0 0 1824 49
<< scnmos >>
rect 84 179 114 263
rect 294 47 324 131
rect 446 47 476 131
rect 560 47 590 131
rect 632 47 662 131
rect 753 47 783 131
rect 831 47 861 131
rect 903 47 933 131
rect 989 47 1019 131
rect 1061 47 1091 131
rect 1259 47 1289 131
rect 1331 47 1361 131
rect 1403 47 1433 131
rect 1601 55 1631 139
rect 1710 55 1740 223
<< scpmoshvt >>
rect 84 483 114 611
rect 283 491 313 619
rect 505 491 535 619
rect 591 491 621 619
rect 690 491 720 619
rect 799 419 849 619
rect 897 419 947 619
rect 1118 335 1168 535
rect 1247 335 1277 463
rect 1361 335 1391 463
rect 1587 367 1617 495
rect 1710 367 1740 619
<< ndiff >>
rect 27 238 84 263
rect 27 204 39 238
rect 73 204 84 238
rect 27 179 84 204
rect 114 238 171 263
rect 114 204 125 238
rect 159 204 171 238
rect 114 179 171 204
rect 1653 211 1710 223
rect 1653 177 1665 211
rect 1699 177 1710 211
rect 1653 139 1710 177
rect 237 104 294 131
rect 237 70 249 104
rect 283 70 294 104
rect 237 47 294 70
rect 324 73 446 131
rect 324 47 381 73
rect 369 39 381 47
rect 415 47 446 73
rect 476 110 560 131
rect 476 76 488 110
rect 522 76 560 110
rect 476 47 560 76
rect 590 47 632 131
rect 662 110 753 131
rect 662 76 708 110
rect 742 76 753 110
rect 662 47 753 76
rect 783 47 831 131
rect 861 47 903 131
rect 933 106 989 131
rect 933 72 944 106
rect 978 72 989 106
rect 933 47 989 72
rect 1019 47 1061 131
rect 1091 110 1148 131
rect 1091 76 1102 110
rect 1136 76 1148 110
rect 1091 47 1148 76
rect 1202 110 1259 131
rect 1202 76 1214 110
rect 1248 76 1259 110
rect 1202 47 1259 76
rect 1289 47 1331 131
rect 1361 47 1403 131
rect 1433 99 1490 131
rect 1433 65 1444 99
rect 1478 65 1490 99
rect 1433 47 1490 65
rect 1544 103 1601 139
rect 1544 69 1556 103
rect 1590 69 1601 103
rect 1544 55 1601 69
rect 1631 101 1710 139
rect 1631 67 1665 101
rect 1699 67 1710 101
rect 1631 55 1710 67
rect 1740 211 1797 223
rect 1740 177 1751 211
rect 1785 177 1797 211
rect 1740 101 1797 177
rect 1740 67 1751 101
rect 1785 67 1797 101
rect 1740 55 1797 67
rect 415 39 427 47
rect 369 27 427 39
<< pdiff >>
rect 27 599 84 611
rect 27 565 39 599
rect 73 565 84 599
rect 27 529 84 565
rect 27 495 39 529
rect 73 495 84 529
rect 27 483 84 495
rect 114 599 171 611
rect 114 565 125 599
rect 159 565 171 599
rect 114 529 171 565
rect 114 495 125 529
rect 159 495 171 529
rect 114 483 171 495
rect 226 568 283 619
rect 226 534 238 568
rect 272 534 283 568
rect 226 491 283 534
rect 313 606 505 619
rect 313 572 338 606
rect 372 572 505 606
rect 313 491 505 572
rect 535 539 591 619
rect 535 505 546 539
rect 580 505 591 539
rect 535 491 591 505
rect 621 491 690 619
rect 720 498 799 619
rect 720 491 754 498
rect 742 464 754 491
rect 788 464 799 498
rect 742 419 799 464
rect 849 419 897 619
rect 947 566 1004 619
rect 1639 607 1710 619
rect 947 532 958 566
rect 992 532 1004 566
rect 947 419 1004 532
rect 1061 381 1118 535
rect 1061 347 1073 381
rect 1107 347 1118 381
rect 1061 335 1118 347
rect 1168 520 1225 535
rect 1168 486 1179 520
rect 1213 486 1225 520
rect 1168 463 1225 486
rect 1168 335 1247 463
rect 1277 451 1361 463
rect 1277 417 1316 451
rect 1350 417 1361 451
rect 1277 381 1361 417
rect 1277 347 1316 381
rect 1350 347 1361 381
rect 1277 335 1361 347
rect 1391 451 1462 463
rect 1391 417 1416 451
rect 1450 417 1462 451
rect 1391 381 1462 417
rect 1391 347 1416 381
rect 1450 347 1462 381
rect 1391 335 1462 347
rect 1639 573 1651 607
rect 1685 573 1710 607
rect 1639 510 1710 573
rect 1639 495 1651 510
rect 1530 483 1587 495
rect 1530 449 1542 483
rect 1576 449 1587 483
rect 1530 413 1587 449
rect 1530 379 1542 413
rect 1576 379 1587 413
rect 1530 367 1587 379
rect 1617 476 1651 495
rect 1685 476 1710 510
rect 1617 413 1710 476
rect 1617 379 1651 413
rect 1685 379 1710 413
rect 1617 367 1710 379
rect 1740 599 1797 619
rect 1740 565 1751 599
rect 1785 565 1797 599
rect 1740 506 1797 565
rect 1740 472 1751 506
rect 1785 472 1797 506
rect 1740 413 1797 472
rect 1740 379 1751 413
rect 1785 379 1797 413
rect 1740 367 1797 379
<< ndiffc >>
rect 39 204 73 238
rect 125 204 159 238
rect 1665 177 1699 211
rect 249 70 283 104
rect 381 39 415 73
rect 488 76 522 110
rect 708 76 742 110
rect 944 72 978 106
rect 1102 76 1136 110
rect 1214 76 1248 110
rect 1444 65 1478 99
rect 1556 69 1590 103
rect 1665 67 1699 101
rect 1751 177 1785 211
rect 1751 67 1785 101
<< pdiffc >>
rect 39 565 73 599
rect 39 495 73 529
rect 125 565 159 599
rect 125 495 159 529
rect 238 534 272 568
rect 338 572 372 606
rect 546 505 580 539
rect 754 464 788 498
rect 958 532 992 566
rect 1073 347 1107 381
rect 1179 486 1213 520
rect 1316 417 1350 451
rect 1316 347 1350 381
rect 1416 417 1450 451
rect 1416 347 1450 381
rect 1651 573 1685 607
rect 1542 449 1576 483
rect 1542 379 1576 413
rect 1651 476 1685 510
rect 1651 379 1685 413
rect 1751 565 1785 599
rect 1751 472 1785 506
rect 1751 379 1785 413
<< poly >>
rect 84 611 114 637
rect 283 619 313 645
rect 505 619 535 645
rect 591 619 621 645
rect 690 619 720 645
rect 799 619 849 645
rect 897 619 947 645
rect 1710 619 1740 645
rect 84 355 114 483
rect 175 375 241 391
rect 175 355 191 375
rect 84 341 191 355
rect 225 341 241 375
rect 84 325 241 341
rect 84 263 114 325
rect 283 223 313 491
rect 505 469 535 491
rect 355 443 535 469
rect 355 409 371 443
rect 405 439 535 443
rect 591 459 621 491
rect 690 459 720 491
rect 591 443 720 459
rect 405 409 421 439
rect 355 393 421 409
rect 591 409 645 443
rect 679 429 720 443
rect 679 409 695 429
rect 1118 557 1617 587
rect 1118 535 1168 557
rect 591 393 695 409
rect 197 207 313 223
rect 84 153 114 179
rect 197 173 213 207
rect 247 187 313 207
rect 372 219 402 393
rect 591 391 621 393
rect 463 375 621 391
rect 799 375 849 419
rect 463 341 479 375
rect 513 341 621 375
rect 737 345 849 375
rect 897 381 947 419
rect 897 365 983 381
rect 897 351 933 365
rect 463 325 621 341
rect 669 315 767 345
rect 917 331 933 351
rect 967 331 983 365
rect 1247 463 1277 489
rect 1361 463 1391 489
rect 917 315 983 331
rect 669 277 699 315
rect 524 261 699 277
rect 809 287 875 303
rect 809 267 825 287
rect 524 227 540 261
rect 574 247 699 261
rect 753 253 825 267
rect 859 253 875 287
rect 574 227 590 247
rect 372 203 438 219
rect 524 211 590 227
rect 247 173 324 187
rect 197 157 324 173
rect 294 131 324 157
rect 372 169 388 203
rect 422 183 438 203
rect 422 169 476 183
rect 372 153 476 169
rect 446 131 476 153
rect 560 131 590 211
rect 632 131 662 247
rect 753 237 875 253
rect 753 131 783 237
rect 917 189 947 315
rect 1118 235 1168 335
rect 1247 303 1277 335
rect 831 159 947 189
rect 989 219 1168 235
rect 989 185 1005 219
rect 1039 205 1168 219
rect 1216 287 1289 303
rect 1216 253 1232 287
rect 1266 253 1289 287
rect 1216 219 1289 253
rect 1361 221 1391 335
rect 1485 299 1515 557
rect 1587 495 1617 557
rect 1587 341 1617 367
rect 1710 329 1740 367
rect 1667 313 1740 329
rect 1485 269 1547 299
rect 1039 185 1091 205
rect 989 169 1091 185
rect 1216 185 1232 219
rect 1266 185 1289 219
rect 1216 169 1289 185
rect 831 131 861 159
rect 903 131 933 159
rect 989 131 1019 169
rect 1061 131 1091 169
rect 1259 131 1289 169
rect 1331 205 1469 221
rect 1331 191 1419 205
rect 1331 131 1361 191
rect 1403 171 1419 191
rect 1453 171 1469 205
rect 1517 215 1547 269
rect 1667 279 1683 313
rect 1717 279 1740 313
rect 1667 263 1740 279
rect 1710 223 1740 263
rect 1517 185 1631 215
rect 1403 155 1469 171
rect 1403 131 1433 155
rect 1601 139 1631 185
rect 294 21 324 47
rect 446 21 476 47
rect 560 21 590 47
rect 632 21 662 47
rect 753 21 783 47
rect 831 21 861 47
rect 903 21 933 47
rect 989 21 1019 47
rect 1061 21 1091 47
rect 1259 21 1289 47
rect 1331 21 1361 47
rect 1403 21 1433 47
rect 1601 29 1631 55
rect 1710 29 1740 55
<< polycont >>
rect 191 341 225 375
rect 371 409 405 443
rect 645 409 679 443
rect 213 173 247 207
rect 479 341 513 375
rect 933 331 967 365
rect 540 227 574 261
rect 825 253 859 287
rect 388 169 422 203
rect 1005 185 1039 219
rect 1232 253 1266 287
rect 1232 185 1266 219
rect 1419 171 1453 205
rect 1683 279 1717 313
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 23 599 73 649
rect 23 565 39 599
rect 23 529 73 565
rect 23 495 39 529
rect 23 479 73 495
rect 107 599 175 615
rect 107 565 125 599
rect 159 565 175 599
rect 107 529 175 565
rect 107 495 125 529
rect 159 495 175 529
rect 107 479 175 495
rect 222 568 288 615
rect 222 534 238 568
rect 272 534 288 568
rect 322 606 388 649
rect 322 572 338 606
rect 372 572 388 606
rect 322 555 388 572
rect 462 581 875 615
rect 222 521 288 534
rect 222 487 421 521
rect 107 291 141 479
rect 355 443 421 487
rect 355 409 371 443
rect 405 409 421 443
rect 355 393 421 409
rect 462 391 496 581
rect 530 539 596 547
rect 530 505 546 539
rect 580 505 596 539
rect 530 489 596 505
rect 175 375 241 391
rect 175 341 191 375
rect 225 359 241 375
rect 462 375 528 391
rect 462 359 479 375
rect 225 341 479 359
rect 513 341 528 375
rect 175 325 528 341
rect 562 359 596 489
rect 630 443 695 581
rect 630 409 645 443
rect 679 409 695 443
rect 630 393 695 409
rect 738 498 804 547
rect 738 464 754 498
rect 788 464 804 498
rect 738 415 804 464
rect 841 449 875 581
rect 942 581 1031 615
rect 942 566 991 581
rect 1025 578 1031 581
rect 1635 607 1701 649
rect 942 532 958 566
rect 1025 547 1229 578
rect 992 544 1229 547
rect 992 532 1031 544
rect 942 483 1031 532
rect 1163 539 1229 544
rect 1635 573 1651 607
rect 1685 573 1701 607
rect 1163 520 1466 539
rect 1163 486 1179 520
rect 1213 505 1466 520
rect 1213 486 1229 505
rect 1163 483 1229 486
rect 1316 451 1366 467
rect 841 417 1316 449
rect 1350 417 1366 451
rect 841 415 1366 417
rect 562 325 658 359
rect 23 238 73 267
rect 23 204 39 238
rect 23 17 73 204
rect 107 261 590 291
rect 107 257 540 261
rect 107 238 159 257
rect 107 204 125 238
rect 524 227 540 257
rect 574 227 590 261
rect 107 175 159 204
rect 197 207 263 223
rect 197 173 213 207
rect 247 173 263 207
rect 197 157 263 173
rect 372 203 438 219
rect 524 211 590 227
rect 372 169 388 203
rect 422 169 438 203
rect 372 157 438 169
rect 297 123 438 157
rect 624 135 658 325
rect 738 203 772 415
rect 841 303 875 415
rect 1316 381 1366 415
rect 917 365 1073 381
rect 917 331 933 365
rect 967 347 1073 365
rect 1107 347 1123 381
rect 967 331 1123 347
rect 917 315 1123 331
rect 809 287 875 303
rect 809 253 825 287
rect 859 253 875 287
rect 809 237 875 253
rect 989 219 1055 235
rect 989 203 1005 219
rect 233 104 331 123
rect 233 70 249 104
rect 283 70 331 104
rect 472 110 658 135
rect 233 51 331 70
rect 365 73 431 89
rect 365 39 381 73
rect 415 39 431 73
rect 472 76 488 110
rect 522 101 658 110
rect 692 185 1005 203
rect 1039 185 1055 219
rect 692 169 1055 185
rect 692 110 758 169
rect 1089 135 1123 315
rect 1177 287 1282 356
rect 1177 253 1232 287
rect 1266 253 1282 287
rect 1177 219 1282 253
rect 1177 185 1232 219
rect 1266 185 1282 219
rect 1177 169 1282 185
rect 1350 347 1366 381
rect 1316 135 1366 347
rect 1400 451 1466 505
rect 1635 510 1701 573
rect 1400 417 1416 451
rect 1450 417 1466 451
rect 1400 381 1466 417
rect 1400 347 1416 381
rect 1450 347 1466 381
rect 1526 483 1592 499
rect 1526 449 1542 483
rect 1576 449 1592 483
rect 1526 413 1592 449
rect 1526 379 1542 413
rect 1576 379 1592 413
rect 1526 363 1592 379
rect 1635 476 1651 510
rect 1685 476 1701 510
rect 1635 413 1701 476
rect 1635 379 1651 413
rect 1685 379 1701 413
rect 1635 363 1701 379
rect 1735 599 1801 615
rect 1735 565 1751 599
rect 1785 565 1801 599
rect 1735 506 1801 565
rect 1735 472 1751 506
rect 1785 472 1801 506
rect 1735 413 1801 472
rect 1735 379 1751 413
rect 1785 379 1801 413
rect 1735 363 1801 379
rect 1400 331 1466 347
rect 1558 329 1592 363
rect 1558 313 1733 329
rect 1403 205 1511 282
rect 1403 171 1419 205
rect 1453 171 1511 205
rect 1403 155 1511 171
rect 1558 279 1683 313
rect 1717 279 1733 313
rect 1558 263 1733 279
rect 522 76 538 101
rect 472 51 538 76
rect 692 76 708 110
rect 742 76 758 110
rect 692 51 758 76
rect 928 106 994 135
rect 928 72 944 106
rect 978 72 994 106
rect 365 17 431 39
rect 928 17 994 72
rect 1086 110 1152 135
rect 1086 76 1102 110
rect 1136 76 1152 110
rect 1086 51 1152 76
rect 1198 110 1366 135
rect 1558 121 1606 263
rect 1767 227 1801 363
rect 1198 76 1214 110
rect 1248 101 1366 110
rect 1248 76 1264 101
rect 1198 51 1264 76
rect 1428 99 1494 121
rect 1428 65 1444 99
rect 1478 65 1494 99
rect 1428 17 1494 65
rect 1540 103 1606 121
rect 1540 69 1556 103
rect 1590 69 1606 103
rect 1540 51 1606 69
rect 1649 211 1699 227
rect 1649 177 1665 211
rect 1649 101 1699 177
rect 1649 67 1665 101
rect 1649 17 1699 67
rect 1735 211 1801 227
rect 1735 177 1751 211
rect 1785 177 1801 211
rect 1735 101 1801 177
rect 1735 67 1751 101
rect 1785 67 1801 101
rect 1735 51 1801 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 991 566 1025 581
rect 991 547 992 566
rect 992 547 1025 566
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 14 581 1810 589
rect 14 547 991 581
rect 1025 547 1810 581
rect 14 535 1810 547
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 srdlxtp_1
flabel comment s 382 318 382 318 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 14 535 1810 589 0 FreeSans 200 0 0 0 KAPWR
port 4 nsew power bidirectional
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1471 168 1505 202 0 FreeSans 340 0 0 0 SLEEP_B
port 3 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 SLEEP_B
port 3 nsew signal input
flabel locali s 1759 94 1793 128 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 1759 168 1793 202 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4950660
string GDS_START 4937416
<< end >>
