magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 13 49 566 157
rect 0 0 672 49
<< scnmos >>
rect 100 47 130 131
rect 205 47 235 131
rect 277 47 307 131
rect 385 47 415 131
rect 457 47 487 131
<< scpmoshvt >>
rect 117 491 147 619
rect 227 491 257 619
rect 313 491 343 619
rect 421 491 451 619
rect 535 491 565 619
<< ndiff >>
rect 39 103 100 131
rect 39 69 55 103
rect 89 69 100 103
rect 39 47 100 69
rect 130 93 205 131
rect 130 59 141 93
rect 175 59 205 93
rect 130 47 205 59
rect 235 47 277 131
rect 307 106 385 131
rect 307 72 318 106
rect 352 72 385 106
rect 307 47 385 72
rect 415 47 457 131
rect 487 106 540 131
rect 487 72 498 106
rect 532 72 540 106
rect 487 47 540 72
<< pdiff >>
rect 60 607 117 619
rect 60 573 68 607
rect 102 573 117 607
rect 60 539 117 573
rect 60 505 68 539
rect 102 505 117 539
rect 60 491 117 505
rect 147 607 227 619
rect 147 573 168 607
rect 202 573 227 607
rect 147 539 227 573
rect 147 505 168 539
rect 202 505 227 539
rect 147 491 227 505
rect 257 607 313 619
rect 257 573 268 607
rect 302 573 313 607
rect 257 539 313 573
rect 257 505 268 539
rect 302 505 313 539
rect 257 491 313 505
rect 343 543 421 619
rect 343 509 368 543
rect 402 509 421 543
rect 343 491 421 509
rect 451 607 535 619
rect 451 573 478 607
rect 512 573 535 607
rect 451 539 535 573
rect 451 505 478 539
rect 512 505 535 539
rect 451 491 535 505
rect 565 607 618 619
rect 565 573 576 607
rect 610 573 618 607
rect 565 539 618 573
rect 565 505 576 539
rect 610 505 618 539
rect 565 491 618 505
<< ndiffc >>
rect 55 69 89 103
rect 141 59 175 93
rect 318 72 352 106
rect 498 72 532 106
<< pdiffc >>
rect 68 573 102 607
rect 68 505 102 539
rect 168 573 202 607
rect 168 505 202 539
rect 268 573 302 607
rect 268 505 302 539
rect 368 509 402 543
rect 478 573 512 607
rect 478 505 512 539
rect 576 573 610 607
rect 576 505 610 539
<< poly >>
rect 117 619 147 645
rect 227 619 257 645
rect 313 619 343 645
rect 421 619 451 645
rect 535 619 565 645
rect 117 289 147 491
rect 227 401 257 491
rect 313 401 343 491
rect 421 411 451 491
rect 535 424 565 491
rect 199 385 265 401
rect 199 351 215 385
rect 249 351 265 385
rect 199 317 265 351
rect 85 273 151 289
rect 85 239 101 273
rect 135 239 151 273
rect 199 283 215 317
rect 249 283 265 317
rect 199 267 265 283
rect 313 385 379 401
rect 313 351 329 385
rect 363 351 379 385
rect 313 317 379 351
rect 421 395 493 411
rect 421 361 443 395
rect 477 361 493 395
rect 421 345 493 361
rect 535 408 625 424
rect 535 374 575 408
rect 609 374 625 408
rect 313 283 329 317
rect 363 297 379 317
rect 363 283 415 297
rect 313 267 415 283
rect 85 205 151 239
rect 85 171 101 205
rect 135 171 151 205
rect 85 155 151 171
rect 100 131 130 155
rect 205 131 235 267
rect 277 203 343 219
rect 277 169 293 203
rect 327 169 343 203
rect 277 153 343 169
rect 277 131 307 153
rect 385 131 415 267
rect 457 131 487 345
rect 535 340 625 374
rect 535 306 575 340
rect 609 306 625 340
rect 535 290 625 306
rect 100 21 130 47
rect 205 21 235 47
rect 277 21 307 47
rect 385 21 415 47
rect 457 21 487 47
<< polycont >>
rect 215 351 249 385
rect 101 239 135 273
rect 215 283 249 317
rect 329 351 363 385
rect 443 361 477 395
rect 575 374 609 408
rect 329 283 363 317
rect 101 171 135 205
rect 293 169 327 203
rect 575 306 609 340
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 17 607 118 615
rect 17 573 68 607
rect 102 573 118 607
rect 17 539 118 573
rect 17 505 68 539
rect 102 505 118 539
rect 17 499 118 505
rect 152 607 218 649
rect 152 573 168 607
rect 202 573 218 607
rect 152 539 218 573
rect 152 505 168 539
rect 202 505 218 539
rect 152 499 218 505
rect 252 607 528 615
rect 252 573 268 607
rect 302 581 478 607
rect 302 573 318 581
rect 252 539 318 573
rect 462 573 478 581
rect 512 573 528 607
rect 252 505 268 539
rect 302 505 318 539
rect 252 501 318 505
rect 352 543 418 547
rect 352 509 368 543
rect 402 509 418 543
rect 17 119 67 499
rect 352 465 418 509
rect 462 539 528 573
rect 462 505 478 539
rect 512 505 528 539
rect 462 489 528 505
rect 564 607 626 649
rect 564 573 576 607
rect 610 573 626 607
rect 564 539 626 573
rect 564 505 576 539
rect 610 505 626 539
rect 564 489 626 505
rect 101 431 418 465
rect 101 273 152 431
rect 559 408 655 438
rect 135 239 152 273
rect 101 205 152 239
rect 199 385 272 397
rect 199 351 215 385
rect 249 351 272 385
rect 199 317 272 351
rect 199 283 215 317
rect 249 283 272 317
rect 199 237 272 283
rect 306 385 379 397
rect 306 351 329 385
rect 363 351 379 385
rect 306 317 379 351
rect 306 283 329 317
rect 363 283 379 317
rect 306 237 379 283
rect 413 395 493 397
rect 413 361 443 395
rect 477 361 493 395
rect 413 237 493 361
rect 559 374 575 408
rect 609 374 655 408
rect 559 340 655 374
rect 559 306 575 340
rect 609 306 655 340
rect 135 189 152 205
rect 559 203 655 306
rect 135 171 243 189
rect 101 155 243 171
rect 277 169 293 203
rect 327 169 655 203
rect 277 156 655 169
rect 209 122 243 155
rect 17 103 95 119
rect 17 69 55 103
rect 89 69 95 103
rect 17 53 95 69
rect 129 93 175 109
rect 129 59 141 93
rect 129 17 175 59
rect 209 106 356 122
rect 209 72 318 106
rect 352 72 356 106
rect 209 56 356 72
rect 482 106 548 122
rect 482 72 498 106
rect 532 72 548 106
rect 482 17 548 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a22o_0
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1139082
string GDS_START 1131472
<< end >>
