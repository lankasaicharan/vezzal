magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4370 1975
<< nwell >>
rect -38 331 3110 704
<< pwell >>
rect 2111 241 2446 263
rect 2111 229 3069 241
rect 905 223 1371 229
rect 1773 223 3069 229
rect 905 191 3069 223
rect 1 160 189 184
rect 368 160 3069 191
rect 1 49 3069 160
rect 0 0 3072 49
<< scnmos >>
rect 80 74 110 158
rect 270 50 300 134
rect 342 50 372 134
rect 474 81 504 165
rect 546 81 576 165
rect 632 81 662 165
rect 991 119 1021 203
rect 1077 119 1107 203
rect 1171 119 1201 203
rect 1243 119 1273 203
rect 1367 69 1397 197
rect 1494 69 1524 197
rect 1675 113 1705 197
rect 1747 113 1777 197
rect 1872 119 1902 203
rect 1944 119 1974 203
rect 2194 69 2224 237
rect 2333 69 2363 237
rect 2608 47 2638 215
rect 2694 47 2724 215
rect 2780 47 2810 215
rect 2866 47 2896 215
rect 2960 47 2990 215
<< scpmoshvt >>
rect 291 463 321 591
rect 377 463 407 591
rect 449 463 479 591
rect 535 463 565 591
rect 629 463 659 591
rect 746 463 776 591
rect 851 463 881 547
rect 975 463 1005 547
rect 1047 463 1077 547
rect 1167 463 1197 547
rect 1422 379 1452 547
rect 1508 379 1538 547
rect 1632 533 1662 617
rect 1750 533 1780 617
rect 1894 533 1924 617
rect 1980 533 2010 617
rect 2194 367 2224 619
rect 2333 367 2363 619
rect 2608 367 2638 619
rect 2694 367 2724 619
rect 2780 367 2810 619
rect 2874 367 2904 619
rect 2960 367 2990 619
<< ndiff >>
rect 27 133 80 158
rect 27 99 35 133
rect 69 99 80 133
rect 27 74 80 99
rect 110 122 163 158
rect 394 157 474 165
rect 394 134 406 157
rect 110 88 121 122
rect 155 88 163 122
rect 110 74 163 88
rect 217 109 270 134
rect 217 75 225 109
rect 259 75 270 109
rect 217 50 270 75
rect 300 50 342 134
rect 372 123 406 134
rect 440 123 474 157
rect 372 81 474 123
rect 504 81 546 165
rect 576 123 632 165
rect 576 89 587 123
rect 621 89 632 123
rect 576 81 632 89
rect 662 129 715 165
rect 662 95 673 129
rect 707 95 715 129
rect 662 81 715 95
rect 372 50 452 81
rect 931 178 991 203
rect 931 144 939 178
rect 973 144 991 178
rect 931 119 991 144
rect 1021 178 1077 203
rect 1021 144 1032 178
rect 1066 144 1077 178
rect 1021 119 1077 144
rect 1107 119 1171 203
rect 1201 119 1243 203
rect 1273 197 1345 203
rect 2137 229 2194 237
rect 1799 197 1872 203
rect 1273 183 1367 197
rect 1273 149 1303 183
rect 1337 149 1367 183
rect 1273 119 1367 149
rect 1295 115 1367 119
rect 1295 81 1303 115
rect 1337 81 1367 115
rect 1295 69 1367 81
rect 1397 185 1494 197
rect 1397 151 1427 185
rect 1461 151 1494 185
rect 1397 117 1494 151
rect 1397 83 1427 117
rect 1461 83 1494 117
rect 1397 69 1494 83
rect 1524 185 1675 197
rect 1524 151 1535 185
rect 1569 170 1675 185
rect 1569 151 1630 170
rect 1524 136 1630 151
rect 1664 136 1675 170
rect 1524 117 1675 136
rect 1524 83 1535 117
rect 1569 113 1675 117
rect 1705 113 1747 197
rect 1777 177 1872 197
rect 1777 143 1807 177
rect 1841 143 1872 177
rect 1777 119 1872 143
rect 1902 119 1944 203
rect 1974 177 2027 203
rect 1974 143 1985 177
rect 2019 143 2027 177
rect 1974 119 2027 143
rect 2137 195 2149 229
rect 2183 195 2194 229
rect 1777 113 1849 119
rect 1569 83 1577 113
rect 1524 69 1577 83
rect 2137 69 2194 195
rect 2224 89 2333 237
rect 2224 69 2251 89
rect 2239 55 2251 69
rect 2285 69 2333 89
rect 2363 229 2420 237
rect 2363 195 2374 229
rect 2408 195 2420 229
rect 2363 69 2420 195
rect 2555 185 2608 215
rect 2555 151 2563 185
rect 2597 151 2608 185
rect 2555 101 2608 151
rect 2285 55 2297 69
rect 2239 47 2297 55
rect 2555 67 2563 101
rect 2597 67 2608 101
rect 2555 47 2608 67
rect 2638 124 2694 215
rect 2638 90 2649 124
rect 2683 90 2694 124
rect 2638 47 2694 90
rect 2724 203 2780 215
rect 2724 169 2735 203
rect 2769 169 2780 203
rect 2724 101 2780 169
rect 2724 67 2735 101
rect 2769 67 2780 101
rect 2724 47 2780 67
rect 2810 173 2866 215
rect 2810 139 2821 173
rect 2855 139 2866 173
rect 2810 89 2866 139
rect 2810 55 2821 89
rect 2855 55 2866 89
rect 2810 47 2866 55
rect 2896 203 2960 215
rect 2896 169 2907 203
rect 2941 169 2960 203
rect 2896 101 2960 169
rect 2896 67 2907 101
rect 2941 67 2960 101
rect 2896 47 2960 67
rect 2990 161 3043 215
rect 2990 127 3001 161
rect 3035 127 3043 161
rect 2990 93 3043 127
rect 2990 59 3001 93
rect 3035 59 3043 93
rect 2990 47 3043 59
<< pdiff >>
rect 238 579 291 591
rect 238 545 246 579
rect 280 545 291 579
rect 238 509 291 545
rect 238 475 246 509
rect 280 475 291 509
rect 238 463 291 475
rect 321 579 377 591
rect 321 545 332 579
rect 366 545 377 579
rect 321 509 377 545
rect 321 475 332 509
rect 366 475 377 509
rect 321 463 377 475
rect 407 463 449 591
rect 479 579 535 591
rect 479 545 490 579
rect 524 545 535 579
rect 479 509 535 545
rect 479 475 490 509
rect 524 475 535 509
rect 479 463 535 475
rect 565 463 629 591
rect 659 571 746 591
rect 659 537 687 571
rect 721 537 746 571
rect 659 463 746 537
rect 776 577 829 591
rect 776 543 787 577
rect 821 547 829 577
rect 1342 561 1400 569
rect 821 543 851 547
rect 776 509 851 543
rect 776 475 787 509
rect 821 475 851 509
rect 776 463 851 475
rect 881 522 975 547
rect 881 488 911 522
rect 945 488 975 522
rect 881 463 975 488
rect 1005 463 1047 547
rect 1077 535 1167 547
rect 1077 501 1090 535
rect 1124 501 1167 535
rect 1077 463 1167 501
rect 1197 522 1250 547
rect 1197 488 1208 522
rect 1242 488 1250 522
rect 1197 463 1250 488
rect 1342 527 1354 561
rect 1388 547 1400 561
rect 1560 547 1632 617
rect 1388 527 1422 547
rect 1342 379 1422 527
rect 1452 421 1508 547
rect 1452 387 1463 421
rect 1497 387 1508 421
rect 1452 379 1508 387
rect 1538 533 1632 547
rect 1662 533 1750 617
rect 1780 605 1894 617
rect 1780 571 1817 605
rect 1851 571 1894 605
rect 1780 533 1894 571
rect 1924 605 1980 617
rect 1924 571 1935 605
rect 1969 571 1980 605
rect 1924 533 1980 571
rect 2010 605 2086 617
rect 2010 571 2044 605
rect 2078 571 2086 605
rect 2010 533 2086 571
rect 1538 493 1610 533
rect 1538 459 1563 493
rect 1597 459 1610 493
rect 1538 425 1610 459
rect 1538 391 1563 425
rect 1597 391 1610 425
rect 1538 379 1610 391
rect 2140 413 2194 619
rect 2140 379 2148 413
rect 2182 379 2194 413
rect 2140 367 2194 379
rect 2224 607 2333 619
rect 2224 573 2235 607
rect 2269 573 2333 607
rect 2224 539 2333 573
rect 2224 505 2288 539
rect 2322 505 2333 539
rect 2224 471 2333 505
rect 2224 437 2288 471
rect 2322 437 2333 471
rect 2224 367 2333 437
rect 2363 584 2416 619
rect 2363 550 2374 584
rect 2408 550 2416 584
rect 2363 367 2416 550
rect 2555 599 2608 619
rect 2555 565 2563 599
rect 2597 565 2608 599
rect 2555 505 2608 565
rect 2555 471 2563 505
rect 2597 471 2608 505
rect 2555 413 2608 471
rect 2555 379 2563 413
rect 2597 379 2608 413
rect 2555 367 2608 379
rect 2638 607 2694 619
rect 2638 573 2649 607
rect 2683 573 2694 607
rect 2638 532 2694 573
rect 2638 498 2649 532
rect 2683 498 2694 532
rect 2638 453 2694 498
rect 2638 419 2649 453
rect 2683 419 2694 453
rect 2638 367 2694 419
rect 2724 599 2780 619
rect 2724 565 2735 599
rect 2769 565 2780 599
rect 2724 505 2780 565
rect 2724 471 2735 505
rect 2769 471 2780 505
rect 2724 413 2780 471
rect 2724 379 2735 413
rect 2769 379 2780 413
rect 2724 367 2780 379
rect 2810 607 2874 619
rect 2810 573 2825 607
rect 2859 573 2874 607
rect 2810 539 2874 573
rect 2810 505 2825 539
rect 2859 505 2874 539
rect 2810 465 2874 505
rect 2810 431 2825 465
rect 2859 431 2874 465
rect 2810 367 2874 431
rect 2904 599 2960 619
rect 2904 565 2915 599
rect 2949 565 2960 599
rect 2904 505 2960 565
rect 2904 471 2915 505
rect 2949 471 2960 505
rect 2904 413 2960 471
rect 2904 379 2915 413
rect 2949 379 2960 413
rect 2904 367 2960 379
rect 2990 607 3043 619
rect 2990 573 3001 607
rect 3035 573 3043 607
rect 2990 539 3043 573
rect 2990 505 3001 539
rect 3035 505 3043 539
rect 2990 465 3043 505
rect 2990 431 3001 465
rect 3035 431 3043 465
rect 2990 367 3043 431
<< ndiffc >>
rect 35 99 69 133
rect 121 88 155 122
rect 225 75 259 109
rect 406 123 440 157
rect 587 89 621 123
rect 673 95 707 129
rect 939 144 973 178
rect 1032 144 1066 178
rect 1303 149 1337 183
rect 1303 81 1337 115
rect 1427 151 1461 185
rect 1427 83 1461 117
rect 1535 151 1569 185
rect 1630 136 1664 170
rect 1535 83 1569 117
rect 1807 143 1841 177
rect 1985 143 2019 177
rect 2149 195 2183 229
rect 2251 55 2285 89
rect 2374 195 2408 229
rect 2563 151 2597 185
rect 2563 67 2597 101
rect 2649 90 2683 124
rect 2735 169 2769 203
rect 2735 67 2769 101
rect 2821 139 2855 173
rect 2821 55 2855 89
rect 2907 169 2941 203
rect 2907 67 2941 101
rect 3001 127 3035 161
rect 3001 59 3035 93
<< pdiffc >>
rect 246 545 280 579
rect 246 475 280 509
rect 332 545 366 579
rect 332 475 366 509
rect 490 545 524 579
rect 490 475 524 509
rect 687 537 721 571
rect 787 543 821 577
rect 787 475 821 509
rect 911 488 945 522
rect 1090 501 1124 535
rect 1208 488 1242 522
rect 1354 527 1388 561
rect 1463 387 1497 421
rect 1817 571 1851 605
rect 1935 571 1969 605
rect 2044 571 2078 605
rect 1563 459 1597 493
rect 1563 391 1597 425
rect 2148 379 2182 413
rect 2235 573 2269 607
rect 2288 505 2322 539
rect 2288 437 2322 471
rect 2374 550 2408 584
rect 2563 565 2597 599
rect 2563 471 2597 505
rect 2563 379 2597 413
rect 2649 573 2683 607
rect 2649 498 2683 532
rect 2649 419 2683 453
rect 2735 565 2769 599
rect 2735 471 2769 505
rect 2735 379 2769 413
rect 2825 573 2859 607
rect 2825 505 2859 539
rect 2825 431 2859 465
rect 2915 565 2949 599
rect 2915 471 2949 505
rect 2915 379 2949 413
rect 3001 573 3035 607
rect 3001 505 3035 539
rect 3001 431 3035 465
<< poly >>
rect 291 591 321 617
rect 377 591 407 617
rect 449 591 479 617
rect 535 591 565 617
rect 629 591 659 617
rect 746 591 776 617
rect 975 615 1538 645
rect 1632 617 1662 643
rect 1750 617 1780 643
rect 1894 617 1924 643
rect 1980 617 2010 643
rect 2194 619 2224 645
rect 2333 619 2363 645
rect 2608 619 2638 645
rect 2694 619 2724 645
rect 2780 619 2810 645
rect 2874 619 2904 645
rect 2960 619 2990 645
rect 851 547 881 573
rect 975 547 1005 615
rect 1047 547 1077 573
rect 1167 547 1197 573
rect 1422 547 1452 573
rect 1508 547 1538 615
rect 291 441 321 463
rect 377 441 407 463
rect 80 411 407 441
rect 80 360 110 411
rect 449 366 479 463
rect 535 420 565 463
rect 80 344 176 360
rect 80 310 126 344
rect 160 310 176 344
rect 80 276 176 310
rect 306 350 479 366
rect 521 404 587 420
rect 521 370 537 404
rect 571 370 587 404
rect 521 354 587 370
rect 629 392 659 463
rect 629 376 695 392
rect 306 316 322 350
rect 356 336 479 350
rect 629 342 645 376
rect 679 342 695 376
rect 356 316 372 336
rect 306 300 372 316
rect 80 242 126 276
rect 160 242 176 276
rect 80 226 176 242
rect 80 158 110 226
rect 234 206 300 222
rect 234 172 250 206
rect 284 172 300 206
rect 234 156 300 172
rect 270 134 300 156
rect 342 134 372 300
rect 629 308 695 342
rect 420 276 504 292
rect 629 288 645 308
rect 420 242 436 276
rect 470 242 504 276
rect 420 226 504 242
rect 474 165 504 226
rect 546 274 645 288
rect 679 274 695 308
rect 546 258 695 274
rect 546 165 576 258
rect 632 165 662 191
rect 80 48 110 74
rect 474 55 504 81
rect 546 55 576 81
rect 632 51 662 81
rect 746 51 776 463
rect 851 376 881 463
rect 851 360 933 376
rect 851 326 883 360
rect 917 326 933 360
rect 851 292 933 326
rect 851 258 883 292
rect 917 258 933 292
rect 851 242 933 258
rect 975 285 1005 463
rect 1047 399 1077 463
rect 1167 441 1197 463
rect 1167 415 1310 441
rect 1167 411 1260 415
rect 1047 383 1119 399
rect 1047 369 1069 383
rect 1053 349 1069 369
rect 1103 363 1119 383
rect 1243 381 1260 411
rect 1294 381 1310 415
rect 1243 365 1310 381
rect 1632 477 1662 533
rect 1750 477 1780 533
rect 1894 501 1924 533
rect 1872 485 1938 501
rect 1632 461 1708 477
rect 1632 427 1658 461
rect 1692 427 1708 461
rect 1632 411 1708 427
rect 1750 461 1830 477
rect 1750 427 1780 461
rect 1814 427 1830 461
rect 1750 411 1830 427
rect 1103 349 1201 363
rect 1053 333 1201 349
rect 975 255 1021 285
rect 991 203 1021 255
rect 1063 275 1129 291
rect 1063 241 1079 275
rect 1113 241 1129 275
rect 1063 225 1129 241
rect 1077 203 1107 225
rect 1171 203 1201 333
rect 1243 203 1273 365
rect 1422 291 1452 379
rect 1508 363 1538 379
rect 1508 347 1758 363
rect 1508 333 1708 347
rect 1508 327 1538 333
rect 1321 275 1452 291
rect 1675 313 1708 333
rect 1742 313 1758 347
rect 1675 297 1758 313
rect 1321 241 1337 275
rect 1371 261 1452 275
rect 1567 269 1633 285
rect 1371 241 1397 261
rect 1567 249 1583 269
rect 1321 225 1397 241
rect 1367 197 1397 225
rect 1494 235 1583 249
rect 1617 235 1633 269
rect 1494 219 1633 235
rect 1494 197 1524 219
rect 1675 197 1705 297
rect 1800 249 1830 411
rect 1747 219 1830 249
rect 1872 451 1888 485
rect 1922 451 1938 485
rect 1872 435 1938 451
rect 1747 197 1777 219
rect 1872 203 1902 435
rect 1980 291 2010 533
rect 2448 410 2514 426
rect 2448 376 2464 410
rect 2498 376 2514 410
rect 1944 275 2010 291
rect 1944 241 1960 275
rect 1994 241 2010 275
rect 1944 225 2010 241
rect 2194 335 2224 367
rect 2194 319 2268 335
rect 2194 285 2218 319
rect 2252 285 2268 319
rect 2194 269 2268 285
rect 2333 322 2363 367
rect 2448 342 2514 376
rect 2448 322 2464 342
rect 2333 308 2464 322
rect 2498 308 2514 342
rect 2333 292 2514 308
rect 2608 303 2638 367
rect 2194 237 2224 269
rect 2333 237 2363 292
rect 2572 287 2638 303
rect 2572 253 2588 287
rect 2622 253 2638 287
rect 2572 237 2638 253
rect 1944 203 1974 225
rect 991 93 1021 119
rect 1077 93 1107 119
rect 1171 93 1201 119
rect 1243 51 1273 119
rect 1675 87 1705 113
rect 270 24 300 50
rect 342 24 372 50
rect 632 21 1273 51
rect 1367 43 1397 69
rect 1494 43 1524 69
rect 1747 51 1777 113
rect 1872 93 1902 119
rect 1944 93 1974 119
rect 2049 87 2115 103
rect 2049 53 2065 87
rect 2099 53 2115 87
rect 2049 51 2115 53
rect 1747 21 2115 51
rect 2194 43 2224 69
rect 2608 215 2638 237
rect 2694 329 2724 367
rect 2780 329 2810 367
rect 2874 329 2904 367
rect 2960 329 2990 367
rect 2694 313 2990 329
rect 2694 279 2710 313
rect 2744 279 2778 313
rect 2812 279 2846 313
rect 2880 279 2914 313
rect 2948 279 2990 313
rect 2694 263 2990 279
rect 2694 215 2724 263
rect 2780 215 2810 263
rect 2866 215 2896 263
rect 2960 215 2990 263
rect 2333 43 2363 69
rect 2608 21 2638 47
rect 2694 21 2724 47
rect 2780 21 2810 47
rect 2866 21 2896 47
rect 2960 21 2990 47
<< polycont >>
rect 126 310 160 344
rect 537 370 571 404
rect 322 316 356 350
rect 645 342 679 376
rect 126 242 160 276
rect 250 172 284 206
rect 436 242 470 276
rect 645 274 679 308
rect 883 326 917 360
rect 883 258 917 292
rect 1069 349 1103 383
rect 1260 381 1294 415
rect 1658 427 1692 461
rect 1780 427 1814 461
rect 1079 241 1113 275
rect 1708 313 1742 347
rect 1337 241 1371 275
rect 1583 235 1617 269
rect 1888 451 1922 485
rect 2464 376 2498 410
rect 1960 241 1994 275
rect 2218 285 2252 319
rect 2464 308 2498 342
rect 2588 253 2622 287
rect 2065 53 2099 87
rect 2710 279 2744 313
rect 2778 279 2812 313
rect 2846 279 2880 313
rect 2914 279 2948 313
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 230 579 290 595
rect 230 545 246 579
rect 280 545 290 579
rect 230 509 290 545
rect 230 475 246 509
rect 280 475 290 509
rect 230 455 290 475
rect 324 579 382 649
rect 324 545 332 579
rect 366 545 382 579
rect 324 509 382 545
rect 324 475 332 509
rect 366 475 382 509
rect 324 459 382 475
rect 474 579 540 595
rect 474 545 490 579
rect 524 545 540 579
rect 474 509 540 545
rect 671 571 737 649
rect 671 537 687 571
rect 721 537 737 571
rect 671 529 737 537
rect 771 577 847 581
rect 771 543 787 577
rect 821 543 847 577
rect 474 475 490 509
rect 524 495 540 509
rect 771 509 847 543
rect 771 495 787 509
rect 524 475 787 495
rect 821 475 847 509
rect 474 459 847 475
rect 31 425 290 455
rect 31 404 571 425
rect 31 386 537 404
rect 31 206 76 386
rect 521 370 537 386
rect 521 354 571 370
rect 605 376 695 425
rect 110 344 176 352
rect 110 310 126 344
rect 160 310 176 344
rect 210 350 465 352
rect 210 316 322 350
rect 356 316 465 350
rect 210 314 465 316
rect 605 342 645 376
rect 679 342 695 376
rect 110 280 176 310
rect 605 308 695 342
rect 110 276 561 280
rect 110 242 126 276
rect 160 242 436 276
rect 470 242 561 276
rect 605 274 645 308
rect 679 274 695 308
rect 605 258 695 274
rect 110 241 561 242
rect 756 213 847 459
rect 881 522 965 555
rect 881 488 911 522
rect 945 488 965 522
rect 1072 535 1140 649
rect 1338 561 1404 649
rect 1801 605 1867 649
rect 1072 501 1090 535
rect 1124 501 1140 535
rect 1072 495 1140 501
rect 1174 522 1248 538
rect 1338 527 1354 561
rect 1388 527 1404 561
rect 1338 525 1404 527
rect 1440 545 1672 579
rect 1801 571 1817 605
rect 1851 571 1867 605
rect 1801 565 1867 571
rect 1919 605 2008 609
rect 1919 571 1935 605
rect 1969 571 2008 605
rect 1919 565 2008 571
rect 881 461 965 488
rect 1174 488 1208 522
rect 1242 488 1248 522
rect 1440 491 1474 545
rect 1638 531 1672 545
rect 1174 472 1248 488
rect 1174 461 1208 472
rect 881 427 1208 461
rect 1282 457 1474 491
rect 1547 493 1604 509
rect 1638 497 1938 531
rect 1547 459 1563 493
rect 1597 459 1604 493
rect 1872 485 1938 497
rect 881 360 929 376
rect 881 326 883 360
rect 917 326 929 360
rect 881 292 929 326
rect 881 258 883 292
rect 917 276 929 292
rect 881 242 895 258
rect 963 276 999 427
rect 1282 426 1316 457
rect 1242 415 1316 426
rect 1547 425 1604 459
rect 1053 383 1208 393
rect 1053 349 1069 383
rect 1103 349 1208 383
rect 1242 381 1260 415
rect 1294 381 1316 415
rect 1242 379 1316 381
rect 1423 421 1513 423
rect 1423 387 1463 421
rect 1497 387 1513 421
rect 1423 380 1513 387
rect 1547 391 1563 425
rect 1597 391 1604 425
rect 1053 345 1208 349
rect 1423 345 1463 380
rect 1547 346 1604 391
rect 1053 333 1463 345
rect 1174 311 1463 333
rect 1077 276 1123 291
rect 963 242 1043 276
rect 881 228 929 242
rect 31 172 250 206
rect 284 172 300 206
rect 581 197 847 213
rect 31 159 300 172
rect 390 194 847 197
rect 390 179 975 194
rect 390 163 615 179
rect 757 178 975 179
rect 31 133 71 159
rect 31 99 35 133
rect 69 99 71 133
rect 390 157 456 163
rect 31 83 71 99
rect 105 122 171 125
rect 105 88 121 122
rect 155 88 171 122
rect 105 17 171 88
rect 209 109 275 125
rect 390 123 406 157
rect 440 123 456 157
rect 671 129 723 145
rect 390 119 456 123
rect 571 123 637 129
rect 209 75 225 109
rect 259 85 275 109
rect 571 89 587 123
rect 621 89 637 123
rect 571 85 637 89
rect 259 75 637 85
rect 209 51 637 75
rect 671 95 673 129
rect 707 95 723 129
rect 757 144 939 178
rect 973 144 975 178
rect 757 128 975 144
rect 1009 191 1043 242
rect 1077 275 1087 276
rect 1077 241 1079 275
rect 1121 242 1123 276
rect 1113 241 1123 242
rect 1077 225 1123 241
rect 1157 275 1387 277
rect 1157 241 1337 275
rect 1371 241 1387 275
rect 1157 233 1387 241
rect 1157 191 1191 233
rect 1009 178 1191 191
rect 1009 144 1032 178
rect 1066 144 1191 178
rect 1009 128 1191 144
rect 1287 183 1353 199
rect 1287 149 1303 183
rect 1337 149 1353 183
rect 671 17 723 95
rect 1287 115 1353 149
rect 1287 81 1303 115
rect 1337 81 1353 115
rect 1287 17 1353 81
rect 1421 185 1463 311
rect 1421 151 1427 185
rect 1461 151 1463 185
rect 1421 117 1463 151
rect 1421 83 1427 117
rect 1461 83 1463 117
rect 1421 67 1463 83
rect 1497 312 1604 346
rect 1638 461 1708 463
rect 1638 427 1658 461
rect 1692 427 1708 461
rect 1638 411 1708 427
rect 1764 461 1830 463
rect 1764 427 1780 461
rect 1814 427 1830 461
rect 1872 451 1888 485
rect 1922 451 1938 485
rect 1872 449 1938 451
rect 1764 415 1830 427
rect 1974 415 2008 565
rect 2042 605 2082 649
rect 2042 571 2044 605
rect 2078 571 2082 605
rect 2042 533 2082 571
rect 2219 607 2322 649
rect 2219 573 2235 607
rect 2269 573 2322 607
rect 2219 539 2322 573
rect 2219 533 2288 539
rect 2286 505 2288 533
rect 1764 411 2008 415
rect 1497 189 1531 312
rect 1638 276 1672 411
rect 1796 381 2008 411
rect 2044 465 2252 499
rect 1706 347 1758 363
rect 1706 313 1708 347
rect 1742 345 1758 347
rect 2044 345 2078 465
rect 1742 313 2078 345
rect 1706 311 2078 313
rect 2133 413 2184 429
rect 2133 379 2148 413
rect 2182 379 2184 413
rect 1706 297 1758 311
rect 1601 269 1672 276
rect 2133 276 2184 379
rect 1567 235 1583 242
rect 1617 235 1672 269
rect 1944 261 1960 275
rect 1708 241 1960 261
rect 1994 241 2097 275
rect 1708 227 2097 241
rect 1708 189 1742 227
rect 1497 185 1742 189
rect 1497 151 1535 185
rect 1569 170 1742 185
rect 1569 151 1630 170
rect 1497 136 1630 151
rect 1664 136 1742 170
rect 1497 117 1742 136
rect 1497 83 1535 117
rect 1569 83 1742 117
rect 1497 79 1742 83
rect 1791 177 1857 193
rect 1791 143 1807 177
rect 1841 143 1857 177
rect 1791 17 1857 143
rect 1969 177 2029 193
rect 1969 143 1985 177
rect 2019 143 2029 177
rect 1969 91 2029 143
rect 2063 159 2097 227
rect 2133 242 2143 276
rect 2177 242 2184 276
rect 2218 335 2252 465
rect 2286 471 2322 505
rect 2286 437 2288 471
rect 2286 421 2322 437
rect 2361 584 2412 600
rect 2361 550 2374 584
rect 2408 550 2412 584
rect 2361 534 2412 550
rect 2548 599 2599 615
rect 2548 565 2563 599
rect 2597 565 2599 599
rect 2361 335 2397 534
rect 2548 505 2599 565
rect 2218 319 2397 335
rect 2252 285 2397 319
rect 2431 410 2514 505
rect 2431 376 2464 410
rect 2498 376 2514 410
rect 2431 342 2514 376
rect 2548 471 2563 505
rect 2597 471 2599 505
rect 2548 413 2599 471
rect 2633 607 2699 649
rect 2633 573 2649 607
rect 2683 573 2699 607
rect 2633 532 2699 573
rect 2633 498 2649 532
rect 2683 498 2699 532
rect 2633 453 2699 498
rect 2633 419 2649 453
rect 2683 419 2699 453
rect 2733 599 2775 615
rect 2733 565 2735 599
rect 2769 565 2775 599
rect 2733 505 2775 565
rect 2733 471 2735 505
rect 2769 471 2775 505
rect 2548 379 2563 413
rect 2597 385 2599 413
rect 2733 413 2775 471
rect 2809 607 2875 649
rect 2809 573 2825 607
rect 2859 573 2875 607
rect 2809 539 2875 573
rect 2809 505 2825 539
rect 2859 505 2875 539
rect 2809 465 2875 505
rect 2809 431 2825 465
rect 2859 431 2875 465
rect 2909 599 2949 615
rect 2909 565 2915 599
rect 2909 505 2949 565
rect 2909 471 2915 505
rect 2597 379 2695 385
rect 2548 351 2695 379
rect 2431 308 2464 342
rect 2498 308 2514 342
rect 2431 305 2514 308
rect 2661 313 2695 351
rect 2733 379 2735 413
rect 2769 397 2775 413
rect 2909 413 2949 471
rect 2985 607 3051 649
rect 2985 573 3001 607
rect 3035 573 3051 607
rect 2985 539 3051 573
rect 2985 505 3001 539
rect 3035 505 3051 539
rect 2985 465 3051 505
rect 2985 431 3001 465
rect 3035 431 3051 465
rect 2909 397 2915 413
rect 2769 379 2915 397
rect 2949 379 3052 397
rect 2733 347 3052 379
rect 2218 269 2397 285
rect 2572 287 2627 303
rect 2572 271 2588 287
rect 2133 233 2184 242
rect 2358 233 2397 269
rect 2460 253 2588 271
rect 2622 253 2627 287
rect 2460 237 2627 253
rect 2661 279 2710 313
rect 2744 279 2778 313
rect 2812 279 2846 313
rect 2880 279 2914 313
rect 2948 279 2964 313
rect 2133 229 2199 233
rect 2133 195 2149 229
rect 2183 195 2199 229
rect 2358 229 2424 233
rect 2358 195 2374 229
rect 2408 195 2424 229
rect 2133 193 2199 195
rect 2460 159 2494 237
rect 2661 203 2695 279
rect 3000 245 3052 347
rect 2063 125 2494 159
rect 2547 185 2695 203
rect 2547 151 2563 185
rect 2597 167 2695 185
rect 2733 211 3052 245
rect 2733 209 2958 211
rect 2733 203 2771 209
rect 2733 169 2735 203
rect 2769 169 2771 203
rect 2905 203 2958 209
rect 2597 151 2599 167
rect 2547 101 2599 151
rect 1969 87 2115 91
rect 1969 53 2065 87
rect 2099 53 2115 87
rect 1969 51 2115 53
rect 2235 89 2301 91
rect 2235 55 2251 89
rect 2285 55 2301 89
rect 2235 17 2301 55
rect 2547 67 2563 101
rect 2597 67 2599 101
rect 2547 51 2599 67
rect 2633 124 2699 133
rect 2633 90 2649 124
rect 2683 90 2699 124
rect 2633 17 2699 90
rect 2733 101 2771 169
rect 2733 67 2735 101
rect 2769 67 2771 101
rect 2733 51 2771 67
rect 2805 173 2871 175
rect 2805 139 2821 173
rect 2855 139 2871 173
rect 2805 89 2871 139
rect 2805 55 2821 89
rect 2855 55 2871 89
rect 2805 17 2871 55
rect 2905 169 2907 203
rect 2941 169 2958 203
rect 2905 101 2958 169
rect 2905 67 2907 101
rect 2941 67 2958 101
rect 2905 51 2958 67
rect 2992 161 3051 177
rect 2992 127 3001 161
rect 3035 127 3051 161
rect 2992 93 3051 127
rect 2992 59 3001 93
rect 3035 59 3051 93
rect 2992 17 3051 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 895 258 917 276
rect 917 258 929 276
rect 895 242 929 258
rect 1087 275 1121 276
rect 1087 242 1113 275
rect 1113 242 1121 275
rect 1567 269 1601 276
rect 1567 242 1583 269
rect 1583 242 1601 269
rect 2143 242 2177 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 683 3072 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 0 617 3072 649
rect 883 276 941 282
rect 883 242 895 276
rect 929 273 941 276
rect 1075 276 1133 282
rect 1075 273 1087 276
rect 929 245 1087 273
rect 929 242 941 245
rect 883 236 941 242
rect 1075 242 1087 245
rect 1121 273 1133 276
rect 1555 276 1613 282
rect 1555 273 1567 276
rect 1121 245 1567 273
rect 1121 242 1133 245
rect 1075 236 1133 242
rect 1555 242 1567 245
rect 1601 273 1613 276
rect 2131 276 2189 282
rect 2131 273 2143 276
rect 1601 245 2143 273
rect 1601 242 1613 245
rect 1555 236 1613 242
rect 2131 242 2143 245
rect 2177 242 2189 276
rect 2131 236 2189 242
rect 0 17 3072 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
rect 0 -49 3072 -17
<< labels >>
flabel pwell s 0 0 3072 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 3072 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfrtp_4
flabel comment s 1812 345 1812 345 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 3072 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 3072 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 2431 316 2465 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2431 390 2465 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2431 464 2465 498 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2911 168 2945 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3072 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3167146
string GDS_START 3145112
<< end >>
