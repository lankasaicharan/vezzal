magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 287 167 657 193
rect 1 49 657 167
rect 0 0 672 49
<< scnmos >>
rect 84 57 114 141
rect 162 57 192 141
rect 370 83 400 167
rect 456 83 486 167
rect 548 83 578 167
<< scpmoshvt >>
rect 95 419 145 619
rect 201 419 251 619
rect 334 419 384 619
rect 440 419 490 619
rect 538 419 588 619
<< ndiff >>
rect 313 142 370 167
rect 27 116 84 141
rect 27 82 39 116
rect 73 82 84 116
rect 27 57 84 82
rect 114 57 162 141
rect 192 116 249 141
rect 192 82 203 116
rect 237 82 249 116
rect 313 108 325 142
rect 359 108 370 142
rect 313 83 370 108
rect 400 142 456 167
rect 400 108 411 142
rect 445 108 456 142
rect 400 83 456 108
rect 486 129 548 167
rect 486 95 497 129
rect 531 95 548 129
rect 486 83 548 95
rect 578 142 631 167
rect 578 108 589 142
rect 623 108 631 142
rect 578 83 631 108
rect 192 57 249 82
<< pdiff >>
rect 36 607 95 619
rect 36 573 48 607
rect 82 573 95 607
rect 36 536 95 573
rect 36 502 48 536
rect 82 502 95 536
rect 36 465 95 502
rect 36 431 48 465
rect 82 431 95 465
rect 36 419 95 431
rect 145 597 201 619
rect 145 563 156 597
rect 190 563 201 597
rect 145 465 201 563
rect 145 431 156 465
rect 190 431 201 465
rect 145 419 201 431
rect 251 607 334 619
rect 251 573 262 607
rect 296 573 334 607
rect 251 473 334 573
rect 251 439 262 473
rect 296 439 334 473
rect 251 419 334 439
rect 384 597 440 619
rect 384 563 395 597
rect 429 563 440 597
rect 384 473 440 563
rect 384 439 395 473
rect 429 439 440 473
rect 384 419 440 439
rect 490 419 538 619
rect 588 607 641 619
rect 588 573 599 607
rect 633 573 641 607
rect 588 536 641 573
rect 588 502 599 536
rect 633 502 641 536
rect 588 465 641 502
rect 588 431 599 465
rect 633 431 641 465
rect 588 419 641 431
<< ndiffc >>
rect 39 82 73 116
rect 203 82 237 116
rect 325 108 359 142
rect 411 108 445 142
rect 497 95 531 129
rect 589 108 623 142
<< pdiffc >>
rect 48 573 82 607
rect 48 502 82 536
rect 48 431 82 465
rect 156 563 190 597
rect 156 431 190 465
rect 262 573 296 607
rect 262 439 296 473
rect 395 563 429 597
rect 395 439 429 473
rect 599 573 633 607
rect 599 502 633 536
rect 599 431 633 465
<< poly >>
rect 95 619 145 645
rect 201 619 251 645
rect 334 619 384 645
rect 440 619 490 645
rect 538 619 588 645
rect 95 379 145 419
rect 44 363 145 379
rect 44 329 60 363
rect 94 329 145 363
rect 44 295 145 329
rect 201 315 251 419
rect 334 387 384 419
rect 301 371 384 387
rect 301 337 317 371
rect 351 337 384 371
rect 301 321 384 337
rect 44 261 60 295
rect 94 261 145 295
rect 44 245 145 261
rect 193 299 259 315
rect 193 265 209 299
rect 243 265 259 299
rect 84 141 114 245
rect 193 231 259 265
rect 193 197 209 231
rect 243 197 259 231
rect 162 167 259 197
rect 354 212 384 321
rect 440 345 490 419
rect 538 393 588 419
rect 548 345 588 393
rect 440 329 506 345
rect 440 295 456 329
rect 490 295 506 329
rect 440 279 506 295
rect 548 329 629 345
rect 548 295 579 329
rect 613 295 629 329
rect 548 279 629 295
rect 354 182 400 212
rect 370 167 400 182
rect 456 167 486 279
rect 548 167 578 279
rect 162 141 192 167
rect 370 57 400 83
rect 456 57 486 83
rect 548 57 578 83
rect 84 31 114 57
rect 162 31 192 57
<< polycont >>
rect 60 329 94 363
rect 317 337 351 371
rect 60 261 94 295
rect 209 265 243 299
rect 209 197 243 231
rect 456 295 490 329
rect 579 295 613 329
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 32 607 98 649
rect 32 573 48 607
rect 82 573 98 607
rect 32 536 98 573
rect 32 502 48 536
rect 82 502 98 536
rect 32 465 98 502
rect 32 431 48 465
rect 82 431 98 465
rect 32 415 98 431
rect 134 597 206 613
rect 134 563 156 597
rect 190 563 206 597
rect 134 465 206 563
rect 134 431 156 465
rect 190 431 206 465
rect 134 387 206 431
rect 246 607 312 649
rect 246 573 262 607
rect 296 573 312 607
rect 246 473 312 573
rect 246 439 262 473
rect 296 439 312 473
rect 246 423 312 439
rect 379 597 445 613
rect 379 563 395 597
rect 429 563 445 597
rect 379 473 445 563
rect 379 439 395 473
rect 429 439 445 473
rect 379 423 445 439
rect 583 607 649 649
rect 583 573 599 607
rect 633 573 649 607
rect 583 536 649 573
rect 583 502 599 536
rect 633 502 649 536
rect 583 465 649 502
rect 583 431 599 465
rect 633 431 649 465
rect 25 363 98 379
rect 25 329 60 363
rect 94 329 98 363
rect 25 295 98 329
rect 25 261 60 295
rect 94 261 98 295
rect 25 236 98 261
rect 134 371 351 387
rect 134 353 317 371
rect 134 145 168 353
rect 301 337 317 353
rect 301 321 351 337
rect 204 299 263 315
rect 204 265 209 299
rect 243 265 263 299
rect 385 285 419 423
rect 583 415 649 431
rect 204 231 263 265
rect 204 197 209 231
rect 243 197 263 231
rect 204 181 263 197
rect 309 251 419 285
rect 453 329 545 356
rect 453 295 456 329
rect 490 295 545 329
rect 23 116 89 145
rect 23 82 39 116
rect 73 82 89 116
rect 134 116 253 145
rect 134 111 203 116
rect 23 17 89 82
rect 187 82 203 111
rect 237 82 253 116
rect 187 53 253 82
rect 309 142 375 251
rect 453 237 545 295
rect 579 329 652 352
rect 613 295 652 329
rect 579 237 652 295
rect 309 108 325 142
rect 359 108 375 142
rect 309 79 375 108
rect 411 169 639 203
rect 411 142 445 169
rect 583 142 639 169
rect 411 92 445 108
rect 481 129 547 135
rect 481 95 497 129
rect 531 95 547 129
rect 481 17 547 95
rect 583 108 589 142
rect 623 108 639 142
rect 583 92 639 108
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2bb2ai_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4079858
string GDS_START 4073182
<< end >>
