magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
rect 863 321 1031 331
<< pwell >>
rect 934 241 1244 249
rect 1 49 1244 241
rect 0 0 1248 49
<< scnmos >>
rect 84 47 114 215
rect 170 47 200 215
rect 270 47 300 215
rect 370 47 400 215
rect 456 47 486 215
rect 542 47 572 215
rect 628 47 658 215
rect 714 47 744 215
rect 1017 55 1047 223
rect 1131 55 1161 223
<< scpmoshvt >>
rect 84 367 114 619
rect 170 367 200 619
rect 270 367 300 619
rect 370 367 400 619
rect 470 367 500 619
rect 584 367 614 619
rect 670 367 700 619
rect 792 367 822 619
rect 1017 367 1047 619
rect 1117 367 1147 619
<< ndiff >>
rect 27 186 84 215
rect 27 152 39 186
rect 73 152 84 186
rect 27 101 84 152
rect 27 67 39 101
rect 73 67 84 101
rect 27 47 84 67
rect 114 178 170 215
rect 114 144 125 178
rect 159 144 170 178
rect 114 47 170 144
rect 200 161 270 215
rect 200 127 225 161
rect 259 127 270 161
rect 200 93 270 127
rect 200 59 225 93
rect 259 59 270 93
rect 200 47 270 59
rect 300 178 370 215
rect 300 144 325 178
rect 359 144 370 178
rect 300 47 370 144
rect 400 203 456 215
rect 400 169 411 203
rect 445 169 456 203
rect 400 101 456 169
rect 400 67 411 101
rect 445 67 456 101
rect 400 47 456 67
rect 486 177 542 215
rect 486 143 497 177
rect 531 143 542 177
rect 486 93 542 143
rect 486 59 497 93
rect 531 59 542 93
rect 486 47 542 59
rect 572 203 628 215
rect 572 169 583 203
rect 617 169 628 203
rect 572 101 628 169
rect 572 67 583 101
rect 617 67 628 101
rect 572 47 628 67
rect 658 105 714 215
rect 658 71 669 105
rect 703 71 714 105
rect 658 47 714 71
rect 744 186 801 215
rect 744 152 755 186
rect 789 152 801 186
rect 744 101 801 152
rect 744 67 755 101
rect 789 67 801 101
rect 960 186 1017 223
rect 960 152 972 186
rect 1006 152 1017 186
rect 960 101 1017 152
rect 744 47 801 67
rect 960 67 972 101
rect 1006 67 1017 101
rect 960 55 1017 67
rect 1047 211 1131 223
rect 1047 177 1072 211
rect 1106 177 1131 211
rect 1047 101 1131 177
rect 1047 67 1072 101
rect 1106 67 1131 101
rect 1047 55 1131 67
rect 1161 211 1218 223
rect 1161 177 1172 211
rect 1206 177 1218 211
rect 1161 101 1218 177
rect 1161 67 1172 101
rect 1206 67 1218 101
rect 1161 55 1218 67
<< pdiff >>
rect 27 599 84 619
rect 27 565 39 599
rect 73 565 84 599
rect 27 506 84 565
rect 27 472 39 506
rect 73 472 84 506
rect 27 413 84 472
rect 27 379 39 413
rect 73 379 84 413
rect 27 367 84 379
rect 114 531 170 619
rect 114 497 125 531
rect 159 497 170 531
rect 114 413 170 497
rect 114 379 125 413
rect 159 379 170 413
rect 114 367 170 379
rect 200 607 270 619
rect 200 573 225 607
rect 259 573 270 607
rect 200 536 270 573
rect 200 502 225 536
rect 259 502 270 536
rect 200 465 270 502
rect 200 431 225 465
rect 259 431 270 465
rect 200 367 270 431
rect 300 547 370 619
rect 300 513 325 547
rect 359 513 370 547
rect 300 413 370 513
rect 300 379 325 413
rect 359 379 370 413
rect 300 367 370 379
rect 400 599 470 619
rect 400 565 425 599
rect 459 565 470 599
rect 400 521 470 565
rect 400 487 425 521
rect 459 487 470 521
rect 400 367 470 487
rect 500 598 584 619
rect 500 564 525 598
rect 559 564 584 598
rect 500 367 584 564
rect 614 599 670 619
rect 614 565 625 599
rect 659 565 670 599
rect 614 521 670 565
rect 614 487 625 521
rect 659 487 670 521
rect 614 367 670 487
rect 700 607 792 619
rect 700 573 725 607
rect 759 573 792 607
rect 700 367 792 573
rect 822 577 879 619
rect 822 543 833 577
rect 867 543 879 577
rect 822 367 879 543
rect 937 403 1017 619
rect 937 369 949 403
rect 983 369 1017 403
rect 937 367 1017 369
rect 1047 581 1117 619
rect 1047 547 1058 581
rect 1092 547 1117 581
rect 1047 367 1117 547
rect 1147 599 1204 619
rect 1147 565 1158 599
rect 1192 565 1204 599
rect 1147 519 1204 565
rect 1147 485 1158 519
rect 1192 485 1204 519
rect 1147 440 1204 485
rect 1147 406 1158 440
rect 1192 406 1204 440
rect 1147 367 1204 406
rect 937 357 995 367
<< ndiffc >>
rect 39 152 73 186
rect 39 67 73 101
rect 125 144 159 178
rect 225 127 259 161
rect 225 59 259 93
rect 325 144 359 178
rect 411 169 445 203
rect 411 67 445 101
rect 497 143 531 177
rect 497 59 531 93
rect 583 169 617 203
rect 583 67 617 101
rect 669 71 703 105
rect 755 152 789 186
rect 755 67 789 101
rect 972 152 1006 186
rect 972 67 1006 101
rect 1072 177 1106 211
rect 1072 67 1106 101
rect 1172 177 1206 211
rect 1172 67 1206 101
<< pdiffc >>
rect 39 565 73 599
rect 39 472 73 506
rect 39 379 73 413
rect 125 497 159 531
rect 125 379 159 413
rect 225 573 259 607
rect 225 502 259 536
rect 225 431 259 465
rect 325 513 359 547
rect 325 379 359 413
rect 425 565 459 599
rect 425 487 459 521
rect 525 564 559 598
rect 625 565 659 599
rect 625 487 659 521
rect 725 573 759 607
rect 833 543 867 577
rect 949 369 983 403
rect 1058 547 1092 581
rect 1158 565 1192 599
rect 1158 485 1192 519
rect 1158 406 1192 440
<< poly >>
rect 84 619 114 645
rect 170 619 200 645
rect 270 619 300 645
rect 370 619 400 645
rect 470 619 500 645
rect 584 619 614 645
rect 670 619 700 645
rect 792 619 822 645
rect 1017 619 1047 645
rect 1117 619 1147 645
rect 84 329 114 367
rect 170 329 200 367
rect 270 329 300 367
rect 370 329 400 367
rect 84 313 400 329
rect 470 345 500 367
rect 584 345 614 367
rect 670 345 700 367
rect 792 345 822 367
rect 470 339 822 345
rect 470 315 954 339
rect 84 279 191 313
rect 225 279 259 313
rect 293 279 327 313
rect 361 279 400 313
rect 792 309 954 315
rect 84 263 400 279
rect 888 303 954 309
rect 888 269 904 303
rect 938 283 954 303
rect 1017 283 1047 367
rect 1117 335 1147 367
rect 938 269 1047 283
rect 1095 319 1161 335
rect 1095 285 1111 319
rect 1145 285 1161 319
rect 1095 269 1161 285
rect 84 215 114 263
rect 170 215 200 263
rect 270 215 300 263
rect 370 215 400 263
rect 456 237 846 267
rect 888 253 1047 269
rect 456 215 486 237
rect 542 215 572 237
rect 628 215 658 237
rect 714 215 744 237
rect 816 202 846 237
rect 1017 223 1047 253
rect 1131 223 1161 269
rect 816 186 905 202
rect 816 152 855 186
rect 889 152 905 186
rect 816 118 905 152
rect 816 84 855 118
rect 889 84 905 118
rect 816 68 905 84
rect 84 21 114 47
rect 170 21 200 47
rect 270 21 300 47
rect 370 21 400 47
rect 456 21 486 47
rect 542 21 572 47
rect 628 21 658 47
rect 714 21 744 47
rect 1017 29 1047 55
rect 1131 29 1161 55
<< polycont >>
rect 191 279 225 313
rect 259 279 293 313
rect 327 279 361 313
rect 904 269 938 303
rect 1111 285 1145 319
rect 855 152 889 186
rect 855 84 889 118
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 23 607 475 615
rect 23 599 225 607
rect 23 565 39 599
rect 73 581 225 599
rect 23 506 73 565
rect 209 573 225 581
rect 259 599 475 607
rect 259 581 425 599
rect 259 573 275 581
rect 23 472 39 506
rect 23 413 73 472
rect 23 379 39 413
rect 23 363 73 379
rect 107 531 175 547
rect 107 497 125 531
rect 159 497 175 531
rect 107 413 175 497
rect 209 536 275 573
rect 409 565 425 581
rect 459 565 475 599
rect 209 502 225 536
rect 259 502 275 536
rect 209 465 275 502
rect 209 431 225 465
rect 259 431 275 465
rect 309 513 325 547
rect 359 513 375 547
rect 107 379 125 413
rect 159 397 175 413
rect 309 413 375 513
rect 409 521 475 565
rect 509 598 575 649
rect 509 564 525 598
rect 559 564 575 598
rect 509 539 575 564
rect 609 599 675 615
rect 609 565 625 599
rect 659 565 675 599
rect 709 607 775 649
rect 709 573 725 607
rect 759 573 775 607
rect 817 577 883 615
rect 609 539 675 565
rect 817 543 833 577
rect 867 543 883 577
rect 817 539 883 543
rect 409 487 425 521
rect 459 505 475 521
rect 609 521 883 539
rect 609 505 625 521
rect 459 487 625 505
rect 659 505 883 521
rect 1042 581 1108 649
rect 1042 547 1058 581
rect 1092 547 1108 581
rect 1042 505 1108 547
rect 1142 599 1229 615
rect 1142 565 1158 599
rect 1192 565 1229 599
rect 1142 519 1229 565
rect 659 487 675 505
rect 409 471 675 487
rect 1142 485 1158 519
rect 1192 485 1229 519
rect 1142 471 1229 485
rect 865 440 1229 471
rect 865 437 1158 440
rect 309 397 325 413
rect 159 379 325 397
rect 359 379 375 413
rect 107 363 375 379
rect 409 403 899 437
rect 1142 406 1158 437
rect 1192 406 1229 440
rect 107 282 141 363
rect 409 329 443 403
rect 933 369 949 403
rect 983 369 1022 403
rect 1142 390 1229 406
rect 933 353 1022 369
rect 25 236 141 282
rect 175 313 443 329
rect 175 279 191 313
rect 225 279 259 313
rect 293 279 327 313
rect 361 295 443 313
rect 888 303 954 319
rect 361 279 377 295
rect 888 282 904 303
rect 175 263 377 279
rect 697 269 904 282
rect 938 269 954 303
rect 107 229 141 236
rect 23 186 73 202
rect 23 152 39 186
rect 23 101 73 152
rect 107 195 375 229
rect 107 178 175 195
rect 107 144 125 178
rect 159 144 175 178
rect 309 178 375 195
rect 107 119 175 144
rect 209 127 225 161
rect 259 127 275 161
rect 23 67 39 101
rect 209 93 275 127
rect 309 144 325 178
rect 359 144 375 178
rect 309 119 375 144
rect 411 227 617 261
rect 697 236 954 269
rect 411 203 445 227
rect 583 203 617 227
rect 209 85 225 93
rect 73 67 225 85
rect 23 59 225 67
rect 259 85 275 93
rect 411 101 445 169
rect 259 67 411 85
rect 259 59 445 67
rect 23 51 445 59
rect 481 177 547 193
rect 481 143 497 177
rect 531 143 547 177
rect 481 93 547 143
rect 481 59 497 93
rect 531 59 547 93
rect 481 17 547 59
rect 988 202 1022 353
rect 1081 319 1161 356
rect 1081 285 1111 319
rect 1145 285 1161 319
rect 1081 269 1161 285
rect 1195 227 1229 390
rect 617 186 805 202
rect 617 169 755 186
rect 583 168 755 169
rect 583 101 617 168
rect 739 152 755 168
rect 789 152 805 186
rect 583 51 617 67
rect 653 105 703 134
rect 653 71 669 105
rect 653 17 703 71
rect 739 101 805 152
rect 739 67 755 101
rect 789 67 805 101
rect 839 186 1022 202
rect 839 152 855 186
rect 889 152 972 186
rect 1006 152 1022 186
rect 839 118 1022 152
rect 839 84 855 118
rect 889 101 1022 118
rect 889 84 972 101
rect 839 68 972 84
rect 739 51 805 67
rect 956 67 972 68
rect 1006 67 1022 101
rect 956 51 1022 67
rect 1056 211 1122 227
rect 1056 177 1072 211
rect 1106 177 1122 211
rect 1056 101 1122 177
rect 1056 67 1072 101
rect 1106 67 1122 101
rect 1056 17 1122 67
rect 1156 211 1229 227
rect 1156 177 1172 211
rect 1206 177 1229 211
rect 1156 101 1229 177
rect 1156 67 1172 101
rect 1206 67 1229 101
rect 1156 51 1229 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ebufn_4
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3440388
string GDS_START 3430938
<< end >>
