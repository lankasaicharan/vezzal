magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2586 1852
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 1 21 1279 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 194 47 224 177
rect 475 47 505 177
rect 579 47 609 177
rect 673 47 703 177
rect 767 47 797 177
rect 875 47 905 177
rect 969 47 999 177
rect 1063 47 1093 177
rect 1167 47 1197 177
<< scpmoshvt >>
rect 81 297 117 497
rect 196 297 232 497
rect 394 309 430 497
rect 488 309 524 497
rect 582 309 618 497
rect 676 309 712 497
rect 877 297 913 497
rect 971 297 1007 497
rect 1065 297 1101 497
rect 1159 297 1195 497
<< ndiff >>
rect 27 106 79 177
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 89 194 177
rect 109 55 129 89
rect 163 55 194 89
rect 109 47 194 55
rect 224 103 286 177
rect 224 69 244 103
rect 278 69 286 103
rect 224 47 286 69
rect 413 129 475 177
rect 413 95 421 129
rect 455 95 475 129
rect 413 47 475 95
rect 505 89 579 177
rect 505 55 525 89
rect 559 55 579 89
rect 505 47 579 55
rect 609 129 673 177
rect 609 95 619 129
rect 653 95 673 129
rect 609 47 673 95
rect 703 89 767 177
rect 703 55 713 89
rect 747 55 767 89
rect 703 47 767 55
rect 797 129 875 177
rect 797 95 819 129
rect 853 95 875 129
rect 797 47 875 95
rect 905 169 969 177
rect 905 135 925 169
rect 959 135 969 169
rect 905 47 969 135
rect 999 89 1063 177
rect 999 55 1019 89
rect 1053 55 1063 89
rect 999 47 1063 55
rect 1093 169 1167 177
rect 1093 135 1113 169
rect 1147 135 1167 169
rect 1093 47 1167 135
rect 1197 89 1253 177
rect 1197 55 1207 89
rect 1241 55 1253 89
rect 1197 47 1253 55
<< pdiff >>
rect 27 477 81 497
rect 27 443 35 477
rect 69 443 81 477
rect 27 409 81 443
rect 27 375 35 409
rect 69 375 81 409
rect 27 297 81 375
rect 117 489 196 497
rect 117 455 137 489
rect 171 455 196 489
rect 117 421 196 455
rect 117 387 137 421
rect 171 387 196 421
rect 117 297 196 387
rect 232 477 286 497
rect 232 443 244 477
rect 278 443 286 477
rect 232 409 286 443
rect 232 375 244 409
rect 278 375 286 409
rect 232 297 286 375
rect 340 477 394 497
rect 340 443 348 477
rect 382 443 394 477
rect 340 309 394 443
rect 430 489 488 497
rect 430 455 442 489
rect 476 455 488 489
rect 430 309 488 455
rect 524 477 582 497
rect 524 443 536 477
rect 570 443 582 477
rect 524 309 582 443
rect 618 489 676 497
rect 618 455 630 489
rect 664 455 676 489
rect 618 309 676 455
rect 712 489 877 497
rect 712 455 742 489
rect 776 455 820 489
rect 854 455 877 489
rect 712 421 877 455
rect 712 387 742 421
rect 776 387 820 421
rect 854 387 877 421
rect 712 309 877 387
rect 729 297 877 309
rect 913 345 971 497
rect 913 311 925 345
rect 959 311 971 345
rect 913 297 971 311
rect 1007 489 1065 497
rect 1007 455 1019 489
rect 1053 455 1065 489
rect 1007 421 1065 455
rect 1007 387 1019 421
rect 1053 387 1065 421
rect 1007 297 1065 387
rect 1101 345 1159 497
rect 1101 311 1113 345
rect 1147 311 1159 345
rect 1101 297 1159 311
rect 1195 489 1253 497
rect 1195 455 1207 489
rect 1241 455 1253 489
rect 1195 421 1253 455
rect 1195 387 1207 421
rect 1241 387 1253 421
rect 1195 297 1253 387
<< ndiffc >>
rect 35 72 69 106
rect 129 55 163 89
rect 244 69 278 103
rect 421 95 455 129
rect 525 55 559 89
rect 619 95 653 129
rect 713 55 747 89
rect 819 95 853 129
rect 925 135 959 169
rect 1019 55 1053 89
rect 1113 135 1147 169
rect 1207 55 1241 89
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 137 455 171 489
rect 137 387 171 421
rect 244 443 278 477
rect 244 375 278 409
rect 348 443 382 477
rect 442 455 476 489
rect 536 443 570 477
rect 630 455 664 489
rect 742 455 776 489
rect 820 455 854 489
rect 742 387 776 421
rect 820 387 854 421
rect 925 311 959 345
rect 1019 455 1053 489
rect 1019 387 1053 421
rect 1113 311 1147 345
rect 1207 455 1241 489
rect 1207 387 1241 421
<< poly >>
rect 81 497 117 523
rect 196 497 232 523
rect 394 497 430 523
rect 488 497 524 523
rect 582 497 618 523
rect 676 497 712 523
rect 877 497 913 523
rect 971 497 1007 523
rect 1065 497 1101 523
rect 1159 497 1195 523
rect 81 282 117 297
rect 196 282 232 297
rect 394 294 430 309
rect 488 294 524 309
rect 582 294 618 309
rect 676 294 712 309
rect 301 282 714 294
rect 877 282 913 297
rect 971 282 1007 297
rect 1065 282 1101 297
rect 1159 282 1195 297
rect 79 265 119 282
rect 79 249 152 265
rect 79 215 98 249
rect 132 215 152 249
rect 79 199 152 215
rect 194 264 714 282
rect 194 252 339 264
rect 875 259 915 282
rect 969 259 1009 282
rect 1063 259 1103 282
rect 1157 259 1197 282
rect 194 249 280 252
rect 194 215 216 249
rect 250 215 280 249
rect 756 249 832 259
rect 756 222 772 249
rect 194 210 280 215
rect 475 215 772 222
rect 806 215 832 249
rect 194 205 276 210
rect 79 177 109 199
rect 194 177 224 205
rect 475 192 832 215
rect 875 249 1197 259
rect 875 215 903 249
rect 937 215 981 249
rect 1015 215 1059 249
rect 1093 215 1137 249
rect 1171 215 1197 249
rect 875 205 1197 215
rect 475 177 505 192
rect 579 177 609 192
rect 673 177 703 192
rect 767 177 797 192
rect 875 177 905 205
rect 969 177 999 205
rect 1063 177 1093 205
rect 1167 177 1197 205
rect 79 21 109 47
rect 194 21 224 47
rect 475 21 505 47
rect 579 21 609 47
rect 673 21 703 47
rect 767 21 797 47
rect 875 21 905 47
rect 969 21 999 47
rect 1063 21 1093 47
rect 1167 21 1197 47
<< polycont >>
rect 98 215 132 249
rect 216 215 250 249
rect 772 215 806 249
rect 903 215 937 249
rect 981 215 1015 249
rect 1059 215 1093 249
rect 1137 215 1171 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 17 477 69 493
rect 17 443 35 477
rect 17 409 69 443
rect 17 375 35 409
rect 17 353 69 375
rect 103 489 196 527
rect 103 455 137 489
rect 171 455 196 489
rect 103 421 196 455
rect 103 387 137 421
rect 171 387 196 421
rect 103 369 196 387
rect 240 477 291 493
rect 240 443 244 477
rect 278 443 291 477
rect 240 409 291 443
rect 240 375 244 409
rect 278 375 291 409
rect 333 477 382 493
rect 333 443 348 477
rect 416 489 492 527
rect 416 455 442 489
rect 476 455 492 489
rect 536 477 570 493
rect 333 421 382 443
rect 614 489 680 527
rect 614 455 630 489
rect 664 455 680 489
rect 724 489 1257 493
rect 724 455 742 489
rect 776 455 820 489
rect 854 455 1019 489
rect 1053 455 1207 489
rect 1241 455 1257 489
rect 536 421 570 443
rect 724 421 1257 455
rect 333 387 742 421
rect 776 387 820 421
rect 854 387 1019 421
rect 1053 387 1207 421
rect 1241 387 1257 421
rect 399 379 1257 387
rect 240 353 291 375
rect 17 255 64 353
rect 17 221 30 255
rect 17 133 64 221
rect 98 249 166 335
rect 240 319 365 353
rect 132 215 166 249
rect 98 153 166 215
rect 200 249 276 285
rect 200 215 216 249
rect 250 215 276 249
rect 200 153 276 215
rect 310 255 365 319
rect 399 311 925 345
rect 959 311 1113 345
rect 1147 311 1267 345
rect 399 289 1267 311
rect 310 249 832 255
rect 310 215 772 249
rect 806 215 832 249
rect 310 205 832 215
rect 866 249 942 255
rect 866 215 903 249
rect 937 221 942 249
rect 976 249 1187 255
rect 976 221 981 249
rect 937 215 981 221
rect 1015 215 1059 249
rect 1093 215 1137 249
rect 1171 215 1187 249
rect 866 205 1187 215
rect 17 106 69 133
rect 310 119 365 205
rect 1221 171 1267 289
rect 17 72 35 106
rect 17 56 69 72
rect 103 89 196 119
rect 103 55 129 89
rect 163 55 196 89
rect 103 17 196 55
rect 240 103 365 119
rect 240 69 244 103
rect 278 69 365 103
rect 240 51 365 69
rect 399 131 865 171
rect 399 129 465 131
rect 399 95 421 129
rect 455 95 465 129
rect 619 129 653 131
rect 399 51 465 95
rect 499 89 575 97
rect 499 55 525 89
rect 559 55 575 89
rect 807 129 865 131
rect 619 55 653 95
rect 687 89 763 97
rect 687 55 713 89
rect 747 55 763 89
rect 499 17 575 55
rect 687 17 763 55
rect 807 95 819 129
rect 853 95 865 129
rect 899 169 1267 171
rect 899 135 925 169
rect 959 135 1113 169
rect 1147 135 1267 169
rect 899 123 1267 135
rect 807 89 865 95
rect 807 55 1019 89
rect 1053 55 1207 89
rect 1241 55 1257 89
rect 807 51 1257 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 30 221 64 255
rect 942 221 976 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 17 255 988 261
rect 17 221 30 255
rect 64 233 942 255
rect 64 221 76 233
rect 17 215 76 221
rect 930 221 942 233
rect 976 221 988 255
rect 930 215 988 221
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 122 153 156 187 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 840 289 874 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 738 289 772 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 636 289 670 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 534 289 568 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 432 289 466 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1225 153 1259 187 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1146 289 1180 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1044 289 1078 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 215 153 249 187 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 122 289 156 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1223 289 1257 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ebufn_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1525902
string GDS_START 1516168
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
