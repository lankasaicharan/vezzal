magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 59 252 637 290
rect 59 49 857 252
rect 0 0 864 49
<< scpmos >>
rect 132 392 168 592
rect 230 392 266 592
rect 320 392 356 592
rect 398 392 434 592
rect 476 392 512 592
rect 742 368 778 592
<< nmoslvt >>
rect 138 136 168 264
rect 210 136 240 264
rect 318 136 348 264
rect 404 136 434 264
rect 528 136 558 264
rect 748 78 778 226
<< ndiff >>
rect 85 235 138 264
rect 85 201 93 235
rect 127 201 138 235
rect 85 136 138 201
rect 168 136 210 264
rect 240 182 318 264
rect 240 148 251 182
rect 285 148 318 182
rect 240 136 318 148
rect 348 234 404 264
rect 348 200 359 234
rect 393 200 404 234
rect 348 136 404 200
rect 434 182 528 264
rect 434 148 483 182
rect 517 148 528 182
rect 434 136 528 148
rect 558 250 611 264
rect 558 216 569 250
rect 603 216 611 250
rect 558 182 611 216
rect 558 148 569 182
rect 603 148 611 182
rect 558 136 611 148
rect 695 214 748 226
rect 695 180 703 214
rect 737 180 748 214
rect 695 124 748 180
rect 695 90 703 124
rect 737 90 748 124
rect 695 78 748 90
rect 778 214 831 226
rect 778 180 789 214
rect 823 180 831 214
rect 778 124 831 180
rect 778 90 789 124
rect 823 90 831 124
rect 778 78 831 90
<< pdiff >>
rect 80 580 132 592
rect 80 546 88 580
rect 122 546 132 580
rect 80 509 132 546
rect 80 475 88 509
rect 122 475 132 509
rect 80 438 132 475
rect 80 404 88 438
rect 122 404 132 438
rect 80 392 132 404
rect 168 580 230 592
rect 168 546 182 580
rect 216 546 230 580
rect 168 512 230 546
rect 168 478 182 512
rect 216 478 230 512
rect 168 392 230 478
rect 266 580 320 592
rect 266 546 276 580
rect 310 546 320 580
rect 266 512 320 546
rect 266 478 276 512
rect 310 478 320 512
rect 266 444 320 478
rect 266 410 276 444
rect 310 410 320 444
rect 266 392 320 410
rect 356 392 398 592
rect 434 392 476 592
rect 512 580 564 592
rect 512 546 522 580
rect 556 546 564 580
rect 512 512 564 546
rect 512 478 522 512
rect 556 478 564 512
rect 512 444 564 478
rect 512 410 522 444
rect 556 410 564 444
rect 512 392 564 410
rect 690 580 742 592
rect 690 546 698 580
rect 732 546 742 580
rect 690 497 742 546
rect 690 463 698 497
rect 732 463 742 497
rect 690 414 742 463
rect 690 380 698 414
rect 732 380 742 414
rect 690 368 742 380
rect 778 580 830 592
rect 778 546 788 580
rect 822 546 830 580
rect 778 497 830 546
rect 778 463 788 497
rect 822 463 830 497
rect 778 414 830 463
rect 778 380 788 414
rect 822 380 830 414
rect 778 368 830 380
<< ndiffc >>
rect 93 201 127 235
rect 251 148 285 182
rect 359 200 393 234
rect 483 148 517 182
rect 569 216 603 250
rect 569 148 603 182
rect 703 180 737 214
rect 703 90 737 124
rect 789 180 823 214
rect 789 90 823 124
<< pdiffc >>
rect 88 546 122 580
rect 88 475 122 509
rect 88 404 122 438
rect 182 546 216 580
rect 182 478 216 512
rect 276 546 310 580
rect 276 478 310 512
rect 276 410 310 444
rect 522 546 556 580
rect 522 478 556 512
rect 522 410 556 444
rect 698 546 732 580
rect 698 463 732 497
rect 698 380 732 414
rect 788 546 822 580
rect 788 463 822 497
rect 788 380 822 414
<< poly >>
rect 132 592 168 618
rect 230 592 266 618
rect 320 592 356 618
rect 398 592 434 618
rect 476 592 512 618
rect 742 592 778 618
rect 132 279 168 392
rect 230 360 266 392
rect 138 264 168 279
rect 210 344 276 360
rect 210 310 226 344
rect 260 310 276 344
rect 210 294 276 310
rect 320 309 356 392
rect 210 264 240 294
rect 318 279 356 309
rect 398 279 434 392
rect 476 360 512 392
rect 476 344 558 360
rect 476 310 505 344
rect 539 310 558 344
rect 742 330 778 368
rect 476 294 558 310
rect 318 264 348 279
rect 404 264 434 279
rect 528 264 558 294
rect 672 314 778 330
rect 672 280 688 314
rect 722 280 778 314
rect 672 264 778 280
rect 748 226 778 264
rect 138 114 168 136
rect 102 98 168 114
rect 210 110 240 136
rect 318 107 348 136
rect 404 107 434 136
rect 528 110 558 136
rect 102 64 118 98
rect 152 64 168 98
rect 102 48 168 64
rect 287 91 353 107
rect 287 57 303 91
rect 337 57 353 91
rect 287 41 353 57
rect 401 91 467 107
rect 401 57 417 91
rect 451 57 467 91
rect 401 41 467 57
rect 748 52 778 78
<< polycont >>
rect 226 310 260 344
rect 505 310 539 344
rect 688 280 722 314
rect 118 64 152 98
rect 303 57 337 91
rect 417 57 451 91
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 72 580 138 596
rect 72 546 88 580
rect 122 546 138 580
rect 72 509 138 546
rect 72 475 88 509
rect 122 475 138 509
rect 72 438 138 475
rect 178 580 220 649
rect 178 546 182 580
rect 216 546 220 580
rect 178 512 220 546
rect 178 478 182 512
rect 216 478 220 512
rect 178 462 220 478
rect 260 580 326 596
rect 260 546 276 580
rect 310 546 326 580
rect 260 512 326 546
rect 260 478 276 512
rect 310 478 326 512
rect 72 404 88 438
rect 122 428 138 438
rect 260 444 326 478
rect 260 428 276 444
rect 122 410 276 428
rect 310 410 326 444
rect 122 404 326 410
rect 72 394 326 404
rect 506 580 572 596
rect 506 546 522 580
rect 556 546 572 580
rect 506 512 572 546
rect 506 478 522 512
rect 556 478 572 512
rect 506 444 572 478
rect 506 410 522 444
rect 556 428 572 444
rect 682 580 732 649
rect 682 546 698 580
rect 682 497 732 546
rect 682 463 698 497
rect 556 410 623 428
rect 506 394 623 410
rect 72 388 138 394
rect 210 344 455 360
rect 210 310 226 344
rect 260 310 455 344
rect 210 300 455 310
rect 489 344 555 360
rect 489 310 505 344
rect 539 310 555 344
rect 489 300 555 310
rect 589 330 623 394
rect 682 414 732 463
rect 682 380 698 414
rect 682 364 732 380
rect 772 580 839 596
rect 772 546 788 580
rect 822 546 839 580
rect 772 497 839 546
rect 772 463 788 497
rect 822 463 839 497
rect 772 414 839 463
rect 772 380 788 414
rect 822 380 839 414
rect 589 314 738 330
rect 589 280 688 314
rect 722 280 738 314
rect 77 266 143 268
rect 589 266 738 280
rect 77 264 738 266
rect 77 250 623 264
rect 77 235 569 250
rect 77 201 93 235
rect 127 234 569 235
rect 127 232 359 234
rect 127 201 143 232
rect 77 168 143 201
rect 343 200 359 232
rect 393 232 569 234
rect 393 200 409 232
rect 219 182 285 198
rect 219 148 251 182
rect 343 168 409 200
rect 603 216 623 250
rect 483 182 535 198
rect 25 98 168 134
rect 25 88 118 98
rect 102 64 118 88
rect 152 64 168 98
rect 102 51 168 64
rect 219 132 285 148
rect 517 148 535 182
rect 219 17 253 132
rect 319 98 359 134
rect 287 91 359 98
rect 287 57 303 91
rect 337 57 359 91
rect 287 51 359 57
rect 401 98 449 134
rect 483 132 535 148
rect 569 182 623 216
rect 603 148 623 182
rect 569 132 623 148
rect 687 214 737 230
rect 687 180 703 214
rect 401 91 467 98
rect 401 57 417 91
rect 451 57 467 91
rect 401 51 467 57
rect 501 17 535 132
rect 687 124 737 180
rect 687 90 703 124
rect 687 17 737 90
rect 772 214 839 380
rect 772 180 789 214
rect 823 180 839 214
rect 772 124 839 180
rect 772 90 789 124
rect 823 90 839 124
rect 772 74 839 90
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2111o_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 51324
string GDS_START 42588
<< end >>
