magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 32 49 881 243
rect 0 0 960 49
<< scnmos >>
rect 111 49 141 217
rect 197 49 227 217
rect 313 49 343 217
rect 399 49 429 217
rect 514 49 544 217
rect 600 49 630 217
rect 686 49 716 217
rect 772 49 802 217
<< scpmoshvt >>
rect 111 367 141 619
rect 183 367 213 619
rect 291 367 321 619
rect 399 367 429 619
rect 514 367 544 619
rect 600 367 630 619
rect 686 367 716 619
rect 772 367 802 619
<< ndiff >>
rect 58 203 111 217
rect 58 169 66 203
rect 100 169 111 203
rect 58 95 111 169
rect 58 61 66 95
rect 100 61 111 95
rect 58 49 111 61
rect 141 205 197 217
rect 141 171 152 205
rect 186 171 197 205
rect 141 101 197 171
rect 141 67 152 101
rect 186 67 197 101
rect 141 49 197 67
rect 227 165 313 217
rect 227 131 254 165
rect 288 131 313 165
rect 227 91 313 131
rect 227 57 254 91
rect 288 57 313 91
rect 227 49 313 57
rect 343 205 399 217
rect 343 171 354 205
rect 388 171 399 205
rect 343 91 399 171
rect 343 57 354 91
rect 388 57 399 91
rect 343 49 399 57
rect 429 165 514 217
rect 429 131 454 165
rect 488 131 514 165
rect 429 91 514 131
rect 429 57 454 91
rect 488 57 514 91
rect 429 49 514 57
rect 544 205 600 217
rect 544 171 555 205
rect 589 171 600 205
rect 544 101 600 171
rect 544 67 555 101
rect 589 67 600 101
rect 544 49 600 67
rect 630 183 686 217
rect 630 149 641 183
rect 675 149 686 183
rect 630 95 686 149
rect 630 61 641 95
rect 675 61 686 95
rect 630 49 686 61
rect 716 205 772 217
rect 716 171 727 205
rect 761 171 772 205
rect 716 101 772 171
rect 716 67 727 101
rect 761 67 772 101
rect 716 49 772 67
rect 802 167 855 217
rect 802 133 813 167
rect 847 133 855 167
rect 802 95 855 133
rect 802 61 813 95
rect 847 61 855 95
rect 802 49 855 61
<< pdiff >>
rect 58 607 111 619
rect 58 573 66 607
rect 100 573 111 607
rect 58 518 111 573
rect 58 484 66 518
rect 100 484 111 518
rect 58 424 111 484
rect 58 390 66 424
rect 100 390 111 424
rect 58 367 111 390
rect 141 367 183 619
rect 213 367 291 619
rect 321 367 399 619
rect 429 607 514 619
rect 429 573 453 607
rect 487 573 514 607
rect 429 496 514 573
rect 429 462 453 496
rect 487 462 514 496
rect 429 367 514 462
rect 544 599 600 619
rect 544 565 555 599
rect 589 565 600 599
rect 544 504 600 565
rect 544 470 555 504
rect 589 470 600 504
rect 544 413 600 470
rect 544 379 555 413
rect 589 379 600 413
rect 544 367 600 379
rect 630 611 686 619
rect 630 577 641 611
rect 675 577 686 611
rect 630 534 686 577
rect 630 500 641 534
rect 675 500 686 534
rect 630 455 686 500
rect 630 421 641 455
rect 675 421 686 455
rect 630 367 686 421
rect 716 599 772 619
rect 716 565 727 599
rect 761 565 772 599
rect 716 504 772 565
rect 716 470 727 504
rect 761 470 772 504
rect 716 413 772 470
rect 716 379 727 413
rect 761 379 772 413
rect 716 367 772 379
rect 802 607 855 619
rect 802 573 813 607
rect 847 573 855 607
rect 802 534 855 573
rect 802 500 813 534
rect 847 500 855 534
rect 802 455 855 500
rect 802 421 813 455
rect 847 421 855 455
rect 802 367 855 421
<< ndiffc >>
rect 66 169 100 203
rect 66 61 100 95
rect 152 171 186 205
rect 152 67 186 101
rect 254 131 288 165
rect 254 57 288 91
rect 354 171 388 205
rect 354 57 388 91
rect 454 131 488 165
rect 454 57 488 91
rect 555 171 589 205
rect 555 67 589 101
rect 641 149 675 183
rect 641 61 675 95
rect 727 171 761 205
rect 727 67 761 101
rect 813 133 847 167
rect 813 61 847 95
<< pdiffc >>
rect 66 573 100 607
rect 66 484 100 518
rect 66 390 100 424
rect 453 573 487 607
rect 453 462 487 496
rect 555 565 589 599
rect 555 470 589 504
rect 555 379 589 413
rect 641 577 675 611
rect 641 500 675 534
rect 641 421 675 455
rect 727 565 761 599
rect 727 470 761 504
rect 727 379 761 413
rect 813 573 847 607
rect 813 500 847 534
rect 813 421 847 455
<< poly >>
rect 111 619 141 645
rect 183 619 213 645
rect 291 619 321 645
rect 399 619 429 645
rect 514 619 544 645
rect 600 619 630 645
rect 686 619 716 645
rect 772 619 802 645
rect 111 308 141 367
rect 41 292 141 308
rect 41 258 57 292
rect 91 258 141 292
rect 183 335 213 367
rect 291 335 321 367
rect 399 335 429 367
rect 514 335 544 367
rect 600 335 630 367
rect 686 335 716 367
rect 772 335 802 367
rect 183 319 249 335
rect 183 285 199 319
rect 233 285 249 319
rect 183 269 249 285
rect 291 319 357 335
rect 291 285 307 319
rect 341 285 357 319
rect 291 269 357 285
rect 399 319 465 335
rect 399 285 415 319
rect 449 285 465 319
rect 399 269 465 285
rect 514 319 852 335
rect 514 285 530 319
rect 564 285 598 319
rect 632 285 666 319
rect 700 285 734 319
rect 768 285 802 319
rect 836 285 852 319
rect 514 269 852 285
rect 41 242 141 258
rect 111 217 141 242
rect 197 217 227 269
rect 313 217 343 269
rect 399 217 429 269
rect 514 217 544 269
rect 600 217 630 269
rect 686 217 716 269
rect 772 217 802 269
rect 111 23 141 49
rect 197 23 227 49
rect 313 23 343 49
rect 399 23 429 49
rect 514 23 544 49
rect 600 23 630 49
rect 686 23 716 49
rect 772 23 802 49
<< polycont >>
rect 57 258 91 292
rect 199 285 233 319
rect 307 285 341 319
rect 415 285 449 319
rect 530 285 564 319
rect 598 285 632 319
rect 666 285 700 319
rect 734 285 768 319
rect 802 285 836 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 50 607 116 615
rect 50 573 66 607
rect 100 573 116 607
rect 50 518 116 573
rect 50 484 66 518
rect 100 484 116 518
rect 50 424 116 484
rect 437 607 503 649
rect 437 573 453 607
rect 487 573 503 607
rect 437 496 503 573
rect 437 462 453 496
rect 487 462 503 496
rect 437 454 503 462
rect 553 599 591 615
rect 553 565 555 599
rect 589 565 591 599
rect 553 504 591 565
rect 553 470 555 504
rect 589 470 591 504
rect 50 390 66 424
rect 100 420 116 424
rect 100 390 519 420
rect 50 386 519 390
rect 17 292 91 352
rect 17 258 57 292
rect 125 319 265 352
rect 125 285 199 319
rect 233 285 265 319
rect 299 319 366 352
rect 299 285 307 319
rect 341 285 366 319
rect 299 269 366 285
rect 400 319 451 352
rect 400 285 415 319
rect 449 285 451 319
rect 400 269 451 285
rect 485 319 519 386
rect 553 413 591 470
rect 625 611 691 649
rect 625 577 641 611
rect 675 577 691 611
rect 625 534 691 577
rect 625 500 641 534
rect 675 500 691 534
rect 625 455 691 500
rect 625 421 641 455
rect 675 421 691 455
rect 725 599 763 615
rect 725 565 727 599
rect 761 565 763 599
rect 725 504 763 565
rect 725 470 727 504
rect 761 470 763 504
rect 553 379 555 413
rect 589 387 591 413
rect 725 413 763 470
rect 797 607 863 649
rect 797 573 813 607
rect 847 573 863 607
rect 797 534 863 573
rect 797 500 813 534
rect 847 500 863 534
rect 797 455 863 500
rect 797 421 813 455
rect 847 421 863 455
rect 725 387 727 413
rect 589 379 727 387
rect 761 387 763 413
rect 761 379 943 387
rect 553 353 943 379
rect 485 285 530 319
rect 564 285 598 319
rect 632 285 666 319
rect 700 285 734 319
rect 768 285 802 319
rect 836 285 852 319
rect 17 242 91 258
rect 485 233 519 285
rect 886 251 943 353
rect 50 203 116 208
rect 50 169 66 203
rect 100 169 116 203
rect 50 95 116 169
rect 50 61 66 95
rect 100 61 116 95
rect 50 17 116 61
rect 150 205 519 233
rect 150 171 152 205
rect 186 199 354 205
rect 186 171 202 199
rect 150 101 202 171
rect 338 171 354 199
rect 388 199 519 205
rect 553 217 943 251
rect 553 205 591 217
rect 388 171 404 199
rect 150 67 152 101
rect 186 67 202 101
rect 150 51 202 67
rect 238 131 254 165
rect 288 131 304 165
rect 238 91 304 131
rect 238 57 254 91
rect 288 57 304 91
rect 238 17 304 57
rect 338 91 404 171
rect 553 171 555 205
rect 589 171 591 205
rect 725 205 770 217
rect 338 57 354 91
rect 388 57 404 91
rect 338 51 404 57
rect 438 131 454 165
rect 488 131 504 165
rect 438 91 504 131
rect 438 57 454 91
rect 488 57 504 91
rect 438 17 504 57
rect 553 101 591 171
rect 553 67 555 101
rect 589 67 591 101
rect 553 51 591 67
rect 625 149 641 183
rect 675 149 691 183
rect 625 95 691 149
rect 625 61 641 95
rect 675 61 691 95
rect 625 17 691 61
rect 725 171 727 205
rect 761 171 770 205
rect 725 101 770 171
rect 725 67 727 101
rect 761 67 770 101
rect 725 51 770 67
rect 804 167 857 183
rect 804 133 813 167
rect 847 133 857 167
rect 804 95 857 133
rect 804 61 813 95
rect 847 61 857 95
rect 891 94 943 217
rect 804 17 857 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or4_4
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 895 94 929 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 287008
string GDS_START 278552
<< end >>
