magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 6 49 1148 241
rect 0 0 1152 49
<< scnmos >>
rect 85 47 115 215
rect 171 47 201 215
rect 257 47 287 215
rect 343 47 373 215
rect 429 47 459 215
rect 515 47 545 215
rect 601 47 631 215
rect 695 47 725 215
rect 781 47 811 215
rect 867 47 897 215
rect 953 47 983 215
rect 1039 47 1069 215
<< scpmoshvt >>
rect 85 367 115 619
rect 171 367 201 619
rect 257 367 287 619
rect 343 367 373 619
rect 429 367 459 619
rect 515 367 545 619
rect 601 367 631 619
rect 687 367 717 619
rect 781 367 811 619
rect 867 367 897 619
rect 953 367 983 619
rect 1039 367 1069 619
<< ndiff >>
rect 32 192 85 215
rect 32 158 40 192
rect 74 158 85 192
rect 32 101 85 158
rect 32 67 40 101
rect 74 67 85 101
rect 32 47 85 67
rect 115 128 171 215
rect 115 94 126 128
rect 160 94 171 128
rect 115 47 171 94
rect 201 171 257 215
rect 201 137 212 171
rect 246 137 257 171
rect 201 103 257 137
rect 201 69 212 103
rect 246 69 257 103
rect 201 47 257 69
rect 287 105 343 215
rect 287 71 298 105
rect 332 71 343 105
rect 287 47 343 71
rect 373 181 429 215
rect 373 147 384 181
rect 418 147 429 181
rect 373 101 429 147
rect 373 67 384 101
rect 418 67 429 101
rect 373 47 429 67
rect 459 105 515 215
rect 459 71 470 105
rect 504 71 515 105
rect 459 47 515 71
rect 545 181 601 215
rect 545 147 556 181
rect 590 147 601 181
rect 545 101 601 147
rect 545 67 556 101
rect 590 67 601 101
rect 545 47 601 67
rect 631 105 695 215
rect 631 71 642 105
rect 676 71 695 105
rect 631 47 695 71
rect 725 181 781 215
rect 725 147 736 181
rect 770 147 781 181
rect 725 101 781 147
rect 725 67 736 101
rect 770 67 781 101
rect 725 47 781 67
rect 811 190 867 215
rect 811 156 822 190
rect 856 156 867 190
rect 811 47 867 156
rect 897 100 953 215
rect 897 66 908 100
rect 942 66 953 100
rect 897 47 953 66
rect 983 190 1039 215
rect 983 156 994 190
rect 1028 156 1039 190
rect 983 47 1039 156
rect 1069 104 1122 215
rect 1069 70 1080 104
rect 1114 70 1122 104
rect 1069 47 1122 70
<< pdiff >>
rect 32 607 85 619
rect 32 573 40 607
rect 74 573 85 607
rect 32 506 85 573
rect 32 472 40 506
rect 74 472 85 506
rect 32 413 85 472
rect 32 379 40 413
rect 74 379 85 413
rect 32 367 85 379
rect 115 599 171 619
rect 115 565 126 599
rect 160 565 171 599
rect 115 504 171 565
rect 115 470 126 504
rect 160 470 171 504
rect 115 413 171 470
rect 115 379 126 413
rect 160 379 171 413
rect 115 367 171 379
rect 201 607 257 619
rect 201 573 212 607
rect 246 573 257 607
rect 201 532 257 573
rect 201 498 212 532
rect 246 498 257 532
rect 201 453 257 498
rect 201 419 212 453
rect 246 419 257 453
rect 201 367 257 419
rect 287 599 343 619
rect 287 565 298 599
rect 332 565 343 599
rect 287 504 343 565
rect 287 470 298 504
rect 332 470 343 504
rect 287 413 343 470
rect 287 379 298 413
rect 332 379 343 413
rect 287 367 343 379
rect 373 537 429 619
rect 373 503 384 537
rect 418 503 429 537
rect 373 434 429 503
rect 373 400 384 434
rect 418 400 429 434
rect 373 367 429 400
rect 459 599 515 619
rect 459 565 470 599
rect 504 565 515 599
rect 459 504 515 565
rect 459 470 470 504
rect 504 470 515 504
rect 459 367 515 470
rect 545 537 601 619
rect 545 503 556 537
rect 590 503 601 537
rect 545 434 601 503
rect 545 400 556 434
rect 590 400 601 434
rect 545 367 601 400
rect 631 599 687 619
rect 631 565 642 599
rect 676 565 687 599
rect 631 504 687 565
rect 631 470 642 504
rect 676 470 687 504
rect 631 367 687 470
rect 717 607 781 619
rect 717 573 732 607
rect 766 573 781 607
rect 717 497 781 573
rect 717 463 732 497
rect 766 463 781 497
rect 717 367 781 463
rect 811 599 867 619
rect 811 565 822 599
rect 856 565 867 599
rect 811 504 867 565
rect 811 470 822 504
rect 856 470 867 504
rect 811 413 867 470
rect 811 379 822 413
rect 856 379 867 413
rect 811 367 867 379
rect 897 607 953 619
rect 897 573 908 607
rect 942 573 953 607
rect 897 532 953 573
rect 897 498 908 532
rect 942 498 953 532
rect 897 455 953 498
rect 897 421 908 455
rect 942 421 953 455
rect 897 367 953 421
rect 983 599 1039 619
rect 983 565 994 599
rect 1028 565 1039 599
rect 983 504 1039 565
rect 983 470 994 504
rect 1028 470 1039 504
rect 983 413 1039 470
rect 983 379 994 413
rect 1028 379 1039 413
rect 983 367 1039 379
rect 1069 607 1122 619
rect 1069 573 1080 607
rect 1114 573 1122 607
rect 1069 532 1122 573
rect 1069 498 1080 532
rect 1114 498 1122 532
rect 1069 455 1122 498
rect 1069 421 1080 455
rect 1114 421 1122 455
rect 1069 367 1122 421
<< ndiffc >>
rect 40 158 74 192
rect 40 67 74 101
rect 126 94 160 128
rect 212 137 246 171
rect 212 69 246 103
rect 298 71 332 105
rect 384 147 418 181
rect 384 67 418 101
rect 470 71 504 105
rect 556 147 590 181
rect 556 67 590 101
rect 642 71 676 105
rect 736 147 770 181
rect 736 67 770 101
rect 822 156 856 190
rect 908 66 942 100
rect 994 156 1028 190
rect 1080 70 1114 104
<< pdiffc >>
rect 40 573 74 607
rect 40 472 74 506
rect 40 379 74 413
rect 126 565 160 599
rect 126 470 160 504
rect 126 379 160 413
rect 212 573 246 607
rect 212 498 246 532
rect 212 419 246 453
rect 298 565 332 599
rect 298 470 332 504
rect 298 379 332 413
rect 384 503 418 537
rect 384 400 418 434
rect 470 565 504 599
rect 470 470 504 504
rect 556 503 590 537
rect 556 400 590 434
rect 642 565 676 599
rect 642 470 676 504
rect 732 573 766 607
rect 732 463 766 497
rect 822 565 856 599
rect 822 470 856 504
rect 822 379 856 413
rect 908 573 942 607
rect 908 498 942 532
rect 908 421 942 455
rect 994 565 1028 599
rect 994 470 1028 504
rect 994 379 1028 413
rect 1080 573 1114 607
rect 1080 498 1114 532
rect 1080 421 1114 455
<< poly >>
rect 85 619 115 645
rect 171 619 201 645
rect 257 619 287 645
rect 343 619 373 645
rect 429 619 459 645
rect 515 619 545 645
rect 601 619 631 645
rect 687 619 717 645
rect 781 619 811 645
rect 867 619 897 645
rect 953 619 983 645
rect 1039 619 1069 645
rect 85 303 115 367
rect 171 303 201 367
rect 257 303 287 367
rect 343 335 373 367
rect 429 335 459 367
rect 515 335 545 367
rect 601 335 631 367
rect 343 319 631 335
rect 25 287 295 303
rect 25 253 41 287
rect 75 253 109 287
rect 143 253 177 287
rect 211 253 245 287
rect 279 253 295 287
rect 25 237 295 253
rect 343 285 415 319
rect 449 285 501 319
rect 535 285 581 319
rect 615 285 631 319
rect 687 303 717 367
rect 781 303 811 367
rect 867 303 897 367
rect 953 303 983 367
rect 1039 303 1069 367
rect 343 269 631 285
rect 85 215 115 237
rect 171 215 201 237
rect 257 215 287 237
rect 343 215 373 269
rect 429 215 459 269
rect 515 215 545 269
rect 601 215 631 269
rect 673 287 739 303
rect 673 253 689 287
rect 723 253 739 287
rect 673 237 739 253
rect 781 287 1069 303
rect 781 253 797 287
rect 831 253 865 287
rect 899 253 933 287
rect 967 253 1001 287
rect 1035 253 1069 287
rect 781 237 1069 253
rect 695 215 725 237
rect 781 215 811 237
rect 867 215 897 237
rect 953 215 983 237
rect 1039 215 1069 237
rect 85 21 115 47
rect 171 21 201 47
rect 257 21 287 47
rect 343 21 373 47
rect 429 21 459 47
rect 515 21 545 47
rect 601 21 631 47
rect 695 21 725 47
rect 781 21 811 47
rect 867 21 897 47
rect 953 21 983 47
rect 1039 21 1069 47
<< polycont >>
rect 41 253 75 287
rect 109 253 143 287
rect 177 253 211 287
rect 245 253 279 287
rect 415 285 449 319
rect 501 285 535 319
rect 581 285 615 319
rect 689 253 723 287
rect 797 253 831 287
rect 865 253 899 287
rect 933 253 967 287
rect 1001 253 1035 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 24 607 81 649
rect 24 573 40 607
rect 74 573 81 607
rect 24 506 81 573
rect 24 472 40 506
rect 74 472 81 506
rect 24 413 81 472
rect 24 379 40 413
rect 74 379 81 413
rect 24 363 81 379
rect 115 599 162 615
rect 115 565 126 599
rect 160 565 162 599
rect 115 504 162 565
rect 115 470 126 504
rect 160 470 162 504
rect 115 413 162 470
rect 196 607 262 649
rect 196 573 212 607
rect 246 573 262 607
rect 196 532 262 573
rect 196 498 212 532
rect 246 498 262 532
rect 196 453 262 498
rect 196 419 212 453
rect 246 419 262 453
rect 296 599 682 615
rect 296 565 298 599
rect 332 581 470 599
rect 332 565 334 581
rect 296 504 334 565
rect 468 565 470 581
rect 504 581 642 599
rect 504 565 506 581
rect 296 470 298 504
rect 332 470 334 504
rect 115 379 126 413
rect 160 385 162 413
rect 296 413 334 470
rect 296 385 298 413
rect 160 379 298 385
rect 332 379 334 413
rect 368 537 434 547
rect 368 503 384 537
rect 418 503 434 537
rect 368 434 434 503
rect 468 504 506 565
rect 640 565 642 581
rect 676 565 682 599
rect 468 470 470 504
rect 504 470 506 504
rect 468 454 506 470
rect 540 537 606 547
rect 540 503 556 537
rect 590 503 606 537
rect 368 400 384 434
rect 418 420 434 434
rect 540 434 606 503
rect 640 504 682 565
rect 640 470 642 504
rect 676 470 682 504
rect 640 454 682 470
rect 716 607 782 649
rect 716 573 732 607
rect 766 573 782 607
rect 716 497 782 573
rect 716 463 732 497
rect 766 463 782 497
rect 716 454 782 463
rect 816 599 858 615
rect 816 565 822 599
rect 856 565 858 599
rect 816 504 858 565
rect 816 470 822 504
rect 856 470 858 504
rect 540 420 556 434
rect 418 400 556 420
rect 590 420 606 434
rect 816 420 858 470
rect 590 413 858 420
rect 892 607 958 649
rect 892 573 908 607
rect 942 573 958 607
rect 892 532 958 573
rect 892 498 908 532
rect 942 498 958 532
rect 892 455 958 498
rect 892 421 908 455
rect 942 421 958 455
rect 892 419 958 421
rect 992 599 1030 615
rect 992 565 994 599
rect 1028 565 1030 599
rect 992 504 1030 565
rect 992 470 994 504
rect 1028 470 1030 504
rect 590 400 822 413
rect 368 386 822 400
rect 115 351 334 379
rect 689 379 822 386
rect 856 385 858 413
rect 992 413 1030 470
rect 1064 607 1130 649
rect 1064 573 1080 607
rect 1114 573 1130 607
rect 1064 532 1130 573
rect 1064 498 1080 532
rect 1114 498 1130 532
rect 1064 455 1130 498
rect 1064 421 1080 455
rect 1114 421 1130 455
rect 992 385 994 413
rect 856 379 994 385
rect 1028 385 1030 413
rect 1028 379 1134 385
rect 399 319 655 352
rect 689 351 1134 379
rect 773 321 1134 351
rect 25 287 365 303
rect 25 253 41 287
rect 75 253 109 287
rect 143 253 177 287
rect 211 253 245 287
rect 279 253 365 287
rect 399 285 415 319
rect 449 285 501 319
rect 535 285 581 319
rect 615 285 655 319
rect 689 287 739 303
rect 25 249 365 253
rect 723 253 739 287
rect 689 249 739 253
rect 25 242 739 249
rect 781 253 797 287
rect 831 253 865 287
rect 899 253 933 287
rect 967 253 1001 287
rect 1035 253 1051 287
rect 781 242 1051 253
rect 284 215 739 242
rect 24 192 250 208
rect 1085 206 1134 321
rect 24 158 40 192
rect 74 181 250 192
rect 820 190 1134 206
rect 74 174 384 181
rect 74 158 76 174
rect 24 101 76 158
rect 210 171 384 174
rect 24 67 40 101
rect 74 67 76 101
rect 24 51 76 67
rect 110 128 176 140
rect 110 94 126 128
rect 160 94 176 128
rect 110 17 176 94
rect 210 137 212 171
rect 246 147 384 171
rect 418 147 556 181
rect 590 147 736 181
rect 770 147 786 181
rect 246 137 248 147
rect 210 103 248 137
rect 210 69 212 103
rect 246 69 248 103
rect 210 51 248 69
rect 282 105 348 113
rect 282 71 298 105
rect 332 71 348 105
rect 282 17 348 71
rect 382 101 420 147
rect 382 67 384 101
rect 418 67 420 101
rect 382 51 420 67
rect 454 105 520 113
rect 454 71 470 105
rect 504 71 520 105
rect 454 17 520 71
rect 554 101 592 147
rect 554 67 556 101
rect 590 67 592 101
rect 554 51 592 67
rect 626 105 692 113
rect 626 71 642 105
rect 676 71 692 105
rect 626 17 692 71
rect 726 106 786 147
rect 820 156 822 190
rect 856 156 994 190
rect 1028 156 1134 190
rect 820 140 1134 156
rect 726 104 1130 106
rect 726 101 1080 104
rect 726 67 736 101
rect 770 100 1080 101
rect 770 67 908 100
rect 726 66 908 67
rect 942 70 1080 100
rect 1114 70 1130 104
rect 942 66 1130 70
rect 726 51 1130 66
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o21ai_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4664720
string GDS_START 4654152
<< end >>
