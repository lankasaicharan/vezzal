magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 3026 1975
<< nwell >>
rect -38 332 1766 704
<< pwell >>
rect 170 49 1678 248
rect 0 0 1728 49
<< scpmos >>
rect 84 392 114 592
rect 174 392 204 592
rect 264 392 294 592
rect 354 392 384 592
rect 594 368 624 592
rect 684 368 714 592
rect 774 368 804 592
rect 864 368 894 592
rect 954 368 984 592
rect 1044 368 1074 592
rect 1134 368 1164 592
rect 1224 368 1254 592
rect 1314 368 1344 592
rect 1404 368 1434 592
rect 1494 368 1524 592
rect 1584 368 1614 592
<< nmoslvt >>
rect 249 74 279 222
rect 335 74 365 222
rect 429 74 459 222
rect 515 74 545 222
rect 601 74 631 222
rect 687 74 717 222
rect 967 74 997 222
rect 1053 74 1083 222
rect 1139 74 1169 222
rect 1225 74 1255 222
rect 1311 74 1341 222
rect 1397 74 1427 222
rect 1483 74 1513 222
rect 1569 74 1599 222
<< ndiff >>
rect 196 190 249 222
rect 196 156 204 190
rect 238 156 249 190
rect 196 122 249 156
rect 196 88 204 122
rect 238 88 249 122
rect 196 74 249 88
rect 279 210 335 222
rect 279 176 290 210
rect 324 176 335 210
rect 279 120 335 176
rect 279 86 290 120
rect 324 86 335 120
rect 279 74 335 86
rect 365 161 429 222
rect 365 127 380 161
rect 414 127 429 161
rect 365 74 429 127
rect 459 192 515 222
rect 459 158 470 192
rect 504 158 515 192
rect 459 120 515 158
rect 459 86 470 120
rect 504 86 515 120
rect 459 74 515 86
rect 545 122 601 222
rect 545 88 556 122
rect 590 88 601 122
rect 545 74 601 88
rect 631 192 687 222
rect 631 158 642 192
rect 676 158 687 192
rect 631 120 687 158
rect 631 86 642 120
rect 676 86 687 120
rect 631 74 687 86
rect 717 122 774 222
rect 717 88 728 122
rect 762 88 774 122
rect 717 74 774 88
rect 914 120 967 222
rect 914 86 922 120
rect 956 86 967 120
rect 914 74 967 86
rect 997 207 1053 222
rect 997 173 1008 207
rect 1042 173 1053 207
rect 997 74 1053 173
rect 1083 120 1139 222
rect 1083 86 1094 120
rect 1128 86 1139 120
rect 1083 74 1139 86
rect 1169 207 1225 222
rect 1169 173 1180 207
rect 1214 173 1225 207
rect 1169 74 1225 173
rect 1255 210 1311 222
rect 1255 176 1266 210
rect 1300 176 1311 210
rect 1255 120 1311 176
rect 1255 86 1266 120
rect 1300 86 1311 120
rect 1255 74 1311 86
rect 1341 152 1397 222
rect 1341 118 1352 152
rect 1386 118 1397 152
rect 1341 74 1397 118
rect 1427 210 1483 222
rect 1427 176 1438 210
rect 1472 176 1483 210
rect 1427 120 1483 176
rect 1427 86 1438 120
rect 1472 86 1483 120
rect 1427 74 1483 86
rect 1513 152 1569 222
rect 1513 118 1524 152
rect 1558 118 1569 152
rect 1513 74 1569 118
rect 1599 210 1652 222
rect 1599 176 1610 210
rect 1644 176 1652 210
rect 1599 120 1652 176
rect 1599 86 1610 120
rect 1644 86 1652 120
rect 1599 74 1652 86
<< pdiff >>
rect 29 580 84 592
rect 29 546 37 580
rect 71 546 84 580
rect 29 509 84 546
rect 29 475 37 509
rect 71 475 84 509
rect 29 438 84 475
rect 29 404 37 438
rect 71 404 84 438
rect 29 392 84 404
rect 114 531 174 592
rect 114 497 127 531
rect 161 497 174 531
rect 114 438 174 497
rect 114 404 127 438
rect 161 404 174 438
rect 114 392 174 404
rect 204 580 264 592
rect 204 546 217 580
rect 251 546 264 580
rect 204 509 264 546
rect 204 475 217 509
rect 251 475 264 509
rect 204 438 264 475
rect 204 404 217 438
rect 251 404 264 438
rect 204 392 264 404
rect 294 580 354 592
rect 294 546 307 580
rect 341 546 354 580
rect 294 512 354 546
rect 294 478 307 512
rect 341 478 354 512
rect 294 392 354 478
rect 384 580 439 592
rect 384 546 397 580
rect 431 546 439 580
rect 384 512 439 546
rect 384 478 397 512
rect 431 478 439 512
rect 384 444 439 478
rect 384 410 397 444
rect 431 410 439 444
rect 384 392 439 410
rect 539 580 594 592
rect 539 546 547 580
rect 581 546 594 580
rect 539 497 594 546
rect 539 463 547 497
rect 581 463 594 497
rect 539 414 594 463
rect 539 380 547 414
rect 581 380 594 414
rect 539 368 594 380
rect 624 531 684 592
rect 624 497 637 531
rect 671 497 684 531
rect 624 414 684 497
rect 624 380 637 414
rect 671 380 684 414
rect 624 368 684 380
rect 714 580 774 592
rect 714 546 727 580
rect 761 546 774 580
rect 714 462 774 546
rect 714 428 727 462
rect 761 428 774 462
rect 714 368 774 428
rect 804 531 864 592
rect 804 497 817 531
rect 851 497 864 531
rect 804 414 864 497
rect 804 380 817 414
rect 851 380 864 414
rect 804 368 864 380
rect 894 580 954 592
rect 894 546 907 580
rect 941 546 954 580
rect 894 510 954 546
rect 894 476 907 510
rect 941 476 954 510
rect 894 440 954 476
rect 894 406 907 440
rect 941 406 954 440
rect 894 368 954 406
rect 984 580 1044 592
rect 984 546 997 580
rect 1031 546 1044 580
rect 984 508 1044 546
rect 984 474 997 508
rect 1031 474 1044 508
rect 984 368 1044 474
rect 1074 580 1134 592
rect 1074 546 1087 580
rect 1121 546 1134 580
rect 1074 510 1134 546
rect 1074 476 1087 510
rect 1121 476 1134 510
rect 1074 440 1134 476
rect 1074 406 1087 440
rect 1121 406 1134 440
rect 1074 368 1134 406
rect 1164 580 1224 592
rect 1164 546 1177 580
rect 1211 546 1224 580
rect 1164 508 1224 546
rect 1164 474 1177 508
rect 1211 474 1224 508
rect 1164 368 1224 474
rect 1254 580 1314 592
rect 1254 546 1267 580
rect 1301 546 1314 580
rect 1254 497 1314 546
rect 1254 463 1267 497
rect 1301 463 1314 497
rect 1254 414 1314 463
rect 1254 380 1267 414
rect 1301 380 1314 414
rect 1254 368 1314 380
rect 1344 580 1404 592
rect 1344 546 1357 580
rect 1391 546 1404 580
rect 1344 508 1404 546
rect 1344 474 1357 508
rect 1391 474 1404 508
rect 1344 368 1404 474
rect 1434 580 1494 592
rect 1434 546 1447 580
rect 1481 546 1494 580
rect 1434 510 1494 546
rect 1434 476 1447 510
rect 1481 476 1494 510
rect 1434 440 1494 476
rect 1434 406 1447 440
rect 1481 406 1494 440
rect 1434 368 1494 406
rect 1524 580 1584 592
rect 1524 546 1537 580
rect 1571 546 1584 580
rect 1524 508 1584 546
rect 1524 474 1537 508
rect 1571 474 1584 508
rect 1524 368 1584 474
rect 1614 580 1669 592
rect 1614 546 1627 580
rect 1661 546 1669 580
rect 1614 510 1669 546
rect 1614 476 1627 510
rect 1661 476 1669 510
rect 1614 440 1669 476
rect 1614 406 1627 440
rect 1661 406 1669 440
rect 1614 368 1669 406
<< ndiffc >>
rect 204 156 238 190
rect 204 88 238 122
rect 290 176 324 210
rect 290 86 324 120
rect 380 127 414 161
rect 470 158 504 192
rect 470 86 504 120
rect 556 88 590 122
rect 642 158 676 192
rect 642 86 676 120
rect 728 88 762 122
rect 922 86 956 120
rect 1008 173 1042 207
rect 1094 86 1128 120
rect 1180 173 1214 207
rect 1266 176 1300 210
rect 1266 86 1300 120
rect 1352 118 1386 152
rect 1438 176 1472 210
rect 1438 86 1472 120
rect 1524 118 1558 152
rect 1610 176 1644 210
rect 1610 86 1644 120
<< pdiffc >>
rect 37 546 71 580
rect 37 475 71 509
rect 37 404 71 438
rect 127 497 161 531
rect 127 404 161 438
rect 217 546 251 580
rect 217 475 251 509
rect 217 404 251 438
rect 307 546 341 580
rect 307 478 341 512
rect 397 546 431 580
rect 397 478 431 512
rect 397 410 431 444
rect 547 546 581 580
rect 547 463 581 497
rect 547 380 581 414
rect 637 497 671 531
rect 637 380 671 414
rect 727 546 761 580
rect 727 428 761 462
rect 817 497 851 531
rect 817 380 851 414
rect 907 546 941 580
rect 907 476 941 510
rect 907 406 941 440
rect 997 546 1031 580
rect 997 474 1031 508
rect 1087 546 1121 580
rect 1087 476 1121 510
rect 1087 406 1121 440
rect 1177 546 1211 580
rect 1177 474 1211 508
rect 1267 546 1301 580
rect 1267 463 1301 497
rect 1267 380 1301 414
rect 1357 546 1391 580
rect 1357 474 1391 508
rect 1447 546 1481 580
rect 1447 476 1481 510
rect 1447 406 1481 440
rect 1537 546 1571 580
rect 1537 474 1571 508
rect 1627 546 1661 580
rect 1627 476 1661 510
rect 1627 406 1661 440
<< poly >>
rect 84 592 114 618
rect 174 592 204 618
rect 264 592 294 618
rect 354 592 384 618
rect 594 592 624 618
rect 684 592 714 618
rect 774 592 804 618
rect 864 592 894 618
rect 954 592 984 618
rect 1044 592 1074 618
rect 1134 592 1164 618
rect 1224 592 1254 618
rect 1314 592 1344 618
rect 1404 592 1434 618
rect 1494 592 1524 618
rect 1584 592 1614 618
rect 84 377 114 392
rect 174 377 204 392
rect 264 377 294 392
rect 354 377 384 392
rect 81 354 117 377
rect 171 354 207 377
rect 25 338 207 354
rect 25 304 41 338
rect 75 304 207 338
rect 261 360 297 377
rect 351 360 387 377
rect 261 344 387 360
rect 594 353 624 368
rect 684 353 714 368
rect 774 353 804 368
rect 864 353 894 368
rect 954 353 984 368
rect 1044 353 1074 368
rect 1134 353 1164 368
rect 1224 353 1254 368
rect 1314 353 1344 368
rect 1404 353 1434 368
rect 1494 353 1524 368
rect 1584 353 1614 368
rect 261 330 337 344
rect 25 270 207 304
rect 321 310 337 330
rect 371 310 387 344
rect 591 310 627 353
rect 681 310 717 353
rect 771 310 807 353
rect 861 310 897 353
rect 321 294 387 310
rect 515 294 897 310
rect 25 236 41 270
rect 75 267 207 270
rect 75 258 279 267
rect 75 236 111 258
rect 177 237 279 258
rect 25 202 111 236
rect 249 222 279 237
rect 335 222 365 294
rect 515 274 531 294
rect 429 260 531 274
rect 565 260 599 294
rect 633 260 667 294
rect 701 280 897 294
rect 951 336 987 353
rect 1041 336 1077 353
rect 1131 336 1167 353
rect 1221 336 1257 353
rect 951 320 1257 336
rect 951 286 967 320
rect 1001 286 1035 320
rect 1069 286 1103 320
rect 1137 286 1171 320
rect 1205 286 1257 320
rect 701 260 717 280
rect 951 270 1257 286
rect 1311 336 1347 353
rect 1401 336 1437 353
rect 1491 336 1527 353
rect 1581 336 1617 353
rect 1311 320 1617 336
rect 1311 286 1363 320
rect 1397 286 1431 320
rect 1465 286 1499 320
rect 1533 286 1567 320
rect 1601 286 1617 320
rect 1311 270 1617 286
rect 429 244 717 260
rect 429 222 459 244
rect 515 222 545 244
rect 601 222 631 244
rect 687 222 717 244
rect 967 222 997 270
rect 1053 222 1083 270
rect 1139 222 1169 270
rect 1225 222 1255 270
rect 1311 222 1341 270
rect 1397 222 1427 270
rect 1483 222 1513 270
rect 1569 222 1599 270
rect 25 168 41 202
rect 75 168 111 202
rect 25 134 111 168
rect 25 100 41 134
rect 75 100 111 134
rect 25 84 111 100
rect 249 48 279 74
rect 335 48 365 74
rect 429 48 459 74
rect 515 48 545 74
rect 601 48 631 74
rect 687 48 717 74
rect 967 48 997 74
rect 1053 48 1083 74
rect 1139 48 1169 74
rect 1225 48 1255 74
rect 1311 48 1341 74
rect 1397 48 1427 74
rect 1483 48 1513 74
rect 1569 48 1599 74
<< polycont >>
rect 41 304 75 338
rect 337 310 371 344
rect 41 236 75 270
rect 531 260 565 294
rect 599 260 633 294
rect 667 260 701 294
rect 967 286 1001 320
rect 1035 286 1069 320
rect 1103 286 1137 320
rect 1171 286 1205 320
rect 1363 286 1397 320
rect 1431 286 1465 320
rect 1499 286 1533 320
rect 1567 286 1601 320
rect 41 168 75 202
rect 41 100 75 134
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 21 581 251 615
rect 21 580 87 581
rect 21 546 37 580
rect 71 546 87 580
rect 217 580 251 581
rect 21 509 87 546
rect 21 475 37 509
rect 71 475 87 509
rect 21 438 87 475
rect 21 404 37 438
rect 71 404 87 438
rect 21 388 87 404
rect 127 531 177 547
rect 161 497 177 531
rect 127 438 177 497
rect 161 404 177 438
rect 25 338 91 354
rect 25 304 41 338
rect 75 304 91 338
rect 25 270 91 304
rect 25 236 41 270
rect 75 236 91 270
rect 25 202 91 236
rect 127 260 177 404
rect 217 509 251 546
rect 217 438 251 475
rect 291 580 341 649
rect 291 546 307 580
rect 291 512 341 546
rect 291 478 307 512
rect 291 462 341 478
rect 381 580 447 596
rect 381 546 397 580
rect 431 546 447 580
rect 381 512 447 546
rect 381 478 397 512
rect 431 478 447 512
rect 381 444 447 478
rect 381 428 397 444
rect 251 410 397 428
rect 431 410 447 444
rect 251 404 447 410
rect 217 394 447 404
rect 531 581 957 615
rect 531 580 597 581
rect 531 546 547 580
rect 581 546 597 580
rect 711 580 777 581
rect 531 497 597 546
rect 531 463 547 497
rect 581 463 597 497
rect 531 414 597 463
rect 217 388 251 394
rect 531 380 547 414
rect 581 380 597 414
rect 531 364 597 380
rect 637 531 671 547
rect 637 414 671 497
rect 711 546 727 580
rect 761 546 777 580
rect 891 580 957 581
rect 711 462 777 546
rect 711 428 727 462
rect 761 428 777 462
rect 711 412 777 428
rect 817 531 851 547
rect 817 414 851 497
rect 637 378 671 380
rect 891 546 907 580
rect 941 546 957 580
rect 891 510 957 546
rect 891 476 907 510
rect 941 476 957 510
rect 891 440 957 476
rect 997 580 1031 649
rect 997 508 1031 546
rect 997 458 1031 474
rect 1071 580 1137 596
rect 1071 546 1087 580
rect 1121 546 1137 580
rect 1071 510 1137 546
rect 1071 476 1087 510
rect 1121 476 1137 510
rect 891 406 907 440
rect 941 424 957 440
rect 1071 440 1137 476
rect 1177 580 1227 649
rect 1211 546 1227 580
rect 1177 508 1227 546
rect 1211 474 1227 508
rect 1177 458 1227 474
rect 1267 580 1301 596
rect 1267 497 1301 546
rect 1071 424 1087 440
rect 941 406 1087 424
rect 1121 424 1137 440
rect 1267 424 1301 463
rect 1341 580 1391 649
rect 1341 546 1357 580
rect 1341 508 1391 546
rect 1341 474 1357 508
rect 1341 458 1391 474
rect 1431 580 1497 596
rect 1431 546 1447 580
rect 1481 546 1497 580
rect 1431 510 1497 546
rect 1431 476 1447 510
rect 1481 476 1497 510
rect 1431 440 1497 476
rect 1537 580 1571 649
rect 1537 508 1571 546
rect 1537 458 1571 474
rect 1611 580 1677 596
rect 1611 546 1627 580
rect 1661 546 1677 580
rect 1611 510 1677 546
rect 1611 476 1627 510
rect 1661 476 1677 510
rect 1431 424 1447 440
rect 1121 414 1447 424
rect 1121 406 1267 414
rect 891 390 1267 406
rect 817 378 851 380
rect 313 344 455 360
rect 637 344 851 378
rect 1301 406 1447 414
rect 1481 424 1497 440
rect 1611 440 1677 476
rect 1611 424 1627 440
rect 1481 406 1627 424
rect 1661 406 1677 440
rect 1301 390 1677 406
rect 1267 364 1301 380
rect 313 310 337 344
rect 371 310 455 344
rect 313 294 455 310
rect 515 294 717 310
rect 515 260 531 294
rect 565 260 599 294
rect 633 260 667 294
rect 701 260 717 294
rect 127 226 717 260
rect 793 226 851 344
rect 889 320 1223 356
rect 889 286 967 320
rect 1001 286 1035 320
rect 1069 286 1103 320
rect 1137 286 1171 320
rect 1205 286 1223 320
rect 889 270 1223 286
rect 1347 320 1703 356
rect 1347 286 1363 320
rect 1397 286 1431 320
rect 1465 286 1499 320
rect 1533 286 1567 320
rect 1601 286 1703 320
rect 1347 270 1703 286
rect 25 168 41 202
rect 75 168 91 202
rect 290 210 324 226
rect 25 134 91 168
rect 25 100 41 134
rect 75 100 91 134
rect 25 84 91 100
rect 188 190 254 192
rect 188 156 204 190
rect 238 156 254 190
rect 188 122 254 156
rect 188 88 204 122
rect 238 88 254 122
rect 188 17 254 88
rect 793 207 1230 226
rect 793 192 1008 207
rect 290 120 324 176
rect 290 70 324 86
rect 360 161 418 177
rect 360 127 380 161
rect 414 127 418 161
rect 360 17 418 127
rect 454 158 470 192
rect 504 158 642 192
rect 676 173 1008 192
rect 1042 173 1180 207
rect 1214 173 1230 207
rect 676 158 1230 173
rect 454 120 504 158
rect 454 86 470 120
rect 454 70 504 86
rect 540 122 606 124
rect 540 88 556 122
rect 590 88 606 122
rect 540 17 606 88
rect 642 120 676 158
rect 992 154 1230 158
rect 1266 210 1660 236
rect 1300 202 1438 210
rect 642 70 676 86
rect 712 122 778 124
rect 712 88 728 122
rect 762 88 778 122
rect 1266 120 1300 176
rect 1422 176 1438 202
rect 1472 202 1610 210
rect 712 17 778 88
rect 906 86 922 120
rect 956 86 1094 120
rect 1128 86 1266 120
rect 906 70 1300 86
rect 1336 152 1386 168
rect 1336 118 1352 152
rect 1336 17 1386 118
rect 1422 120 1472 176
rect 1594 176 1610 202
rect 1644 176 1660 210
rect 1422 86 1438 120
rect 1422 70 1472 86
rect 1508 152 1558 168
rect 1508 118 1524 152
rect 1508 17 1558 118
rect 1594 120 1660 176
rect 1594 86 1610 120
rect 1644 86 1660 120
rect 1594 70 1660 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a2bb2oi_4
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 1927830
string GDS_START 1913258
<< end >>
