magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3794 1975
<< nwell >>
rect -38 371 2534 704
rect -38 331 231 371
rect 485 331 2534 371
<< pwell >>
rect 338 279 443 329
rect 338 257 915 279
rect 1813 273 2172 289
rect 1813 257 2453 273
rect 338 241 1133 257
rect 3 217 1133 241
rect 1711 217 2453 257
rect 3 49 2453 217
rect 0 0 2496 49
<< scnmos >>
rect 86 47 116 215
rect 226 87 256 215
rect 439 73 469 201
rect 525 73 555 201
rect 665 125 695 253
rect 804 125 834 253
rect 1004 63 1034 231
rect 1146 63 1176 191
rect 1232 63 1262 191
rect 1470 63 1500 191
rect 1608 63 1638 191
rect 1787 63 1817 231
rect 1896 135 1926 263
rect 2036 135 2066 263
rect 2168 119 2198 247
rect 2340 79 2370 247
<< scpmoshvt >>
rect 86 367 116 619
rect 242 407 272 607
rect 442 407 472 575
rect 528 407 558 575
rect 660 379 690 547
rect 798 379 828 547
rect 1004 367 1034 619
rect 1122 389 1152 589
rect 1231 389 1261 557
rect 1475 389 1505 557
rect 1584 389 1614 589
rect 1744 367 1774 619
rect 1939 395 1969 563
rect 2025 395 2055 563
rect 2243 419 2273 619
rect 2383 367 2413 619
<< ndiff >>
rect 364 291 417 303
rect 364 257 373 291
rect 407 257 417 291
rect 29 203 86 215
rect 29 169 41 203
rect 75 169 86 203
rect 29 103 86 169
rect 29 69 41 103
rect 75 69 86 103
rect 29 47 86 69
rect 116 120 226 215
rect 116 86 127 120
rect 161 87 226 120
rect 256 181 310 215
rect 256 147 267 181
rect 301 147 310 181
rect 256 87 310 147
rect 364 201 417 257
rect 608 241 665 253
rect 608 207 620 241
rect 654 207 665 241
rect 608 201 665 207
rect 161 86 173 87
rect 116 47 173 86
rect 364 73 439 201
rect 469 119 525 201
rect 469 85 480 119
rect 514 85 525 119
rect 469 73 525 85
rect 555 173 665 201
rect 555 139 620 173
rect 654 139 665 173
rect 555 125 665 139
rect 695 179 804 253
rect 695 145 706 179
rect 740 145 804 179
rect 695 125 804 145
rect 834 241 889 253
rect 834 207 846 241
rect 880 207 889 241
rect 834 173 889 207
rect 834 139 846 173
rect 880 139 889 173
rect 834 125 889 139
rect 555 73 605 125
rect 949 184 1004 231
rect 949 150 959 184
rect 993 150 1004 184
rect 949 109 1004 150
rect 949 75 959 109
rect 993 75 1004 109
rect 949 63 1004 75
rect 1034 191 1107 231
rect 1839 231 1896 263
rect 1737 191 1787 231
rect 1034 111 1146 191
rect 1034 77 1061 111
rect 1095 77 1146 111
rect 1034 63 1146 77
rect 1176 179 1232 191
rect 1176 145 1187 179
rect 1221 145 1232 179
rect 1176 109 1232 145
rect 1176 75 1187 109
rect 1221 75 1232 109
rect 1176 63 1232 75
rect 1262 135 1470 191
rect 1262 101 1289 135
rect 1323 101 1470 135
rect 1262 63 1470 101
rect 1500 140 1608 191
rect 1500 106 1563 140
rect 1597 106 1608 140
rect 1500 63 1608 106
rect 1638 136 1787 191
rect 1638 102 1665 136
rect 1699 102 1787 136
rect 1638 63 1787 102
rect 1817 225 1896 231
rect 1817 191 1851 225
rect 1885 191 1896 225
rect 1817 135 1896 191
rect 1926 213 2036 263
rect 1926 179 1991 213
rect 2025 179 2036 213
rect 1926 135 2036 179
rect 2066 247 2146 263
rect 2066 245 2168 247
rect 2066 211 2100 245
rect 2134 211 2168 245
rect 2066 173 2168 211
rect 2066 139 2100 173
rect 2134 139 2168 173
rect 2066 135 2168 139
rect 1817 63 1867 135
rect 2088 119 2168 135
rect 2198 199 2340 247
rect 2198 165 2279 199
rect 2313 165 2340 199
rect 2198 125 2340 165
rect 2198 119 2279 125
rect 2267 91 2279 119
rect 2313 91 2340 125
rect 2267 79 2340 91
rect 2370 199 2427 247
rect 2370 165 2381 199
rect 2415 165 2427 199
rect 2370 125 2427 165
rect 2370 91 2381 125
rect 2415 91 2427 125
rect 2370 79 2427 91
<< pdiff >>
rect 29 597 86 619
rect 29 563 41 597
rect 75 563 86 597
rect 29 519 86 563
rect 29 485 41 519
rect 75 485 86 519
rect 29 442 86 485
rect 29 408 41 442
rect 75 408 86 442
rect 29 367 86 408
rect 116 607 173 619
rect 116 573 127 607
rect 161 573 242 607
rect 116 534 242 573
rect 116 500 127 534
rect 161 500 242 534
rect 116 461 242 500
rect 116 427 127 461
rect 161 427 242 461
rect 116 407 242 427
rect 272 494 329 607
rect 272 460 283 494
rect 317 460 329 494
rect 272 407 329 460
rect 385 455 442 575
rect 385 421 397 455
rect 431 421 442 455
rect 385 407 442 421
rect 472 527 528 575
rect 472 493 483 527
rect 517 493 528 527
rect 472 453 528 493
rect 472 419 483 453
rect 517 419 528 453
rect 472 407 528 419
rect 558 547 638 575
rect 558 527 660 547
rect 558 493 592 527
rect 626 493 660 527
rect 558 425 660 493
rect 558 407 592 425
rect 116 367 173 407
rect 580 391 592 407
rect 626 391 660 425
rect 580 379 660 391
rect 690 523 798 547
rect 690 489 701 523
rect 735 489 798 523
rect 690 379 798 489
rect 828 527 887 547
rect 828 493 841 527
rect 875 493 887 527
rect 828 425 887 493
rect 828 391 841 425
rect 875 391 887 425
rect 828 379 887 391
rect 947 427 1004 619
rect 947 393 959 427
rect 993 393 1004 427
rect 947 367 1004 393
rect 1034 607 1091 619
rect 1034 573 1045 607
rect 1079 589 1091 607
rect 1687 607 1744 619
rect 1687 589 1699 607
rect 1079 573 1122 589
rect 1034 389 1122 573
rect 1152 557 1209 589
rect 1527 557 1584 589
rect 1152 435 1231 557
rect 1152 401 1163 435
rect 1197 401 1231 435
rect 1152 389 1231 401
rect 1261 527 1475 557
rect 1261 493 1321 527
rect 1355 493 1475 527
rect 1261 442 1475 493
rect 1261 408 1321 442
rect 1355 408 1475 442
rect 1261 389 1475 408
rect 1505 527 1584 557
rect 1505 493 1539 527
rect 1573 493 1584 527
rect 1505 435 1584 493
rect 1505 401 1539 435
rect 1573 401 1584 435
rect 1505 389 1584 401
rect 1614 573 1699 589
rect 1733 573 1744 607
rect 1614 522 1744 573
rect 1614 488 1699 522
rect 1733 488 1744 522
rect 1614 438 1744 488
rect 1614 404 1699 438
rect 1733 404 1744 438
rect 1614 389 1744 404
rect 1034 367 1091 389
rect 1687 367 1744 389
rect 1774 597 1829 619
rect 1774 563 1785 597
rect 1819 563 1829 597
rect 2077 597 2133 609
rect 2077 563 2088 597
rect 2122 563 2133 597
rect 1774 517 1829 563
rect 1774 483 1785 517
rect 1819 483 1829 517
rect 1774 438 1829 483
rect 1774 404 1785 438
rect 1819 404 1829 438
rect 1774 367 1829 404
rect 1883 527 1939 563
rect 1883 493 1894 527
rect 1928 493 1939 527
rect 1883 395 1939 493
rect 1969 441 2025 563
rect 1969 407 1980 441
rect 2014 407 2025 441
rect 1969 395 2025 407
rect 2055 395 2133 563
rect 2187 509 2243 619
rect 2187 475 2198 509
rect 2232 475 2243 509
rect 2187 419 2243 475
rect 2273 607 2383 619
rect 2273 573 2338 607
rect 2372 573 2383 607
rect 2273 514 2383 573
rect 2273 480 2338 514
rect 2372 480 2383 514
rect 2273 421 2383 480
rect 2273 419 2338 421
rect 2326 387 2338 419
rect 2372 387 2383 421
rect 2326 367 2383 387
rect 2413 597 2469 619
rect 2413 563 2424 597
rect 2458 563 2469 597
rect 2413 505 2469 563
rect 2413 471 2424 505
rect 2458 471 2469 505
rect 2413 413 2469 471
rect 2413 379 2424 413
rect 2458 379 2469 413
rect 2413 367 2469 379
<< ndiffc >>
rect 373 257 407 291
rect 41 169 75 203
rect 41 69 75 103
rect 127 86 161 120
rect 267 147 301 181
rect 620 207 654 241
rect 480 85 514 119
rect 620 139 654 173
rect 706 145 740 179
rect 846 207 880 241
rect 846 139 880 173
rect 959 150 993 184
rect 959 75 993 109
rect 1061 77 1095 111
rect 1187 145 1221 179
rect 1187 75 1221 109
rect 1289 101 1323 135
rect 1563 106 1597 140
rect 1665 102 1699 136
rect 1851 191 1885 225
rect 1991 179 2025 213
rect 2100 211 2134 245
rect 2100 139 2134 173
rect 2279 165 2313 199
rect 2279 91 2313 125
rect 2381 165 2415 199
rect 2381 91 2415 125
<< pdiffc >>
rect 41 563 75 597
rect 41 485 75 519
rect 41 408 75 442
rect 127 573 161 607
rect 127 500 161 534
rect 127 427 161 461
rect 283 460 317 494
rect 397 421 431 455
rect 483 493 517 527
rect 483 419 517 453
rect 592 493 626 527
rect 592 391 626 425
rect 701 489 735 523
rect 841 493 875 527
rect 841 391 875 425
rect 959 393 993 427
rect 1045 573 1079 607
rect 1163 401 1197 435
rect 1321 493 1355 527
rect 1321 408 1355 442
rect 1539 493 1573 527
rect 1539 401 1573 435
rect 1699 573 1733 607
rect 1699 488 1733 522
rect 1699 404 1733 438
rect 1785 563 1819 597
rect 2088 563 2122 597
rect 1785 483 1819 517
rect 1785 404 1819 438
rect 1894 493 1928 527
rect 1980 407 2014 441
rect 2198 475 2232 509
rect 2338 573 2372 607
rect 2338 480 2372 514
rect 2338 387 2372 421
rect 2424 563 2458 597
rect 2424 471 2458 505
rect 2424 379 2458 413
<< poly >>
rect 86 619 116 645
rect 242 607 272 633
rect 528 615 828 645
rect 1004 619 1034 645
rect 1744 619 1774 645
rect 2243 619 2273 645
rect 2383 619 2413 645
rect 442 575 472 601
rect 528 575 558 615
rect 798 599 828 615
rect 660 547 690 573
rect 798 569 932 599
rect 798 547 828 569
rect 242 375 272 407
rect 86 335 116 367
rect 206 359 272 375
rect 86 319 158 335
rect 86 285 108 319
rect 142 285 158 319
rect 86 269 158 285
rect 206 325 222 359
rect 256 325 272 359
rect 206 291 272 325
rect 442 305 472 407
rect 528 381 558 407
rect 660 341 690 379
rect 798 353 828 379
rect 660 325 756 341
rect 660 305 706 325
rect 86 215 116 269
rect 206 257 222 291
rect 256 257 272 291
rect 206 241 272 257
rect 226 215 256 241
rect 439 291 706 305
rect 740 291 756 325
rect 439 275 756 291
rect 902 334 932 569
rect 1122 589 1152 615
rect 1584 589 1614 615
rect 1231 557 1261 583
rect 1475 557 1505 583
rect 1004 334 1034 367
rect 902 318 1034 334
rect 1122 319 1152 389
rect 1231 357 1261 389
rect 1475 367 1505 389
rect 902 284 948 318
rect 982 284 1034 318
rect 439 201 469 275
rect 665 253 695 275
rect 804 253 834 279
rect 902 268 1034 284
rect 525 201 555 227
rect 226 61 256 87
rect 665 99 695 125
rect 439 47 469 73
rect 525 51 555 73
rect 804 51 834 125
rect 904 51 934 268
rect 1004 231 1034 268
rect 1076 303 1152 319
rect 1076 269 1092 303
rect 1126 269 1152 303
rect 1218 341 1284 357
rect 1218 307 1234 341
rect 1268 307 1284 341
rect 1218 291 1284 307
rect 1398 337 1505 367
rect 1398 279 1428 337
rect 1584 313 1614 389
rect 1939 563 1969 589
rect 2025 563 2055 589
rect 1076 253 1152 269
rect 1122 243 1152 253
rect 1362 263 1428 279
rect 1362 243 1378 263
rect 1122 213 1176 243
rect 1146 191 1176 213
rect 1232 229 1378 243
rect 1412 229 1428 263
rect 1232 213 1428 229
rect 1470 273 1536 289
rect 1584 283 1679 313
rect 1744 283 1774 367
rect 1939 315 1969 395
rect 2025 363 2055 395
rect 2243 387 2273 419
rect 2207 371 2273 387
rect 1896 285 1969 315
rect 2021 347 2087 363
rect 2207 351 2223 371
rect 2021 313 2037 347
rect 2071 313 2087 347
rect 2021 297 2087 313
rect 2168 337 2223 351
rect 2257 337 2273 371
rect 2168 321 2273 337
rect 2383 335 2413 367
rect 1470 239 1486 273
rect 1520 239 1536 273
rect 1470 223 1536 239
rect 1608 266 1817 283
rect 1608 232 1665 266
rect 1699 253 1817 266
rect 1896 263 1926 285
rect 2036 263 2066 297
rect 1699 232 1715 253
rect 1232 191 1262 213
rect 1470 191 1500 223
rect 1608 216 1715 232
rect 1787 231 1817 253
rect 1608 191 1638 216
rect 2168 247 2198 321
rect 2322 319 2413 335
rect 2322 285 2338 319
rect 2372 285 2413 319
rect 2322 269 2413 285
rect 2340 247 2370 269
rect 1896 113 1926 135
rect 1889 97 1955 113
rect 2036 109 2066 135
rect 1889 63 1905 97
rect 1939 63 1955 97
rect 2168 93 2198 119
rect 86 21 116 47
rect 525 21 934 51
rect 1004 37 1034 63
rect 1146 37 1176 63
rect 1232 37 1262 63
rect 1470 37 1500 63
rect 1608 37 1638 63
rect 1787 37 1817 63
rect 1889 47 1955 63
rect 2340 53 2370 79
<< polycont >>
rect 108 285 142 319
rect 222 325 256 359
rect 222 257 256 291
rect 706 291 740 325
rect 948 284 982 318
rect 1092 269 1126 303
rect 1234 307 1268 341
rect 1378 229 1412 263
rect 2037 313 2071 347
rect 2223 337 2257 371
rect 1486 239 1520 273
rect 1665 232 1699 266
rect 2338 285 2372 319
rect 1905 63 1939 97
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 22 597 75 613
rect 22 563 41 597
rect 22 519 75 563
rect 22 485 41 519
rect 22 442 75 485
rect 22 408 41 442
rect 111 607 177 649
rect 111 573 127 607
rect 161 573 177 607
rect 111 534 177 573
rect 111 500 127 534
rect 161 500 177 534
rect 111 461 177 500
rect 111 427 127 461
rect 161 427 177 461
rect 111 411 177 427
rect 213 579 735 613
rect 22 392 75 408
rect 22 233 56 392
rect 213 375 247 579
rect 283 527 533 543
rect 283 509 483 527
rect 283 494 333 509
rect 317 460 333 494
rect 467 493 483 509
rect 517 493 533 527
rect 283 411 333 460
rect 381 455 431 473
rect 381 421 397 455
rect 197 359 272 375
rect 92 319 161 356
rect 92 285 108 319
rect 142 285 161 319
rect 92 269 161 285
rect 197 325 222 359
rect 256 325 272 359
rect 381 356 431 421
rect 197 291 272 325
rect 313 350 431 356
rect 313 316 319 350
rect 353 316 431 350
rect 313 310 431 316
rect 197 257 222 291
rect 256 257 272 291
rect 197 241 272 257
rect 357 291 431 310
rect 357 257 373 291
rect 407 257 431 291
rect 357 241 431 257
rect 467 453 533 493
rect 467 419 483 453
rect 517 419 533 453
rect 197 233 231 241
rect 22 203 231 233
rect 467 205 533 419
rect 576 527 654 543
rect 576 493 592 527
rect 626 493 654 527
rect 576 426 654 493
rect 701 523 735 579
rect 701 462 735 489
rect 771 579 993 613
rect 771 426 805 579
rect 576 425 805 426
rect 576 391 592 425
rect 626 392 805 425
rect 841 527 896 543
rect 875 493 896 527
rect 841 425 896 493
rect 959 521 993 579
rect 1029 607 1095 649
rect 1029 573 1045 607
rect 1079 573 1095 607
rect 1029 557 1095 573
rect 1233 579 1663 613
rect 1233 521 1269 579
rect 959 487 1269 521
rect 626 391 654 392
rect 576 375 654 391
rect 620 241 654 375
rect 875 391 896 425
rect 841 356 896 391
rect 943 427 1009 451
rect 943 393 959 427
rect 993 404 1009 427
rect 1163 435 1197 451
rect 993 393 1127 404
rect 943 370 1127 393
rect 793 350 896 356
rect 690 325 756 341
rect 690 291 706 325
rect 740 291 756 325
rect 793 316 799 350
rect 833 316 896 350
rect 793 310 896 316
rect 690 274 756 291
rect 690 240 810 274
rect 22 169 41 203
rect 75 199 231 203
rect 75 169 91 199
rect 22 103 91 169
rect 22 69 41 103
rect 75 69 91 103
rect 22 53 91 69
rect 127 120 161 163
rect 127 17 161 86
rect 197 87 231 199
rect 267 181 584 205
rect 301 171 584 181
rect 301 147 317 171
rect 267 123 317 147
rect 464 119 514 135
rect 464 87 480 119
rect 197 85 480 87
rect 197 53 514 85
rect 550 87 584 171
rect 620 173 654 207
rect 620 123 654 139
rect 690 179 740 204
rect 690 145 706 179
rect 690 87 740 145
rect 550 53 740 87
rect 776 87 810 240
rect 846 241 896 310
rect 880 207 896 241
rect 932 318 1031 334
rect 932 284 948 318
rect 982 284 1031 318
rect 932 236 1031 284
rect 1076 303 1127 370
rect 1076 269 1092 303
rect 1126 269 1127 303
rect 846 173 896 207
rect 1076 200 1127 269
rect 880 139 896 173
rect 846 123 896 139
rect 943 184 1127 200
rect 943 150 959 184
rect 993 166 1127 184
rect 1163 195 1197 401
rect 1233 341 1269 487
rect 1233 307 1234 341
rect 1268 307 1269 341
rect 1233 291 1269 307
rect 1305 527 1371 543
rect 1305 493 1321 527
rect 1355 493 1371 527
rect 1305 442 1371 493
rect 1305 408 1321 442
rect 1355 408 1371 442
rect 1305 392 1371 408
rect 1163 179 1237 195
rect 993 150 1009 166
rect 943 109 1009 150
rect 1163 145 1187 179
rect 1221 145 1237 179
rect 1305 177 1339 392
rect 1375 350 1415 356
rect 1409 316 1415 350
rect 1375 279 1415 316
rect 1453 349 1487 579
rect 1523 527 1593 543
rect 1523 493 1539 527
rect 1573 493 1593 527
rect 1523 435 1593 493
rect 1523 401 1539 435
rect 1573 401 1593 435
rect 1523 385 1593 401
rect 1453 315 1523 349
rect 1375 263 1428 279
rect 1375 229 1378 263
rect 1412 229 1428 263
rect 1375 213 1428 229
rect 1470 273 1523 315
rect 1470 239 1486 273
rect 1520 239 1523 273
rect 1470 223 1523 239
rect 1559 187 1593 385
rect 1629 352 1663 579
rect 1699 607 1733 649
rect 1699 522 1733 573
rect 1699 438 1733 488
rect 1699 388 1733 404
rect 1769 597 2302 613
rect 1769 563 1785 597
rect 1819 579 2088 597
rect 1819 563 1858 579
rect 1769 517 1858 563
rect 2072 563 2088 579
rect 2122 579 2302 597
rect 2122 563 2138 579
rect 2072 547 2138 563
rect 1769 483 1785 517
rect 1819 483 1858 517
rect 1769 438 1858 483
rect 1894 527 1944 543
rect 1928 511 1944 527
rect 2182 511 2232 543
rect 1928 509 2232 511
rect 1928 493 2198 509
rect 1894 477 2198 493
rect 2123 475 2198 477
rect 2123 441 2232 475
rect 1769 404 1785 438
rect 1819 404 1858 438
rect 1769 388 1858 404
rect 1629 318 1785 352
rect 1649 266 1715 282
rect 1649 232 1665 266
rect 1699 232 1715 266
rect 1649 216 1715 232
rect 943 87 959 109
rect 776 75 959 87
rect 993 75 1009 109
rect 776 53 1009 75
rect 1045 111 1111 130
rect 1045 77 1061 111
rect 1095 77 1111 111
rect 1045 17 1111 77
rect 1163 109 1237 145
rect 1163 75 1187 109
rect 1221 75 1237 109
rect 1163 59 1237 75
rect 1273 135 1511 177
rect 1273 101 1289 135
rect 1323 101 1511 135
rect 1273 88 1511 101
rect 1547 140 1613 187
rect 1547 106 1563 140
rect 1597 106 1613 140
rect 1273 59 1339 88
rect 1547 59 1613 106
rect 1649 136 1715 180
rect 1649 102 1665 136
rect 1699 102 1715 136
rect 1649 17 1715 102
rect 1751 113 1785 318
rect 1824 267 1858 388
rect 1951 407 1980 441
rect 2014 407 2030 441
rect 1824 225 1901 267
rect 1951 261 1985 407
rect 2021 350 2087 363
rect 2021 347 2047 350
rect 2021 313 2037 347
rect 2081 316 2087 350
rect 2071 313 2087 316
rect 2021 297 2087 313
rect 2123 261 2157 441
rect 2268 405 2302 579
rect 2207 371 2302 405
rect 2338 607 2388 649
rect 2372 573 2388 607
rect 2338 514 2388 573
rect 2372 480 2388 514
rect 2338 421 2388 480
rect 2372 387 2388 421
rect 2338 371 2388 387
rect 2424 597 2474 613
rect 2458 563 2474 597
rect 2424 505 2474 563
rect 2458 471 2474 505
rect 2424 413 2474 471
rect 2458 379 2474 413
rect 2207 337 2223 371
rect 2257 337 2273 371
rect 2207 321 2273 337
rect 2322 319 2388 335
rect 2322 285 2338 319
rect 2372 285 2388 319
rect 1951 227 2041 261
rect 1824 191 1851 225
rect 1885 191 1901 225
rect 1824 149 1901 191
rect 1991 213 2041 227
rect 2025 179 2041 213
rect 1751 97 1955 113
rect 1751 63 1905 97
rect 1939 63 1955 97
rect 1751 53 1955 63
rect 1991 87 2041 179
rect 2084 245 2157 261
rect 2084 211 2100 245
rect 2134 211 2157 245
rect 2084 173 2157 211
rect 2084 139 2100 173
rect 2134 139 2157 173
rect 2084 123 2157 139
rect 2193 251 2388 285
rect 2193 87 2227 251
rect 2424 215 2474 379
rect 1991 53 2227 87
rect 2263 199 2329 215
rect 2263 165 2279 199
rect 2313 165 2329 199
rect 2263 125 2329 165
rect 2263 91 2279 125
rect 2313 91 2329 125
rect 2263 17 2329 91
rect 2365 199 2474 215
rect 2365 165 2381 199
rect 2415 165 2474 199
rect 2365 125 2474 165
rect 2365 91 2381 125
rect 2415 91 2474 125
rect 2365 75 2474 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 319 316 353 350
rect 799 316 833 350
rect 1375 316 1409 350
rect 2047 347 2081 350
rect 2047 316 2071 347
rect 2071 316 2081 347
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 683 2496 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2496 683
rect 0 617 2496 649
rect 307 350 365 356
rect 307 316 319 350
rect 353 347 365 350
rect 787 350 845 356
rect 787 347 799 350
rect 353 319 799 347
rect 353 316 365 319
rect 307 310 365 316
rect 787 316 799 319
rect 833 347 845 350
rect 1363 350 1421 356
rect 1363 347 1375 350
rect 833 319 1375 347
rect 833 316 845 319
rect 787 310 845 316
rect 1363 316 1375 319
rect 1409 347 1421 350
rect 2035 350 2093 356
rect 2035 347 2047 350
rect 1409 319 2047 347
rect 1409 316 1421 319
rect 1363 310 1421 316
rect 2035 316 2047 319
rect 2081 316 2093 350
rect 2035 310 2093 316
rect 0 17 2496 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
rect 0 -49 2496 -17
<< labels >>
flabel pwell s 0 0 2496 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2496 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fahcin_1
flabel metal1 s 0 617 2496 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2496 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 2431 94 2465 128 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2431 168 2465 202 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2431 242 2465 276 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2431 316 2465 350 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2431 390 2465 424 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2431 464 2465 498 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2431 538 2465 572 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1279 94 1313 128 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 1375 94 1409 128 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 1471 94 1505 128 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2496 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5747574
string GDS_START 5729436
<< end >>
