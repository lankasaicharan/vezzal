magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
<< pwell >>
rect 1021 236 1349 281
rect 56 157 1349 236
rect 56 49 1631 157
rect 0 0 1632 49
<< scnmos >>
rect 135 126 165 210
rect 243 126 273 210
rect 315 126 345 210
rect 423 126 453 210
rect 495 126 525 210
rect 586 126 616 210
rect 658 126 688 210
rect 744 126 774 210
rect 816 126 846 210
rect 1154 171 1184 255
rect 1240 171 1270 255
rect 1436 47 1466 131
rect 1522 47 1552 131
<< scpmoshvt >>
rect 112 463 142 547
rect 243 463 273 547
rect 315 463 345 547
rect 401 463 431 547
rect 473 463 503 547
rect 617 463 647 547
rect 689 463 719 547
rect 775 463 805 547
rect 847 463 877 547
rect 1154 463 1184 547
rect 1240 463 1270 547
rect 1436 527 1466 611
rect 1522 527 1552 611
<< ndiff >>
rect 82 198 135 210
rect 82 164 90 198
rect 124 164 135 198
rect 82 126 135 164
rect 165 172 243 210
rect 165 138 192 172
rect 226 138 243 172
rect 165 126 243 138
rect 273 126 315 210
rect 345 175 423 210
rect 345 141 378 175
rect 412 141 423 175
rect 345 126 423 141
rect 453 126 495 210
rect 525 168 586 210
rect 525 134 541 168
rect 575 134 586 168
rect 525 126 586 134
rect 616 126 658 210
rect 688 180 744 210
rect 688 146 699 180
rect 733 146 744 180
rect 688 126 744 146
rect 774 126 816 210
rect 846 172 899 210
rect 846 138 857 172
rect 891 138 899 172
rect 846 126 899 138
rect 1047 243 1154 255
rect 1047 209 1055 243
rect 1089 209 1154 243
rect 1047 171 1154 209
rect 1184 243 1240 255
rect 1184 209 1195 243
rect 1229 209 1240 243
rect 1184 171 1240 209
rect 1270 217 1323 255
rect 1270 183 1281 217
rect 1315 183 1323 217
rect 1270 171 1323 183
rect 1383 103 1436 131
rect 1383 69 1391 103
rect 1425 69 1436 103
rect 1383 47 1436 69
rect 1466 93 1522 131
rect 1466 59 1477 93
rect 1511 59 1522 93
rect 1466 47 1522 59
rect 1552 119 1605 131
rect 1552 85 1563 119
rect 1597 85 1605 119
rect 1552 47 1605 85
<< pdiff >>
rect 59 509 112 547
rect 59 475 67 509
rect 101 475 112 509
rect 59 463 112 475
rect 142 535 243 547
rect 142 501 153 535
rect 187 501 243 535
rect 142 463 243 501
rect 273 463 315 547
rect 345 509 401 547
rect 345 475 356 509
rect 390 475 401 509
rect 345 463 401 475
rect 431 463 473 547
rect 503 539 617 547
rect 503 505 515 539
rect 549 505 617 539
rect 503 463 617 505
rect 647 463 689 547
rect 719 509 775 547
rect 719 475 730 509
rect 764 475 775 509
rect 719 463 775 475
rect 805 463 847 547
rect 877 535 957 547
rect 877 501 915 535
rect 949 501 957 535
rect 877 463 957 501
rect 1047 509 1154 547
rect 1047 475 1055 509
rect 1089 475 1154 509
rect 1047 463 1154 475
rect 1184 509 1240 547
rect 1184 475 1195 509
rect 1229 475 1240 509
rect 1184 463 1240 475
rect 1270 535 1323 547
rect 1270 501 1281 535
rect 1315 501 1323 535
rect 1270 463 1323 501
rect 1383 573 1436 611
rect 1383 539 1391 573
rect 1425 539 1436 573
rect 1383 527 1436 539
rect 1466 599 1522 611
rect 1466 565 1477 599
rect 1511 565 1522 599
rect 1466 527 1522 565
rect 1552 573 1605 611
rect 1552 539 1563 573
rect 1597 539 1605 573
rect 1552 527 1605 539
<< ndiffc >>
rect 90 164 124 198
rect 192 138 226 172
rect 378 141 412 175
rect 541 134 575 168
rect 699 146 733 180
rect 857 138 891 172
rect 1055 209 1089 243
rect 1195 209 1229 243
rect 1281 183 1315 217
rect 1391 69 1425 103
rect 1477 59 1511 93
rect 1563 85 1597 119
<< pdiffc >>
rect 67 475 101 509
rect 153 501 187 535
rect 356 475 390 509
rect 515 505 549 539
rect 730 475 764 509
rect 915 501 949 535
rect 1055 475 1089 509
rect 1195 475 1229 509
rect 1281 501 1315 535
rect 1391 539 1425 573
rect 1477 565 1511 599
rect 1563 539 1597 573
<< poly >>
rect 315 615 1002 645
rect 112 547 142 573
rect 243 547 273 573
rect 315 547 345 615
rect 401 547 431 573
rect 473 547 503 573
rect 617 547 647 573
rect 689 547 719 573
rect 775 547 805 615
rect 847 547 877 573
rect 112 262 142 463
rect 243 431 273 463
rect 315 437 345 463
rect 207 415 273 431
rect 207 381 223 415
rect 257 381 273 415
rect 207 347 273 381
rect 401 366 431 463
rect 207 313 223 347
rect 257 313 273 347
rect 207 297 273 313
rect 112 232 165 262
rect 135 210 165 232
rect 243 210 273 297
rect 315 350 431 366
rect 315 316 331 350
rect 365 336 431 350
rect 473 412 503 463
rect 617 412 647 463
rect 473 396 539 412
rect 473 362 489 396
rect 523 362 539 396
rect 365 316 381 336
rect 315 282 381 316
rect 315 248 331 282
rect 365 248 381 282
rect 473 328 539 362
rect 473 294 489 328
rect 523 294 539 328
rect 473 278 539 294
rect 581 396 647 412
rect 581 362 597 396
rect 631 362 647 396
rect 581 328 647 362
rect 581 294 597 328
rect 631 294 647 328
rect 689 376 719 463
rect 775 437 805 463
rect 689 360 774 376
rect 689 326 705 360
rect 739 326 774 360
rect 689 310 774 326
rect 581 278 647 294
rect 315 232 381 248
rect 315 210 345 232
rect 423 210 453 236
rect 495 210 525 278
rect 586 210 616 278
rect 658 210 688 236
rect 744 210 774 310
rect 847 298 877 463
rect 847 282 913 298
rect 847 262 863 282
rect 816 248 863 262
rect 897 248 913 282
rect 816 232 913 248
rect 816 210 846 232
rect 135 103 165 126
rect 69 87 165 103
rect 243 100 273 126
rect 315 100 345 126
rect 69 53 85 87
rect 119 53 165 87
rect 69 52 165 53
rect 423 52 453 126
rect 495 100 525 126
rect 586 100 616 126
rect 658 52 688 126
rect 744 100 774 126
rect 816 100 846 126
rect 972 52 1002 615
rect 1154 615 1368 645
rect 1154 547 1184 615
rect 1240 547 1270 573
rect 1338 505 1368 615
rect 1436 611 1466 637
rect 1522 611 1552 637
rect 1436 505 1466 527
rect 1338 475 1466 505
rect 1154 437 1184 463
rect 1240 427 1270 463
rect 1240 411 1335 427
rect 1240 389 1285 411
rect 1154 377 1285 389
rect 1319 377 1335 411
rect 1154 359 1335 377
rect 1154 255 1184 359
rect 1395 307 1425 475
rect 1522 372 1552 527
rect 1240 277 1425 307
rect 1240 255 1270 277
rect 1359 271 1425 277
rect 1359 237 1375 271
rect 1409 237 1425 271
rect 1473 356 1552 372
rect 1473 322 1489 356
rect 1523 322 1552 356
rect 1473 288 1552 322
rect 1473 254 1489 288
rect 1523 254 1552 288
rect 1473 238 1552 254
rect 1359 203 1425 237
rect 1154 103 1184 171
rect 1240 145 1270 171
rect 1359 169 1375 203
rect 1409 183 1425 203
rect 1409 169 1466 183
rect 1359 153 1466 169
rect 1436 131 1466 153
rect 1522 131 1552 238
rect 69 22 1002 52
rect 1118 87 1184 103
rect 1118 53 1134 87
rect 1168 53 1184 87
rect 1118 37 1184 53
rect 1436 21 1466 47
rect 1522 21 1552 47
<< polycont >>
rect 223 381 257 415
rect 223 313 257 347
rect 331 316 365 350
rect 489 362 523 396
rect 331 248 365 282
rect 489 294 523 328
rect 597 362 631 396
rect 597 294 631 328
rect 705 326 739 360
rect 863 248 897 282
rect 85 53 119 87
rect 1285 377 1319 411
rect 1375 237 1409 271
rect 1489 322 1523 356
rect 1489 254 1523 288
rect 1375 169 1409 203
rect 1134 53 1168 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 149 535 187 649
rect 63 509 105 525
rect 63 475 67 509
rect 101 475 105 509
rect 149 501 153 535
rect 149 485 187 501
rect 63 261 105 475
rect 223 415 257 572
rect 499 539 565 649
rect 352 509 401 525
rect 352 475 356 509
rect 390 475 401 509
rect 499 505 515 539
rect 549 505 565 539
rect 601 549 879 583
rect 352 469 401 475
rect 601 469 635 549
rect 714 509 809 513
rect 714 475 730 509
rect 764 475 809 509
rect 714 471 809 475
rect 352 435 635 469
rect 223 347 257 381
rect 223 297 257 313
rect 304 350 365 366
rect 304 316 331 350
rect 304 282 365 316
rect 304 261 331 282
rect 63 248 331 261
rect 63 227 365 248
rect 63 198 140 227
rect 63 164 90 198
rect 124 164 140 198
rect 176 172 242 176
rect 176 138 192 172
rect 226 138 242 172
rect 31 87 65 128
rect 31 53 85 87
rect 119 53 135 87
rect 176 17 242 138
rect 304 89 338 227
rect 401 191 435 435
rect 473 362 489 396
rect 523 362 545 396
rect 473 328 545 362
rect 473 294 489 328
rect 523 294 545 328
rect 581 362 597 396
rect 631 362 647 396
rect 775 379 809 471
rect 845 449 879 549
rect 915 535 949 649
rect 1473 599 1515 649
rect 915 485 949 501
rect 985 561 1319 595
rect 985 449 1019 561
rect 845 415 1019 449
rect 1055 509 1089 525
rect 1055 379 1089 475
rect 581 328 647 362
rect 581 294 597 328
rect 631 294 647 328
rect 705 360 739 376
rect 705 254 739 326
rect 374 175 435 191
rect 374 141 378 175
rect 412 141 435 175
rect 374 125 435 141
rect 471 220 739 254
rect 775 345 1089 379
rect 471 89 505 220
rect 775 184 809 345
rect 863 282 929 298
rect 897 248 929 282
rect 863 232 929 248
rect 1051 243 1089 345
rect 1051 209 1055 243
rect 1051 193 1089 209
rect 304 55 505 89
rect 541 168 579 184
rect 575 134 579 168
rect 683 180 809 184
rect 683 146 699 180
rect 733 146 809 180
rect 683 142 809 146
rect 853 172 895 188
rect 541 17 579 134
rect 853 138 857 172
rect 891 138 895 172
rect 853 17 895 138
rect 1125 157 1159 561
rect 1277 535 1319 561
rect 1195 509 1233 525
rect 1229 475 1233 509
rect 1277 501 1281 535
rect 1315 501 1319 535
rect 1277 485 1319 501
rect 1387 573 1429 589
rect 1387 539 1391 573
rect 1425 539 1429 573
rect 1473 565 1477 599
rect 1511 565 1515 599
rect 1473 549 1515 565
rect 1559 573 1601 589
rect 1195 341 1233 475
rect 1387 411 1429 539
rect 1269 377 1285 411
rect 1319 377 1429 411
rect 1559 539 1563 573
rect 1597 539 1601 573
rect 1489 356 1523 372
rect 1195 322 1489 341
rect 1195 307 1523 322
rect 1195 243 1233 307
rect 1489 288 1523 307
rect 1229 209 1233 243
rect 1359 237 1375 271
rect 1409 237 1425 271
rect 1489 238 1523 254
rect 1195 193 1233 209
rect 1277 217 1319 233
rect 1277 183 1281 217
rect 1315 183 1319 217
rect 1277 157 1319 183
rect 1359 203 1425 237
rect 1359 169 1375 203
rect 1409 169 1425 203
rect 1359 168 1425 169
rect 1125 123 1319 157
rect 1559 119 1601 539
rect 1387 103 1429 119
rect 1387 87 1391 103
rect 1118 53 1134 87
rect 1168 69 1391 87
rect 1425 69 1429 103
rect 1168 53 1429 69
rect 1477 93 1515 109
rect 1511 59 1515 93
rect 1559 85 1563 119
rect 1597 85 1601 119
rect 1559 69 1601 85
rect 1477 17 1515 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux4_m
flabel comment s 1167 281 1167 281 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 1375 168 1409 202 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1548504
string GDS_START 1536338
<< end >>
