magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1586 1975
<< nwell >>
rect -38 331 326 704
<< pwell >>
rect 3 49 269 263
rect 0 0 288 49
<< scnmos >>
rect 82 69 112 237
rect 160 69 190 237
<< scpmoshvt >>
rect 82 367 112 619
rect 168 367 198 619
<< ndiff >>
rect 29 208 82 237
rect 29 174 37 208
rect 71 174 82 208
rect 29 115 82 174
rect 29 81 37 115
rect 71 81 82 115
rect 29 69 82 81
rect 112 69 160 237
rect 190 208 243 237
rect 190 174 201 208
rect 235 174 243 208
rect 190 122 243 174
rect 190 88 201 122
rect 235 88 243 122
rect 190 69 243 88
<< pdiff >>
rect 29 607 82 619
rect 29 573 37 607
rect 71 573 82 607
rect 29 515 82 573
rect 29 481 37 515
rect 71 481 82 515
rect 29 418 82 481
rect 29 384 37 418
rect 71 384 82 418
rect 29 367 82 384
rect 112 599 168 619
rect 112 565 123 599
rect 157 565 168 599
rect 112 508 168 565
rect 112 474 123 508
rect 157 474 168 508
rect 112 413 168 474
rect 112 379 123 413
rect 157 379 168 413
rect 112 367 168 379
rect 198 607 251 619
rect 198 573 209 607
rect 243 573 251 607
rect 198 523 251 573
rect 198 489 209 523
rect 243 489 251 523
rect 198 434 251 489
rect 198 400 209 434
rect 243 400 251 434
rect 198 367 251 400
<< ndiffc >>
rect 37 174 71 208
rect 37 81 71 115
rect 201 174 235 208
rect 201 88 235 122
<< pdiffc >>
rect 37 573 71 607
rect 37 481 71 515
rect 37 384 71 418
rect 123 565 157 599
rect 123 474 157 508
rect 123 379 157 413
rect 209 573 243 607
rect 209 489 243 523
rect 209 400 243 434
<< poly >>
rect 82 619 112 645
rect 168 619 198 645
rect 82 325 112 367
rect 33 309 112 325
rect 33 275 49 309
rect 83 275 112 309
rect 168 325 198 367
rect 168 309 247 325
rect 168 289 197 309
rect 33 259 112 275
rect 82 237 112 259
rect 160 275 197 289
rect 231 275 247 309
rect 160 259 247 275
rect 160 237 190 259
rect 82 43 112 69
rect 160 43 190 69
<< polycont >>
rect 49 275 83 309
rect 197 275 231 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 21 607 87 649
rect 21 573 37 607
rect 71 573 87 607
rect 21 515 87 573
rect 21 481 37 515
rect 71 481 87 515
rect 21 418 87 481
rect 21 384 37 418
rect 71 384 87 418
rect 121 599 163 615
rect 121 565 123 599
rect 157 565 163 599
rect 121 508 163 565
rect 121 474 123 508
rect 157 474 163 508
rect 121 413 163 474
rect 121 379 123 413
rect 157 379 163 413
rect 197 607 259 649
rect 197 573 209 607
rect 243 573 259 607
rect 197 523 259 573
rect 197 489 209 523
rect 243 489 259 523
rect 197 434 259 489
rect 197 400 209 434
rect 243 400 259 434
rect 197 384 259 400
rect 17 309 87 350
rect 17 275 49 309
rect 83 275 87 309
rect 17 242 87 275
rect 121 208 163 379
rect 197 309 271 350
rect 231 275 271 309
rect 197 242 271 275
rect 21 174 37 208
rect 71 174 87 208
rect 21 115 87 174
rect 21 81 37 115
rect 71 81 87 115
rect 21 17 87 81
rect 121 174 201 208
rect 235 174 251 208
rect 121 122 251 174
rect 121 88 201 122
rect 235 88 251 122
rect 121 72 251 88
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
<< metal1 >>
rect 0 683 288 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 288 683
rect 0 617 288 649
rect 0 17 288 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 288 17
rect 0 -49 288 -17
<< labels >>
flabel pwell s 0 0 288 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 288 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2_1
flabel metal1 s 0 617 288 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 288 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 288 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5696964
string GDS_START 5692300
<< end >>
