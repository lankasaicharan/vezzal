magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3506 1975
<< nwell >>
rect -38 332 2246 704
rect 496 313 1735 332
<< pwell >>
rect 1 49 2207 248
rect 0 0 2208 49
<< scpmos >>
rect 83 368 119 592
rect 183 368 219 592
rect 283 368 319 592
rect 373 368 409 592
rect 481 368 517 592
rect 582 349 618 573
rect 672 349 708 573
rect 772 349 808 573
rect 864 349 900 573
rect 954 349 990 573
rect 1078 349 1114 573
rect 1168 349 1204 573
rect 1258 349 1294 573
rect 1350 349 1386 573
rect 1440 349 1476 573
rect 1601 349 1637 573
rect 1819 424 1855 592
rect 1909 424 1945 592
rect 1999 424 2035 592
rect 2089 424 2125 592
<< nmoslvt >>
rect 98 74 128 222
rect 184 74 214 222
rect 289 74 319 222
rect 384 74 414 222
rect 492 74 522 222
rect 582 74 612 222
rect 678 74 708 222
rect 778 74 808 222
rect 864 74 894 222
rect 964 74 994 222
rect 1064 74 1094 222
rect 1162 74 1192 222
rect 1264 74 1294 222
rect 1350 74 1380 222
rect 1516 74 1546 222
rect 1607 74 1637 222
rect 1826 74 1856 222
rect 2094 74 2124 222
<< ndiff >>
rect 27 210 98 222
rect 27 176 39 210
rect 73 176 98 210
rect 27 120 98 176
rect 27 86 39 120
rect 73 86 98 120
rect 27 74 98 86
rect 128 210 184 222
rect 128 176 139 210
rect 173 176 184 210
rect 128 120 184 176
rect 128 86 139 120
rect 173 86 184 120
rect 128 74 184 86
rect 214 127 289 222
rect 214 93 239 127
rect 273 93 289 127
rect 214 74 289 93
rect 319 202 384 222
rect 319 168 339 202
rect 373 168 384 202
rect 319 120 384 168
rect 319 86 339 120
rect 373 86 384 120
rect 319 74 384 86
rect 414 127 492 222
rect 414 93 439 127
rect 473 93 492 127
rect 414 74 492 93
rect 522 201 582 222
rect 522 167 533 201
rect 567 167 582 201
rect 522 120 582 167
rect 522 86 533 120
rect 567 86 582 120
rect 522 74 582 86
rect 612 133 678 222
rect 612 99 633 133
rect 667 99 678 133
rect 612 74 678 99
rect 708 201 778 222
rect 708 167 719 201
rect 753 167 778 201
rect 708 120 778 167
rect 708 86 719 120
rect 753 86 778 120
rect 708 74 778 86
rect 808 133 864 222
rect 808 99 819 133
rect 853 99 864 133
rect 808 74 864 99
rect 894 201 964 222
rect 894 167 919 201
rect 953 167 964 201
rect 894 120 964 167
rect 894 86 919 120
rect 953 86 964 120
rect 894 74 964 86
rect 994 133 1064 222
rect 994 99 1019 133
rect 1053 99 1064 133
rect 994 74 1064 99
rect 1094 210 1162 222
rect 1094 176 1105 210
rect 1139 176 1162 210
rect 1094 120 1162 176
rect 1094 86 1105 120
rect 1139 86 1162 120
rect 1094 74 1162 86
rect 1192 210 1264 222
rect 1192 176 1205 210
rect 1239 176 1264 210
rect 1192 120 1264 176
rect 1192 86 1205 120
rect 1239 86 1264 120
rect 1192 74 1264 86
rect 1294 195 1350 222
rect 1294 161 1305 195
rect 1339 161 1350 195
rect 1294 120 1350 161
rect 1294 86 1305 120
rect 1339 86 1350 120
rect 1294 74 1350 86
rect 1380 120 1516 222
rect 1380 86 1391 120
rect 1425 86 1471 120
rect 1505 86 1516 120
rect 1380 74 1516 86
rect 1546 195 1607 222
rect 1546 161 1557 195
rect 1591 161 1607 195
rect 1546 120 1607 161
rect 1546 86 1557 120
rect 1591 86 1607 120
rect 1546 74 1607 86
rect 1637 120 1826 222
rect 1637 86 1648 120
rect 1682 86 1716 120
rect 1750 86 1826 120
rect 1637 74 1826 86
rect 1856 184 1913 222
rect 1856 150 1867 184
rect 1901 150 1913 184
rect 1856 74 1913 150
rect 2023 188 2094 222
rect 2023 154 2049 188
rect 2083 154 2094 188
rect 2023 120 2094 154
rect 2023 86 2049 120
rect 2083 86 2094 120
rect 2023 74 2094 86
rect 2124 210 2181 222
rect 2124 176 2135 210
rect 2169 176 2181 210
rect 2124 120 2181 176
rect 2124 86 2135 120
rect 2169 86 2181 120
rect 2124 74 2181 86
<< pdiff >>
rect 1005 615 1063 627
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 183 592
rect 119 546 139 580
rect 173 546 183 580
rect 119 512 183 546
rect 119 478 139 512
rect 173 478 183 512
rect 119 368 183 478
rect 219 580 283 592
rect 219 546 239 580
rect 273 546 283 580
rect 219 368 283 546
rect 319 580 373 592
rect 319 546 329 580
rect 363 546 373 580
rect 319 512 373 546
rect 319 478 329 512
rect 363 478 373 512
rect 319 368 373 478
rect 409 580 481 592
rect 409 546 433 580
rect 467 546 481 580
rect 409 368 481 546
rect 517 573 567 592
rect 1005 581 1017 615
rect 1051 581 1063 615
rect 1005 573 1063 581
rect 1753 580 1819 592
rect 517 528 582 573
rect 517 494 527 528
rect 561 494 582 528
rect 517 368 582 494
rect 532 349 582 368
rect 618 531 672 573
rect 618 497 628 531
rect 662 497 672 531
rect 618 463 672 497
rect 618 429 628 463
rect 662 429 672 463
rect 618 395 672 429
rect 618 361 628 395
rect 662 361 672 395
rect 618 349 672 361
rect 708 561 772 573
rect 708 527 728 561
rect 762 527 772 561
rect 708 469 772 527
rect 708 435 728 469
rect 762 435 772 469
rect 708 349 772 435
rect 808 561 864 573
rect 808 527 818 561
rect 852 527 864 561
rect 808 481 864 527
rect 808 447 818 481
rect 852 447 864 481
rect 808 401 864 447
rect 808 367 818 401
rect 852 367 864 401
rect 808 349 864 367
rect 900 531 954 573
rect 900 497 910 531
rect 944 497 954 531
rect 900 463 954 497
rect 900 429 910 463
rect 944 429 954 463
rect 900 395 954 429
rect 900 361 910 395
rect 944 361 954 395
rect 900 349 954 361
rect 990 349 1078 573
rect 1114 547 1168 573
rect 1114 513 1124 547
rect 1158 513 1168 547
rect 1114 349 1168 513
rect 1204 395 1258 573
rect 1204 361 1214 395
rect 1248 361 1258 395
rect 1204 349 1258 361
rect 1294 547 1350 573
rect 1294 513 1305 547
rect 1339 513 1350 547
rect 1294 349 1350 513
rect 1386 403 1440 573
rect 1386 369 1396 403
rect 1430 369 1440 403
rect 1386 349 1440 369
rect 1476 547 1601 573
rect 1476 513 1486 547
rect 1520 513 1557 547
rect 1591 513 1601 547
rect 1476 463 1601 513
rect 1476 429 1557 463
rect 1591 429 1601 463
rect 1476 349 1601 429
rect 1637 561 1699 573
rect 1637 527 1648 561
rect 1682 527 1699 561
rect 1637 463 1699 527
rect 1637 429 1648 463
rect 1682 429 1699 463
rect 1637 349 1699 429
rect 1753 546 1774 580
rect 1808 546 1819 580
rect 1753 508 1819 546
rect 1753 474 1774 508
rect 1808 474 1819 508
rect 1753 424 1819 474
rect 1855 580 1909 592
rect 1855 546 1865 580
rect 1899 546 1909 580
rect 1855 470 1909 546
rect 1855 436 1865 470
rect 1899 436 1909 470
rect 1855 424 1909 436
rect 1945 580 1999 592
rect 1945 546 1955 580
rect 1989 546 1999 580
rect 1945 470 1999 546
rect 1945 436 1955 470
rect 1989 436 1999 470
rect 1945 424 1999 436
rect 2035 580 2089 592
rect 2035 546 2045 580
rect 2079 546 2089 580
rect 2035 470 2089 546
rect 2035 436 2045 470
rect 2079 436 2089 470
rect 2035 424 2089 436
rect 2125 580 2181 592
rect 2125 546 2135 580
rect 2169 546 2181 580
rect 2125 496 2181 546
rect 2125 462 2135 496
rect 2169 462 2181 496
rect 2125 424 2181 462
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 176 173 210
rect 139 86 173 120
rect 239 93 273 127
rect 339 168 373 202
rect 339 86 373 120
rect 439 93 473 127
rect 533 167 567 201
rect 533 86 567 120
rect 633 99 667 133
rect 719 167 753 201
rect 719 86 753 120
rect 819 99 853 133
rect 919 167 953 201
rect 919 86 953 120
rect 1019 99 1053 133
rect 1105 176 1139 210
rect 1105 86 1139 120
rect 1205 176 1239 210
rect 1205 86 1239 120
rect 1305 161 1339 195
rect 1305 86 1339 120
rect 1391 86 1425 120
rect 1471 86 1505 120
rect 1557 161 1591 195
rect 1557 86 1591 120
rect 1648 86 1682 120
rect 1716 86 1750 120
rect 1867 150 1901 184
rect 2049 154 2083 188
rect 2049 86 2083 120
rect 2135 176 2169 210
rect 2135 86 2169 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 546 173 580
rect 139 478 173 512
rect 239 546 273 580
rect 329 546 363 580
rect 329 478 363 512
rect 433 546 467 580
rect 1017 581 1051 615
rect 527 494 561 528
rect 628 497 662 531
rect 628 429 662 463
rect 628 361 662 395
rect 728 527 762 561
rect 728 435 762 469
rect 818 527 852 561
rect 818 447 852 481
rect 818 367 852 401
rect 910 497 944 531
rect 910 429 944 463
rect 910 361 944 395
rect 1124 513 1158 547
rect 1214 361 1248 395
rect 1305 513 1339 547
rect 1396 369 1430 403
rect 1486 513 1520 547
rect 1557 513 1591 547
rect 1557 429 1591 463
rect 1648 527 1682 561
rect 1648 429 1682 463
rect 1774 546 1808 580
rect 1774 474 1808 508
rect 1865 546 1899 580
rect 1865 436 1899 470
rect 1955 546 1989 580
rect 1955 436 1989 470
rect 2045 546 2079 580
rect 2045 436 2079 470
rect 2135 546 2169 580
rect 2135 462 2169 496
<< poly >>
rect 83 592 119 618
rect 183 592 219 618
rect 283 592 319 618
rect 373 592 409 618
rect 481 592 517 618
rect 582 573 618 599
rect 672 573 708 599
rect 772 573 808 599
rect 864 573 900 599
rect 954 573 990 599
rect 1078 573 1114 599
rect 1168 573 1204 599
rect 1258 573 1294 599
rect 1350 573 1386 599
rect 1440 573 1476 599
rect 1601 573 1637 599
rect 1819 592 1855 618
rect 1909 592 1945 618
rect 1999 592 2035 618
rect 2089 592 2125 618
rect 83 330 119 368
rect 53 314 119 330
rect 53 280 69 314
rect 103 294 119 314
rect 183 310 219 368
rect 283 310 319 368
rect 373 310 409 368
rect 481 310 517 368
rect 1819 372 1855 424
rect 1909 372 1945 424
rect 1819 356 1945 372
rect 582 317 618 349
rect 672 317 708 349
rect 772 317 808 349
rect 183 294 522 310
rect 103 280 128 294
rect 183 280 313 294
rect 53 264 128 280
rect 98 222 128 264
rect 184 260 313 280
rect 347 260 381 294
rect 415 260 449 294
rect 483 260 522 294
rect 184 244 522 260
rect 184 222 214 244
rect 289 222 319 244
rect 384 222 414 244
rect 492 222 522 244
rect 582 301 808 317
rect 582 267 598 301
rect 632 267 666 301
rect 700 267 734 301
rect 768 267 808 301
rect 582 251 808 267
rect 582 222 612 251
rect 678 222 708 251
rect 778 222 808 251
rect 864 317 900 349
rect 954 317 990 349
rect 1078 317 1114 349
rect 864 301 1114 317
rect 864 267 885 301
rect 919 267 953 301
rect 987 267 1021 301
rect 1055 267 1114 301
rect 1168 281 1204 349
rect 1258 281 1294 349
rect 1350 311 1386 349
rect 1440 311 1476 349
rect 1350 295 1559 311
rect 1350 281 1373 295
rect 864 251 1114 267
rect 1162 261 1373 281
rect 1407 261 1441 295
rect 1475 261 1509 295
rect 1543 261 1559 295
rect 1162 251 1559 261
rect 864 222 894 251
rect 964 222 994 251
rect 1064 222 1094 251
rect 1162 222 1192 251
rect 1264 222 1294 251
rect 1350 245 1559 251
rect 1601 307 1637 349
rect 1819 322 1835 356
rect 1869 342 1945 356
rect 1999 356 2035 424
rect 2089 356 2125 424
rect 1869 322 1885 342
rect 1709 307 1775 310
rect 1601 294 1775 307
rect 1819 306 1885 322
rect 1999 340 2125 356
rect 1999 306 2041 340
rect 2075 326 2125 340
rect 2075 306 2124 326
rect 1601 260 1725 294
rect 1759 260 1775 294
rect 1350 222 1380 245
rect 1516 222 1546 245
rect 1601 244 1775 260
rect 1607 222 1637 244
rect 1826 222 1856 306
rect 1999 290 2124 306
rect 2094 222 2124 290
rect 98 48 128 74
rect 184 48 214 74
rect 289 48 319 74
rect 384 48 414 74
rect 492 48 522 74
rect 582 48 612 74
rect 678 48 708 74
rect 778 48 808 74
rect 864 48 894 74
rect 964 48 994 74
rect 1064 48 1094 74
rect 1162 48 1192 74
rect 1264 48 1294 74
rect 1350 48 1380 74
rect 1516 48 1546 74
rect 1607 48 1637 74
rect 1826 48 1856 74
rect 2094 48 2124 74
<< polycont >>
rect 69 280 103 314
rect 313 260 347 294
rect 381 260 415 294
rect 449 260 483 294
rect 598 267 632 301
rect 666 267 700 301
rect 734 267 768 301
rect 885 267 919 301
rect 953 267 987 301
rect 1021 267 1055 301
rect 1373 261 1407 295
rect 1441 261 1475 295
rect 1509 261 1543 295
rect 1835 322 1869 356
rect 2041 306 2075 340
rect 1725 260 1759 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 497 89 546
rect 23 463 39 497
rect 73 463 89 497
rect 123 580 189 596
rect 123 546 139 580
rect 173 546 189 580
rect 223 580 289 649
rect 223 546 239 580
rect 273 546 289 580
rect 329 580 379 596
rect 363 546 379 580
rect 413 580 487 649
rect 413 546 433 580
rect 467 546 487 580
rect 527 581 778 615
rect 123 512 189 546
rect 329 512 379 546
rect 527 528 577 581
rect 712 561 778 581
rect 123 478 139 512
rect 173 478 329 512
rect 363 494 527 512
rect 561 494 577 528
rect 363 478 577 494
rect 612 531 678 547
rect 612 497 628 531
rect 662 497 678 531
rect 23 444 89 463
rect 612 463 678 497
rect 612 444 628 463
rect 23 429 628 444
rect 662 429 678 463
rect 23 414 678 429
rect 712 527 728 561
rect 762 527 778 561
rect 712 469 778 527
rect 712 435 728 469
rect 762 435 778 469
rect 712 419 778 435
rect 818 581 1017 615
rect 1051 581 1698 615
rect 818 561 852 581
rect 1641 561 1698 581
rect 818 481 852 527
rect 23 380 39 414
rect 73 410 678 414
rect 73 380 89 410
rect 23 364 89 380
rect 612 395 678 410
rect 217 342 578 376
rect 612 361 628 395
rect 662 385 678 395
rect 818 401 852 447
rect 662 367 818 385
rect 662 361 852 367
rect 612 351 852 361
rect 894 531 1124 547
rect 894 497 910 531
rect 944 513 1124 531
rect 1158 513 1305 547
rect 1339 513 1486 547
rect 1520 513 1557 547
rect 1591 513 1607 547
rect 944 497 960 513
rect 894 463 960 497
rect 894 429 910 463
rect 944 429 960 463
rect 894 395 960 429
rect 894 361 910 395
rect 944 361 960 395
rect 894 351 960 361
rect 1037 445 1514 479
rect 217 330 263 342
rect 53 314 263 330
rect 53 280 69 314
rect 103 280 263 314
rect 544 317 578 342
rect 1037 317 1071 445
rect 53 264 263 280
rect 297 294 499 308
rect 297 260 313 294
rect 347 260 381 294
rect 415 260 449 294
rect 483 260 499 294
rect 297 236 499 260
rect 544 301 784 317
rect 544 267 598 301
rect 632 267 666 301
rect 700 267 734 301
rect 768 267 784 301
rect 544 251 784 267
rect 869 301 1071 317
rect 869 267 885 301
rect 919 267 953 301
rect 987 267 1021 301
rect 1055 267 1071 301
rect 1198 403 1446 411
rect 1198 395 1396 403
rect 1198 361 1214 395
rect 1248 369 1396 395
rect 1430 369 1446 403
rect 1248 361 1446 369
rect 1198 345 1446 361
rect 1480 379 1514 445
rect 1552 463 1607 513
rect 1552 429 1557 463
rect 1591 429 1607 463
rect 1552 413 1607 429
rect 1641 527 1648 561
rect 1682 527 1698 561
rect 1641 463 1698 527
rect 1758 580 1824 649
rect 1758 546 1774 580
rect 1808 546 1824 580
rect 1758 508 1824 546
rect 1758 474 1774 508
rect 1808 474 1824 508
rect 1860 580 1915 596
rect 1860 546 1865 580
rect 1899 546 1915 580
rect 1641 429 1648 463
rect 1682 429 1698 463
rect 1860 470 1915 546
rect 1860 440 1865 470
rect 1641 413 1698 429
rect 1741 436 1865 440
rect 1899 436 1915 470
rect 1741 406 1915 436
rect 1955 580 1989 649
rect 1955 470 1989 546
rect 1955 420 1989 436
rect 2029 580 2079 596
rect 2029 546 2045 580
rect 2029 470 2079 546
rect 2029 436 2045 470
rect 2119 580 2185 649
rect 2119 546 2135 580
rect 2169 546 2185 580
rect 2119 496 2185 546
rect 2119 462 2135 496
rect 2169 462 2185 496
rect 2119 458 2185 462
rect 2029 424 2079 436
rect 1741 379 1775 406
rect 2029 390 2185 424
rect 1480 345 1775 379
rect 1198 294 1264 345
rect 1357 295 1675 311
rect 869 251 1071 267
rect 1105 260 1323 294
rect 23 210 89 226
rect 23 176 39 210
rect 73 176 89 210
rect 23 120 89 176
rect 23 86 39 120
rect 73 86 89 120
rect 23 17 89 86
rect 123 210 189 226
rect 1105 217 1155 260
rect 123 176 139 210
rect 173 202 189 210
rect 533 210 1155 217
rect 533 202 1105 210
rect 173 176 339 202
rect 123 168 339 176
rect 373 201 1105 202
rect 373 168 533 201
rect 123 120 189 168
rect 123 86 139 120
rect 173 86 189 120
rect 123 70 189 86
rect 223 127 289 134
rect 223 93 239 127
rect 273 93 289 127
rect 223 17 289 93
rect 323 120 389 168
rect 567 183 719 201
rect 567 167 583 183
rect 323 86 339 120
rect 373 86 389 120
rect 323 70 389 86
rect 423 127 489 134
rect 423 93 439 127
rect 473 93 489 127
rect 423 17 489 93
rect 533 120 583 167
rect 753 183 919 201
rect 753 167 769 183
rect 567 86 583 120
rect 533 70 583 86
rect 617 133 683 149
rect 617 99 633 133
rect 667 99 683 133
rect 617 17 683 99
rect 719 120 769 167
rect 903 167 919 183
rect 953 183 1105 201
rect 953 167 969 183
rect 753 86 769 120
rect 719 70 769 86
rect 803 133 869 149
rect 803 99 819 133
rect 853 99 869 133
rect 803 17 869 99
rect 903 120 969 167
rect 1139 176 1155 210
rect 903 86 919 120
rect 953 86 969 120
rect 903 70 969 86
rect 1003 133 1069 149
rect 1003 99 1019 133
rect 1053 99 1069 133
rect 1003 17 1069 99
rect 1105 120 1155 176
rect 1139 86 1155 120
rect 1105 70 1155 86
rect 1189 210 1255 226
rect 1189 176 1205 210
rect 1239 176 1255 210
rect 1189 120 1255 176
rect 1189 86 1205 120
rect 1239 86 1255 120
rect 1189 17 1255 86
rect 1289 211 1323 260
rect 1357 261 1373 295
rect 1407 261 1441 295
rect 1475 261 1509 295
rect 1543 261 1675 295
rect 1357 245 1675 261
rect 1289 195 1607 211
rect 1289 161 1305 195
rect 1339 177 1557 195
rect 1339 161 1355 177
rect 1289 120 1355 161
rect 1541 161 1557 177
rect 1591 161 1607 195
rect 1641 204 1675 245
rect 1709 294 1775 345
rect 1819 356 1991 372
rect 1819 322 1835 356
rect 1869 322 1991 356
rect 1819 306 1991 322
rect 2025 340 2091 356
rect 2025 306 2041 340
rect 2075 306 2091 340
rect 1709 260 1725 294
rect 1759 272 1775 294
rect 2025 290 2091 306
rect 1759 260 1917 272
rect 1709 238 1917 260
rect 2151 256 2185 390
rect 1641 170 1818 204
rect 1289 86 1305 120
rect 1339 86 1355 120
rect 1289 70 1355 86
rect 1389 120 1507 136
rect 1389 86 1391 120
rect 1425 86 1471 120
rect 1505 86 1507 120
rect 1389 17 1507 86
rect 1541 120 1607 161
rect 1541 86 1557 120
rect 1591 86 1607 120
rect 1541 70 1607 86
rect 1641 120 1750 136
rect 1641 86 1648 120
rect 1682 86 1716 120
rect 1641 17 1750 86
rect 1784 85 1818 170
rect 1852 184 1917 238
rect 1852 150 1867 184
rect 1901 150 1917 184
rect 1852 134 1917 150
rect 1951 222 2185 256
rect 1951 85 1985 222
rect 2133 210 2185 222
rect 1784 51 1985 85
rect 2019 154 2049 188
rect 2083 154 2099 188
rect 2019 120 2099 154
rect 2019 86 2049 120
rect 2083 86 2099 120
rect 2019 17 2099 86
rect 2133 176 2135 210
rect 2169 176 2185 210
rect 2133 120 2185 176
rect 2133 86 2135 120
rect 2169 86 2185 120
rect 2133 70 2185 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4bb_4
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1567 94 1601 128 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1567 168 1601 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 1309274
string GDS_START 1293910
<< end >>
