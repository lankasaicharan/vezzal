magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 1 49 863 241
rect 0 0 864 49
<< scnmos >>
rect 80 131 110 215
rect 178 47 208 215
rect 368 131 398 215
rect 466 47 496 215
rect 656 131 686 215
rect 754 47 784 215
<< scpmoshvt >>
rect 80 367 110 451
rect 178 367 208 619
rect 368 367 398 451
rect 466 367 496 619
rect 656 367 686 451
rect 754 367 784 619
<< ndiff >>
rect 27 190 80 215
rect 27 156 35 190
rect 69 156 80 190
rect 27 131 80 156
rect 110 161 178 215
rect 110 131 133 161
rect 125 127 133 131
rect 167 127 178 161
rect 125 93 178 127
rect 125 59 133 93
rect 167 59 178 93
rect 125 47 178 59
rect 208 199 261 215
rect 208 165 219 199
rect 253 165 261 199
rect 208 101 261 165
rect 315 190 368 215
rect 315 156 323 190
rect 357 156 368 190
rect 315 131 368 156
rect 398 161 466 215
rect 398 131 421 161
rect 413 127 421 131
rect 455 127 466 161
rect 208 67 219 101
rect 253 67 261 101
rect 208 47 261 67
rect 413 93 466 127
rect 413 59 421 93
rect 455 59 466 93
rect 413 47 466 59
rect 496 199 549 215
rect 496 165 507 199
rect 541 165 549 199
rect 496 101 549 165
rect 603 190 656 215
rect 603 156 611 190
rect 645 156 656 190
rect 603 131 656 156
rect 686 161 754 215
rect 686 131 709 161
rect 701 127 709 131
rect 743 127 754 161
rect 496 67 507 101
rect 541 67 549 101
rect 496 47 549 67
rect 701 93 754 127
rect 701 59 709 93
rect 743 59 754 93
rect 701 47 754 59
rect 784 199 837 215
rect 784 165 795 199
rect 829 165 837 199
rect 784 101 837 165
rect 784 67 795 101
rect 829 67 837 101
rect 784 47 837 67
<< pdiff >>
rect 125 607 178 619
rect 125 573 133 607
rect 167 573 178 607
rect 125 516 178 573
rect 125 482 133 516
rect 167 482 178 516
rect 125 451 178 482
rect 27 429 80 451
rect 27 395 35 429
rect 69 395 80 429
rect 27 367 80 395
rect 110 367 178 451
rect 208 599 261 619
rect 208 565 219 599
rect 253 565 261 599
rect 208 510 261 565
rect 208 476 219 510
rect 253 476 261 510
rect 413 607 466 619
rect 413 573 421 607
rect 455 573 466 607
rect 413 516 466 573
rect 413 482 421 516
rect 455 482 466 516
rect 208 417 261 476
rect 413 451 466 482
rect 208 383 219 417
rect 253 383 261 417
rect 208 367 261 383
rect 315 429 368 451
rect 315 395 323 429
rect 357 395 368 429
rect 315 367 368 395
rect 398 367 466 451
rect 496 599 549 619
rect 496 565 507 599
rect 541 565 549 599
rect 496 510 549 565
rect 496 476 507 510
rect 541 476 549 510
rect 701 607 754 619
rect 701 573 709 607
rect 743 573 754 607
rect 701 516 754 573
rect 701 482 709 516
rect 743 482 754 516
rect 496 417 549 476
rect 701 451 754 482
rect 496 383 507 417
rect 541 383 549 417
rect 496 367 549 383
rect 603 429 656 451
rect 603 395 611 429
rect 645 395 656 429
rect 603 367 656 395
rect 686 367 754 451
rect 784 599 837 619
rect 784 565 795 599
rect 829 565 837 599
rect 784 510 837 565
rect 784 476 795 510
rect 829 476 837 510
rect 784 417 837 476
rect 784 383 795 417
rect 829 383 837 417
rect 784 367 837 383
<< ndiffc >>
rect 35 156 69 190
rect 133 127 167 161
rect 133 59 167 93
rect 219 165 253 199
rect 323 156 357 190
rect 421 127 455 161
rect 219 67 253 101
rect 421 59 455 93
rect 507 165 541 199
rect 611 156 645 190
rect 709 127 743 161
rect 507 67 541 101
rect 709 59 743 93
rect 795 165 829 199
rect 795 67 829 101
<< pdiffc >>
rect 133 573 167 607
rect 133 482 167 516
rect 35 395 69 429
rect 219 565 253 599
rect 219 476 253 510
rect 421 573 455 607
rect 421 482 455 516
rect 219 383 253 417
rect 323 395 357 429
rect 507 565 541 599
rect 507 476 541 510
rect 709 573 743 607
rect 709 482 743 516
rect 507 383 541 417
rect 611 395 645 429
rect 795 565 829 599
rect 795 476 829 510
rect 795 383 829 417
<< poly >>
rect 178 619 208 645
rect 466 619 496 645
rect 754 619 784 645
rect 80 451 110 477
rect 368 451 398 477
rect 656 451 686 477
rect 80 321 110 367
rect 178 321 208 367
rect 368 321 398 367
rect 466 321 496 367
rect 656 321 686 367
rect 754 321 784 367
rect 44 305 110 321
rect 44 271 60 305
rect 94 271 110 305
rect 44 255 110 271
rect 80 215 110 255
rect 152 305 218 321
rect 152 271 168 305
rect 202 271 218 305
rect 152 252 218 271
rect 332 305 398 321
rect 332 271 348 305
rect 382 271 398 305
rect 332 255 398 271
rect 178 215 208 252
rect 368 215 398 255
rect 440 305 506 321
rect 440 271 456 305
rect 490 271 506 305
rect 440 252 506 271
rect 620 305 686 321
rect 620 271 636 305
rect 670 271 686 305
rect 620 255 686 271
rect 466 215 496 252
rect 656 215 686 255
rect 728 305 794 321
rect 728 271 744 305
rect 778 271 794 305
rect 728 252 794 271
rect 754 215 784 252
rect 80 105 110 131
rect 368 105 398 131
rect 656 105 686 131
rect 178 21 208 47
rect 466 21 496 47
rect 754 21 784 47
<< polycont >>
rect 60 271 94 305
rect 168 271 202 305
rect 348 271 382 305
rect 456 271 490 305
rect 636 271 670 305
rect 744 271 778 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 117 607 176 649
rect 117 573 133 607
rect 167 573 176 607
rect 117 516 176 573
rect 117 482 133 516
rect 167 482 176 516
rect 117 466 176 482
rect 212 599 270 615
rect 212 565 219 599
rect 253 565 270 599
rect 212 510 270 565
rect 212 476 219 510
rect 253 476 270 510
rect 19 432 85 445
rect 19 429 178 432
rect 19 395 35 429
rect 69 395 178 429
rect 19 387 178 395
rect 20 305 110 353
rect 20 271 60 305
rect 94 271 110 305
rect 20 263 110 271
rect 144 321 178 387
rect 212 424 270 476
rect 405 607 464 649
rect 405 573 421 607
rect 455 573 464 607
rect 405 516 464 573
rect 405 482 421 516
rect 455 482 464 516
rect 405 466 464 482
rect 500 599 558 615
rect 500 565 507 599
rect 541 565 558 599
rect 500 510 558 565
rect 500 476 507 510
rect 541 476 558 510
rect 212 383 219 424
rect 253 383 270 424
rect 212 367 270 383
rect 307 432 373 445
rect 307 429 466 432
rect 307 395 323 429
rect 357 395 466 429
rect 307 379 466 395
rect 236 321 270 367
rect 432 321 466 379
rect 500 424 558 476
rect 693 607 752 649
rect 693 573 709 607
rect 743 573 752 607
rect 693 516 752 573
rect 693 482 709 516
rect 743 482 752 516
rect 693 466 752 482
rect 788 599 847 615
rect 788 565 795 599
rect 829 565 847 599
rect 788 510 847 565
rect 788 476 795 510
rect 829 476 847 510
rect 500 383 507 424
rect 541 383 558 424
rect 500 367 558 383
rect 595 432 661 445
rect 595 429 754 432
rect 595 395 611 429
rect 645 395 754 429
rect 595 379 754 395
rect 524 321 558 367
rect 720 321 754 379
rect 788 424 847 476
rect 788 383 795 424
rect 829 383 847 424
rect 788 367 847 383
rect 144 305 202 321
rect 144 271 168 305
rect 144 255 202 271
rect 236 305 398 321
rect 236 271 348 305
rect 382 271 398 305
rect 236 263 398 271
rect 432 305 490 321
rect 432 271 456 305
rect 144 229 178 255
rect 19 195 178 229
rect 236 215 270 263
rect 432 255 490 271
rect 524 305 686 321
rect 524 271 636 305
rect 670 271 686 305
rect 524 263 686 271
rect 720 305 778 321
rect 720 271 744 305
rect 432 229 466 255
rect 217 199 270 215
rect 19 190 78 195
rect 19 156 35 190
rect 69 156 78 190
rect 217 165 219 199
rect 253 165 270 199
rect 19 140 78 156
rect 117 127 133 161
rect 167 127 183 161
rect 117 93 183 127
rect 117 59 133 93
rect 167 59 183 93
rect 117 17 183 59
rect 217 101 270 165
rect 307 195 466 229
rect 524 215 558 263
rect 720 255 778 271
rect 720 229 754 255
rect 505 199 558 215
rect 307 190 366 195
rect 307 156 323 190
rect 357 156 366 190
rect 505 165 507 199
rect 541 165 558 199
rect 307 140 366 156
rect 217 67 219 101
rect 253 67 270 101
rect 217 51 270 67
rect 405 127 421 161
rect 455 127 471 161
rect 405 93 471 127
rect 405 59 421 93
rect 455 59 471 93
rect 405 17 471 59
rect 505 101 558 165
rect 595 195 754 229
rect 812 215 847 367
rect 793 199 847 215
rect 595 190 654 195
rect 595 156 611 190
rect 645 156 654 190
rect 793 165 795 199
rect 829 165 847 199
rect 595 140 654 156
rect 505 67 507 101
rect 541 67 558 101
rect 505 51 558 67
rect 693 127 709 161
rect 743 127 759 161
rect 693 93 759 127
rect 693 59 709 93
rect 743 59 759 93
rect 693 17 759 59
rect 793 101 847 165
rect 793 67 795 101
rect 829 67 847 101
rect 793 51 847 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 219 417 253 424
rect 219 390 253 417
rect 507 417 541 424
rect 507 390 541 417
rect 795 417 829 424
rect 795 390 829 417
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 192 464 841 498
rect 192 424 265 430
rect 192 390 219 424
rect 253 390 265 424
rect 192 384 265 390
rect 480 424 553 430
rect 480 390 507 424
rect 541 390 553 424
rect 480 384 553 390
rect 768 424 841 464
rect 768 390 795 424
rect 829 390 841 424
rect 768 384 841 390
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlymetal6s6s_1
flabel metal1 s 192 464 841 498 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4582924
string GDS_START 4575084
<< end >>
