magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -2403 -11413 16394 11152
<< dnwell >>
rect 13147 4289 13273 4326
rect 13147 3073 15054 4289
rect 13147 -56 15031 3073
<< nwell >>
rect 13067 8723 15134 8773
rect 1099 7312 4519 8647
rect 1099 7164 4511 7312
rect 14947 4339 15053 4362
rect 14825 4326 15053 4339
rect -238 1344 1092 1944
rect 13067 2949 13353 4326
rect 14825 2949 15134 4326
rect 13067 2779 15134 2949
rect 13067 150 13353 2779
rect 14825 150 15134 2779
rect 13067 -136 15134 150
<< pwell >>
rect 774 8731 4799 8817
rect 774 7104 860 8731
rect 774 7018 4757 7104
rect -900 6062 951 6792
rect 4385 5805 4757 7018
rect 4041 4242 4757 5805
rect 4041 4042 8318 4242
rect 4041 3951 9482 4042
rect 3838 3646 9482 3951
rect 3838 -22 4966 3646
rect 11483 2718 12391 3070
rect 11815 2176 12391 2718
rect 13413 4113 14641 4199
rect 13413 3347 14605 4113
rect 13413 3208 14606 3347
rect 13526 3009 14606 3208
rect 5273 819 8672 1119
rect 8011 -70 10609 -36
rect 11288 -70 12864 905
rect 7537 -102 12864 -70
rect 5709 -241 12864 -102
rect 13413 210 14765 2718
rect 12251 -1021 12823 -241
<< mvnmos >>
rect 13603 3415 13703 4015
rect 13875 3415 13975 4015
rect 14151 3415 14251 4015
rect 14423 3415 14523 4015
rect 13608 3237 13708 3321
rect 13880 3237 13980 3321
rect 14152 3237 14252 3321
rect 14424 3237 14524 3321
rect 13608 3035 13708 3119
rect 13880 3035 13980 3119
rect 14152 3035 14252 3119
rect 14424 3035 14524 3119
rect 13630 2428 14630 2528
rect 13630 2272 14630 2372
rect 13630 2116 14630 2216
rect 13630 1960 14630 2060
rect 13630 1804 14630 1904
rect 13630 1648 14630 1748
rect 13630 1492 14630 1592
rect 13630 1336 14630 1436
rect 13630 1180 14630 1280
rect 13630 1024 14630 1124
rect 13630 868 14630 968
rect 13630 712 14630 812
rect 13630 556 14630 656
rect 13630 400 14630 500
<< mvpmos >>
rect 1282 8327 4282 8427
rect 1282 8171 4282 8271
rect 1282 8015 4282 8115
rect 1282 7859 4282 7959
rect 1282 7703 4282 7803
rect 1282 7547 4282 7647
rect 1282 7391 4282 7491
<< mvndiff >>
rect 13547 3937 13603 4015
rect 13547 3903 13558 3937
rect 13592 3903 13603 3937
rect 13547 3869 13603 3903
rect 13547 3835 13558 3869
rect 13592 3835 13603 3869
rect 13547 3801 13603 3835
rect 13547 3767 13558 3801
rect 13592 3767 13603 3801
rect 13547 3733 13603 3767
rect 13547 3699 13558 3733
rect 13592 3699 13603 3733
rect 13547 3665 13603 3699
rect 13547 3631 13558 3665
rect 13592 3631 13603 3665
rect 13547 3597 13603 3631
rect 13547 3563 13558 3597
rect 13592 3563 13603 3597
rect 13547 3529 13603 3563
rect 13547 3495 13558 3529
rect 13592 3495 13603 3529
rect 13547 3461 13603 3495
rect 13547 3427 13558 3461
rect 13592 3427 13603 3461
rect 13547 3415 13603 3427
rect 13703 3937 13759 4015
rect 13703 3903 13714 3937
rect 13748 3903 13759 3937
rect 13703 3869 13759 3903
rect 13703 3835 13714 3869
rect 13748 3835 13759 3869
rect 13703 3801 13759 3835
rect 13703 3767 13714 3801
rect 13748 3767 13759 3801
rect 13703 3733 13759 3767
rect 13703 3699 13714 3733
rect 13748 3699 13759 3733
rect 13703 3665 13759 3699
rect 13703 3631 13714 3665
rect 13748 3631 13759 3665
rect 13703 3597 13759 3631
rect 13703 3563 13714 3597
rect 13748 3563 13759 3597
rect 13703 3529 13759 3563
rect 13703 3495 13714 3529
rect 13748 3495 13759 3529
rect 13703 3461 13759 3495
rect 13703 3427 13714 3461
rect 13748 3427 13759 3461
rect 13703 3415 13759 3427
rect 13819 3937 13875 4015
rect 13819 3903 13830 3937
rect 13864 3903 13875 3937
rect 13819 3869 13875 3903
rect 13819 3835 13830 3869
rect 13864 3835 13875 3869
rect 13819 3801 13875 3835
rect 13819 3767 13830 3801
rect 13864 3767 13875 3801
rect 13819 3733 13875 3767
rect 13819 3699 13830 3733
rect 13864 3699 13875 3733
rect 13819 3665 13875 3699
rect 13819 3631 13830 3665
rect 13864 3631 13875 3665
rect 13819 3597 13875 3631
rect 13819 3563 13830 3597
rect 13864 3563 13875 3597
rect 13819 3529 13875 3563
rect 13819 3495 13830 3529
rect 13864 3495 13875 3529
rect 13819 3461 13875 3495
rect 13819 3427 13830 3461
rect 13864 3427 13875 3461
rect 13819 3415 13875 3427
rect 13975 3937 14031 4015
rect 13975 3903 13986 3937
rect 14020 3903 14031 3937
rect 13975 3869 14031 3903
rect 13975 3835 13986 3869
rect 14020 3835 14031 3869
rect 13975 3801 14031 3835
rect 13975 3767 13986 3801
rect 14020 3767 14031 3801
rect 13975 3733 14031 3767
rect 13975 3699 13986 3733
rect 14020 3699 14031 3733
rect 13975 3665 14031 3699
rect 13975 3631 13986 3665
rect 14020 3631 14031 3665
rect 13975 3597 14031 3631
rect 13975 3563 13986 3597
rect 14020 3563 14031 3597
rect 13975 3529 14031 3563
rect 13975 3495 13986 3529
rect 14020 3495 14031 3529
rect 13975 3461 14031 3495
rect 13975 3427 13986 3461
rect 14020 3427 14031 3461
rect 13975 3415 14031 3427
rect 14095 3937 14151 4015
rect 14095 3903 14106 3937
rect 14140 3903 14151 3937
rect 14095 3869 14151 3903
rect 14095 3835 14106 3869
rect 14140 3835 14151 3869
rect 14095 3801 14151 3835
rect 14095 3767 14106 3801
rect 14140 3767 14151 3801
rect 14095 3733 14151 3767
rect 14095 3699 14106 3733
rect 14140 3699 14151 3733
rect 14095 3665 14151 3699
rect 14095 3631 14106 3665
rect 14140 3631 14151 3665
rect 14095 3597 14151 3631
rect 14095 3563 14106 3597
rect 14140 3563 14151 3597
rect 14095 3529 14151 3563
rect 14095 3495 14106 3529
rect 14140 3495 14151 3529
rect 14095 3461 14151 3495
rect 14095 3427 14106 3461
rect 14140 3427 14151 3461
rect 14095 3415 14151 3427
rect 14251 3937 14307 4015
rect 14251 3903 14262 3937
rect 14296 3903 14307 3937
rect 14251 3869 14307 3903
rect 14251 3835 14262 3869
rect 14296 3835 14307 3869
rect 14251 3801 14307 3835
rect 14251 3767 14262 3801
rect 14296 3767 14307 3801
rect 14251 3733 14307 3767
rect 14251 3699 14262 3733
rect 14296 3699 14307 3733
rect 14251 3665 14307 3699
rect 14251 3631 14262 3665
rect 14296 3631 14307 3665
rect 14251 3597 14307 3631
rect 14251 3563 14262 3597
rect 14296 3563 14307 3597
rect 14251 3529 14307 3563
rect 14251 3495 14262 3529
rect 14296 3495 14307 3529
rect 14251 3461 14307 3495
rect 14251 3427 14262 3461
rect 14296 3427 14307 3461
rect 14251 3415 14307 3427
rect 14367 3937 14423 4015
rect 14367 3903 14378 3937
rect 14412 3903 14423 3937
rect 14367 3869 14423 3903
rect 14367 3835 14378 3869
rect 14412 3835 14423 3869
rect 14367 3801 14423 3835
rect 14367 3767 14378 3801
rect 14412 3767 14423 3801
rect 14367 3733 14423 3767
rect 14367 3699 14378 3733
rect 14412 3699 14423 3733
rect 14367 3665 14423 3699
rect 14367 3631 14378 3665
rect 14412 3631 14423 3665
rect 14367 3597 14423 3631
rect 14367 3563 14378 3597
rect 14412 3563 14423 3597
rect 14367 3529 14423 3563
rect 14367 3495 14378 3529
rect 14412 3495 14423 3529
rect 14367 3461 14423 3495
rect 14367 3427 14378 3461
rect 14412 3427 14423 3461
rect 14367 3415 14423 3427
rect 14523 3937 14579 4015
rect 14523 3903 14534 3937
rect 14568 3903 14579 3937
rect 14523 3869 14579 3903
rect 14523 3835 14534 3869
rect 14568 3835 14579 3869
rect 14523 3801 14579 3835
rect 14523 3767 14534 3801
rect 14568 3767 14579 3801
rect 14523 3733 14579 3767
rect 14523 3699 14534 3733
rect 14568 3699 14579 3733
rect 14523 3665 14579 3699
rect 14523 3631 14534 3665
rect 14568 3631 14579 3665
rect 14523 3597 14579 3631
rect 14523 3563 14534 3597
rect 14568 3563 14579 3597
rect 14523 3529 14579 3563
rect 14523 3495 14534 3529
rect 14568 3495 14579 3529
rect 14523 3461 14579 3495
rect 14523 3427 14534 3461
rect 14568 3427 14579 3461
rect 14523 3415 14579 3427
rect 13552 3309 13608 3321
rect 13552 3275 13563 3309
rect 13597 3275 13608 3309
rect 13552 3237 13608 3275
rect 13708 3309 13764 3321
rect 13708 3275 13719 3309
rect 13753 3275 13764 3309
rect 13708 3237 13764 3275
rect 13824 3309 13880 3321
rect 13824 3275 13835 3309
rect 13869 3275 13880 3309
rect 13824 3237 13880 3275
rect 13980 3309 14036 3321
rect 13980 3275 13991 3309
rect 14025 3275 14036 3309
rect 13980 3237 14036 3275
rect 14096 3309 14152 3321
rect 14096 3275 14107 3309
rect 14141 3275 14152 3309
rect 14096 3237 14152 3275
rect 14252 3309 14308 3321
rect 14252 3275 14263 3309
rect 14297 3275 14308 3309
rect 14252 3237 14308 3275
rect 14368 3309 14424 3321
rect 14368 3275 14379 3309
rect 14413 3275 14424 3309
rect 14368 3237 14424 3275
rect 14524 3309 14580 3321
rect 14524 3275 14535 3309
rect 14569 3275 14580 3309
rect 14524 3237 14580 3275
rect 13552 3081 13608 3119
rect 13552 3047 13563 3081
rect 13597 3047 13608 3081
rect 13552 3035 13608 3047
rect 13708 3081 13764 3119
rect 13708 3047 13719 3081
rect 13753 3047 13764 3081
rect 13708 3035 13764 3047
rect 13824 3081 13880 3119
rect 13824 3047 13835 3081
rect 13869 3047 13880 3081
rect 13824 3035 13880 3047
rect 13980 3081 14036 3119
rect 13980 3047 13991 3081
rect 14025 3047 14036 3081
rect 13980 3035 14036 3047
rect 14096 3081 14152 3119
rect 14096 3047 14107 3081
rect 14141 3047 14152 3081
rect 14096 3035 14152 3047
rect 14252 3081 14308 3119
rect 14252 3047 14263 3081
rect 14297 3047 14308 3081
rect 14252 3035 14308 3047
rect 14368 3081 14424 3119
rect 14368 3047 14379 3081
rect 14413 3047 14424 3081
rect 14368 3035 14424 3047
rect 14524 3081 14580 3119
rect 14524 3047 14535 3081
rect 14569 3047 14580 3081
rect 14524 3035 14580 3047
rect 13630 2573 14630 2584
rect 13630 2539 13700 2573
rect 13734 2539 13768 2573
rect 13802 2539 13836 2573
rect 13870 2539 13904 2573
rect 13938 2539 13972 2573
rect 14006 2539 14040 2573
rect 14074 2539 14108 2573
rect 14142 2539 14176 2573
rect 14210 2539 14244 2573
rect 14278 2539 14312 2573
rect 14346 2539 14380 2573
rect 14414 2539 14448 2573
rect 14482 2539 14516 2573
rect 14550 2539 14584 2573
rect 14618 2539 14630 2573
rect 13630 2528 14630 2539
rect 13630 2417 14630 2428
rect 13630 2383 13700 2417
rect 13734 2383 13768 2417
rect 13802 2383 13836 2417
rect 13870 2383 13904 2417
rect 13938 2383 13972 2417
rect 14006 2383 14040 2417
rect 14074 2383 14108 2417
rect 14142 2383 14176 2417
rect 14210 2383 14244 2417
rect 14278 2383 14312 2417
rect 14346 2383 14380 2417
rect 14414 2383 14448 2417
rect 14482 2383 14516 2417
rect 14550 2383 14584 2417
rect 14618 2383 14630 2417
rect 13630 2372 14630 2383
rect 13630 2261 14630 2272
rect 13630 2227 13700 2261
rect 13734 2227 13768 2261
rect 13802 2227 13836 2261
rect 13870 2227 13904 2261
rect 13938 2227 13972 2261
rect 14006 2227 14040 2261
rect 14074 2227 14108 2261
rect 14142 2227 14176 2261
rect 14210 2227 14244 2261
rect 14278 2227 14312 2261
rect 14346 2227 14380 2261
rect 14414 2227 14448 2261
rect 14482 2227 14516 2261
rect 14550 2227 14584 2261
rect 14618 2227 14630 2261
rect 13630 2216 14630 2227
rect 13630 2105 14630 2116
rect 13630 2071 13700 2105
rect 13734 2071 13768 2105
rect 13802 2071 13836 2105
rect 13870 2071 13904 2105
rect 13938 2071 13972 2105
rect 14006 2071 14040 2105
rect 14074 2071 14108 2105
rect 14142 2071 14176 2105
rect 14210 2071 14244 2105
rect 14278 2071 14312 2105
rect 14346 2071 14380 2105
rect 14414 2071 14448 2105
rect 14482 2071 14516 2105
rect 14550 2071 14584 2105
rect 14618 2071 14630 2105
rect 13630 2060 14630 2071
rect 13630 1949 14630 1960
rect 13630 1915 13700 1949
rect 13734 1915 13768 1949
rect 13802 1915 13836 1949
rect 13870 1915 13904 1949
rect 13938 1915 13972 1949
rect 14006 1915 14040 1949
rect 14074 1915 14108 1949
rect 14142 1915 14176 1949
rect 14210 1915 14244 1949
rect 14278 1915 14312 1949
rect 14346 1915 14380 1949
rect 14414 1915 14448 1949
rect 14482 1915 14516 1949
rect 14550 1915 14584 1949
rect 14618 1915 14630 1949
rect 13630 1904 14630 1915
rect 13630 1793 14630 1804
rect 13630 1759 13700 1793
rect 13734 1759 13768 1793
rect 13802 1759 13836 1793
rect 13870 1759 13904 1793
rect 13938 1759 13972 1793
rect 14006 1759 14040 1793
rect 14074 1759 14108 1793
rect 14142 1759 14176 1793
rect 14210 1759 14244 1793
rect 14278 1759 14312 1793
rect 14346 1759 14380 1793
rect 14414 1759 14448 1793
rect 14482 1759 14516 1793
rect 14550 1759 14584 1793
rect 14618 1759 14630 1793
rect 13630 1748 14630 1759
rect 13630 1637 14630 1648
rect 13630 1603 13700 1637
rect 13734 1603 13768 1637
rect 13802 1603 13836 1637
rect 13870 1603 13904 1637
rect 13938 1603 13972 1637
rect 14006 1603 14040 1637
rect 14074 1603 14108 1637
rect 14142 1603 14176 1637
rect 14210 1603 14244 1637
rect 14278 1603 14312 1637
rect 14346 1603 14380 1637
rect 14414 1603 14448 1637
rect 14482 1603 14516 1637
rect 14550 1603 14584 1637
rect 14618 1603 14630 1637
rect 13630 1592 14630 1603
rect 13630 1481 14630 1492
rect 13630 1447 13700 1481
rect 13734 1447 13768 1481
rect 13802 1447 13836 1481
rect 13870 1447 13904 1481
rect 13938 1447 13972 1481
rect 14006 1447 14040 1481
rect 14074 1447 14108 1481
rect 14142 1447 14176 1481
rect 14210 1447 14244 1481
rect 14278 1447 14312 1481
rect 14346 1447 14380 1481
rect 14414 1447 14448 1481
rect 14482 1447 14516 1481
rect 14550 1447 14584 1481
rect 14618 1447 14630 1481
rect 13630 1436 14630 1447
rect 13630 1325 14630 1336
rect 13630 1291 13700 1325
rect 13734 1291 13768 1325
rect 13802 1291 13836 1325
rect 13870 1291 13904 1325
rect 13938 1291 13972 1325
rect 14006 1291 14040 1325
rect 14074 1291 14108 1325
rect 14142 1291 14176 1325
rect 14210 1291 14244 1325
rect 14278 1291 14312 1325
rect 14346 1291 14380 1325
rect 14414 1291 14448 1325
rect 14482 1291 14516 1325
rect 14550 1291 14584 1325
rect 14618 1291 14630 1325
rect 13630 1280 14630 1291
rect 13630 1169 14630 1180
rect 13630 1135 13700 1169
rect 13734 1135 13768 1169
rect 13802 1135 13836 1169
rect 13870 1135 13904 1169
rect 13938 1135 13972 1169
rect 14006 1135 14040 1169
rect 14074 1135 14108 1169
rect 14142 1135 14176 1169
rect 14210 1135 14244 1169
rect 14278 1135 14312 1169
rect 14346 1135 14380 1169
rect 14414 1135 14448 1169
rect 14482 1135 14516 1169
rect 14550 1135 14584 1169
rect 14618 1135 14630 1169
rect 13630 1124 14630 1135
rect 13630 1013 14630 1024
rect 13630 979 13700 1013
rect 13734 979 13768 1013
rect 13802 979 13836 1013
rect 13870 979 13904 1013
rect 13938 979 13972 1013
rect 14006 979 14040 1013
rect 14074 979 14108 1013
rect 14142 979 14176 1013
rect 14210 979 14244 1013
rect 14278 979 14312 1013
rect 14346 979 14380 1013
rect 14414 979 14448 1013
rect 14482 979 14516 1013
rect 14550 979 14584 1013
rect 14618 979 14630 1013
rect 13630 968 14630 979
rect 13630 857 14630 868
rect 13630 823 13700 857
rect 13734 823 13768 857
rect 13802 823 13836 857
rect 13870 823 13904 857
rect 13938 823 13972 857
rect 14006 823 14040 857
rect 14074 823 14108 857
rect 14142 823 14176 857
rect 14210 823 14244 857
rect 14278 823 14312 857
rect 14346 823 14380 857
rect 14414 823 14448 857
rect 14482 823 14516 857
rect 14550 823 14584 857
rect 14618 823 14630 857
rect 13630 812 14630 823
rect 13630 701 14630 712
rect 13630 667 13700 701
rect 13734 667 13768 701
rect 13802 667 13836 701
rect 13870 667 13904 701
rect 13938 667 13972 701
rect 14006 667 14040 701
rect 14074 667 14108 701
rect 14142 667 14176 701
rect 14210 667 14244 701
rect 14278 667 14312 701
rect 14346 667 14380 701
rect 14414 667 14448 701
rect 14482 667 14516 701
rect 14550 667 14584 701
rect 14618 667 14630 701
rect 13630 656 14630 667
rect 13630 545 14630 556
rect 13630 511 13700 545
rect 13734 511 13768 545
rect 13802 511 13836 545
rect 13870 511 13904 545
rect 13938 511 13972 545
rect 14006 511 14040 545
rect 14074 511 14108 545
rect 14142 511 14176 545
rect 14210 511 14244 545
rect 14278 511 14312 545
rect 14346 511 14380 545
rect 14414 511 14448 545
rect 14482 511 14516 545
rect 14550 511 14584 545
rect 14618 511 14630 545
rect 13630 500 14630 511
rect 13630 389 14630 400
rect 13630 355 13700 389
rect 13734 355 13768 389
rect 13802 355 13836 389
rect 13870 355 13904 389
rect 13938 355 13972 389
rect 14006 355 14040 389
rect 14074 355 14108 389
rect 14142 355 14176 389
rect 14210 355 14244 389
rect 14278 355 14312 389
rect 14346 355 14380 389
rect 14414 355 14448 389
rect 14482 355 14516 389
rect 14550 355 14584 389
rect 14618 355 14630 389
rect 13630 344 14630 355
<< mvpdiff >>
rect 1282 8472 4282 8483
rect 1282 8438 1294 8472
rect 1328 8438 1362 8472
rect 1396 8438 1430 8472
rect 1464 8438 1498 8472
rect 1532 8438 1566 8472
rect 1600 8438 1634 8472
rect 1668 8438 1702 8472
rect 1736 8438 1770 8472
rect 1804 8438 1838 8472
rect 1872 8438 1906 8472
rect 1940 8438 1974 8472
rect 2008 8438 2042 8472
rect 2076 8438 2110 8472
rect 2144 8438 2178 8472
rect 2212 8438 2246 8472
rect 2280 8438 2314 8472
rect 2348 8438 2382 8472
rect 2416 8438 2450 8472
rect 2484 8438 2518 8472
rect 2552 8438 2586 8472
rect 2620 8438 2654 8472
rect 2688 8438 2722 8472
rect 2756 8438 2790 8472
rect 2824 8438 2858 8472
rect 2892 8438 2926 8472
rect 2960 8438 2994 8472
rect 3028 8438 3062 8472
rect 3096 8438 3130 8472
rect 3164 8438 3198 8472
rect 3232 8438 3266 8472
rect 3300 8438 3334 8472
rect 3368 8438 3402 8472
rect 3436 8438 3470 8472
rect 3504 8438 3538 8472
rect 3572 8438 3606 8472
rect 3640 8438 3674 8472
rect 3708 8438 3742 8472
rect 3776 8438 3810 8472
rect 3844 8438 3878 8472
rect 3912 8438 3946 8472
rect 3980 8438 4014 8472
rect 4048 8438 4082 8472
rect 4116 8438 4150 8472
rect 4184 8438 4218 8472
rect 4252 8438 4282 8472
rect 1282 8427 4282 8438
rect 1282 8316 4282 8327
rect 1282 8282 1294 8316
rect 1328 8282 1362 8316
rect 1396 8282 1430 8316
rect 1464 8282 1498 8316
rect 1532 8282 1566 8316
rect 1600 8282 1634 8316
rect 1668 8282 1702 8316
rect 1736 8282 1770 8316
rect 1804 8282 1838 8316
rect 1872 8282 1906 8316
rect 1940 8282 1974 8316
rect 2008 8282 2042 8316
rect 2076 8282 2110 8316
rect 2144 8282 2178 8316
rect 2212 8282 2246 8316
rect 2280 8282 2314 8316
rect 2348 8282 2382 8316
rect 2416 8282 2450 8316
rect 2484 8282 2518 8316
rect 2552 8282 2586 8316
rect 2620 8282 2654 8316
rect 2688 8282 2722 8316
rect 2756 8282 2790 8316
rect 2824 8282 2858 8316
rect 2892 8282 2926 8316
rect 2960 8282 2994 8316
rect 3028 8282 3062 8316
rect 3096 8282 3130 8316
rect 3164 8282 3198 8316
rect 3232 8282 3266 8316
rect 3300 8282 3334 8316
rect 3368 8282 3402 8316
rect 3436 8282 3470 8316
rect 3504 8282 3538 8316
rect 3572 8282 3606 8316
rect 3640 8282 3674 8316
rect 3708 8282 3742 8316
rect 3776 8282 3810 8316
rect 3844 8282 3878 8316
rect 3912 8282 3946 8316
rect 3980 8282 4014 8316
rect 4048 8282 4082 8316
rect 4116 8282 4150 8316
rect 4184 8282 4218 8316
rect 4252 8282 4282 8316
rect 1282 8271 4282 8282
rect 1282 8160 4282 8171
rect 1282 8126 1294 8160
rect 1328 8126 1362 8160
rect 1396 8126 1430 8160
rect 1464 8126 1498 8160
rect 1532 8126 1566 8160
rect 1600 8126 1634 8160
rect 1668 8126 1702 8160
rect 1736 8126 1770 8160
rect 1804 8126 1838 8160
rect 1872 8126 1906 8160
rect 1940 8126 1974 8160
rect 2008 8126 2042 8160
rect 2076 8126 2110 8160
rect 2144 8126 2178 8160
rect 2212 8126 2246 8160
rect 2280 8126 2314 8160
rect 2348 8126 2382 8160
rect 2416 8126 2450 8160
rect 2484 8126 2518 8160
rect 2552 8126 2586 8160
rect 2620 8126 2654 8160
rect 2688 8126 2722 8160
rect 2756 8126 2790 8160
rect 2824 8126 2858 8160
rect 2892 8126 2926 8160
rect 2960 8126 2994 8160
rect 3028 8126 3062 8160
rect 3096 8126 3130 8160
rect 3164 8126 3198 8160
rect 3232 8126 3266 8160
rect 3300 8126 3334 8160
rect 3368 8126 3402 8160
rect 3436 8126 3470 8160
rect 3504 8126 3538 8160
rect 3572 8126 3606 8160
rect 3640 8126 3674 8160
rect 3708 8126 3742 8160
rect 3776 8126 3810 8160
rect 3844 8126 3878 8160
rect 3912 8126 3946 8160
rect 3980 8126 4014 8160
rect 4048 8126 4082 8160
rect 4116 8126 4150 8160
rect 4184 8126 4218 8160
rect 4252 8126 4282 8160
rect 1282 8115 4282 8126
rect 1282 8004 4282 8015
rect 1282 7970 1294 8004
rect 1328 7970 1362 8004
rect 1396 7970 1430 8004
rect 1464 7970 1498 8004
rect 1532 7970 1566 8004
rect 1600 7970 1634 8004
rect 1668 7970 1702 8004
rect 1736 7970 1770 8004
rect 1804 7970 1838 8004
rect 1872 7970 1906 8004
rect 1940 7970 1974 8004
rect 2008 7970 2042 8004
rect 2076 7970 2110 8004
rect 2144 7970 2178 8004
rect 2212 7970 2246 8004
rect 2280 7970 2314 8004
rect 2348 7970 2382 8004
rect 2416 7970 2450 8004
rect 2484 7970 2518 8004
rect 2552 7970 2586 8004
rect 2620 7970 2654 8004
rect 2688 7970 2722 8004
rect 2756 7970 2790 8004
rect 2824 7970 2858 8004
rect 2892 7970 2926 8004
rect 2960 7970 2994 8004
rect 3028 7970 3062 8004
rect 3096 7970 3130 8004
rect 3164 7970 3198 8004
rect 3232 7970 3266 8004
rect 3300 7970 3334 8004
rect 3368 7970 3402 8004
rect 3436 7970 3470 8004
rect 3504 7970 3538 8004
rect 3572 7970 3606 8004
rect 3640 7970 3674 8004
rect 3708 7970 3742 8004
rect 3776 7970 3810 8004
rect 3844 7970 3878 8004
rect 3912 7970 3946 8004
rect 3980 7970 4014 8004
rect 4048 7970 4082 8004
rect 4116 7970 4150 8004
rect 4184 7970 4218 8004
rect 4252 7970 4282 8004
rect 1282 7959 4282 7970
rect 1282 7848 4282 7859
rect 1282 7814 1294 7848
rect 1328 7814 1362 7848
rect 1396 7814 1430 7848
rect 1464 7814 1498 7848
rect 1532 7814 1566 7848
rect 1600 7814 1634 7848
rect 1668 7814 1702 7848
rect 1736 7814 1770 7848
rect 1804 7814 1838 7848
rect 1872 7814 1906 7848
rect 1940 7814 1974 7848
rect 2008 7814 2042 7848
rect 2076 7814 2110 7848
rect 2144 7814 2178 7848
rect 2212 7814 2246 7848
rect 2280 7814 2314 7848
rect 2348 7814 2382 7848
rect 2416 7814 2450 7848
rect 2484 7814 2518 7848
rect 2552 7814 2586 7848
rect 2620 7814 2654 7848
rect 2688 7814 2722 7848
rect 2756 7814 2790 7848
rect 2824 7814 2858 7848
rect 2892 7814 2926 7848
rect 2960 7814 2994 7848
rect 3028 7814 3062 7848
rect 3096 7814 3130 7848
rect 3164 7814 3198 7848
rect 3232 7814 3266 7848
rect 3300 7814 3334 7848
rect 3368 7814 3402 7848
rect 3436 7814 3470 7848
rect 3504 7814 3538 7848
rect 3572 7814 3606 7848
rect 3640 7814 3674 7848
rect 3708 7814 3742 7848
rect 3776 7814 3810 7848
rect 3844 7814 3878 7848
rect 3912 7814 3946 7848
rect 3980 7814 4014 7848
rect 4048 7814 4082 7848
rect 4116 7814 4150 7848
rect 4184 7814 4218 7848
rect 4252 7814 4282 7848
rect 1282 7803 4282 7814
rect 1282 7692 4282 7703
rect 1282 7658 1294 7692
rect 1328 7658 1362 7692
rect 1396 7658 1430 7692
rect 1464 7658 1498 7692
rect 1532 7658 1566 7692
rect 1600 7658 1634 7692
rect 1668 7658 1702 7692
rect 1736 7658 1770 7692
rect 1804 7658 1838 7692
rect 1872 7658 1906 7692
rect 1940 7658 1974 7692
rect 2008 7658 2042 7692
rect 2076 7658 2110 7692
rect 2144 7658 2178 7692
rect 2212 7658 2246 7692
rect 2280 7658 2314 7692
rect 2348 7658 2382 7692
rect 2416 7658 2450 7692
rect 2484 7658 2518 7692
rect 2552 7658 2586 7692
rect 2620 7658 2654 7692
rect 2688 7658 2722 7692
rect 2756 7658 2790 7692
rect 2824 7658 2858 7692
rect 2892 7658 2926 7692
rect 2960 7658 2994 7692
rect 3028 7658 3062 7692
rect 3096 7658 3130 7692
rect 3164 7658 3198 7692
rect 3232 7658 3266 7692
rect 3300 7658 3334 7692
rect 3368 7658 3402 7692
rect 3436 7658 3470 7692
rect 3504 7658 3538 7692
rect 3572 7658 3606 7692
rect 3640 7658 3674 7692
rect 3708 7658 3742 7692
rect 3776 7658 3810 7692
rect 3844 7658 3878 7692
rect 3912 7658 3946 7692
rect 3980 7658 4014 7692
rect 4048 7658 4082 7692
rect 4116 7658 4150 7692
rect 4184 7658 4218 7692
rect 4252 7658 4282 7692
rect 1282 7647 4282 7658
rect 1282 7536 4282 7547
rect 1282 7502 1294 7536
rect 1328 7502 1362 7536
rect 1396 7502 1430 7536
rect 1464 7502 1498 7536
rect 1532 7502 1566 7536
rect 1600 7502 1634 7536
rect 1668 7502 1702 7536
rect 1736 7502 1770 7536
rect 1804 7502 1838 7536
rect 1872 7502 1906 7536
rect 1940 7502 1974 7536
rect 2008 7502 2042 7536
rect 2076 7502 2110 7536
rect 2144 7502 2178 7536
rect 2212 7502 2246 7536
rect 2280 7502 2314 7536
rect 2348 7502 2382 7536
rect 2416 7502 2450 7536
rect 2484 7502 2518 7536
rect 2552 7502 2586 7536
rect 2620 7502 2654 7536
rect 2688 7502 2722 7536
rect 2756 7502 2790 7536
rect 2824 7502 2858 7536
rect 2892 7502 2926 7536
rect 2960 7502 2994 7536
rect 3028 7502 3062 7536
rect 3096 7502 3130 7536
rect 3164 7502 3198 7536
rect 3232 7502 3266 7536
rect 3300 7502 3334 7536
rect 3368 7502 3402 7536
rect 3436 7502 3470 7536
rect 3504 7502 3538 7536
rect 3572 7502 3606 7536
rect 3640 7502 3674 7536
rect 3708 7502 3742 7536
rect 3776 7502 3810 7536
rect 3844 7502 3878 7536
rect 3912 7502 3946 7536
rect 3980 7502 4014 7536
rect 4048 7502 4082 7536
rect 4116 7502 4150 7536
rect 4184 7502 4218 7536
rect 4252 7502 4282 7536
rect 1282 7491 4282 7502
rect 1282 7380 4282 7391
rect 1282 7346 1294 7380
rect 1328 7346 1362 7380
rect 1396 7346 1430 7380
rect 1464 7346 1498 7380
rect 1532 7346 1566 7380
rect 1600 7346 1634 7380
rect 1668 7346 1702 7380
rect 1736 7346 1770 7380
rect 1804 7346 1838 7380
rect 1872 7346 1906 7380
rect 1940 7346 1974 7380
rect 2008 7346 2042 7380
rect 2076 7346 2110 7380
rect 2144 7346 2178 7380
rect 2212 7346 2246 7380
rect 2280 7346 2314 7380
rect 2348 7346 2382 7380
rect 2416 7346 2450 7380
rect 2484 7346 2518 7380
rect 2552 7346 2586 7380
rect 2620 7346 2654 7380
rect 2688 7346 2722 7380
rect 2756 7346 2790 7380
rect 2824 7346 2858 7380
rect 2892 7346 2926 7380
rect 2960 7346 2994 7380
rect 3028 7346 3062 7380
rect 3096 7346 3130 7380
rect 3164 7346 3198 7380
rect 3232 7346 3266 7380
rect 3300 7346 3334 7380
rect 3368 7346 3402 7380
rect 3436 7346 3470 7380
rect 3504 7346 3538 7380
rect 3572 7346 3606 7380
rect 3640 7346 3674 7380
rect 3708 7346 3742 7380
rect 3776 7346 3810 7380
rect 3844 7346 3878 7380
rect 3912 7346 3946 7380
rect 3980 7346 4014 7380
rect 4048 7346 4082 7380
rect 4116 7346 4150 7380
rect 4184 7346 4218 7380
rect 4252 7346 4282 7380
rect 1282 7335 4282 7346
<< mvndiffc >>
rect 13558 3903 13592 3937
rect 13558 3835 13592 3869
rect 13558 3767 13592 3801
rect 13558 3699 13592 3733
rect 13558 3631 13592 3665
rect 13558 3563 13592 3597
rect 13558 3495 13592 3529
rect 13558 3427 13592 3461
rect 13714 3903 13748 3937
rect 13714 3835 13748 3869
rect 13714 3767 13748 3801
rect 13714 3699 13748 3733
rect 13714 3631 13748 3665
rect 13714 3563 13748 3597
rect 13714 3495 13748 3529
rect 13714 3427 13748 3461
rect 13830 3903 13864 3937
rect 13830 3835 13864 3869
rect 13830 3767 13864 3801
rect 13830 3699 13864 3733
rect 13830 3631 13864 3665
rect 13830 3563 13864 3597
rect 13830 3495 13864 3529
rect 13830 3427 13864 3461
rect 13986 3903 14020 3937
rect 13986 3835 14020 3869
rect 13986 3767 14020 3801
rect 13986 3699 14020 3733
rect 13986 3631 14020 3665
rect 13986 3563 14020 3597
rect 13986 3495 14020 3529
rect 13986 3427 14020 3461
rect 14106 3903 14140 3937
rect 14106 3835 14140 3869
rect 14106 3767 14140 3801
rect 14106 3699 14140 3733
rect 14106 3631 14140 3665
rect 14106 3563 14140 3597
rect 14106 3495 14140 3529
rect 14106 3427 14140 3461
rect 14262 3903 14296 3937
rect 14262 3835 14296 3869
rect 14262 3767 14296 3801
rect 14262 3699 14296 3733
rect 14262 3631 14296 3665
rect 14262 3563 14296 3597
rect 14262 3495 14296 3529
rect 14262 3427 14296 3461
rect 14378 3903 14412 3937
rect 14378 3835 14412 3869
rect 14378 3767 14412 3801
rect 14378 3699 14412 3733
rect 14378 3631 14412 3665
rect 14378 3563 14412 3597
rect 14378 3495 14412 3529
rect 14378 3427 14412 3461
rect 14534 3903 14568 3937
rect 14534 3835 14568 3869
rect 14534 3767 14568 3801
rect 14534 3699 14568 3733
rect 14534 3631 14568 3665
rect 14534 3563 14568 3597
rect 14534 3495 14568 3529
rect 14534 3427 14568 3461
rect 13563 3275 13597 3309
rect 13719 3275 13753 3309
rect 13835 3275 13869 3309
rect 13991 3275 14025 3309
rect 14107 3275 14141 3309
rect 14263 3275 14297 3309
rect 14379 3275 14413 3309
rect 14535 3275 14569 3309
rect 13563 3047 13597 3081
rect 13719 3047 13753 3081
rect 13835 3047 13869 3081
rect 13991 3047 14025 3081
rect 14107 3047 14141 3081
rect 14263 3047 14297 3081
rect 14379 3047 14413 3081
rect 14535 3047 14569 3081
rect 13700 2539 13734 2573
rect 13768 2539 13802 2573
rect 13836 2539 13870 2573
rect 13904 2539 13938 2573
rect 13972 2539 14006 2573
rect 14040 2539 14074 2573
rect 14108 2539 14142 2573
rect 14176 2539 14210 2573
rect 14244 2539 14278 2573
rect 14312 2539 14346 2573
rect 14380 2539 14414 2573
rect 14448 2539 14482 2573
rect 14516 2539 14550 2573
rect 14584 2539 14618 2573
rect 13700 2383 13734 2417
rect 13768 2383 13802 2417
rect 13836 2383 13870 2417
rect 13904 2383 13938 2417
rect 13972 2383 14006 2417
rect 14040 2383 14074 2417
rect 14108 2383 14142 2417
rect 14176 2383 14210 2417
rect 14244 2383 14278 2417
rect 14312 2383 14346 2417
rect 14380 2383 14414 2417
rect 14448 2383 14482 2417
rect 14516 2383 14550 2417
rect 14584 2383 14618 2417
rect 13700 2227 13734 2261
rect 13768 2227 13802 2261
rect 13836 2227 13870 2261
rect 13904 2227 13938 2261
rect 13972 2227 14006 2261
rect 14040 2227 14074 2261
rect 14108 2227 14142 2261
rect 14176 2227 14210 2261
rect 14244 2227 14278 2261
rect 14312 2227 14346 2261
rect 14380 2227 14414 2261
rect 14448 2227 14482 2261
rect 14516 2227 14550 2261
rect 14584 2227 14618 2261
rect 13700 2071 13734 2105
rect 13768 2071 13802 2105
rect 13836 2071 13870 2105
rect 13904 2071 13938 2105
rect 13972 2071 14006 2105
rect 14040 2071 14074 2105
rect 14108 2071 14142 2105
rect 14176 2071 14210 2105
rect 14244 2071 14278 2105
rect 14312 2071 14346 2105
rect 14380 2071 14414 2105
rect 14448 2071 14482 2105
rect 14516 2071 14550 2105
rect 14584 2071 14618 2105
rect 13700 1915 13734 1949
rect 13768 1915 13802 1949
rect 13836 1915 13870 1949
rect 13904 1915 13938 1949
rect 13972 1915 14006 1949
rect 14040 1915 14074 1949
rect 14108 1915 14142 1949
rect 14176 1915 14210 1949
rect 14244 1915 14278 1949
rect 14312 1915 14346 1949
rect 14380 1915 14414 1949
rect 14448 1915 14482 1949
rect 14516 1915 14550 1949
rect 14584 1915 14618 1949
rect 13700 1759 13734 1793
rect 13768 1759 13802 1793
rect 13836 1759 13870 1793
rect 13904 1759 13938 1793
rect 13972 1759 14006 1793
rect 14040 1759 14074 1793
rect 14108 1759 14142 1793
rect 14176 1759 14210 1793
rect 14244 1759 14278 1793
rect 14312 1759 14346 1793
rect 14380 1759 14414 1793
rect 14448 1759 14482 1793
rect 14516 1759 14550 1793
rect 14584 1759 14618 1793
rect 13700 1603 13734 1637
rect 13768 1603 13802 1637
rect 13836 1603 13870 1637
rect 13904 1603 13938 1637
rect 13972 1603 14006 1637
rect 14040 1603 14074 1637
rect 14108 1603 14142 1637
rect 14176 1603 14210 1637
rect 14244 1603 14278 1637
rect 14312 1603 14346 1637
rect 14380 1603 14414 1637
rect 14448 1603 14482 1637
rect 14516 1603 14550 1637
rect 14584 1603 14618 1637
rect 13700 1447 13734 1481
rect 13768 1447 13802 1481
rect 13836 1447 13870 1481
rect 13904 1447 13938 1481
rect 13972 1447 14006 1481
rect 14040 1447 14074 1481
rect 14108 1447 14142 1481
rect 14176 1447 14210 1481
rect 14244 1447 14278 1481
rect 14312 1447 14346 1481
rect 14380 1447 14414 1481
rect 14448 1447 14482 1481
rect 14516 1447 14550 1481
rect 14584 1447 14618 1481
rect 13700 1291 13734 1325
rect 13768 1291 13802 1325
rect 13836 1291 13870 1325
rect 13904 1291 13938 1325
rect 13972 1291 14006 1325
rect 14040 1291 14074 1325
rect 14108 1291 14142 1325
rect 14176 1291 14210 1325
rect 14244 1291 14278 1325
rect 14312 1291 14346 1325
rect 14380 1291 14414 1325
rect 14448 1291 14482 1325
rect 14516 1291 14550 1325
rect 14584 1291 14618 1325
rect 13700 1135 13734 1169
rect 13768 1135 13802 1169
rect 13836 1135 13870 1169
rect 13904 1135 13938 1169
rect 13972 1135 14006 1169
rect 14040 1135 14074 1169
rect 14108 1135 14142 1169
rect 14176 1135 14210 1169
rect 14244 1135 14278 1169
rect 14312 1135 14346 1169
rect 14380 1135 14414 1169
rect 14448 1135 14482 1169
rect 14516 1135 14550 1169
rect 14584 1135 14618 1169
rect 13700 979 13734 1013
rect 13768 979 13802 1013
rect 13836 979 13870 1013
rect 13904 979 13938 1013
rect 13972 979 14006 1013
rect 14040 979 14074 1013
rect 14108 979 14142 1013
rect 14176 979 14210 1013
rect 14244 979 14278 1013
rect 14312 979 14346 1013
rect 14380 979 14414 1013
rect 14448 979 14482 1013
rect 14516 979 14550 1013
rect 14584 979 14618 1013
rect 13700 823 13734 857
rect 13768 823 13802 857
rect 13836 823 13870 857
rect 13904 823 13938 857
rect 13972 823 14006 857
rect 14040 823 14074 857
rect 14108 823 14142 857
rect 14176 823 14210 857
rect 14244 823 14278 857
rect 14312 823 14346 857
rect 14380 823 14414 857
rect 14448 823 14482 857
rect 14516 823 14550 857
rect 14584 823 14618 857
rect 13700 667 13734 701
rect 13768 667 13802 701
rect 13836 667 13870 701
rect 13904 667 13938 701
rect 13972 667 14006 701
rect 14040 667 14074 701
rect 14108 667 14142 701
rect 14176 667 14210 701
rect 14244 667 14278 701
rect 14312 667 14346 701
rect 14380 667 14414 701
rect 14448 667 14482 701
rect 14516 667 14550 701
rect 14584 667 14618 701
rect 13700 511 13734 545
rect 13768 511 13802 545
rect 13836 511 13870 545
rect 13904 511 13938 545
rect 13972 511 14006 545
rect 14040 511 14074 545
rect 14108 511 14142 545
rect 14176 511 14210 545
rect 14244 511 14278 545
rect 14312 511 14346 545
rect 14380 511 14414 545
rect 14448 511 14482 545
rect 14516 511 14550 545
rect 14584 511 14618 545
rect 13700 355 13734 389
rect 13768 355 13802 389
rect 13836 355 13870 389
rect 13904 355 13938 389
rect 13972 355 14006 389
rect 14040 355 14074 389
rect 14108 355 14142 389
rect 14176 355 14210 389
rect 14244 355 14278 389
rect 14312 355 14346 389
rect 14380 355 14414 389
rect 14448 355 14482 389
rect 14516 355 14550 389
rect 14584 355 14618 389
<< mvpdiffc >>
rect 1294 8438 1328 8472
rect 1362 8438 1396 8472
rect 1430 8438 1464 8472
rect 1498 8438 1532 8472
rect 1566 8438 1600 8472
rect 1634 8438 1668 8472
rect 1702 8438 1736 8472
rect 1770 8438 1804 8472
rect 1838 8438 1872 8472
rect 1906 8438 1940 8472
rect 1974 8438 2008 8472
rect 2042 8438 2076 8472
rect 2110 8438 2144 8472
rect 2178 8438 2212 8472
rect 2246 8438 2280 8472
rect 2314 8438 2348 8472
rect 2382 8438 2416 8472
rect 2450 8438 2484 8472
rect 2518 8438 2552 8472
rect 2586 8438 2620 8472
rect 2654 8438 2688 8472
rect 2722 8438 2756 8472
rect 2790 8438 2824 8472
rect 2858 8438 2892 8472
rect 2926 8438 2960 8472
rect 2994 8438 3028 8472
rect 3062 8438 3096 8472
rect 3130 8438 3164 8472
rect 3198 8438 3232 8472
rect 3266 8438 3300 8472
rect 3334 8438 3368 8472
rect 3402 8438 3436 8472
rect 3470 8438 3504 8472
rect 3538 8438 3572 8472
rect 3606 8438 3640 8472
rect 3674 8438 3708 8472
rect 3742 8438 3776 8472
rect 3810 8438 3844 8472
rect 3878 8438 3912 8472
rect 3946 8438 3980 8472
rect 4014 8438 4048 8472
rect 4082 8438 4116 8472
rect 4150 8438 4184 8472
rect 4218 8438 4252 8472
rect 1294 8282 1328 8316
rect 1362 8282 1396 8316
rect 1430 8282 1464 8316
rect 1498 8282 1532 8316
rect 1566 8282 1600 8316
rect 1634 8282 1668 8316
rect 1702 8282 1736 8316
rect 1770 8282 1804 8316
rect 1838 8282 1872 8316
rect 1906 8282 1940 8316
rect 1974 8282 2008 8316
rect 2042 8282 2076 8316
rect 2110 8282 2144 8316
rect 2178 8282 2212 8316
rect 2246 8282 2280 8316
rect 2314 8282 2348 8316
rect 2382 8282 2416 8316
rect 2450 8282 2484 8316
rect 2518 8282 2552 8316
rect 2586 8282 2620 8316
rect 2654 8282 2688 8316
rect 2722 8282 2756 8316
rect 2790 8282 2824 8316
rect 2858 8282 2892 8316
rect 2926 8282 2960 8316
rect 2994 8282 3028 8316
rect 3062 8282 3096 8316
rect 3130 8282 3164 8316
rect 3198 8282 3232 8316
rect 3266 8282 3300 8316
rect 3334 8282 3368 8316
rect 3402 8282 3436 8316
rect 3470 8282 3504 8316
rect 3538 8282 3572 8316
rect 3606 8282 3640 8316
rect 3674 8282 3708 8316
rect 3742 8282 3776 8316
rect 3810 8282 3844 8316
rect 3878 8282 3912 8316
rect 3946 8282 3980 8316
rect 4014 8282 4048 8316
rect 4082 8282 4116 8316
rect 4150 8282 4184 8316
rect 4218 8282 4252 8316
rect 1294 8126 1328 8160
rect 1362 8126 1396 8160
rect 1430 8126 1464 8160
rect 1498 8126 1532 8160
rect 1566 8126 1600 8160
rect 1634 8126 1668 8160
rect 1702 8126 1736 8160
rect 1770 8126 1804 8160
rect 1838 8126 1872 8160
rect 1906 8126 1940 8160
rect 1974 8126 2008 8160
rect 2042 8126 2076 8160
rect 2110 8126 2144 8160
rect 2178 8126 2212 8160
rect 2246 8126 2280 8160
rect 2314 8126 2348 8160
rect 2382 8126 2416 8160
rect 2450 8126 2484 8160
rect 2518 8126 2552 8160
rect 2586 8126 2620 8160
rect 2654 8126 2688 8160
rect 2722 8126 2756 8160
rect 2790 8126 2824 8160
rect 2858 8126 2892 8160
rect 2926 8126 2960 8160
rect 2994 8126 3028 8160
rect 3062 8126 3096 8160
rect 3130 8126 3164 8160
rect 3198 8126 3232 8160
rect 3266 8126 3300 8160
rect 3334 8126 3368 8160
rect 3402 8126 3436 8160
rect 3470 8126 3504 8160
rect 3538 8126 3572 8160
rect 3606 8126 3640 8160
rect 3674 8126 3708 8160
rect 3742 8126 3776 8160
rect 3810 8126 3844 8160
rect 3878 8126 3912 8160
rect 3946 8126 3980 8160
rect 4014 8126 4048 8160
rect 4082 8126 4116 8160
rect 4150 8126 4184 8160
rect 4218 8126 4252 8160
rect 1294 7970 1328 8004
rect 1362 7970 1396 8004
rect 1430 7970 1464 8004
rect 1498 7970 1532 8004
rect 1566 7970 1600 8004
rect 1634 7970 1668 8004
rect 1702 7970 1736 8004
rect 1770 7970 1804 8004
rect 1838 7970 1872 8004
rect 1906 7970 1940 8004
rect 1974 7970 2008 8004
rect 2042 7970 2076 8004
rect 2110 7970 2144 8004
rect 2178 7970 2212 8004
rect 2246 7970 2280 8004
rect 2314 7970 2348 8004
rect 2382 7970 2416 8004
rect 2450 7970 2484 8004
rect 2518 7970 2552 8004
rect 2586 7970 2620 8004
rect 2654 7970 2688 8004
rect 2722 7970 2756 8004
rect 2790 7970 2824 8004
rect 2858 7970 2892 8004
rect 2926 7970 2960 8004
rect 2994 7970 3028 8004
rect 3062 7970 3096 8004
rect 3130 7970 3164 8004
rect 3198 7970 3232 8004
rect 3266 7970 3300 8004
rect 3334 7970 3368 8004
rect 3402 7970 3436 8004
rect 3470 7970 3504 8004
rect 3538 7970 3572 8004
rect 3606 7970 3640 8004
rect 3674 7970 3708 8004
rect 3742 7970 3776 8004
rect 3810 7970 3844 8004
rect 3878 7970 3912 8004
rect 3946 7970 3980 8004
rect 4014 7970 4048 8004
rect 4082 7970 4116 8004
rect 4150 7970 4184 8004
rect 4218 7970 4252 8004
rect 1294 7814 1328 7848
rect 1362 7814 1396 7848
rect 1430 7814 1464 7848
rect 1498 7814 1532 7848
rect 1566 7814 1600 7848
rect 1634 7814 1668 7848
rect 1702 7814 1736 7848
rect 1770 7814 1804 7848
rect 1838 7814 1872 7848
rect 1906 7814 1940 7848
rect 1974 7814 2008 7848
rect 2042 7814 2076 7848
rect 2110 7814 2144 7848
rect 2178 7814 2212 7848
rect 2246 7814 2280 7848
rect 2314 7814 2348 7848
rect 2382 7814 2416 7848
rect 2450 7814 2484 7848
rect 2518 7814 2552 7848
rect 2586 7814 2620 7848
rect 2654 7814 2688 7848
rect 2722 7814 2756 7848
rect 2790 7814 2824 7848
rect 2858 7814 2892 7848
rect 2926 7814 2960 7848
rect 2994 7814 3028 7848
rect 3062 7814 3096 7848
rect 3130 7814 3164 7848
rect 3198 7814 3232 7848
rect 3266 7814 3300 7848
rect 3334 7814 3368 7848
rect 3402 7814 3436 7848
rect 3470 7814 3504 7848
rect 3538 7814 3572 7848
rect 3606 7814 3640 7848
rect 3674 7814 3708 7848
rect 3742 7814 3776 7848
rect 3810 7814 3844 7848
rect 3878 7814 3912 7848
rect 3946 7814 3980 7848
rect 4014 7814 4048 7848
rect 4082 7814 4116 7848
rect 4150 7814 4184 7848
rect 4218 7814 4252 7848
rect 1294 7658 1328 7692
rect 1362 7658 1396 7692
rect 1430 7658 1464 7692
rect 1498 7658 1532 7692
rect 1566 7658 1600 7692
rect 1634 7658 1668 7692
rect 1702 7658 1736 7692
rect 1770 7658 1804 7692
rect 1838 7658 1872 7692
rect 1906 7658 1940 7692
rect 1974 7658 2008 7692
rect 2042 7658 2076 7692
rect 2110 7658 2144 7692
rect 2178 7658 2212 7692
rect 2246 7658 2280 7692
rect 2314 7658 2348 7692
rect 2382 7658 2416 7692
rect 2450 7658 2484 7692
rect 2518 7658 2552 7692
rect 2586 7658 2620 7692
rect 2654 7658 2688 7692
rect 2722 7658 2756 7692
rect 2790 7658 2824 7692
rect 2858 7658 2892 7692
rect 2926 7658 2960 7692
rect 2994 7658 3028 7692
rect 3062 7658 3096 7692
rect 3130 7658 3164 7692
rect 3198 7658 3232 7692
rect 3266 7658 3300 7692
rect 3334 7658 3368 7692
rect 3402 7658 3436 7692
rect 3470 7658 3504 7692
rect 3538 7658 3572 7692
rect 3606 7658 3640 7692
rect 3674 7658 3708 7692
rect 3742 7658 3776 7692
rect 3810 7658 3844 7692
rect 3878 7658 3912 7692
rect 3946 7658 3980 7692
rect 4014 7658 4048 7692
rect 4082 7658 4116 7692
rect 4150 7658 4184 7692
rect 4218 7658 4252 7692
rect 1294 7502 1328 7536
rect 1362 7502 1396 7536
rect 1430 7502 1464 7536
rect 1498 7502 1532 7536
rect 1566 7502 1600 7536
rect 1634 7502 1668 7536
rect 1702 7502 1736 7536
rect 1770 7502 1804 7536
rect 1838 7502 1872 7536
rect 1906 7502 1940 7536
rect 1974 7502 2008 7536
rect 2042 7502 2076 7536
rect 2110 7502 2144 7536
rect 2178 7502 2212 7536
rect 2246 7502 2280 7536
rect 2314 7502 2348 7536
rect 2382 7502 2416 7536
rect 2450 7502 2484 7536
rect 2518 7502 2552 7536
rect 2586 7502 2620 7536
rect 2654 7502 2688 7536
rect 2722 7502 2756 7536
rect 2790 7502 2824 7536
rect 2858 7502 2892 7536
rect 2926 7502 2960 7536
rect 2994 7502 3028 7536
rect 3062 7502 3096 7536
rect 3130 7502 3164 7536
rect 3198 7502 3232 7536
rect 3266 7502 3300 7536
rect 3334 7502 3368 7536
rect 3402 7502 3436 7536
rect 3470 7502 3504 7536
rect 3538 7502 3572 7536
rect 3606 7502 3640 7536
rect 3674 7502 3708 7536
rect 3742 7502 3776 7536
rect 3810 7502 3844 7536
rect 3878 7502 3912 7536
rect 3946 7502 3980 7536
rect 4014 7502 4048 7536
rect 4082 7502 4116 7536
rect 4150 7502 4184 7536
rect 4218 7502 4252 7536
rect 1294 7346 1328 7380
rect 1362 7346 1396 7380
rect 1430 7346 1464 7380
rect 1498 7346 1532 7380
rect 1566 7346 1600 7380
rect 1634 7346 1668 7380
rect 1702 7346 1736 7380
rect 1770 7346 1804 7380
rect 1838 7346 1872 7380
rect 1906 7346 1940 7380
rect 1974 7346 2008 7380
rect 2042 7346 2076 7380
rect 2110 7346 2144 7380
rect 2178 7346 2212 7380
rect 2246 7346 2280 7380
rect 2314 7346 2348 7380
rect 2382 7346 2416 7380
rect 2450 7346 2484 7380
rect 2518 7346 2552 7380
rect 2586 7346 2620 7380
rect 2654 7346 2688 7380
rect 2722 7346 2756 7380
rect 2790 7346 2824 7380
rect 2858 7346 2892 7380
rect 2926 7346 2960 7380
rect 2994 7346 3028 7380
rect 3062 7346 3096 7380
rect 3130 7346 3164 7380
rect 3198 7346 3232 7380
rect 3266 7346 3300 7380
rect 3334 7346 3368 7380
rect 3402 7346 3436 7380
rect 3470 7346 3504 7380
rect 3538 7346 3572 7380
rect 3606 7346 3640 7380
rect 3674 7346 3708 7380
rect 3742 7346 3776 7380
rect 3810 7346 3844 7380
rect 3878 7346 3912 7380
rect 3946 7346 3980 7380
rect 4014 7346 4048 7380
rect 4082 7346 4116 7380
rect 4150 7346 4184 7380
rect 4218 7346 4252 7380
<< psubdiff >>
rect 8037 -96 8071 -62
rect 8105 -96 8119 -62
rect 10501 -96 10515 -62
rect 10549 -96 10583 -62
rect 7563 -128 8119 -96
rect 5735 -140 8119 -128
rect 10501 -140 11128 -96
rect 5735 -174 5769 -140
rect 5803 -174 5838 -140
rect 5872 -174 5907 -140
rect 5941 -174 5976 -140
rect 6010 -174 6045 -140
rect 6079 -174 6114 -140
rect 6148 -174 6183 -140
rect 6217 -174 6252 -140
rect 6286 -174 6321 -140
rect 6355 -174 6390 -140
rect 6424 -174 6459 -140
rect 6493 -174 6528 -140
rect 6562 -174 6597 -140
rect 6631 -174 6666 -140
rect 6700 -174 6735 -140
rect 6769 -174 6804 -140
rect 6838 -174 6873 -140
rect 6907 -174 6942 -140
rect 6976 -174 7011 -140
rect 7045 -174 7080 -140
rect 7114 -174 7149 -140
rect 7183 -174 7218 -140
rect 7252 -174 7287 -140
rect 7321 -174 7356 -140
rect 7390 -174 7425 -140
rect 7459 -174 7494 -140
rect 7528 -174 7563 -140
rect 7597 -174 7632 -140
rect 7666 -174 7701 -140
rect 7735 -174 7770 -140
rect 7804 -174 7839 -140
rect 7873 -174 7908 -140
rect 7942 -174 7977 -140
rect 8011 -174 8046 -140
rect 8080 -174 8115 -140
rect 10532 -174 10566 -140
rect 10600 -174 10634 -140
rect 10668 -174 10702 -140
rect 10736 -174 10770 -140
rect 10804 -174 10838 -140
rect 10872 -174 10906 -140
rect 10940 -174 10974 -140
rect 11008 -174 11042 -140
rect 11076 -174 11110 -140
rect 5735 -191 8119 -174
rect 10501 -191 11128 -174
rect 5735 -215 12838 -191
rect 12277 -255 12797 -215
rect 12277 -289 12316 -255
rect 12350 -289 12384 -255
rect 12418 -289 12452 -255
rect 12486 -289 12520 -255
rect 12554 -289 12588 -255
rect 12622 -289 12656 -255
rect 12690 -289 12724 -255
rect 12758 -289 12797 -255
rect 12277 -325 12797 -289
rect 12277 -359 12316 -325
rect 12350 -359 12384 -325
rect 12418 -359 12452 -325
rect 12486 -359 12520 -325
rect 12554 -359 12588 -325
rect 12622 -359 12656 -325
rect 12690 -359 12724 -325
rect 12758 -359 12797 -325
rect 12277 -395 12797 -359
rect 12277 -429 12316 -395
rect 12350 -429 12384 -395
rect 12418 -429 12452 -395
rect 12486 -429 12520 -395
rect 12554 -429 12588 -395
rect 12622 -429 12656 -395
rect 12690 -429 12724 -395
rect 12758 -429 12797 -395
rect 12277 -465 12797 -429
rect 12277 -499 12316 -465
rect 12350 -499 12384 -465
rect 12418 -499 12452 -465
rect 12486 -499 12520 -465
rect 12554 -499 12588 -465
rect 12622 -499 12656 -465
rect 12690 -499 12724 -465
rect 12758 -499 12797 -465
rect 12277 -535 12797 -499
rect 12277 -569 12316 -535
rect 12350 -569 12384 -535
rect 12418 -569 12452 -535
rect 12486 -569 12520 -535
rect 12554 -569 12588 -535
rect 12622 -569 12656 -535
rect 12690 -569 12724 -535
rect 12758 -569 12797 -535
rect 12277 -606 12797 -569
rect 12277 -640 12316 -606
rect 12350 -640 12384 -606
rect 12418 -640 12452 -606
rect 12486 -640 12520 -606
rect 12554 -640 12588 -606
rect 12622 -640 12656 -606
rect 12690 -640 12724 -606
rect 12758 -640 12797 -606
rect 12277 -677 12797 -640
rect 12277 -711 12316 -677
rect 12350 -711 12384 -677
rect 12418 -711 12452 -677
rect 12486 -711 12520 -677
rect 12554 -711 12588 -677
rect 12622 -711 12656 -677
rect 12690 -711 12724 -677
rect 12758 -711 12797 -677
rect 12277 -748 12797 -711
rect 12277 -782 12316 -748
rect 12350 -782 12384 -748
rect 12418 -782 12452 -748
rect 12486 -782 12520 -748
rect 12554 -782 12588 -748
rect 12622 -782 12656 -748
rect 12690 -782 12724 -748
rect 12758 -782 12797 -748
rect 12277 -819 12797 -782
rect 12277 -853 12316 -819
rect 12350 -853 12384 -819
rect 12418 -853 12452 -819
rect 12486 -853 12520 -819
rect 12554 -853 12588 -819
rect 12622 -853 12656 -819
rect 12690 -853 12724 -819
rect 12758 -853 12797 -819
rect 12277 -890 12797 -853
rect 12277 -924 12316 -890
rect 12350 -924 12384 -890
rect 12418 -924 12452 -890
rect 12486 -924 12520 -890
rect 12554 -924 12588 -890
rect 12622 -924 12656 -890
rect 12690 -924 12724 -890
rect 12758 -924 12797 -890
rect 12277 -961 12797 -924
rect 12277 -995 12316 -961
rect 12350 -995 12384 -961
rect 12418 -995 12452 -961
rect 12486 -995 12520 -961
rect 12554 -995 12588 -961
rect 12622 -995 12656 -961
rect 12690 -995 12724 -961
rect 12758 -995 12797 -961
<< mvpsubdiff >>
rect 800 8767 907 8791
rect 834 8757 907 8767
rect 941 8757 975 8791
rect 1009 8757 1043 8791
rect 1077 8757 1111 8791
rect 1145 8757 1179 8791
rect 1213 8757 1247 8791
rect 1281 8757 1315 8791
rect 1349 8757 1383 8791
rect 1417 8757 1451 8791
rect 1485 8757 1519 8791
rect 1553 8757 1587 8791
rect 1621 8757 1655 8791
rect 1689 8757 1723 8791
rect 1757 8757 1791 8791
rect 1825 8757 1859 8791
rect 1893 8757 1927 8791
rect 1961 8757 1995 8791
rect 2029 8757 2063 8791
rect 2097 8757 2131 8791
rect 2165 8757 2199 8791
rect 2233 8757 2267 8791
rect 2301 8757 2335 8791
rect 2369 8757 2403 8791
rect 2437 8757 2471 8791
rect 2505 8757 2539 8791
rect 2573 8757 2607 8791
rect 2641 8757 2675 8791
rect 2709 8757 2743 8791
rect 2777 8757 2811 8791
rect 2845 8757 2879 8791
rect 2913 8757 2947 8791
rect 2981 8757 3015 8791
rect 3049 8757 3083 8791
rect 3117 8757 3151 8791
rect 3185 8757 3219 8791
rect 3253 8757 3287 8791
rect 3321 8757 3355 8791
rect 3389 8757 3423 8791
rect 3457 8757 3491 8791
rect 3525 8757 3559 8791
rect 3593 8757 3627 8791
rect 3661 8757 3695 8791
rect 3729 8757 3763 8791
rect 3797 8757 3831 8791
rect 3865 8757 3899 8791
rect 3933 8757 3967 8791
rect 4001 8757 4035 8791
rect 4069 8757 4103 8791
rect 4137 8757 4171 8791
rect 4205 8757 4239 8791
rect 4273 8757 4307 8791
rect 4341 8757 4375 8791
rect 4409 8757 4443 8791
rect 4477 8757 4511 8791
rect 4545 8757 4579 8791
rect 4613 8757 4647 8791
rect 4681 8757 4715 8791
rect 4749 8757 4773 8791
rect 800 8699 834 8733
rect 800 8631 834 8665
rect 800 8563 834 8597
rect 800 8495 834 8529
rect 800 8427 834 8461
rect 800 8359 834 8393
rect 800 8291 834 8325
rect 800 8223 834 8257
rect 800 8155 834 8189
rect 800 8087 834 8121
rect 800 8019 834 8053
rect 800 7951 834 7985
rect 800 7883 834 7917
rect 800 7815 834 7849
rect 800 7747 834 7781
rect 800 7679 834 7713
rect 800 7611 834 7645
rect 800 7543 834 7577
rect 800 7475 834 7509
rect 800 7407 834 7441
rect 800 7339 834 7373
rect 800 7271 834 7305
rect 800 7203 834 7237
rect 800 7078 834 7169
rect 800 7044 841 7078
rect 875 7044 909 7078
rect 943 7044 977 7078
rect 1011 7044 1045 7078
rect 1079 7044 1113 7078
rect 1147 7044 1181 7078
rect 1215 7044 1249 7078
rect 1283 7044 1317 7078
rect 1351 7044 1385 7078
rect 1419 7044 1453 7078
rect 1487 7044 1521 7078
rect 1555 7044 1589 7078
rect 1623 7044 1657 7078
rect 1691 7044 1725 7078
rect 1759 7044 1793 7078
rect 1827 7044 1861 7078
rect 1895 7044 1929 7078
rect 1963 7044 1997 7078
rect 2031 7044 2065 7078
rect 2099 7044 2133 7078
rect 2167 7044 2201 7078
rect 2235 7044 2269 7078
rect 2303 7044 2337 7078
rect 2371 7044 2405 7078
rect 2439 7044 2473 7078
rect 2507 7044 2541 7078
rect 2575 7044 2609 7078
rect 2643 7044 2677 7078
rect 2711 7044 2745 7078
rect 2779 7044 2813 7078
rect 2847 7044 2881 7078
rect 2915 7044 2949 7078
rect 2983 7044 3017 7078
rect 3051 7044 3085 7078
rect 3119 7044 3153 7078
rect 3187 7044 3221 7078
rect 3255 7044 3289 7078
rect 3323 7044 3357 7078
rect 3391 7044 3425 7078
rect 3459 7044 3493 7078
rect 3527 7044 3561 7078
rect 3595 7044 3629 7078
rect 3663 7044 3697 7078
rect 3731 7044 3765 7078
rect 3799 7044 3833 7078
rect 3867 7044 3901 7078
rect 3935 7044 3969 7078
rect 4003 7044 4037 7078
rect 4071 7044 4105 7078
rect 4139 7044 4173 7078
rect 4207 7044 4241 7078
rect 4275 7044 4309 7078
rect 4343 7044 4377 7078
rect 4411 7044 4445 7078
rect 4479 7044 4513 7078
rect 4547 7044 4581 7078
rect 4615 7044 4649 7078
rect 4683 7044 4731 7078
rect 4411 7007 4731 7044
rect 4411 6973 4446 7007
rect 4480 6973 4518 7007
rect 4552 6973 4590 7007
rect 4624 6973 4662 7007
rect 4696 6973 4731 7007
rect 4411 6939 4731 6973
rect 4411 6905 4446 6939
rect 4480 6905 4518 6939
rect 4552 6905 4590 6939
rect 4624 6905 4662 6939
rect 4696 6905 4731 6939
rect 4411 6871 4731 6905
rect 4411 6837 4446 6871
rect 4480 6837 4518 6871
rect 4552 6837 4590 6871
rect 4624 6837 4662 6871
rect 4696 6837 4731 6871
rect 4411 6803 4731 6837
rect 4411 6769 4446 6803
rect 4480 6769 4518 6803
rect 4552 6769 4590 6803
rect 4624 6769 4662 6803
rect 4696 6769 4731 6803
rect -874 6759 925 6766
rect -874 6725 -850 6759
rect -816 6725 -781 6759
rect -747 6725 -712 6759
rect -678 6725 -643 6759
rect -609 6725 -574 6759
rect -540 6725 -505 6759
rect -471 6725 -436 6759
rect -402 6725 -367 6759
rect -333 6725 -298 6759
rect -264 6725 -229 6759
rect -195 6725 -160 6759
rect -126 6725 -91 6759
rect -57 6725 -22 6759
rect 12 6725 47 6759
rect 81 6725 116 6759
rect 150 6725 185 6759
rect 219 6725 254 6759
rect 288 6725 323 6759
rect 357 6725 391 6759
rect 425 6725 459 6759
rect 493 6725 527 6759
rect 561 6725 595 6759
rect 629 6725 663 6759
rect 697 6725 731 6759
rect 765 6725 799 6759
rect 833 6725 867 6759
rect 901 6725 925 6759
rect -874 6689 925 6725
rect -874 6655 -850 6689
rect -816 6655 -781 6689
rect -747 6655 -712 6689
rect -678 6655 -643 6689
rect -609 6655 -574 6689
rect -540 6655 -505 6689
rect -471 6655 -436 6689
rect -402 6655 -367 6689
rect -333 6655 -298 6689
rect -264 6655 -229 6689
rect -195 6655 -160 6689
rect -126 6655 -91 6689
rect -57 6655 -22 6689
rect 12 6655 47 6689
rect 81 6655 116 6689
rect 150 6655 185 6689
rect 219 6655 254 6689
rect 288 6655 323 6689
rect 357 6655 391 6689
rect 425 6655 459 6689
rect 493 6655 527 6689
rect 561 6655 595 6689
rect 629 6655 663 6689
rect 697 6655 731 6689
rect 765 6655 799 6689
rect 833 6655 867 6689
rect 901 6655 925 6689
rect -874 6619 925 6655
rect -874 6585 -850 6619
rect -816 6585 -781 6619
rect -747 6585 -712 6619
rect -678 6585 -643 6619
rect -609 6585 -574 6619
rect -540 6585 -505 6619
rect -471 6585 -436 6619
rect -402 6585 -367 6619
rect -333 6585 -298 6619
rect -264 6585 -229 6619
rect -195 6585 -160 6619
rect -126 6585 -91 6619
rect -57 6585 -22 6619
rect 12 6585 47 6619
rect 81 6585 116 6619
rect 150 6585 185 6619
rect 219 6585 254 6619
rect 288 6585 323 6619
rect 357 6585 391 6619
rect 425 6585 459 6619
rect 493 6585 527 6619
rect 561 6585 595 6619
rect 629 6585 663 6619
rect 697 6585 731 6619
rect 765 6585 799 6619
rect 833 6585 867 6619
rect 901 6585 925 6619
rect -874 6549 925 6585
rect -874 6515 -850 6549
rect -816 6515 -781 6549
rect -747 6515 -712 6549
rect -678 6515 -643 6549
rect -609 6515 -574 6549
rect -540 6515 -505 6549
rect -471 6515 -436 6549
rect -402 6515 -367 6549
rect -333 6515 -298 6549
rect -264 6515 -229 6549
rect -195 6515 -160 6549
rect -126 6515 -91 6549
rect -57 6515 -22 6549
rect 12 6515 47 6549
rect 81 6515 116 6549
rect 150 6515 185 6549
rect 219 6515 254 6549
rect 288 6515 323 6549
rect 357 6515 391 6549
rect 425 6515 459 6549
rect 493 6515 527 6549
rect 561 6515 595 6549
rect 629 6515 663 6549
rect 697 6515 731 6549
rect 765 6515 799 6549
rect 833 6515 867 6549
rect 901 6515 925 6549
rect -874 6479 925 6515
rect -874 6445 -850 6479
rect -816 6445 -781 6479
rect -747 6445 -712 6479
rect -678 6445 -643 6479
rect -609 6445 -574 6479
rect -540 6445 -505 6479
rect -471 6445 -436 6479
rect -402 6445 -367 6479
rect -333 6445 -298 6479
rect -264 6445 -229 6479
rect -195 6445 -160 6479
rect -126 6445 -91 6479
rect -57 6445 -22 6479
rect 12 6445 47 6479
rect 81 6445 116 6479
rect 150 6445 185 6479
rect 219 6445 254 6479
rect 288 6445 323 6479
rect 357 6445 391 6479
rect 425 6445 459 6479
rect 493 6445 527 6479
rect 561 6445 595 6479
rect 629 6445 663 6479
rect 697 6445 731 6479
rect 765 6445 799 6479
rect 833 6445 867 6479
rect 901 6445 925 6479
rect -874 6409 925 6445
rect -874 6375 -850 6409
rect -816 6375 -781 6409
rect -747 6375 -712 6409
rect -678 6375 -643 6409
rect -609 6375 -574 6409
rect -540 6375 -505 6409
rect -471 6375 -436 6409
rect -402 6375 -367 6409
rect -333 6375 -298 6409
rect -264 6375 -229 6409
rect -195 6375 -160 6409
rect -126 6375 -91 6409
rect -57 6375 -22 6409
rect 12 6375 47 6409
rect 81 6375 116 6409
rect 150 6375 185 6409
rect 219 6375 254 6409
rect 288 6375 323 6409
rect 357 6375 391 6409
rect 425 6375 459 6409
rect 493 6375 527 6409
rect 561 6375 595 6409
rect 629 6375 663 6409
rect 697 6375 731 6409
rect 765 6375 799 6409
rect 833 6375 867 6409
rect 901 6375 925 6409
rect -874 6339 925 6375
rect -874 6305 -850 6339
rect -816 6305 -781 6339
rect -747 6305 -712 6339
rect -678 6305 -643 6339
rect -609 6305 -574 6339
rect -540 6305 -505 6339
rect -471 6305 -436 6339
rect -402 6305 -367 6339
rect -333 6305 -298 6339
rect -264 6305 -229 6339
rect -195 6305 -160 6339
rect -126 6305 -91 6339
rect -57 6305 -22 6339
rect 12 6305 47 6339
rect 81 6305 116 6339
rect 150 6305 185 6339
rect 219 6305 254 6339
rect 288 6305 323 6339
rect 357 6305 391 6339
rect 425 6305 459 6339
rect 493 6305 527 6339
rect 561 6305 595 6339
rect 629 6305 663 6339
rect 697 6305 731 6339
rect 765 6305 799 6339
rect 833 6305 867 6339
rect 901 6305 925 6339
rect -874 6269 925 6305
rect -874 6235 -850 6269
rect -816 6235 -781 6269
rect -747 6235 -712 6269
rect -678 6235 -643 6269
rect -609 6235 -574 6269
rect -540 6235 -505 6269
rect -471 6235 -436 6269
rect -402 6235 -367 6269
rect -333 6235 -298 6269
rect -264 6235 -229 6269
rect -195 6235 -160 6269
rect -126 6235 -91 6269
rect -57 6235 -22 6269
rect 12 6235 47 6269
rect 81 6235 116 6269
rect 150 6235 185 6269
rect 219 6235 254 6269
rect 288 6235 323 6269
rect 357 6235 391 6269
rect 425 6235 459 6269
rect 493 6235 527 6269
rect 561 6235 595 6269
rect 629 6235 663 6269
rect 697 6235 731 6269
rect 765 6235 799 6269
rect 833 6235 867 6269
rect 901 6235 925 6269
rect -874 6199 925 6235
rect -874 6165 -850 6199
rect -816 6165 -781 6199
rect -747 6165 -712 6199
rect -678 6165 -643 6199
rect -609 6165 -574 6199
rect -540 6165 -505 6199
rect -471 6165 -436 6199
rect -402 6165 -367 6199
rect -333 6165 -298 6199
rect -264 6165 -229 6199
rect -195 6165 -160 6199
rect -126 6165 -91 6199
rect -57 6165 -22 6199
rect 12 6165 47 6199
rect 81 6165 116 6199
rect 150 6165 185 6199
rect 219 6165 254 6199
rect 288 6165 323 6199
rect 357 6165 391 6199
rect 425 6165 459 6199
rect 493 6165 527 6199
rect 561 6165 595 6199
rect 629 6165 663 6199
rect 697 6165 731 6199
rect 765 6165 799 6199
rect 833 6165 867 6199
rect 901 6165 925 6199
rect -874 6129 925 6165
rect -874 6095 -850 6129
rect -816 6095 -781 6129
rect -747 6095 -712 6129
rect -678 6095 -643 6129
rect -609 6095 -574 6129
rect -540 6095 -505 6129
rect -471 6095 -436 6129
rect -402 6095 -367 6129
rect -333 6095 -298 6129
rect -264 6095 -229 6129
rect -195 6095 -160 6129
rect -126 6095 -91 6129
rect -57 6095 -22 6129
rect 12 6095 47 6129
rect 81 6095 116 6129
rect 150 6095 185 6129
rect 219 6095 254 6129
rect 288 6095 323 6129
rect 357 6095 391 6129
rect 425 6095 459 6129
rect 493 6095 527 6129
rect 561 6095 595 6129
rect 629 6095 663 6129
rect 697 6095 731 6129
rect 765 6095 799 6129
rect 833 6095 867 6129
rect 901 6095 925 6129
rect -874 6088 925 6095
rect 4411 6735 4731 6769
rect 4411 6701 4446 6735
rect 4480 6701 4518 6735
rect 4552 6701 4590 6735
rect 4624 6701 4662 6735
rect 4696 6701 4731 6735
rect 4411 6667 4731 6701
rect 4411 6633 4446 6667
rect 4480 6633 4518 6667
rect 4552 6633 4590 6667
rect 4624 6633 4662 6667
rect 4696 6633 4731 6667
rect 4411 6599 4731 6633
rect 4411 6565 4446 6599
rect 4480 6565 4518 6599
rect 4552 6565 4590 6599
rect 4624 6565 4662 6599
rect 4696 6565 4731 6599
rect 4411 6531 4731 6565
rect 4411 6497 4446 6531
rect 4480 6497 4518 6531
rect 4552 6497 4590 6531
rect 4624 6497 4662 6531
rect 4696 6497 4731 6531
rect 4411 6463 4731 6497
rect 4411 6429 4446 6463
rect 4480 6429 4518 6463
rect 4552 6429 4590 6463
rect 4624 6429 4662 6463
rect 4696 6429 4731 6463
rect 4411 6395 4731 6429
rect 4411 6361 4446 6395
rect 4480 6361 4518 6395
rect 4552 6361 4590 6395
rect 4624 6361 4662 6395
rect 4696 6361 4731 6395
rect 4411 6327 4731 6361
rect 4411 6293 4446 6327
rect 4480 6293 4518 6327
rect 4552 6293 4590 6327
rect 4624 6293 4662 6327
rect 4696 6293 4731 6327
rect 4411 6259 4731 6293
rect 4411 6225 4446 6259
rect 4480 6225 4518 6259
rect 4552 6225 4590 6259
rect 4624 6225 4662 6259
rect 4696 6225 4731 6259
rect 4411 6191 4731 6225
rect 4411 6157 4446 6191
rect 4480 6157 4518 6191
rect 4552 6157 4590 6191
rect 4624 6157 4662 6191
rect 4696 6157 4731 6191
rect 4411 6123 4731 6157
rect 4411 6089 4446 6123
rect 4480 6089 4518 6123
rect 4552 6089 4590 6123
rect 4624 6089 4662 6123
rect 4696 6089 4731 6123
rect 4411 6055 4731 6089
rect 4411 6021 4446 6055
rect 4480 6021 4518 6055
rect 4552 6021 4590 6055
rect 4624 6021 4662 6055
rect 4696 6021 4731 6055
rect 4411 5987 4731 6021
rect 4411 5953 4446 5987
rect 4480 5953 4518 5987
rect 4552 5953 4590 5987
rect 4624 5953 4662 5987
rect 4696 5953 4731 5987
rect 4411 5919 4731 5953
rect 4411 5885 4446 5919
rect 4480 5885 4518 5919
rect 4552 5885 4590 5919
rect 4624 5885 4662 5919
rect 4696 5885 4731 5919
rect 4411 5850 4731 5885
rect 4411 5816 4446 5850
rect 4480 5816 4518 5850
rect 4552 5816 4590 5850
rect 4624 5816 4662 5850
rect 4696 5816 4731 5850
rect 4411 5779 4731 5816
rect 4067 5745 4102 5779
rect 4136 5745 4172 5779
rect 4206 5745 4242 5779
rect 4276 5745 4312 5779
rect 4346 5745 4382 5779
rect 4416 5745 4452 5779
rect 4486 5745 4522 5779
rect 4556 5745 4592 5779
rect 4626 5745 4662 5779
rect 4696 5745 4731 5779
rect 4067 5710 4731 5745
rect 4067 5676 4102 5710
rect 4136 5676 4172 5710
rect 4206 5676 4242 5710
rect 4276 5676 4312 5710
rect 4346 5676 4382 5710
rect 4416 5676 4452 5710
rect 4486 5676 4522 5710
rect 4556 5676 4592 5710
rect 4626 5676 4662 5710
rect 4696 5676 4731 5710
rect 4067 5641 4731 5676
rect 4067 5607 4102 5641
rect 4136 5607 4172 5641
rect 4206 5607 4242 5641
rect 4276 5607 4312 5641
rect 4346 5607 4382 5641
rect 4416 5607 4452 5641
rect 4486 5607 4522 5641
rect 4556 5607 4592 5641
rect 4626 5607 4662 5641
rect 4696 5607 4731 5641
rect 4067 5572 4731 5607
rect 4067 5538 4102 5572
rect 4136 5538 4172 5572
rect 4206 5538 4242 5572
rect 4276 5538 4312 5572
rect 4346 5538 4382 5572
rect 4416 5538 4452 5572
rect 4486 5538 4522 5572
rect 4556 5538 4592 5572
rect 4626 5538 4662 5572
rect 4696 5538 4731 5572
rect 4067 5503 4731 5538
rect 4067 5469 4102 5503
rect 4136 5469 4172 5503
rect 4206 5469 4242 5503
rect 4276 5469 4312 5503
rect 4346 5469 4382 5503
rect 4416 5469 4452 5503
rect 4486 5469 4522 5503
rect 4556 5469 4592 5503
rect 4626 5469 4662 5503
rect 4696 5469 4731 5503
rect 4067 5434 4731 5469
rect 4067 5400 4102 5434
rect 4136 5400 4172 5434
rect 4206 5400 4242 5434
rect 4276 5400 4312 5434
rect 4346 5400 4382 5434
rect 4416 5400 4452 5434
rect 4486 5400 4522 5434
rect 4556 5400 4592 5434
rect 4626 5400 4662 5434
rect 4696 5400 4731 5434
rect 4067 5365 4731 5400
rect 4067 5331 4102 5365
rect 4136 5331 4172 5365
rect 4206 5331 4242 5365
rect 4276 5331 4312 5365
rect 4346 5331 4382 5365
rect 4416 5331 4452 5365
rect 4486 5331 4522 5365
rect 4556 5331 4592 5365
rect 4626 5331 4662 5365
rect 4696 5331 4731 5365
rect 4067 5296 4731 5331
rect 4067 5262 4102 5296
rect 4136 5262 4172 5296
rect 4206 5262 4242 5296
rect 4276 5262 4312 5296
rect 4346 5262 4382 5296
rect 4416 5262 4452 5296
rect 4486 5262 4522 5296
rect 4556 5262 4592 5296
rect 4626 5262 4662 5296
rect 4696 5262 4731 5296
rect 4067 5227 4731 5262
rect 4067 5193 4102 5227
rect 4136 5193 4172 5227
rect 4206 5193 4242 5227
rect 4276 5193 4312 5227
rect 4346 5193 4382 5227
rect 4416 5193 4452 5227
rect 4486 5193 4522 5227
rect 4556 5193 4592 5227
rect 4626 5193 4662 5227
rect 4696 5193 4731 5227
rect 4067 5158 4731 5193
rect 4067 5124 4102 5158
rect 4136 5124 4172 5158
rect 4206 5124 4242 5158
rect 4276 5124 4312 5158
rect 4346 5124 4382 5158
rect 4416 5124 4452 5158
rect 4486 5124 4522 5158
rect 4556 5124 4592 5158
rect 4626 5124 4662 5158
rect 4696 5124 4731 5158
rect 4067 5089 4731 5124
rect 4067 5055 4102 5089
rect 4136 5055 4172 5089
rect 4206 5055 4242 5089
rect 4276 5055 4312 5089
rect 4346 5055 4382 5089
rect 4416 5055 4452 5089
rect 4486 5055 4522 5089
rect 4556 5055 4592 5089
rect 4626 5055 4662 5089
rect 4696 5055 4731 5089
rect 4067 5019 4731 5055
rect 4067 4985 4102 5019
rect 4136 4985 4172 5019
rect 4206 4985 4242 5019
rect 4276 4985 4312 5019
rect 4346 4985 4382 5019
rect 4416 4985 4452 5019
rect 4486 4985 4522 5019
rect 4556 4985 4592 5019
rect 4626 4985 4662 5019
rect 4696 4985 4731 5019
rect 4067 4949 4731 4985
rect 4067 4915 4102 4949
rect 4136 4915 4172 4949
rect 4206 4915 4242 4949
rect 4276 4915 4312 4949
rect 4346 4915 4382 4949
rect 4416 4915 4452 4949
rect 4486 4915 4522 4949
rect 4556 4915 4592 4949
rect 4626 4915 4662 4949
rect 4696 4915 4731 4949
rect 4067 4879 4731 4915
rect 4067 4845 4102 4879
rect 4136 4845 4172 4879
rect 4206 4845 4242 4879
rect 4276 4845 4312 4879
rect 4346 4845 4382 4879
rect 4416 4845 4452 4879
rect 4486 4845 4522 4879
rect 4556 4845 4592 4879
rect 4626 4845 4662 4879
rect 4696 4845 4731 4879
rect 4067 4809 4731 4845
rect 4067 4775 4102 4809
rect 4136 4775 4172 4809
rect 4206 4775 4242 4809
rect 4276 4775 4312 4809
rect 4346 4775 4382 4809
rect 4416 4775 4452 4809
rect 4486 4775 4522 4809
rect 4556 4775 4592 4809
rect 4626 4775 4662 4809
rect 4696 4775 4731 4809
rect 4067 4739 4731 4775
rect 4067 4705 4102 4739
rect 4136 4705 4172 4739
rect 4206 4705 4242 4739
rect 4276 4705 4312 4739
rect 4346 4705 4382 4739
rect 4416 4705 4452 4739
rect 4486 4705 4522 4739
rect 4556 4705 4592 4739
rect 4626 4705 4662 4739
rect 4696 4705 4731 4739
rect 4067 4669 4731 4705
rect 4067 4635 4102 4669
rect 4136 4635 4172 4669
rect 4206 4635 4242 4669
rect 4276 4635 4312 4669
rect 4346 4635 4382 4669
rect 4416 4635 4452 4669
rect 4486 4635 4522 4669
rect 4556 4635 4592 4669
rect 4626 4635 4662 4669
rect 4696 4635 4731 4669
rect 4067 4599 4731 4635
rect 4067 4565 4102 4599
rect 4136 4565 4172 4599
rect 4206 4565 4242 4599
rect 4276 4565 4312 4599
rect 4346 4565 4382 4599
rect 4416 4565 4452 4599
rect 4486 4565 4522 4599
rect 4556 4565 4592 4599
rect 4626 4565 4662 4599
rect 4696 4565 4731 4599
rect 4067 4529 4731 4565
rect 4067 4495 4102 4529
rect 4136 4495 4172 4529
rect 4206 4495 4242 4529
rect 4276 4495 4312 4529
rect 4346 4495 4382 4529
rect 4416 4495 4452 4529
rect 4486 4495 4522 4529
rect 4556 4495 4592 4529
rect 4626 4495 4662 4529
rect 4696 4495 4731 4529
rect 4067 4459 4731 4495
rect 4067 4425 4102 4459
rect 4136 4425 4172 4459
rect 4206 4425 4242 4459
rect 4276 4425 4312 4459
rect 4346 4425 4382 4459
rect 4416 4425 4452 4459
rect 4486 4425 4522 4459
rect 4556 4425 4592 4459
rect 4626 4425 4662 4459
rect 4696 4425 4731 4459
rect 4067 4389 4731 4425
rect 4067 4355 4102 4389
rect 4136 4355 4172 4389
rect 4206 4355 4242 4389
rect 4276 4355 4312 4389
rect 4346 4355 4382 4389
rect 4416 4355 4452 4389
rect 4486 4355 4522 4389
rect 4556 4355 4592 4389
rect 4626 4355 4662 4389
rect 4696 4355 4731 4389
rect 4067 4319 4731 4355
rect 4067 4285 4102 4319
rect 4136 4285 4172 4319
rect 4206 4285 4242 4319
rect 4276 4285 4312 4319
rect 4346 4285 4382 4319
rect 4416 4285 4452 4319
rect 4486 4285 4522 4319
rect 4556 4285 4592 4319
rect 4626 4285 4662 4319
rect 4696 4285 4731 4319
rect 4067 4249 4731 4285
rect 4067 4215 4102 4249
rect 4136 4215 4172 4249
rect 4206 4215 4242 4249
rect 4276 4215 4312 4249
rect 4346 4215 4382 4249
rect 4416 4215 4452 4249
rect 4486 4215 4522 4249
rect 4556 4215 4592 4249
rect 4626 4215 4662 4249
rect 4696 4216 4731 4249
rect 4696 4215 8292 4216
rect 4067 4182 8292 4215
rect 4067 4179 4731 4182
rect 4067 4145 4102 4179
rect 4136 4145 4172 4179
rect 4206 4145 4242 4179
rect 4276 4145 4312 4179
rect 4346 4145 4382 4179
rect 4416 4145 4452 4179
rect 4486 4145 4522 4179
rect 4556 4145 4592 4179
rect 4626 4145 4662 4179
rect 4696 4148 4731 4179
rect 4765 4148 4801 4182
rect 4835 4148 4871 4182
rect 4905 4148 4941 4182
rect 4975 4148 5011 4182
rect 5045 4148 5081 4182
rect 5115 4148 5151 4182
rect 5185 4148 5221 4182
rect 5255 4148 5291 4182
rect 5325 4148 5360 4182
rect 5394 4148 5429 4182
rect 5463 4148 5498 4182
rect 5532 4148 5567 4182
rect 5601 4148 5636 4182
rect 5670 4148 5705 4182
rect 5739 4148 5774 4182
rect 5808 4148 5843 4182
rect 5877 4148 5912 4182
rect 5946 4148 5981 4182
rect 6015 4148 6050 4182
rect 6084 4148 6119 4182
rect 6153 4148 6188 4182
rect 6222 4148 6257 4182
rect 6291 4148 6326 4182
rect 6360 4148 6395 4182
rect 6429 4148 6464 4182
rect 6498 4148 6533 4182
rect 6567 4148 6602 4182
rect 6636 4148 6671 4182
rect 6705 4148 6740 4182
rect 6774 4148 6809 4182
rect 6843 4148 6878 4182
rect 6912 4148 6947 4182
rect 6981 4148 7016 4182
rect 7050 4148 7085 4182
rect 7119 4148 7154 4182
rect 7188 4148 7223 4182
rect 7257 4148 7292 4182
rect 7326 4148 7361 4182
rect 7395 4148 7430 4182
rect 7464 4148 7499 4182
rect 7533 4148 7568 4182
rect 7602 4148 7637 4182
rect 7671 4148 7706 4182
rect 7740 4148 7775 4182
rect 7809 4148 7844 4182
rect 7878 4148 7913 4182
rect 7947 4148 7982 4182
rect 8016 4148 8051 4182
rect 8085 4148 8120 4182
rect 8154 4148 8189 4182
rect 8223 4148 8258 4182
rect 4696 4145 8292 4148
rect 4067 4109 8292 4145
rect 4067 4075 4102 4109
rect 4136 4075 4172 4109
rect 4206 4075 4242 4109
rect 4276 4075 4312 4109
rect 4346 4075 4382 4109
rect 4416 4075 4452 4109
rect 4486 4075 4522 4109
rect 4556 4075 4592 4109
rect 4626 4075 4662 4109
rect 4696 4084 8292 4109
rect 4696 4075 4731 4084
rect 4067 4050 4731 4075
rect 4765 4050 4801 4084
rect 4835 4050 4871 4084
rect 4905 4050 4941 4084
rect 4975 4050 5011 4084
rect 5045 4050 5081 4084
rect 5115 4050 5151 4084
rect 5185 4050 5221 4084
rect 5255 4050 5291 4084
rect 5325 4050 5360 4084
rect 5394 4050 5429 4084
rect 5463 4050 5498 4084
rect 5532 4050 5567 4084
rect 5601 4050 5636 4084
rect 5670 4050 5705 4084
rect 5739 4050 5774 4084
rect 5808 4050 5843 4084
rect 5877 4050 5912 4084
rect 5946 4050 5981 4084
rect 6015 4050 6050 4084
rect 6084 4050 6119 4084
rect 6153 4050 6188 4084
rect 6222 4050 6257 4084
rect 6291 4050 6326 4084
rect 6360 4050 6395 4084
rect 6429 4050 6464 4084
rect 6498 4050 6533 4084
rect 6567 4050 6602 4084
rect 6636 4050 6671 4084
rect 6705 4050 6740 4084
rect 6774 4050 6809 4084
rect 6843 4050 6878 4084
rect 6912 4050 6947 4084
rect 6981 4050 7016 4084
rect 7050 4050 7085 4084
rect 7119 4050 7154 4084
rect 7188 4050 7223 4084
rect 7257 4050 7292 4084
rect 7326 4050 7361 4084
rect 7395 4050 7430 4084
rect 7464 4050 7499 4084
rect 7533 4050 7568 4084
rect 7602 4050 7637 4084
rect 7671 4050 7706 4084
rect 7740 4050 7775 4084
rect 7809 4050 7844 4084
rect 7878 4050 7913 4084
rect 7947 4050 7982 4084
rect 8016 4050 8051 4084
rect 8085 4050 8120 4084
rect 8154 4050 8189 4084
rect 8223 4050 8258 4084
rect 4067 4039 8292 4050
rect 4067 4005 4102 4039
rect 4136 4005 4172 4039
rect 4206 4005 4242 4039
rect 4276 4005 4312 4039
rect 4346 4005 4382 4039
rect 4416 4005 4452 4039
rect 4486 4005 4522 4039
rect 4556 4005 4592 4039
rect 4626 4005 4662 4039
rect 4696 4016 8292 4039
rect 4696 4013 9456 4016
rect 4696 4005 4974 4013
rect 4067 3979 4974 4005
rect 5008 3979 5043 4013
rect 5077 3979 5112 4013
rect 5146 3979 5181 4013
rect 5215 3979 5250 4013
rect 5284 3979 5319 4013
rect 5353 3979 5388 4013
rect 5422 3979 5457 4013
rect 5491 3979 5526 4013
rect 5560 3979 5595 4013
rect 5629 3979 5664 4013
rect 5698 3979 5733 4013
rect 5767 3979 5802 4013
rect 5836 3979 5871 4013
rect 5905 3979 5940 4013
rect 5974 3979 6009 4013
rect 6043 3979 6078 4013
rect 6112 3979 6147 4013
rect 6181 3979 6216 4013
rect 6250 3979 6285 4013
rect 6319 3979 6354 4013
rect 6388 3979 6423 4013
rect 6457 3979 6492 4013
rect 6526 3979 6561 4013
rect 6595 3979 6630 4013
rect 6664 3979 6699 4013
rect 6733 3979 6768 4013
rect 6802 3979 6837 4013
rect 6871 3979 6906 4013
rect 6940 3979 6975 4013
rect 7009 3979 7044 4013
rect 7078 3979 7113 4013
rect 7147 3979 7182 4013
rect 7216 3979 7251 4013
rect 7285 3979 7320 4013
rect 7354 3979 7389 4013
rect 7423 3979 7458 4013
rect 7492 3979 7527 4013
rect 7561 3979 7596 4013
rect 7630 3979 7665 4013
rect 7699 3979 7734 4013
rect 7768 3979 7803 4013
rect 7837 3979 7872 4013
rect 7906 3979 7941 4013
rect 7975 3979 8010 4013
rect 8044 3979 8079 4013
rect 8113 3979 8148 4013
rect 8182 3979 8217 4013
rect 8251 3979 8286 4013
rect 8320 3979 8355 4013
rect 8389 3979 8424 4013
rect 8458 3979 8493 4013
rect 8527 3979 8562 4013
rect 8596 3979 8631 4013
rect 8665 3979 8700 4013
rect 8734 3979 8769 4013
rect 8803 3979 8838 4013
rect 8872 3979 8907 4013
rect 8941 3979 8976 4013
rect 9010 3979 9045 4013
rect 9079 3979 9114 4013
rect 9148 3979 9183 4013
rect 9217 3979 9252 4013
rect 9286 3979 9320 4013
rect 9354 3979 9388 4013
rect 9422 3979 9456 4013
rect 4067 3969 9456 3979
rect 4067 3935 4102 3969
rect 4136 3935 4172 3969
rect 4206 3935 4242 3969
rect 4276 3935 4312 3969
rect 4346 3935 4382 3969
rect 4416 3935 4452 3969
rect 4486 3935 4522 3969
rect 4556 3935 4592 3969
rect 4626 3935 4662 3969
rect 4696 3937 9456 3969
rect 4696 3935 4974 3937
rect 4067 3925 4974 3935
rect 3864 3903 4974 3925
rect 5008 3903 5043 3937
rect 5077 3903 5112 3937
rect 5146 3903 5181 3937
rect 5215 3903 5250 3937
rect 5284 3903 5319 3937
rect 5353 3903 5388 3937
rect 5422 3903 5457 3937
rect 5491 3903 5526 3937
rect 5560 3903 5595 3937
rect 5629 3903 5664 3937
rect 5698 3903 5733 3937
rect 5767 3903 5802 3937
rect 5836 3903 5871 3937
rect 5905 3903 5940 3937
rect 5974 3903 6009 3937
rect 6043 3903 6078 3937
rect 6112 3903 6147 3937
rect 6181 3903 6216 3937
rect 6250 3903 6285 3937
rect 6319 3903 6354 3937
rect 6388 3903 6423 3937
rect 6457 3903 6492 3937
rect 6526 3903 6561 3937
rect 6595 3903 6630 3937
rect 6664 3903 6699 3937
rect 6733 3903 6768 3937
rect 6802 3903 6837 3937
rect 6871 3903 6906 3937
rect 6940 3903 6975 3937
rect 7009 3903 7044 3937
rect 7078 3903 7113 3937
rect 7147 3903 7182 3937
rect 7216 3903 7251 3937
rect 7285 3903 7320 3937
rect 7354 3903 7389 3937
rect 7423 3903 7458 3937
rect 7492 3903 7527 3937
rect 7561 3903 7596 3937
rect 7630 3903 7665 3937
rect 7699 3903 7734 3937
rect 7768 3903 7803 3937
rect 7837 3903 7872 3937
rect 7906 3903 7941 3937
rect 7975 3903 8010 3937
rect 8044 3903 8079 3937
rect 8113 3903 8148 3937
rect 8182 3903 8217 3937
rect 8251 3903 8286 3937
rect 8320 3903 8355 3937
rect 8389 3903 8424 3937
rect 8458 3903 8493 3937
rect 8527 3903 8562 3937
rect 8596 3903 8631 3937
rect 8665 3903 8700 3937
rect 8734 3903 8769 3937
rect 8803 3903 8838 3937
rect 8872 3903 8907 3937
rect 8941 3903 8976 3937
rect 9010 3903 9045 3937
rect 9079 3903 9114 3937
rect 9148 3903 9183 3937
rect 9217 3903 9252 3937
rect 9286 3903 9320 3937
rect 9354 3903 9388 3937
rect 9422 3903 9456 3937
rect 3864 3901 9456 3903
rect 3864 2167 3875 3901
rect 4929 3861 9456 3901
rect 4929 3827 4974 3861
rect 5008 3827 5043 3861
rect 5077 3827 5112 3861
rect 5146 3827 5181 3861
rect 5215 3827 5250 3861
rect 5284 3827 5319 3861
rect 5353 3827 5388 3861
rect 5422 3827 5457 3861
rect 5491 3827 5526 3861
rect 5560 3827 5595 3861
rect 5629 3827 5664 3861
rect 5698 3827 5733 3861
rect 5767 3827 5802 3861
rect 5836 3827 5871 3861
rect 5905 3827 5940 3861
rect 5974 3827 6009 3861
rect 6043 3827 6078 3861
rect 6112 3827 6147 3861
rect 6181 3827 6216 3861
rect 6250 3827 6285 3861
rect 6319 3827 6354 3861
rect 6388 3827 6423 3861
rect 6457 3827 6492 3861
rect 6526 3827 6561 3861
rect 6595 3827 6630 3861
rect 6664 3827 6699 3861
rect 6733 3827 6768 3861
rect 6802 3827 6837 3861
rect 6871 3827 6906 3861
rect 6940 3827 6975 3861
rect 7009 3827 7044 3861
rect 7078 3827 7113 3861
rect 7147 3827 7182 3861
rect 7216 3827 7251 3861
rect 7285 3827 7320 3861
rect 7354 3827 7389 3861
rect 7423 3827 7458 3861
rect 7492 3827 7527 3861
rect 7561 3827 7596 3861
rect 7630 3827 7665 3861
rect 7699 3827 7734 3861
rect 7768 3827 7803 3861
rect 7837 3827 7872 3861
rect 7906 3827 7941 3861
rect 7975 3827 8010 3861
rect 8044 3827 8079 3861
rect 8113 3827 8148 3861
rect 8182 3827 8217 3861
rect 8251 3827 8286 3861
rect 8320 3827 8355 3861
rect 8389 3827 8424 3861
rect 8458 3827 8493 3861
rect 8527 3827 8562 3861
rect 8596 3827 8631 3861
rect 8665 3827 8700 3861
rect 8734 3827 8769 3861
rect 8803 3827 8838 3861
rect 8872 3827 8907 3861
rect 8941 3827 8976 3861
rect 9010 3827 9045 3861
rect 9079 3827 9114 3861
rect 9148 3827 9183 3861
rect 9217 3827 9252 3861
rect 9286 3827 9320 3861
rect 9354 3827 9388 3861
rect 9422 3827 9456 3861
rect 4929 3785 9456 3827
rect 4929 3751 4974 3785
rect 5008 3751 5043 3785
rect 5077 3751 5112 3785
rect 5146 3751 5181 3785
rect 5215 3751 5250 3785
rect 5284 3751 5319 3785
rect 5353 3751 5388 3785
rect 5422 3751 5457 3785
rect 5491 3751 5526 3785
rect 5560 3751 5595 3785
rect 5629 3751 5664 3785
rect 5698 3751 5733 3785
rect 5767 3751 5802 3785
rect 5836 3751 5871 3785
rect 5905 3751 5940 3785
rect 5974 3751 6009 3785
rect 6043 3751 6078 3785
rect 6112 3751 6147 3785
rect 6181 3751 6216 3785
rect 6250 3751 6285 3785
rect 6319 3751 6354 3785
rect 6388 3751 6423 3785
rect 6457 3751 6492 3785
rect 6526 3751 6561 3785
rect 6595 3751 6630 3785
rect 6664 3751 6699 3785
rect 6733 3751 6768 3785
rect 6802 3751 6837 3785
rect 6871 3751 6906 3785
rect 6940 3751 6975 3785
rect 7009 3751 7044 3785
rect 7078 3751 7113 3785
rect 7147 3751 7182 3785
rect 7216 3751 7251 3785
rect 7285 3751 7320 3785
rect 7354 3751 7389 3785
rect 7423 3751 7458 3785
rect 7492 3751 7527 3785
rect 7561 3751 7596 3785
rect 7630 3751 7665 3785
rect 7699 3751 7734 3785
rect 7768 3751 7803 3785
rect 7837 3751 7872 3785
rect 7906 3751 7941 3785
rect 7975 3751 8010 3785
rect 8044 3751 8079 3785
rect 8113 3751 8148 3785
rect 8182 3751 8217 3785
rect 8251 3751 8286 3785
rect 8320 3751 8355 3785
rect 8389 3751 8424 3785
rect 8458 3751 8493 3785
rect 8527 3751 8562 3785
rect 8596 3751 8631 3785
rect 8665 3751 8700 3785
rect 8734 3751 8769 3785
rect 8803 3751 8838 3785
rect 8872 3751 8907 3785
rect 8941 3751 8976 3785
rect 9010 3751 9045 3785
rect 9079 3751 9114 3785
rect 9148 3751 9183 3785
rect 9217 3751 9252 3785
rect 9286 3751 9320 3785
rect 9354 3751 9388 3785
rect 9422 3751 9456 3785
rect 4929 3709 9456 3751
rect 4929 3675 4974 3709
rect 5008 3675 5043 3709
rect 5077 3675 5112 3709
rect 5146 3675 5181 3709
rect 5215 3675 5250 3709
rect 5284 3675 5319 3709
rect 5353 3675 5388 3709
rect 5422 3675 5457 3709
rect 5491 3675 5526 3709
rect 5560 3675 5595 3709
rect 5629 3675 5664 3709
rect 5698 3675 5733 3709
rect 5767 3675 5802 3709
rect 5836 3675 5871 3709
rect 5905 3675 5940 3709
rect 5974 3675 6009 3709
rect 6043 3675 6078 3709
rect 6112 3675 6147 3709
rect 6181 3675 6216 3709
rect 6250 3675 6285 3709
rect 6319 3675 6354 3709
rect 6388 3675 6423 3709
rect 6457 3675 6492 3709
rect 6526 3675 6561 3709
rect 6595 3675 6630 3709
rect 6664 3675 6699 3709
rect 6733 3675 6768 3709
rect 6802 3675 6837 3709
rect 6871 3675 6906 3709
rect 6940 3675 6975 3709
rect 7009 3675 7044 3709
rect 7078 3675 7113 3709
rect 7147 3675 7182 3709
rect 7216 3675 7251 3709
rect 7285 3675 7320 3709
rect 7354 3675 7389 3709
rect 7423 3675 7458 3709
rect 7492 3675 7527 3709
rect 7561 3675 7596 3709
rect 7630 3675 7665 3709
rect 7699 3675 7734 3709
rect 7768 3675 7803 3709
rect 7837 3675 7872 3709
rect 7906 3675 7941 3709
rect 7975 3675 8010 3709
rect 8044 3675 8079 3709
rect 8113 3675 8148 3709
rect 8182 3675 8217 3709
rect 8251 3675 8286 3709
rect 8320 3675 8355 3709
rect 8389 3675 8424 3709
rect 8458 3675 8493 3709
rect 8527 3675 8562 3709
rect 8596 3675 8631 3709
rect 8665 3675 8700 3709
rect 8734 3675 8769 3709
rect 8803 3675 8838 3709
rect 8872 3675 8907 3709
rect 8941 3675 8976 3709
rect 9010 3675 9045 3709
rect 9079 3675 9114 3709
rect 9148 3675 9183 3709
rect 9217 3675 9252 3709
rect 9286 3675 9320 3709
rect 9354 3675 9388 3709
rect 9422 3675 9456 3709
rect 4929 3672 9456 3675
rect 4929 2167 4940 3672
rect 13439 4139 13507 4173
rect 13541 4139 13575 4173
rect 13609 4139 13643 4173
rect 13677 4139 13711 4173
rect 13745 4139 13779 4173
rect 13813 4139 13847 4173
rect 13881 4139 13915 4173
rect 13949 4139 13983 4173
rect 14017 4139 14051 4173
rect 14085 4139 14119 4173
rect 14153 4139 14187 4173
rect 14221 4139 14255 4173
rect 14289 4139 14323 4173
rect 14357 4139 14391 4173
rect 14425 4139 14459 4173
rect 14493 4139 14527 4173
rect 14561 4139 14615 4173
rect 13439 4050 13473 4139
rect 13439 3982 13473 4016
rect 13439 3914 13473 3948
rect 13439 3846 13473 3880
rect 13439 3778 13473 3812
rect 13439 3710 13473 3744
rect 13439 3642 13473 3676
rect 13439 3574 13473 3608
rect 13439 3506 13473 3540
rect 13439 3438 13473 3472
rect 13439 3370 13473 3404
rect 13439 3302 13473 3336
rect 13439 3234 13473 3268
rect 11509 3043 12365 3044
rect 11509 3009 11543 3043
rect 11577 3009 11612 3043
rect 11646 3009 11681 3043
rect 11715 3009 11750 3043
rect 11784 3009 11819 3043
rect 11853 3009 11888 3043
rect 11922 3009 11957 3043
rect 11991 3009 12025 3043
rect 12059 3009 12093 3043
rect 12127 3009 12161 3043
rect 12195 3009 12229 3043
rect 12263 3009 12297 3043
rect 12331 3009 12365 3043
rect 11509 2955 12365 3009
rect 11509 2921 11543 2955
rect 11577 2921 11612 2955
rect 11646 2921 11681 2955
rect 11715 2921 11750 2955
rect 11784 2921 11819 2955
rect 11853 2921 11888 2955
rect 11922 2921 11957 2955
rect 11991 2921 12025 2955
rect 12059 2921 12093 2955
rect 12127 2921 12161 2955
rect 12195 2921 12229 2955
rect 12263 2921 12297 2955
rect 12331 2921 12365 2955
rect 11509 2867 12365 2921
rect 11509 2833 11543 2867
rect 11577 2833 11612 2867
rect 11646 2833 11681 2867
rect 11715 2833 11750 2867
rect 11784 2833 11819 2867
rect 11853 2833 11888 2867
rect 11922 2833 11957 2867
rect 11991 2833 12025 2867
rect 12059 2833 12093 2867
rect 12127 2833 12161 2867
rect 12195 2833 12229 2867
rect 12263 2833 12297 2867
rect 12331 2833 12365 2867
rect 11509 2779 12365 2833
rect 11509 2745 11543 2779
rect 11577 2745 11612 2779
rect 11646 2745 11681 2779
rect 11715 2745 11750 2779
rect 11784 2745 11819 2779
rect 11853 2745 11888 2779
rect 11922 2745 11957 2779
rect 11991 2745 12025 2779
rect 12059 2745 12093 2779
rect 12127 2745 12161 2779
rect 12195 2745 12229 2779
rect 12263 2745 12297 2779
rect 12331 2745 12365 2779
rect 11509 2744 12365 2745
rect 11841 2710 12365 2744
rect 11875 2676 11911 2710
rect 11945 2676 11981 2710
rect 12015 2676 12051 2710
rect 12085 2676 12121 2710
rect 12155 2676 12191 2710
rect 12225 2676 12261 2710
rect 12295 2676 12331 2710
rect 11841 2637 12365 2676
rect 11875 2603 11911 2637
rect 11945 2603 11981 2637
rect 12015 2603 12051 2637
rect 12085 2603 12121 2637
rect 12155 2603 12191 2637
rect 12225 2603 12261 2637
rect 12295 2603 12331 2637
rect 11841 2564 12365 2603
rect 11875 2530 11911 2564
rect 11945 2530 11981 2564
rect 12015 2530 12051 2564
rect 12085 2530 12121 2564
rect 12155 2530 12191 2564
rect 12225 2530 12261 2564
rect 12295 2530 12331 2564
rect 11841 2491 12365 2530
rect 11875 2457 11911 2491
rect 11945 2457 11981 2491
rect 12015 2457 12051 2491
rect 12085 2457 12121 2491
rect 12155 2457 12191 2491
rect 12225 2457 12261 2491
rect 12295 2457 12331 2491
rect 11841 2418 12365 2457
rect 11875 2384 11911 2418
rect 11945 2384 11981 2418
rect 12015 2384 12051 2418
rect 12085 2384 12121 2418
rect 12155 2384 12191 2418
rect 12225 2384 12261 2418
rect 12295 2384 12331 2418
rect 11841 2344 12365 2384
rect 11875 2310 11911 2344
rect 11945 2310 11981 2344
rect 12015 2310 12051 2344
rect 12085 2310 12121 2344
rect 12155 2310 12191 2344
rect 12225 2310 12261 2344
rect 12295 2310 12331 2344
rect 11841 2270 12365 2310
rect 11875 2236 11911 2270
rect 11945 2236 11981 2270
rect 12015 2236 12051 2270
rect 12085 2236 12121 2270
rect 12155 2236 12191 2270
rect 12225 2236 12261 2270
rect 12295 2236 12331 2270
rect 11841 2202 12365 2236
rect 3864 2132 4940 2167
rect 3864 2098 3875 2132
rect 3909 2098 3943 2132
rect 3977 2098 4011 2132
rect 4045 2098 4079 2132
rect 4113 2098 4147 2132
rect 4181 2098 4215 2132
rect 4249 2098 4283 2132
rect 4317 2098 4351 2132
rect 4385 2098 4419 2132
rect 4453 2098 4487 2132
rect 4521 2098 4555 2132
rect 4589 2098 4623 2132
rect 4657 2098 4691 2132
rect 4725 2098 4759 2132
rect 4793 2098 4827 2132
rect 4861 2098 4895 2132
rect 4929 2098 4940 2132
rect 3864 2063 4940 2098
rect 3864 2029 3875 2063
rect 3909 2029 3943 2063
rect 3977 2029 4011 2063
rect 4045 2029 4079 2063
rect 4113 2029 4147 2063
rect 4181 2029 4215 2063
rect 4249 2029 4283 2063
rect 4317 2029 4351 2063
rect 4385 2029 4419 2063
rect 4453 2029 4487 2063
rect 4521 2029 4555 2063
rect 4589 2029 4623 2063
rect 4657 2029 4691 2063
rect 4725 2029 4759 2063
rect 4793 2029 4827 2063
rect 4861 2029 4895 2063
rect 4929 2029 4940 2063
rect 3864 1994 4940 2029
rect 3864 1960 3875 1994
rect 3909 1960 3943 1994
rect 3977 1960 4011 1994
rect 4045 1960 4079 1994
rect 4113 1960 4147 1994
rect 4181 1960 4215 1994
rect 4249 1960 4283 1994
rect 4317 1960 4351 1994
rect 4385 1960 4419 1994
rect 4453 1960 4487 1994
rect 4521 1960 4555 1994
rect 4589 1960 4623 1994
rect 4657 1960 4691 1994
rect 4725 1960 4759 1994
rect 4793 1960 4827 1994
rect 4861 1960 4895 1994
rect 4929 1960 4940 1994
rect 3864 1925 4940 1960
rect 3864 1891 3875 1925
rect 3909 1891 3943 1925
rect 3977 1891 4011 1925
rect 4045 1891 4079 1925
rect 4113 1891 4147 1925
rect 4181 1891 4215 1925
rect 4249 1891 4283 1925
rect 4317 1891 4351 1925
rect 4385 1891 4419 1925
rect 4453 1891 4487 1925
rect 4521 1891 4555 1925
rect 4589 1891 4623 1925
rect 4657 1891 4691 1925
rect 4725 1891 4759 1925
rect 4793 1891 4827 1925
rect 4861 1891 4895 1925
rect 4929 1891 4940 1925
rect 3864 1856 4940 1891
rect 3864 1822 3875 1856
rect 3909 1822 3943 1856
rect 3977 1822 4011 1856
rect 4045 1822 4079 1856
rect 4113 1822 4147 1856
rect 4181 1822 4215 1856
rect 4249 1822 4283 1856
rect 4317 1822 4351 1856
rect 4385 1822 4419 1856
rect 4453 1822 4487 1856
rect 4521 1822 4555 1856
rect 4589 1822 4623 1856
rect 4657 1822 4691 1856
rect 4725 1822 4759 1856
rect 4793 1822 4827 1856
rect 4861 1822 4895 1856
rect 4929 1822 4940 1856
rect 3864 1787 4940 1822
rect 3864 1753 3875 1787
rect 3909 1753 3943 1787
rect 3977 1753 4011 1787
rect 4045 1753 4079 1787
rect 4113 1753 4147 1787
rect 4181 1753 4215 1787
rect 4249 1753 4283 1787
rect 4317 1753 4351 1787
rect 4385 1753 4419 1787
rect 4453 1753 4487 1787
rect 4521 1753 4555 1787
rect 4589 1753 4623 1787
rect 4657 1753 4691 1787
rect 4725 1753 4759 1787
rect 4793 1753 4827 1787
rect 4861 1753 4895 1787
rect 4929 1753 4940 1787
rect 3864 1718 4940 1753
rect 3864 1684 3875 1718
rect 3909 1684 3943 1718
rect 3977 1684 4011 1718
rect 4045 1684 4079 1718
rect 4113 1684 4147 1718
rect 4181 1684 4215 1718
rect 4249 1684 4283 1718
rect 4317 1684 4351 1718
rect 4385 1684 4419 1718
rect 4453 1684 4487 1718
rect 4521 1684 4555 1718
rect 4589 1684 4623 1718
rect 4657 1684 4691 1718
rect 4725 1684 4759 1718
rect 4793 1684 4827 1718
rect 4861 1684 4895 1718
rect 4929 1684 4940 1718
rect 3864 1649 4940 1684
rect 3864 1615 3875 1649
rect 3909 1615 3943 1649
rect 3977 1615 4011 1649
rect 4045 1615 4079 1649
rect 4113 1615 4147 1649
rect 4181 1615 4215 1649
rect 4249 1615 4283 1649
rect 4317 1615 4351 1649
rect 4385 1615 4419 1649
rect 4453 1615 4487 1649
rect 4521 1615 4555 1649
rect 4589 1615 4623 1649
rect 4657 1615 4691 1649
rect 4725 1615 4759 1649
rect 4793 1615 4827 1649
rect 4861 1615 4895 1649
rect 4929 1615 4940 1649
rect 3864 1580 4940 1615
rect 3864 1546 3875 1580
rect 3909 1546 3943 1580
rect 3977 1546 4011 1580
rect 4045 1546 4079 1580
rect 4113 1546 4147 1580
rect 4181 1546 4215 1580
rect 4249 1546 4283 1580
rect 4317 1546 4351 1580
rect 4385 1546 4419 1580
rect 4453 1546 4487 1580
rect 4521 1546 4555 1580
rect 4589 1546 4623 1580
rect 4657 1546 4691 1580
rect 4725 1546 4759 1580
rect 4793 1546 4827 1580
rect 4861 1546 4895 1580
rect 4929 1546 4940 1580
rect 3864 1511 4940 1546
rect 3864 1477 3875 1511
rect 3909 1477 3943 1511
rect 3977 1477 4011 1511
rect 4045 1477 4079 1511
rect 4113 1477 4147 1511
rect 4181 1477 4215 1511
rect 4249 1477 4283 1511
rect 4317 1477 4351 1511
rect 4385 1477 4419 1511
rect 4453 1477 4487 1511
rect 4521 1477 4555 1511
rect 4589 1477 4623 1511
rect 4657 1477 4691 1511
rect 4725 1477 4759 1511
rect 4793 1477 4827 1511
rect 4861 1477 4895 1511
rect 4929 1477 4940 1511
rect 3864 1442 4940 1477
rect 3864 1408 3875 1442
rect 3909 1408 3943 1442
rect 3977 1408 4011 1442
rect 4045 1408 4079 1442
rect 4113 1408 4147 1442
rect 4181 1408 4215 1442
rect 4249 1408 4283 1442
rect 4317 1408 4351 1442
rect 4385 1408 4419 1442
rect 4453 1408 4487 1442
rect 4521 1408 4555 1442
rect 4589 1408 4623 1442
rect 4657 1408 4691 1442
rect 4725 1408 4759 1442
rect 4793 1408 4827 1442
rect 4861 1408 4895 1442
rect 4929 1408 4940 1442
rect 3864 1373 4940 1408
rect 3864 1339 3875 1373
rect 3909 1339 3943 1373
rect 3977 1339 4011 1373
rect 4045 1339 4079 1373
rect 4113 1339 4147 1373
rect 4181 1339 4215 1373
rect 4249 1339 4283 1373
rect 4317 1339 4351 1373
rect 4385 1339 4419 1373
rect 4453 1339 4487 1373
rect 4521 1339 4555 1373
rect 4589 1339 4623 1373
rect 4657 1339 4691 1373
rect 4725 1339 4759 1373
rect 4793 1339 4827 1373
rect 4861 1339 4895 1373
rect 4929 1339 4940 1373
rect 3864 1304 4940 1339
rect 3864 1270 3875 1304
rect 3909 1270 3943 1304
rect 3977 1270 4011 1304
rect 4045 1270 4079 1304
rect 4113 1270 4147 1304
rect 4181 1270 4215 1304
rect 4249 1270 4283 1304
rect 4317 1270 4351 1304
rect 4385 1270 4419 1304
rect 4453 1270 4487 1304
rect 4521 1270 4555 1304
rect 4589 1270 4623 1304
rect 4657 1270 4691 1304
rect 4725 1270 4759 1304
rect 4793 1270 4827 1304
rect 4861 1270 4895 1304
rect 4929 1270 4940 1304
rect 3864 1235 4940 1270
rect 3864 1201 3875 1235
rect 3909 1201 3943 1235
rect 3977 1201 4011 1235
rect 4045 1201 4079 1235
rect 4113 1201 4147 1235
rect 4181 1201 4215 1235
rect 4249 1201 4283 1235
rect 4317 1201 4351 1235
rect 4385 1201 4419 1235
rect 4453 1201 4487 1235
rect 4521 1201 4555 1235
rect 4589 1201 4623 1235
rect 4657 1201 4691 1235
rect 4725 1201 4759 1235
rect 4793 1201 4827 1235
rect 4861 1201 4895 1235
rect 4929 1201 4940 1235
rect 3864 1166 4940 1201
rect 3864 1132 3875 1166
rect 3909 1132 3943 1166
rect 3977 1132 4011 1166
rect 4045 1132 4079 1166
rect 4113 1132 4147 1166
rect 4181 1132 4215 1166
rect 4249 1132 4283 1166
rect 4317 1132 4351 1166
rect 4385 1132 4419 1166
rect 4453 1132 4487 1166
rect 4521 1132 4555 1166
rect 4589 1132 4623 1166
rect 4657 1132 4691 1166
rect 4725 1132 4759 1166
rect 4793 1132 4827 1166
rect 4861 1132 4895 1166
rect 4929 1132 4940 1166
rect 3864 1097 4940 1132
rect 3864 1063 3875 1097
rect 3909 1063 3943 1097
rect 3977 1063 4011 1097
rect 4045 1063 4079 1097
rect 4113 1063 4147 1097
rect 4181 1063 4215 1097
rect 4249 1063 4283 1097
rect 4317 1063 4351 1097
rect 4385 1063 4419 1097
rect 4453 1063 4487 1097
rect 4521 1063 4555 1097
rect 4589 1063 4623 1097
rect 4657 1063 4691 1097
rect 4725 1063 4759 1097
rect 4793 1063 4827 1097
rect 4861 1063 4895 1097
rect 4929 1063 4940 1097
rect 3864 1028 4940 1063
rect 3864 994 3875 1028
rect 3909 994 3943 1028
rect 3977 994 4011 1028
rect 4045 994 4079 1028
rect 4113 994 4147 1028
rect 4181 994 4215 1028
rect 4249 994 4283 1028
rect 4317 994 4351 1028
rect 4385 994 4419 1028
rect 4453 994 4487 1028
rect 4521 994 4555 1028
rect 4589 994 4623 1028
rect 4657 994 4691 1028
rect 4725 994 4759 1028
rect 4793 994 4827 1028
rect 4861 994 4895 1028
rect 4929 994 4940 1028
rect 3864 959 4940 994
rect 3864 925 3875 959
rect 3909 925 3943 959
rect 3977 925 4011 959
rect 4045 925 4079 959
rect 4113 925 4147 959
rect 4181 925 4215 959
rect 4249 925 4283 959
rect 4317 925 4351 959
rect 4385 925 4419 959
rect 4453 925 4487 959
rect 4521 925 4555 959
rect 4589 925 4623 959
rect 4657 925 4691 959
rect 4725 925 4759 959
rect 4793 925 4827 959
rect 4861 925 4895 959
rect 4929 925 4940 959
rect 3864 890 4940 925
rect 3864 856 3875 890
rect 3909 856 3943 890
rect 3977 856 4011 890
rect 4045 856 4079 890
rect 4113 856 4147 890
rect 4181 856 4215 890
rect 4249 856 4283 890
rect 4317 856 4351 890
rect 4385 856 4419 890
rect 4453 856 4487 890
rect 4521 856 4555 890
rect 4589 856 4623 890
rect 4657 856 4691 890
rect 4725 856 4759 890
rect 4793 856 4827 890
rect 4861 856 4895 890
rect 4929 856 4940 890
rect 3864 821 4940 856
rect 5299 1058 8646 1093
rect 5333 1024 5369 1058
rect 5403 1024 5438 1058
rect 5472 1024 5507 1058
rect 5541 1024 5576 1058
rect 5610 1024 5645 1058
rect 5679 1024 5714 1058
rect 5748 1024 5783 1058
rect 5817 1024 5852 1058
rect 5886 1024 5921 1058
rect 5955 1024 5990 1058
rect 6024 1024 6059 1058
rect 6093 1024 6128 1058
rect 6162 1024 6197 1058
rect 6231 1024 6266 1058
rect 6300 1024 6335 1058
rect 6369 1024 6404 1058
rect 6438 1024 6473 1058
rect 6507 1024 6542 1058
rect 6576 1024 6611 1058
rect 6645 1024 6680 1058
rect 6714 1024 6749 1058
rect 6783 1024 6818 1058
rect 6852 1024 6887 1058
rect 6921 1024 6956 1058
rect 6990 1024 7025 1058
rect 7059 1024 7094 1058
rect 7128 1024 7163 1058
rect 7197 1024 7232 1058
rect 7266 1024 7301 1058
rect 7335 1024 7370 1058
rect 7404 1024 7439 1058
rect 7473 1024 7508 1058
rect 7542 1024 7577 1058
rect 7611 1024 7646 1058
rect 7680 1024 7715 1058
rect 7749 1024 7784 1058
rect 7818 1024 7853 1058
rect 7887 1024 7922 1058
rect 7956 1024 7991 1058
rect 8025 1024 8060 1058
rect 8094 1024 8129 1058
rect 8163 1024 8198 1058
rect 8232 1024 8267 1058
rect 8301 1024 8336 1058
rect 8370 1024 8405 1058
rect 8439 1024 8474 1058
rect 8508 1024 8543 1058
rect 8577 1024 8612 1058
rect 5299 986 8646 1024
rect 5333 952 5369 986
rect 5403 952 5438 986
rect 5472 952 5507 986
rect 5541 952 5576 986
rect 5610 952 5645 986
rect 5679 952 5714 986
rect 5748 952 5783 986
rect 5817 952 5852 986
rect 5886 952 5921 986
rect 5955 952 5990 986
rect 6024 952 6059 986
rect 6093 952 6128 986
rect 6162 952 6197 986
rect 6231 952 6266 986
rect 6300 952 6335 986
rect 6369 952 6404 986
rect 6438 952 6473 986
rect 6507 952 6542 986
rect 6576 952 6611 986
rect 6645 952 6680 986
rect 6714 952 6749 986
rect 6783 952 6818 986
rect 6852 952 6887 986
rect 6921 952 6956 986
rect 6990 952 7025 986
rect 7059 952 7094 986
rect 7128 952 7163 986
rect 7197 952 7232 986
rect 7266 952 7301 986
rect 7335 952 7370 986
rect 7404 952 7439 986
rect 7473 952 7508 986
rect 7542 952 7577 986
rect 7611 952 7646 986
rect 7680 952 7715 986
rect 7749 952 7784 986
rect 7818 952 7853 986
rect 7887 952 7922 986
rect 7956 952 7991 986
rect 8025 952 8060 986
rect 8094 952 8129 986
rect 8163 952 8198 986
rect 8232 952 8267 986
rect 8301 952 8336 986
rect 8370 952 8405 986
rect 8439 952 8474 986
rect 8508 952 8543 986
rect 8577 952 8612 986
rect 5299 914 8646 952
rect 5333 880 5369 914
rect 5403 880 5438 914
rect 5472 880 5507 914
rect 5541 880 5576 914
rect 5610 880 5645 914
rect 5679 880 5714 914
rect 5748 880 5783 914
rect 5817 880 5852 914
rect 5886 880 5921 914
rect 5955 880 5990 914
rect 6024 880 6059 914
rect 6093 880 6128 914
rect 6162 880 6197 914
rect 6231 880 6266 914
rect 6300 880 6335 914
rect 6369 880 6404 914
rect 6438 880 6473 914
rect 6507 880 6542 914
rect 6576 880 6611 914
rect 6645 880 6680 914
rect 6714 880 6749 914
rect 6783 880 6818 914
rect 6852 880 6887 914
rect 6921 880 6956 914
rect 6990 880 7025 914
rect 7059 880 7094 914
rect 7128 880 7163 914
rect 7197 880 7232 914
rect 7266 880 7301 914
rect 7335 880 7370 914
rect 7404 880 7439 914
rect 7473 880 7508 914
rect 7542 880 7577 914
rect 7611 880 7646 914
rect 7680 880 7715 914
rect 7749 880 7784 914
rect 7818 880 7853 914
rect 7887 880 7922 914
rect 7956 880 7991 914
rect 8025 880 8060 914
rect 8094 880 8129 914
rect 8163 880 8198 914
rect 8232 880 8267 914
rect 8301 880 8336 914
rect 8370 880 8405 914
rect 8439 880 8474 914
rect 8508 880 8543 914
rect 8577 880 8612 914
rect 5299 845 8646 880
rect 3864 787 3875 821
rect 3909 787 3943 821
rect 3977 787 4011 821
rect 4045 787 4079 821
rect 4113 787 4147 821
rect 4181 787 4215 821
rect 4249 787 4283 821
rect 4317 787 4351 821
rect 4385 787 4419 821
rect 4453 787 4487 821
rect 4521 787 4555 821
rect 4589 787 4623 821
rect 4657 787 4691 821
rect 4725 787 4759 821
rect 4793 787 4827 821
rect 4861 787 4895 821
rect 4929 787 4940 821
rect 3864 752 4940 787
rect 3864 718 3875 752
rect 3909 718 3943 752
rect 3977 718 4011 752
rect 4045 718 4079 752
rect 4113 718 4147 752
rect 4181 718 4215 752
rect 4249 718 4283 752
rect 4317 718 4351 752
rect 4385 718 4419 752
rect 4453 718 4487 752
rect 4521 718 4555 752
rect 4589 718 4623 752
rect 4657 718 4691 752
rect 4725 718 4759 752
rect 4793 718 4827 752
rect 4861 718 4895 752
rect 4929 718 4940 752
rect 3864 683 4940 718
rect 3864 649 3875 683
rect 3909 649 3943 683
rect 3977 649 4011 683
rect 4045 649 4079 683
rect 4113 649 4147 683
rect 4181 649 4215 683
rect 4249 649 4283 683
rect 4317 649 4351 683
rect 4385 649 4419 683
rect 4453 649 4487 683
rect 4521 649 4555 683
rect 4589 649 4623 683
rect 4657 649 4691 683
rect 4725 649 4759 683
rect 4793 649 4827 683
rect 4861 649 4895 683
rect 4929 649 4940 683
rect 3864 614 4940 649
rect 3864 580 3875 614
rect 3909 580 3943 614
rect 3977 580 4011 614
rect 4045 580 4079 614
rect 4113 580 4147 614
rect 4181 580 4215 614
rect 4249 580 4283 614
rect 4317 580 4351 614
rect 4385 580 4419 614
rect 4453 580 4487 614
rect 4521 580 4555 614
rect 4589 580 4623 614
rect 4657 580 4691 614
rect 4725 580 4759 614
rect 4793 580 4827 614
rect 4861 580 4895 614
rect 4929 580 4940 614
rect 3864 545 4940 580
rect 3864 511 3875 545
rect 3909 511 3943 545
rect 3977 511 4011 545
rect 4045 511 4079 545
rect 4113 511 4147 545
rect 4181 511 4215 545
rect 4249 511 4283 545
rect 4317 511 4351 545
rect 4385 511 4419 545
rect 4453 511 4487 545
rect 4521 511 4555 545
rect 4589 511 4623 545
rect 4657 511 4691 545
rect 4725 511 4759 545
rect 4793 511 4827 545
rect 4861 511 4895 545
rect 4929 511 4940 545
rect 3864 476 4940 511
rect 3864 442 3875 476
rect 3909 442 3943 476
rect 3977 442 4011 476
rect 4045 442 4079 476
rect 4113 442 4147 476
rect 4181 442 4215 476
rect 4249 442 4283 476
rect 4317 442 4351 476
rect 4385 442 4419 476
rect 4453 442 4487 476
rect 4521 442 4555 476
rect 4589 442 4623 476
rect 4657 442 4691 476
rect 4725 442 4759 476
rect 4793 442 4827 476
rect 4861 442 4895 476
rect 4929 442 4940 476
rect 3864 407 4940 442
rect 3864 373 3875 407
rect 3909 373 3943 407
rect 3977 373 4011 407
rect 4045 373 4079 407
rect 4113 373 4147 407
rect 4181 373 4215 407
rect 4249 373 4283 407
rect 4317 373 4351 407
rect 4385 373 4419 407
rect 4453 373 4487 407
rect 4521 373 4555 407
rect 4589 373 4623 407
rect 4657 373 4691 407
rect 4725 373 4759 407
rect 4793 373 4827 407
rect 4861 373 4895 407
rect 4929 373 4940 407
rect 3864 338 4940 373
rect 3864 304 3875 338
rect 3909 304 3943 338
rect 3977 304 4011 338
rect 4045 304 4079 338
rect 4113 304 4147 338
rect 4181 304 4215 338
rect 4249 304 4283 338
rect 4317 304 4351 338
rect 4385 304 4419 338
rect 4453 304 4487 338
rect 4521 304 4555 338
rect 4589 304 4623 338
rect 4657 304 4691 338
rect 4725 304 4759 338
rect 4793 304 4827 338
rect 4861 304 4895 338
rect 4929 304 4940 338
rect 3864 269 4940 304
rect 3864 235 3875 269
rect 3909 235 3943 269
rect 3977 235 4011 269
rect 4045 235 4079 269
rect 4113 235 4147 269
rect 4181 235 4215 269
rect 4249 235 4283 269
rect 4317 235 4351 269
rect 4385 235 4419 269
rect 4453 235 4487 269
rect 4521 235 4555 269
rect 4589 235 4623 269
rect 4657 235 4691 269
rect 4725 235 4759 269
rect 4793 235 4827 269
rect 4861 235 4895 269
rect 4929 235 4940 269
rect 3864 200 4940 235
rect 3864 166 3875 200
rect 3909 166 3943 200
rect 3977 166 4011 200
rect 4045 166 4079 200
rect 4113 166 4147 200
rect 4181 166 4215 200
rect 4249 166 4283 200
rect 4317 166 4351 200
rect 4385 166 4419 200
rect 4453 166 4487 200
rect 4521 166 4555 200
rect 4589 166 4623 200
rect 4657 166 4691 200
rect 4725 166 4759 200
rect 4793 166 4827 200
rect 4861 166 4895 200
rect 4929 166 4940 200
rect 3864 131 4940 166
rect 3864 97 3875 131
rect 3909 97 3943 131
rect 3977 97 4011 131
rect 4045 97 4079 131
rect 4113 97 4147 131
rect 4181 97 4215 131
rect 4249 97 4283 131
rect 4317 97 4351 131
rect 4385 97 4419 131
rect 4453 97 4487 131
rect 4521 97 4555 131
rect 4589 97 4623 131
rect 4657 97 4691 131
rect 4725 97 4759 131
rect 4793 97 4827 131
rect 4861 97 4895 131
rect 4929 97 4940 131
rect 3864 62 4940 97
rect 3864 28 3875 62
rect 3909 28 3943 62
rect 3977 28 4011 62
rect 4045 28 4079 62
rect 4113 28 4147 62
rect 4181 28 4215 62
rect 4249 28 4283 62
rect 4317 28 4351 62
rect 4385 28 4419 62
rect 4453 28 4487 62
rect 4521 28 4555 62
rect 4589 28 4623 62
rect 4657 28 4691 62
rect 4725 28 4759 62
rect 4793 28 4827 62
rect 4861 28 4895 62
rect 4929 28 4940 62
rect 3864 4 4940 28
rect 11314 839 12838 879
rect 11348 805 11385 839
rect 11419 805 11456 839
rect 11490 805 11527 839
rect 11561 805 11598 839
rect 11632 805 11669 839
rect 11703 805 11740 839
rect 11774 805 11811 839
rect 11845 805 11882 839
rect 11916 805 11953 839
rect 11987 805 12024 839
rect 12058 805 12095 839
rect 12129 805 12166 839
rect 12200 805 12237 839
rect 12271 805 12308 839
rect 12342 805 12379 839
rect 12413 805 12450 839
rect 12484 805 12521 839
rect 12555 805 12592 839
rect 12626 805 12663 839
rect 12697 805 12734 839
rect 12768 805 12804 839
rect 11314 769 12838 805
rect 11348 735 11385 769
rect 11419 735 11456 769
rect 11490 735 11527 769
rect 11561 735 11598 769
rect 11632 735 11669 769
rect 11703 735 11740 769
rect 11774 735 11811 769
rect 11845 735 11882 769
rect 11916 735 11953 769
rect 11987 735 12024 769
rect 12058 735 12095 769
rect 12129 735 12166 769
rect 12200 735 12237 769
rect 12271 735 12308 769
rect 12342 735 12379 769
rect 12413 735 12450 769
rect 12484 735 12521 769
rect 12555 735 12592 769
rect 12626 735 12663 769
rect 12697 735 12734 769
rect 12768 735 12804 769
rect 11314 699 12838 735
rect 11348 665 11385 699
rect 11419 665 11456 699
rect 11490 665 11527 699
rect 11561 665 11598 699
rect 11632 665 11669 699
rect 11703 665 11740 699
rect 11774 665 11811 699
rect 11845 665 11882 699
rect 11916 665 11953 699
rect 11987 665 12024 699
rect 12058 665 12095 699
rect 12129 665 12166 699
rect 12200 665 12237 699
rect 12271 665 12308 699
rect 12342 665 12379 699
rect 12413 665 12450 699
rect 12484 665 12521 699
rect 12555 665 12592 699
rect 12626 665 12663 699
rect 12697 665 12734 699
rect 12768 665 12804 699
rect 11314 629 12838 665
rect 11348 595 11385 629
rect 11419 595 11456 629
rect 11490 595 11527 629
rect 11561 595 11598 629
rect 11632 595 11669 629
rect 11703 595 11740 629
rect 11774 595 11811 629
rect 11845 595 11882 629
rect 11916 595 11953 629
rect 11987 595 12024 629
rect 12058 595 12095 629
rect 12129 595 12166 629
rect 12200 595 12237 629
rect 12271 595 12308 629
rect 12342 595 12379 629
rect 12413 595 12450 629
rect 12484 595 12521 629
rect 12555 595 12592 629
rect 12626 595 12663 629
rect 12697 595 12734 629
rect 12768 595 12804 629
rect 11314 559 12838 595
rect 11348 525 11385 559
rect 11419 525 11456 559
rect 11490 525 11527 559
rect 11561 525 11598 559
rect 11632 525 11669 559
rect 11703 525 11740 559
rect 11774 525 11811 559
rect 11845 525 11882 559
rect 11916 525 11953 559
rect 11987 525 12024 559
rect 12058 525 12095 559
rect 12129 525 12166 559
rect 12200 525 12237 559
rect 12271 525 12308 559
rect 12342 525 12379 559
rect 12413 525 12450 559
rect 12484 525 12521 559
rect 12555 525 12592 559
rect 12626 525 12663 559
rect 12697 525 12734 559
rect 12768 525 12804 559
rect 11314 489 12838 525
rect 11348 455 11385 489
rect 11419 455 11456 489
rect 11490 455 11527 489
rect 11561 455 11598 489
rect 11632 455 11669 489
rect 11703 455 11740 489
rect 11774 455 11811 489
rect 11845 455 11882 489
rect 11916 455 11953 489
rect 11987 455 12024 489
rect 12058 455 12095 489
rect 12129 455 12166 489
rect 12200 455 12237 489
rect 12271 455 12308 489
rect 12342 455 12379 489
rect 12413 455 12450 489
rect 12484 455 12521 489
rect 12555 455 12592 489
rect 12626 455 12663 489
rect 12697 455 12734 489
rect 12768 455 12804 489
rect 11314 419 12838 455
rect 11348 385 11385 419
rect 11419 385 11456 419
rect 11490 385 11527 419
rect 11561 385 11598 419
rect 11632 385 11669 419
rect 11703 385 11740 419
rect 11774 385 11811 419
rect 11845 385 11882 419
rect 11916 385 11953 419
rect 11987 385 12024 419
rect 12058 385 12095 419
rect 12129 385 12166 419
rect 12200 385 12237 419
rect 12271 385 12308 419
rect 12342 385 12379 419
rect 12413 385 12450 419
rect 12484 385 12521 419
rect 12555 385 12592 419
rect 12626 385 12663 419
rect 12697 385 12734 419
rect 12768 385 12804 419
rect 11314 349 12838 385
rect 11348 315 11385 349
rect 11419 315 11456 349
rect 11490 315 11527 349
rect 11561 315 11598 349
rect 11632 315 11669 349
rect 11703 315 11740 349
rect 11774 315 11811 349
rect 11845 315 11882 349
rect 11916 315 11953 349
rect 11987 315 12024 349
rect 12058 315 12095 349
rect 12129 315 12166 349
rect 12200 315 12237 349
rect 12271 315 12308 349
rect 12342 315 12379 349
rect 12413 315 12450 349
rect 12484 315 12521 349
rect 12555 315 12592 349
rect 12626 315 12663 349
rect 12697 315 12734 349
rect 12768 315 12804 349
rect 11314 279 12838 315
rect 11348 245 11385 279
rect 11419 245 11456 279
rect 11490 245 11527 279
rect 11561 245 11598 279
rect 11632 245 11669 279
rect 11703 245 11740 279
rect 11774 245 11811 279
rect 11845 245 11882 279
rect 11916 245 11953 279
rect 11987 245 12024 279
rect 12058 245 12095 279
rect 12129 245 12166 279
rect 12200 245 12237 279
rect 12271 245 12308 279
rect 12342 245 12379 279
rect 12413 245 12450 279
rect 12484 245 12521 279
rect 12555 245 12592 279
rect 12626 245 12663 279
rect 12697 245 12734 279
rect 12768 245 12804 279
rect 11314 209 12838 245
rect 11348 175 11385 209
rect 11419 175 11456 209
rect 11490 175 11527 209
rect 11561 175 11598 209
rect 11632 175 11669 209
rect 11703 175 11740 209
rect 11774 175 11811 209
rect 11845 175 11882 209
rect 11916 175 11953 209
rect 11987 175 12024 209
rect 12058 175 12095 209
rect 12129 175 12166 209
rect 12200 175 12237 209
rect 12271 175 12308 209
rect 12342 175 12379 209
rect 12413 175 12450 209
rect 12484 175 12521 209
rect 12555 175 12592 209
rect 12626 175 12663 209
rect 12697 175 12734 209
rect 12768 175 12804 209
rect 11314 139 12838 175
rect 11348 105 11385 139
rect 11419 105 11456 139
rect 11490 105 11527 139
rect 11561 105 11598 139
rect 11632 105 11669 139
rect 11703 105 11740 139
rect 11774 105 11811 139
rect 11845 105 11882 139
rect 11916 105 11953 139
rect 11987 105 12024 139
rect 12058 105 12095 139
rect 12129 105 12166 139
rect 12200 105 12237 139
rect 12271 105 12308 139
rect 12342 105 12379 139
rect 12413 105 12450 139
rect 12484 105 12521 139
rect 12555 105 12592 139
rect 12626 105 12663 139
rect 12697 105 12734 139
rect 12768 105 12804 139
rect 11314 69 12838 105
rect 11348 35 11385 69
rect 11419 35 11456 69
rect 11490 35 11527 69
rect 11561 35 11598 69
rect 11632 35 11669 69
rect 11703 35 11740 69
rect 11774 35 11811 69
rect 11845 35 11882 69
rect 11916 35 11953 69
rect 11987 35 12024 69
rect 12058 35 12095 69
rect 12129 35 12166 69
rect 12200 35 12237 69
rect 12271 35 12308 69
rect 12342 35 12379 69
rect 12413 35 12450 69
rect 12484 35 12521 69
rect 12555 35 12592 69
rect 12626 35 12663 69
rect 12697 35 12734 69
rect 12768 35 12804 69
rect 11314 -1 12838 35
rect 11348 -35 11385 -1
rect 11419 -35 11456 -1
rect 11490 -35 11527 -1
rect 11561 -35 11598 -1
rect 11632 -35 11669 -1
rect 11703 -35 11740 -1
rect 11774 -35 11811 -1
rect 11845 -35 11882 -1
rect 11916 -35 11953 -1
rect 11987 -35 12024 -1
rect 12058 -35 12095 -1
rect 12129 -35 12166 -1
rect 12200 -35 12237 -1
rect 12271 -35 12308 -1
rect 12342 -35 12379 -1
rect 12413 -35 12450 -1
rect 12484 -35 12521 -1
rect 12555 -35 12592 -1
rect 12626 -35 12663 -1
rect 12697 -35 12734 -1
rect 12768 -35 12804 -1
rect 13439 2658 13507 2692
rect 13541 2658 13575 2692
rect 13609 2658 13643 2692
rect 13677 2658 13711 2692
rect 13745 2658 13779 2692
rect 13813 2658 13847 2692
rect 13881 2658 13915 2692
rect 13949 2658 13983 2692
rect 14017 2658 14051 2692
rect 14085 2658 14119 2692
rect 14153 2658 14187 2692
rect 14221 2658 14255 2692
rect 14289 2658 14323 2692
rect 14357 2658 14391 2692
rect 14425 2658 14459 2692
rect 14493 2658 14527 2692
rect 14561 2658 14595 2692
rect 14629 2658 14739 2692
rect 13439 2588 13473 2658
rect 14705 2624 14739 2658
rect 13439 2520 13473 2554
rect 14705 2556 14739 2590
rect 13439 2452 13473 2486
rect 13439 2384 13473 2418
rect 13439 2316 13473 2350
rect 13439 2248 13473 2282
rect 13439 2180 13473 2214
rect 13439 2112 13473 2146
rect 13439 2044 13473 2078
rect 13439 1976 13473 2010
rect 13439 1908 13473 1942
rect 13439 1840 13473 1874
rect 13439 1772 13473 1806
rect 13439 1704 13473 1738
rect 13439 1562 13473 1670
rect 13439 1494 13473 1528
rect 13439 1426 13473 1460
rect 13439 1358 13473 1392
rect 13439 1290 13473 1324
rect 13439 1222 13473 1256
rect 13439 1154 13473 1188
rect 13439 1086 13473 1120
rect 13439 1018 13473 1052
rect 13439 950 13473 984
rect 13439 882 13473 916
rect 13439 814 13473 848
rect 13439 746 13473 780
rect 13439 678 13473 712
rect 13439 610 13473 644
rect 13439 542 13473 576
rect 13439 474 13473 508
rect 13439 406 13473 440
rect 14705 2488 14739 2522
rect 14705 2420 14739 2454
rect 14705 2352 14739 2386
rect 14705 2284 14739 2318
rect 14705 2216 14739 2250
rect 14705 2148 14739 2182
rect 14705 2080 14739 2114
rect 14705 2012 14739 2046
rect 14705 1944 14739 1978
rect 14705 1876 14739 1910
rect 14705 1808 14739 1842
rect 14705 1740 14739 1774
rect 14705 1672 14739 1706
rect 14705 1604 14739 1638
rect 14705 1536 14739 1570
rect 14705 1468 14739 1502
rect 14705 1400 14739 1434
rect 14705 1332 14739 1366
rect 14705 1264 14739 1298
rect 14705 1196 14739 1230
rect 14705 1128 14739 1162
rect 14705 1060 14739 1094
rect 14705 992 14739 1026
rect 14705 924 14739 958
rect 14705 856 14739 890
rect 14705 788 14739 822
rect 14705 720 14739 754
rect 14705 652 14739 686
rect 14705 584 14739 618
rect 14705 516 14739 550
rect 14705 448 14739 482
rect 13439 338 13473 372
rect 14705 380 14739 414
rect 13439 270 13473 304
rect 14705 270 14739 346
rect 13439 236 13549 270
rect 13583 236 13617 270
rect 13651 236 13685 270
rect 13719 236 13753 270
rect 13787 236 13821 270
rect 13855 236 13889 270
rect 13923 236 13957 270
rect 13991 236 14025 270
rect 14059 236 14093 270
rect 14127 236 14161 270
rect 14195 236 14229 270
rect 14263 236 14297 270
rect 14331 236 14365 270
rect 14399 236 14433 270
rect 14467 236 14501 270
rect 14535 236 14569 270
rect 14603 236 14637 270
rect 14671 236 14739 270
rect 8119 -96 8141 -62
rect 8175 -96 8211 -62
rect 8245 -96 8281 -62
rect 8315 -96 8351 -62
rect 8385 -96 8421 -62
rect 8455 -96 8491 -62
rect 8525 -96 8561 -62
rect 8595 -96 8631 -62
rect 8665 -96 8701 -62
rect 8735 -96 8771 -62
rect 8805 -96 8841 -62
rect 8875 -96 8911 -62
rect 8945 -96 8981 -62
rect 9015 -96 9051 -62
rect 9085 -96 9121 -62
rect 9155 -96 9191 -62
rect 9225 -96 9261 -62
rect 9295 -96 9331 -62
rect 9365 -96 9401 -62
rect 9435 -96 9471 -62
rect 9505 -96 9541 -62
rect 9575 -96 9611 -62
rect 9645 -96 9681 -62
rect 9715 -96 9751 -62
rect 9785 -96 9821 -62
rect 9855 -96 9891 -62
rect 9925 -96 9961 -62
rect 9995 -96 10031 -62
rect 10065 -96 10101 -62
rect 10135 -96 10170 -62
rect 10204 -96 10239 -62
rect 10273 -96 10308 -62
rect 10342 -96 10377 -62
rect 10411 -96 10446 -62
rect 10480 -96 10501 -62
rect 11314 -71 12838 -35
rect 8119 -140 10501 -96
rect 11128 -105 11314 -96
rect 11348 -105 11385 -71
rect 11419 -105 11456 -71
rect 11490 -105 11527 -71
rect 11561 -105 11598 -71
rect 11632 -105 11669 -71
rect 11703 -105 11740 -71
rect 11774 -105 11811 -71
rect 11845 -105 11882 -71
rect 11916 -105 11953 -71
rect 11987 -105 12024 -71
rect 12058 -105 12095 -71
rect 12129 -105 12166 -71
rect 12200 -105 12237 -71
rect 12271 -105 12308 -71
rect 12342 -105 12379 -71
rect 12413 -105 12450 -71
rect 12484 -105 12521 -71
rect 12555 -105 12592 -71
rect 12626 -105 12663 -71
rect 12697 -105 12734 -71
rect 12768 -105 12804 -71
rect 11128 -140 12838 -105
rect 8149 -174 8184 -140
rect 8218 -174 8253 -140
rect 8287 -174 8322 -140
rect 8356 -174 8390 -140
rect 8424 -174 8458 -140
rect 8492 -174 8526 -140
rect 8560 -174 8594 -140
rect 8628 -174 8662 -140
rect 8696 -174 8730 -140
rect 8764 -174 8798 -140
rect 8832 -174 8866 -140
rect 8900 -174 8934 -140
rect 8968 -174 9002 -140
rect 9036 -174 9070 -140
rect 9104 -174 9138 -140
rect 9172 -174 9206 -140
rect 9240 -174 9274 -140
rect 9308 -174 9342 -140
rect 9376 -174 9410 -140
rect 9444 -174 9478 -140
rect 9512 -174 9546 -140
rect 9580 -174 9614 -140
rect 9648 -174 9682 -140
rect 9716 -174 9750 -140
rect 9784 -174 9818 -140
rect 9852 -174 9886 -140
rect 9920 -174 9954 -140
rect 9988 -174 10022 -140
rect 10056 -174 10090 -140
rect 10124 -174 10158 -140
rect 10192 -174 10226 -140
rect 10260 -174 10294 -140
rect 10328 -174 10362 -140
rect 10396 -174 10430 -140
rect 10464 -174 10498 -140
rect 11144 -174 11178 -140
rect 11212 -174 11246 -140
rect 11280 -141 12838 -140
rect 11280 -174 11314 -141
rect 8119 -191 10501 -174
rect 11128 -175 11314 -174
rect 11348 -175 11385 -141
rect 11419 -175 11456 -141
rect 11490 -175 11527 -141
rect 11561 -175 11598 -141
rect 11632 -175 11669 -141
rect 11703 -175 11740 -141
rect 11774 -175 11811 -141
rect 11845 -175 11882 -141
rect 11916 -175 11953 -141
rect 11987 -175 12024 -141
rect 12058 -175 12095 -141
rect 12129 -175 12166 -141
rect 12200 -175 12237 -141
rect 12271 -175 12308 -141
rect 12342 -175 12379 -141
rect 12413 -175 12450 -141
rect 12484 -175 12521 -141
rect 12555 -175 12592 -141
rect 12626 -175 12663 -141
rect 12697 -175 12734 -141
rect 12768 -175 12804 -141
rect 11128 -191 12838 -175
<< mvnsubdiff >>
rect 1166 8579 4444 8580
rect 1166 8545 1234 8579
rect 1268 8545 1302 8579
rect 1336 8545 1370 8579
rect 1404 8545 1438 8579
rect 1472 8545 1506 8579
rect 1540 8545 1574 8579
rect 1608 8545 1642 8579
rect 1676 8545 1710 8579
rect 1744 8545 1778 8579
rect 1812 8545 1846 8579
rect 1880 8545 1914 8579
rect 1948 8545 1982 8579
rect 2016 8545 2050 8579
rect 2084 8545 2118 8579
rect 2152 8545 2186 8579
rect 2220 8545 2254 8579
rect 2288 8545 2322 8579
rect 2356 8545 2390 8579
rect 2424 8545 2458 8579
rect 2492 8545 2526 8579
rect 2560 8545 2594 8579
rect 2628 8545 2662 8579
rect 2696 8545 2730 8579
rect 2764 8545 2798 8579
rect 2832 8545 2866 8579
rect 2900 8545 2934 8579
rect 2968 8545 3002 8579
rect 3036 8545 3070 8579
rect 3104 8545 3138 8579
rect 3172 8545 3206 8579
rect 3240 8545 3274 8579
rect 3308 8545 3342 8579
rect 3376 8545 3410 8579
rect 3444 8545 3478 8579
rect 3512 8545 3546 8579
rect 3580 8545 3614 8579
rect 3648 8545 3682 8579
rect 3716 8545 3750 8579
rect 3784 8545 3818 8579
rect 3852 8545 3886 8579
rect 3920 8545 3954 8579
rect 3988 8545 4022 8579
rect 4056 8545 4090 8579
rect 4124 8545 4158 8579
rect 4192 8545 4226 8579
rect 4260 8545 4294 8579
rect 4328 8545 4444 8579
rect 1166 8544 4444 8545
rect 1166 8489 1202 8544
rect 1166 8455 1167 8489
rect 1201 8455 1202 8489
rect 4408 8512 4444 8544
rect 1166 8421 1202 8455
rect 4408 8478 4409 8512
rect 4443 8478 4444 8512
rect 4408 8444 4444 8478
rect 1166 8387 1167 8421
rect 1201 8387 1202 8421
rect 1166 8353 1202 8387
rect 1166 8319 1167 8353
rect 1201 8319 1202 8353
rect 1166 8285 1202 8319
rect 1166 8251 1167 8285
rect 1201 8251 1202 8285
rect 1166 8217 1202 8251
rect 1166 8183 1167 8217
rect 1201 8183 1202 8217
rect 1166 8149 1202 8183
rect 1166 8115 1167 8149
rect 1201 8115 1202 8149
rect 1166 8081 1202 8115
rect 1166 8047 1167 8081
rect 1201 8047 1202 8081
rect 1166 8013 1202 8047
rect 1166 7979 1167 8013
rect 1201 7979 1202 8013
rect 1166 7945 1202 7979
rect 1166 7911 1167 7945
rect 1201 7911 1202 7945
rect 1166 7877 1202 7911
rect 1166 7843 1167 7877
rect 1201 7843 1202 7877
rect 1166 7809 1202 7843
rect 1166 7775 1167 7809
rect 1201 7775 1202 7809
rect 1166 7741 1202 7775
rect 1166 7707 1167 7741
rect 1201 7707 1202 7741
rect 1166 7673 1202 7707
rect 1166 7639 1167 7673
rect 1201 7639 1202 7673
rect 1166 7605 1202 7639
rect 1166 7571 1167 7605
rect 1201 7571 1202 7605
rect 1166 7537 1202 7571
rect 1166 7503 1167 7537
rect 1201 7503 1202 7537
rect 1166 7469 1202 7503
rect 1166 7435 1167 7469
rect 1201 7435 1202 7469
rect 1166 7401 1202 7435
rect 1166 7367 1167 7401
rect 1201 7367 1202 7401
rect 4408 8410 4409 8444
rect 4443 8410 4444 8444
rect 4408 8376 4444 8410
rect 4408 8342 4409 8376
rect 4443 8342 4444 8376
rect 4408 8308 4444 8342
rect 4408 8274 4409 8308
rect 4443 8274 4444 8308
rect 4408 8240 4444 8274
rect 4408 8206 4409 8240
rect 4443 8206 4444 8240
rect 4408 8172 4444 8206
rect 4408 8138 4409 8172
rect 4443 8138 4444 8172
rect 4408 8104 4444 8138
rect 4408 8070 4409 8104
rect 4443 8070 4444 8104
rect 4408 8036 4444 8070
rect 4408 8002 4409 8036
rect 4443 8002 4444 8036
rect 4408 7968 4444 8002
rect 4408 7934 4409 7968
rect 4443 7934 4444 7968
rect 4408 7900 4444 7934
rect 4408 7866 4409 7900
rect 4443 7866 4444 7900
rect 4408 7832 4444 7866
rect 4408 7798 4409 7832
rect 4443 7798 4444 7832
rect 4408 7764 4444 7798
rect 4408 7730 4409 7764
rect 4443 7730 4444 7764
rect 4408 7696 4444 7730
rect 4408 7662 4409 7696
rect 4443 7662 4444 7696
rect 4408 7628 4444 7662
rect 4408 7594 4409 7628
rect 4443 7594 4444 7628
rect 4408 7560 4444 7594
rect 4408 7526 4409 7560
rect 4443 7526 4444 7560
rect 4408 7492 4444 7526
rect 4408 7458 4409 7492
rect 4443 7458 4444 7492
rect 4408 7424 4444 7458
rect 1166 7333 1202 7367
rect 4408 7390 4409 7424
rect 4443 7390 4444 7424
rect 4408 7356 4444 7390
rect 1166 7299 1167 7333
rect 1201 7299 1202 7333
rect 1166 7267 1202 7299
rect 4408 7322 4409 7356
rect 4443 7322 4444 7356
rect 4408 7267 4444 7322
rect 1166 7266 4444 7267
rect 1166 7232 1291 7266
rect 1325 7232 1359 7266
rect 1393 7232 1427 7266
rect 1461 7232 1495 7266
rect 1529 7232 1622 7266
rect 1656 7232 1690 7266
rect 1724 7232 1758 7266
rect 1792 7232 1826 7266
rect 1860 7232 1894 7266
rect 1928 7232 1962 7266
rect 1996 7232 2030 7266
rect 2064 7232 2098 7266
rect 2132 7232 2166 7266
rect 2200 7232 2234 7266
rect 2268 7232 2302 7266
rect 2336 7232 2370 7266
rect 2404 7232 2438 7266
rect 2472 7232 2506 7266
rect 2540 7232 2574 7266
rect 2608 7232 2642 7266
rect 2676 7232 2710 7266
rect 2744 7232 2778 7266
rect 2812 7232 2846 7266
rect 2880 7232 2914 7266
rect 2948 7232 2982 7266
rect 3016 7232 3050 7266
rect 3084 7232 3118 7266
rect 3152 7232 3186 7266
rect 3220 7232 3254 7266
rect 3288 7232 3322 7266
rect 3356 7232 3390 7266
rect 3424 7232 3458 7266
rect 3492 7232 3526 7266
rect 3560 7232 3594 7266
rect 3628 7232 3662 7266
rect 3696 7232 3730 7266
rect 3764 7232 3798 7266
rect 3832 7232 3866 7266
rect 3900 7232 3934 7266
rect 3968 7232 4002 7266
rect 4036 7232 4070 7266
rect 4104 7232 4138 7266
rect 4172 7232 4206 7266
rect 4240 7232 4274 7266
rect 4308 7232 4342 7266
rect 4376 7232 4444 7266
rect 1166 7231 4444 7232
rect 13193 4240 13227 4326
rect 13193 4172 13227 4206
rect 14983 4302 15017 4326
rect 14983 4234 15017 4268
rect 13193 4104 13227 4138
rect 13193 4036 13227 4070
rect 13193 3968 13227 4002
rect 13193 3900 13227 3934
rect 13193 3832 13227 3866
rect 13193 3764 13227 3798
rect 13193 3696 13227 3730
rect 13193 3628 13227 3662
rect 13193 3560 13227 3594
rect 13193 3492 13227 3526
rect 13193 3424 13227 3458
rect 13193 3356 13227 3390
rect 13193 3288 13227 3322
rect 13193 3220 13227 3254
rect 14983 4166 15017 4200
rect 14983 4098 15017 4132
rect 14983 4030 15017 4064
rect 14983 3962 15017 3996
rect 14983 3894 15017 3928
rect 14983 3826 15017 3860
rect 14983 3758 15017 3792
rect 14983 3690 15017 3724
rect 14983 3622 15017 3656
rect 14983 3554 15017 3588
rect 14983 3486 15017 3520
rect 14983 3418 15017 3452
rect 14983 3350 15017 3384
rect 14983 3282 15017 3316
rect 13193 3152 13227 3186
rect 14983 3214 15017 3248
rect 14983 3146 15017 3180
rect 13193 3084 13227 3118
rect 13193 3016 13227 3050
rect 14983 3078 15017 3112
rect 14983 3010 15017 3044
rect 13193 2948 13227 2982
rect 13193 2883 13227 2914
rect 14983 2942 15017 2976
rect 14983 2883 15017 2908
rect 13193 2881 15017 2883
rect 13193 2880 13261 2881
rect 13227 2847 13261 2880
rect 13295 2847 13330 2881
rect 13364 2847 13399 2881
rect 13433 2847 13468 2881
rect 13502 2847 13537 2881
rect 13571 2847 13606 2881
rect 13640 2847 13675 2881
rect 13709 2847 13744 2881
rect 13778 2847 13813 2881
rect 13847 2847 13882 2881
rect 13916 2847 13951 2881
rect 13985 2847 14020 2881
rect 14054 2847 14089 2881
rect 14123 2847 14158 2881
rect 14192 2847 14227 2881
rect 14261 2847 14296 2881
rect 14330 2847 14365 2881
rect 14399 2847 14434 2881
rect 14468 2847 14503 2881
rect 14537 2847 14572 2881
rect 14606 2847 14641 2881
rect 14675 2847 14710 2881
rect 14744 2847 14779 2881
rect 14813 2847 14847 2881
rect 14881 2847 14915 2881
rect 14949 2874 15017 2881
rect 14949 2847 14983 2874
rect 13227 2846 14983 2847
rect 13193 2845 14983 2846
rect 13193 2812 13227 2845
rect 13193 2744 13227 2778
rect 13193 2676 13227 2710
rect 14983 2806 15017 2840
rect 14983 2738 15017 2772
rect 13193 2608 13227 2642
rect 13193 2540 13227 2574
rect 13193 2472 13227 2506
rect 13193 2404 13227 2438
rect 13193 2336 13227 2370
rect 13193 2268 13227 2302
rect 13193 2200 13227 2234
rect 13193 2132 13227 2166
rect 13193 2064 13227 2098
rect 13193 1996 13227 2030
rect 13193 1928 13227 1962
rect 13193 1860 13227 1894
rect 13193 1792 13227 1826
rect 13193 1724 13227 1758
rect 13193 1656 13227 1690
rect 13193 1588 13227 1622
rect 13193 1520 13227 1554
rect 13193 1452 13227 1486
rect 13193 1384 13227 1418
rect 13193 1316 13227 1350
rect 13193 1248 13227 1282
rect 13193 1180 13227 1214
rect 13193 1112 13227 1146
rect 13193 1044 13227 1078
rect 13193 976 13227 1010
rect 13193 908 13227 942
rect 13193 840 13227 874
rect 13193 772 13227 806
rect 13193 704 13227 738
rect 13193 636 13227 670
rect 13193 568 13227 602
rect 13193 500 13227 534
rect 13193 432 13227 466
rect 13193 364 13227 398
rect 13193 296 13227 330
rect 13193 228 13227 262
rect 14983 2670 15017 2704
rect 14983 2602 15017 2636
rect 14983 2534 15017 2568
rect 14983 2466 15017 2500
rect 14983 2398 15017 2432
rect 14983 2330 15017 2364
rect 14983 2262 15017 2296
rect 14983 2194 15017 2228
rect 14983 2126 15017 2160
rect 14983 2058 15017 2092
rect 14983 1990 15017 2024
rect 14983 1922 15017 1956
rect 14983 1854 15017 1888
rect 14983 1786 15017 1820
rect 14983 1718 15017 1752
rect 14983 1650 15017 1684
rect 14983 1582 15017 1616
rect 14983 1514 15017 1548
rect 14983 1446 15017 1480
rect 14983 1378 15017 1412
rect 14983 1310 15017 1344
rect 14983 1242 15017 1276
rect 14983 1174 15017 1208
rect 14983 1106 15017 1140
rect 14983 1038 15017 1072
rect 14983 970 15017 1004
rect 14983 902 15017 936
rect 14983 834 15017 868
rect 14983 766 15017 800
rect 14983 698 15017 732
rect 14983 630 15017 664
rect 14983 562 15017 596
rect 14983 494 15017 528
rect 14983 426 15017 460
rect 14983 358 15017 392
rect 14983 290 15017 324
rect 13193 160 13227 194
rect 13193 92 13227 126
rect 13193 24 13227 58
rect 14983 222 15017 256
rect 14983 154 15017 188
rect 14983 86 15017 120
rect 14983 24 15017 52
rect 13193 -10 13283 24
rect 13317 -10 13351 24
rect 13385 -10 13419 24
rect 13453 -10 13487 24
rect 13521 -10 13555 24
rect 13589 -10 13623 24
rect 13657 -10 13691 24
rect 13725 -10 13759 24
rect 13793 -10 13827 24
rect 13861 -10 13895 24
rect 13929 -10 13963 24
rect 13997 -10 14031 24
rect 14065 -10 14099 24
rect 14133 -10 14167 24
rect 14201 -10 14235 24
rect 14269 -10 14303 24
rect 14337 -10 14371 24
rect 14405 -10 14439 24
rect 14473 -10 14507 24
rect 14541 -10 14575 24
rect 14609 -10 14643 24
rect 14677 -10 14711 24
rect 14745 -10 14779 24
rect 14813 -10 14847 24
rect 14881 -10 14915 24
rect 14949 -10 15017 24
<< psubdiffcont >>
rect 4731 8757 4749 8766
rect 8071 -96 8105 -62
rect 10515 -96 10549 -62
rect 5769 -174 5803 -140
rect 5838 -174 5872 -140
rect 5907 -174 5941 -140
rect 5976 -174 6010 -140
rect 6045 -174 6079 -140
rect 6114 -174 6148 -140
rect 6183 -174 6217 -140
rect 6252 -174 6286 -140
rect 6321 -174 6355 -140
rect 6390 -174 6424 -140
rect 6459 -174 6493 -140
rect 6528 -174 6562 -140
rect 6597 -174 6631 -140
rect 6666 -174 6700 -140
rect 6735 -174 6769 -140
rect 6804 -174 6838 -140
rect 6873 -174 6907 -140
rect 6942 -174 6976 -140
rect 7011 -174 7045 -140
rect 7080 -174 7114 -140
rect 7149 -174 7183 -140
rect 7218 -174 7252 -140
rect 7287 -174 7321 -140
rect 7356 -174 7390 -140
rect 7425 -174 7459 -140
rect 7494 -174 7528 -140
rect 7563 -174 7597 -140
rect 7632 -174 7666 -140
rect 7701 -174 7735 -140
rect 7770 -174 7804 -140
rect 7839 -174 7873 -140
rect 7908 -174 7942 -140
rect 7977 -174 8011 -140
rect 8046 -174 8080 -140
rect 8115 -174 8119 -140
rect 10501 -174 10532 -140
rect 10566 -174 10600 -140
rect 10634 -174 10668 -140
rect 10702 -174 10736 -140
rect 10770 -174 10804 -140
rect 10838 -174 10872 -140
rect 10906 -174 10940 -140
rect 10974 -174 11008 -140
rect 11042 -174 11076 -140
rect 11110 -174 11128 -140
rect 12316 -289 12350 -255
rect 12384 -289 12418 -255
rect 12452 -289 12486 -255
rect 12520 -289 12554 -255
rect 12588 -289 12622 -255
rect 12656 -289 12690 -255
rect 12724 -289 12758 -255
rect 12316 -359 12350 -325
rect 12384 -359 12418 -325
rect 12452 -359 12486 -325
rect 12520 -359 12554 -325
rect 12588 -359 12622 -325
rect 12656 -359 12690 -325
rect 12724 -359 12758 -325
rect 12316 -429 12350 -395
rect 12384 -429 12418 -395
rect 12452 -429 12486 -395
rect 12520 -429 12554 -395
rect 12588 -429 12622 -395
rect 12656 -429 12690 -395
rect 12724 -429 12758 -395
rect 12316 -499 12350 -465
rect 12384 -499 12418 -465
rect 12452 -499 12486 -465
rect 12520 -499 12554 -465
rect 12588 -499 12622 -465
rect 12656 -499 12690 -465
rect 12724 -499 12758 -465
rect 12316 -569 12350 -535
rect 12384 -569 12418 -535
rect 12452 -569 12486 -535
rect 12520 -569 12554 -535
rect 12588 -569 12622 -535
rect 12656 -569 12690 -535
rect 12724 -569 12758 -535
rect 12316 -640 12350 -606
rect 12384 -640 12418 -606
rect 12452 -640 12486 -606
rect 12520 -640 12554 -606
rect 12588 -640 12622 -606
rect 12656 -640 12690 -606
rect 12724 -640 12758 -606
rect 12316 -711 12350 -677
rect 12384 -711 12418 -677
rect 12452 -711 12486 -677
rect 12520 -711 12554 -677
rect 12588 -711 12622 -677
rect 12656 -711 12690 -677
rect 12724 -711 12758 -677
rect 12316 -782 12350 -748
rect 12384 -782 12418 -748
rect 12452 -782 12486 -748
rect 12520 -782 12554 -748
rect 12588 -782 12622 -748
rect 12656 -782 12690 -748
rect 12724 -782 12758 -748
rect 12316 -853 12350 -819
rect 12384 -853 12418 -819
rect 12452 -853 12486 -819
rect 12520 -853 12554 -819
rect 12588 -853 12622 -819
rect 12656 -853 12690 -819
rect 12724 -853 12758 -819
rect 12316 -924 12350 -890
rect 12384 -924 12418 -890
rect 12452 -924 12486 -890
rect 12520 -924 12554 -890
rect 12588 -924 12622 -890
rect 12656 -924 12690 -890
rect 12724 -924 12758 -890
rect 12316 -995 12350 -961
rect 12384 -995 12418 -961
rect 12452 -995 12486 -961
rect 12520 -995 12554 -961
rect 12588 -995 12622 -961
rect 12656 -995 12690 -961
rect 12724 -995 12758 -961
<< mvpsubdiffcont >>
rect 800 8733 834 8767
rect 907 8757 941 8791
rect 975 8757 1009 8791
rect 1043 8757 1077 8791
rect 1111 8757 1145 8791
rect 1179 8757 1213 8791
rect 1247 8757 1281 8791
rect 1315 8757 1349 8791
rect 1383 8757 1417 8791
rect 1451 8757 1485 8791
rect 1519 8757 1553 8791
rect 1587 8757 1621 8791
rect 1655 8757 1689 8791
rect 1723 8757 1757 8791
rect 1791 8757 1825 8791
rect 1859 8757 1893 8791
rect 1927 8757 1961 8791
rect 1995 8757 2029 8791
rect 2063 8757 2097 8791
rect 2131 8757 2165 8791
rect 2199 8757 2233 8791
rect 2267 8757 2301 8791
rect 2335 8757 2369 8791
rect 2403 8757 2437 8791
rect 2471 8757 2505 8791
rect 2539 8757 2573 8791
rect 2607 8757 2641 8791
rect 2675 8757 2709 8791
rect 2743 8757 2777 8791
rect 2811 8757 2845 8791
rect 2879 8757 2913 8791
rect 2947 8757 2981 8791
rect 3015 8757 3049 8791
rect 3083 8757 3117 8791
rect 3151 8757 3185 8791
rect 3219 8757 3253 8791
rect 3287 8757 3321 8791
rect 3355 8757 3389 8791
rect 3423 8757 3457 8791
rect 3491 8757 3525 8791
rect 3559 8757 3593 8791
rect 3627 8757 3661 8791
rect 3695 8757 3729 8791
rect 3763 8757 3797 8791
rect 3831 8757 3865 8791
rect 3899 8757 3933 8791
rect 3967 8757 4001 8791
rect 4035 8757 4069 8791
rect 4103 8757 4137 8791
rect 4171 8757 4205 8791
rect 4239 8757 4273 8791
rect 4307 8757 4341 8791
rect 4375 8757 4409 8791
rect 4443 8757 4477 8791
rect 4511 8757 4545 8791
rect 4579 8757 4613 8791
rect 4647 8757 4681 8791
rect 4715 8766 4749 8791
rect 4715 8757 4731 8766
rect 800 8665 834 8699
rect 800 8597 834 8631
rect 800 8529 834 8563
rect 800 8461 834 8495
rect 800 8393 834 8427
rect 800 8325 834 8359
rect 800 8257 834 8291
rect 800 8189 834 8223
rect 800 8121 834 8155
rect 800 8053 834 8087
rect 800 7985 834 8019
rect 800 7917 834 7951
rect 800 7849 834 7883
rect 800 7781 834 7815
rect 800 7713 834 7747
rect 800 7645 834 7679
rect 800 7577 834 7611
rect 800 7509 834 7543
rect 800 7441 834 7475
rect 800 7373 834 7407
rect 800 7305 834 7339
rect 800 7237 834 7271
rect 800 7169 834 7203
rect 841 7044 875 7078
rect 909 7044 943 7078
rect 977 7044 1011 7078
rect 1045 7044 1079 7078
rect 1113 7044 1147 7078
rect 1181 7044 1215 7078
rect 1249 7044 1283 7078
rect 1317 7044 1351 7078
rect 1385 7044 1419 7078
rect 1453 7044 1487 7078
rect 1521 7044 1555 7078
rect 1589 7044 1623 7078
rect 1657 7044 1691 7078
rect 1725 7044 1759 7078
rect 1793 7044 1827 7078
rect 1861 7044 1895 7078
rect 1929 7044 1963 7078
rect 1997 7044 2031 7078
rect 2065 7044 2099 7078
rect 2133 7044 2167 7078
rect 2201 7044 2235 7078
rect 2269 7044 2303 7078
rect 2337 7044 2371 7078
rect 2405 7044 2439 7078
rect 2473 7044 2507 7078
rect 2541 7044 2575 7078
rect 2609 7044 2643 7078
rect 2677 7044 2711 7078
rect 2745 7044 2779 7078
rect 2813 7044 2847 7078
rect 2881 7044 2915 7078
rect 2949 7044 2983 7078
rect 3017 7044 3051 7078
rect 3085 7044 3119 7078
rect 3153 7044 3187 7078
rect 3221 7044 3255 7078
rect 3289 7044 3323 7078
rect 3357 7044 3391 7078
rect 3425 7044 3459 7078
rect 3493 7044 3527 7078
rect 3561 7044 3595 7078
rect 3629 7044 3663 7078
rect 3697 7044 3731 7078
rect 3765 7044 3799 7078
rect 3833 7044 3867 7078
rect 3901 7044 3935 7078
rect 3969 7044 4003 7078
rect 4037 7044 4071 7078
rect 4105 7044 4139 7078
rect 4173 7044 4207 7078
rect 4241 7044 4275 7078
rect 4309 7044 4343 7078
rect 4377 7044 4411 7078
rect 4445 7044 4479 7078
rect 4513 7044 4547 7078
rect 4581 7044 4615 7078
rect 4649 7044 4683 7078
rect 4446 6973 4480 7007
rect 4518 6973 4552 7007
rect 4590 6973 4624 7007
rect 4662 6973 4696 7007
rect 4446 6905 4480 6939
rect 4518 6905 4552 6939
rect 4590 6905 4624 6939
rect 4662 6905 4696 6939
rect 4446 6837 4480 6871
rect 4518 6837 4552 6871
rect 4590 6837 4624 6871
rect 4662 6837 4696 6871
rect 4446 6769 4480 6803
rect 4518 6769 4552 6803
rect 4590 6769 4624 6803
rect 4662 6769 4696 6803
rect -850 6725 -816 6759
rect -781 6725 -747 6759
rect -712 6725 -678 6759
rect -643 6725 -609 6759
rect -574 6725 -540 6759
rect -505 6725 -471 6759
rect -436 6725 -402 6759
rect -367 6725 -333 6759
rect -298 6725 -264 6759
rect -229 6725 -195 6759
rect -160 6725 -126 6759
rect -91 6725 -57 6759
rect -22 6725 12 6759
rect 47 6725 81 6759
rect 116 6725 150 6759
rect 185 6725 219 6759
rect 254 6725 288 6759
rect 323 6725 357 6759
rect 391 6725 425 6759
rect 459 6725 493 6759
rect 527 6725 561 6759
rect 595 6725 629 6759
rect 663 6725 697 6759
rect 731 6725 765 6759
rect 799 6725 833 6759
rect 867 6725 901 6759
rect -850 6655 -816 6689
rect -781 6655 -747 6689
rect -712 6655 -678 6689
rect -643 6655 -609 6689
rect -574 6655 -540 6689
rect -505 6655 -471 6689
rect -436 6655 -402 6689
rect -367 6655 -333 6689
rect -298 6655 -264 6689
rect -229 6655 -195 6689
rect -160 6655 -126 6689
rect -91 6655 -57 6689
rect -22 6655 12 6689
rect 47 6655 81 6689
rect 116 6655 150 6689
rect 185 6655 219 6689
rect 254 6655 288 6689
rect 323 6655 357 6689
rect 391 6655 425 6689
rect 459 6655 493 6689
rect 527 6655 561 6689
rect 595 6655 629 6689
rect 663 6655 697 6689
rect 731 6655 765 6689
rect 799 6655 833 6689
rect 867 6655 901 6689
rect -850 6585 -816 6619
rect -781 6585 -747 6619
rect -712 6585 -678 6619
rect -643 6585 -609 6619
rect -574 6585 -540 6619
rect -505 6585 -471 6619
rect -436 6585 -402 6619
rect -367 6585 -333 6619
rect -298 6585 -264 6619
rect -229 6585 -195 6619
rect -160 6585 -126 6619
rect -91 6585 -57 6619
rect -22 6585 12 6619
rect 47 6585 81 6619
rect 116 6585 150 6619
rect 185 6585 219 6619
rect 254 6585 288 6619
rect 323 6585 357 6619
rect 391 6585 425 6619
rect 459 6585 493 6619
rect 527 6585 561 6619
rect 595 6585 629 6619
rect 663 6585 697 6619
rect 731 6585 765 6619
rect 799 6585 833 6619
rect 867 6585 901 6619
rect -850 6515 -816 6549
rect -781 6515 -747 6549
rect -712 6515 -678 6549
rect -643 6515 -609 6549
rect -574 6515 -540 6549
rect -505 6515 -471 6549
rect -436 6515 -402 6549
rect -367 6515 -333 6549
rect -298 6515 -264 6549
rect -229 6515 -195 6549
rect -160 6515 -126 6549
rect -91 6515 -57 6549
rect -22 6515 12 6549
rect 47 6515 81 6549
rect 116 6515 150 6549
rect 185 6515 219 6549
rect 254 6515 288 6549
rect 323 6515 357 6549
rect 391 6515 425 6549
rect 459 6515 493 6549
rect 527 6515 561 6549
rect 595 6515 629 6549
rect 663 6515 697 6549
rect 731 6515 765 6549
rect 799 6515 833 6549
rect 867 6515 901 6549
rect -850 6445 -816 6479
rect -781 6445 -747 6479
rect -712 6445 -678 6479
rect -643 6445 -609 6479
rect -574 6445 -540 6479
rect -505 6445 -471 6479
rect -436 6445 -402 6479
rect -367 6445 -333 6479
rect -298 6445 -264 6479
rect -229 6445 -195 6479
rect -160 6445 -126 6479
rect -91 6445 -57 6479
rect -22 6445 12 6479
rect 47 6445 81 6479
rect 116 6445 150 6479
rect 185 6445 219 6479
rect 254 6445 288 6479
rect 323 6445 357 6479
rect 391 6445 425 6479
rect 459 6445 493 6479
rect 527 6445 561 6479
rect 595 6445 629 6479
rect 663 6445 697 6479
rect 731 6445 765 6479
rect 799 6445 833 6479
rect 867 6445 901 6479
rect -850 6375 -816 6409
rect -781 6375 -747 6409
rect -712 6375 -678 6409
rect -643 6375 -609 6409
rect -574 6375 -540 6409
rect -505 6375 -471 6409
rect -436 6375 -402 6409
rect -367 6375 -333 6409
rect -298 6375 -264 6409
rect -229 6375 -195 6409
rect -160 6375 -126 6409
rect -91 6375 -57 6409
rect -22 6375 12 6409
rect 47 6375 81 6409
rect 116 6375 150 6409
rect 185 6375 219 6409
rect 254 6375 288 6409
rect 323 6375 357 6409
rect 391 6375 425 6409
rect 459 6375 493 6409
rect 527 6375 561 6409
rect 595 6375 629 6409
rect 663 6375 697 6409
rect 731 6375 765 6409
rect 799 6375 833 6409
rect 867 6375 901 6409
rect -850 6305 -816 6339
rect -781 6305 -747 6339
rect -712 6305 -678 6339
rect -643 6305 -609 6339
rect -574 6305 -540 6339
rect -505 6305 -471 6339
rect -436 6305 -402 6339
rect -367 6305 -333 6339
rect -298 6305 -264 6339
rect -229 6305 -195 6339
rect -160 6305 -126 6339
rect -91 6305 -57 6339
rect -22 6305 12 6339
rect 47 6305 81 6339
rect 116 6305 150 6339
rect 185 6305 219 6339
rect 254 6305 288 6339
rect 323 6305 357 6339
rect 391 6305 425 6339
rect 459 6305 493 6339
rect 527 6305 561 6339
rect 595 6305 629 6339
rect 663 6305 697 6339
rect 731 6305 765 6339
rect 799 6305 833 6339
rect 867 6305 901 6339
rect -850 6235 -816 6269
rect -781 6235 -747 6269
rect -712 6235 -678 6269
rect -643 6235 -609 6269
rect -574 6235 -540 6269
rect -505 6235 -471 6269
rect -436 6235 -402 6269
rect -367 6235 -333 6269
rect -298 6235 -264 6269
rect -229 6235 -195 6269
rect -160 6235 -126 6269
rect -91 6235 -57 6269
rect -22 6235 12 6269
rect 47 6235 81 6269
rect 116 6235 150 6269
rect 185 6235 219 6269
rect 254 6235 288 6269
rect 323 6235 357 6269
rect 391 6235 425 6269
rect 459 6235 493 6269
rect 527 6235 561 6269
rect 595 6235 629 6269
rect 663 6235 697 6269
rect 731 6235 765 6269
rect 799 6235 833 6269
rect 867 6235 901 6269
rect -850 6165 -816 6199
rect -781 6165 -747 6199
rect -712 6165 -678 6199
rect -643 6165 -609 6199
rect -574 6165 -540 6199
rect -505 6165 -471 6199
rect -436 6165 -402 6199
rect -367 6165 -333 6199
rect -298 6165 -264 6199
rect -229 6165 -195 6199
rect -160 6165 -126 6199
rect -91 6165 -57 6199
rect -22 6165 12 6199
rect 47 6165 81 6199
rect 116 6165 150 6199
rect 185 6165 219 6199
rect 254 6165 288 6199
rect 323 6165 357 6199
rect 391 6165 425 6199
rect 459 6165 493 6199
rect 527 6165 561 6199
rect 595 6165 629 6199
rect 663 6165 697 6199
rect 731 6165 765 6199
rect 799 6165 833 6199
rect 867 6165 901 6199
rect -850 6095 -816 6129
rect -781 6095 -747 6129
rect -712 6095 -678 6129
rect -643 6095 -609 6129
rect -574 6095 -540 6129
rect -505 6095 -471 6129
rect -436 6095 -402 6129
rect -367 6095 -333 6129
rect -298 6095 -264 6129
rect -229 6095 -195 6129
rect -160 6095 -126 6129
rect -91 6095 -57 6129
rect -22 6095 12 6129
rect 47 6095 81 6129
rect 116 6095 150 6129
rect 185 6095 219 6129
rect 254 6095 288 6129
rect 323 6095 357 6129
rect 391 6095 425 6129
rect 459 6095 493 6129
rect 527 6095 561 6129
rect 595 6095 629 6129
rect 663 6095 697 6129
rect 731 6095 765 6129
rect 799 6095 833 6129
rect 867 6095 901 6129
rect 4446 6701 4480 6735
rect 4518 6701 4552 6735
rect 4590 6701 4624 6735
rect 4662 6701 4696 6735
rect 4446 6633 4480 6667
rect 4518 6633 4552 6667
rect 4590 6633 4624 6667
rect 4662 6633 4696 6667
rect 4446 6565 4480 6599
rect 4518 6565 4552 6599
rect 4590 6565 4624 6599
rect 4662 6565 4696 6599
rect 4446 6497 4480 6531
rect 4518 6497 4552 6531
rect 4590 6497 4624 6531
rect 4662 6497 4696 6531
rect 4446 6429 4480 6463
rect 4518 6429 4552 6463
rect 4590 6429 4624 6463
rect 4662 6429 4696 6463
rect 4446 6361 4480 6395
rect 4518 6361 4552 6395
rect 4590 6361 4624 6395
rect 4662 6361 4696 6395
rect 4446 6293 4480 6327
rect 4518 6293 4552 6327
rect 4590 6293 4624 6327
rect 4662 6293 4696 6327
rect 4446 6225 4480 6259
rect 4518 6225 4552 6259
rect 4590 6225 4624 6259
rect 4662 6225 4696 6259
rect 4446 6157 4480 6191
rect 4518 6157 4552 6191
rect 4590 6157 4624 6191
rect 4662 6157 4696 6191
rect 4446 6089 4480 6123
rect 4518 6089 4552 6123
rect 4590 6089 4624 6123
rect 4662 6089 4696 6123
rect 4446 6021 4480 6055
rect 4518 6021 4552 6055
rect 4590 6021 4624 6055
rect 4662 6021 4696 6055
rect 4446 5953 4480 5987
rect 4518 5953 4552 5987
rect 4590 5953 4624 5987
rect 4662 5953 4696 5987
rect 4446 5885 4480 5919
rect 4518 5885 4552 5919
rect 4590 5885 4624 5919
rect 4662 5885 4696 5919
rect 4446 5816 4480 5850
rect 4518 5816 4552 5850
rect 4590 5816 4624 5850
rect 4662 5816 4696 5850
rect 4102 5745 4136 5779
rect 4172 5745 4206 5779
rect 4242 5745 4276 5779
rect 4312 5745 4346 5779
rect 4382 5745 4416 5779
rect 4452 5745 4486 5779
rect 4522 5745 4556 5779
rect 4592 5745 4626 5779
rect 4662 5745 4696 5779
rect 4102 5676 4136 5710
rect 4172 5676 4206 5710
rect 4242 5676 4276 5710
rect 4312 5676 4346 5710
rect 4382 5676 4416 5710
rect 4452 5676 4486 5710
rect 4522 5676 4556 5710
rect 4592 5676 4626 5710
rect 4662 5676 4696 5710
rect 4102 5607 4136 5641
rect 4172 5607 4206 5641
rect 4242 5607 4276 5641
rect 4312 5607 4346 5641
rect 4382 5607 4416 5641
rect 4452 5607 4486 5641
rect 4522 5607 4556 5641
rect 4592 5607 4626 5641
rect 4662 5607 4696 5641
rect 4102 5538 4136 5572
rect 4172 5538 4206 5572
rect 4242 5538 4276 5572
rect 4312 5538 4346 5572
rect 4382 5538 4416 5572
rect 4452 5538 4486 5572
rect 4522 5538 4556 5572
rect 4592 5538 4626 5572
rect 4662 5538 4696 5572
rect 4102 5469 4136 5503
rect 4172 5469 4206 5503
rect 4242 5469 4276 5503
rect 4312 5469 4346 5503
rect 4382 5469 4416 5503
rect 4452 5469 4486 5503
rect 4522 5469 4556 5503
rect 4592 5469 4626 5503
rect 4662 5469 4696 5503
rect 4102 5400 4136 5434
rect 4172 5400 4206 5434
rect 4242 5400 4276 5434
rect 4312 5400 4346 5434
rect 4382 5400 4416 5434
rect 4452 5400 4486 5434
rect 4522 5400 4556 5434
rect 4592 5400 4626 5434
rect 4662 5400 4696 5434
rect 4102 5331 4136 5365
rect 4172 5331 4206 5365
rect 4242 5331 4276 5365
rect 4312 5331 4346 5365
rect 4382 5331 4416 5365
rect 4452 5331 4486 5365
rect 4522 5331 4556 5365
rect 4592 5331 4626 5365
rect 4662 5331 4696 5365
rect 4102 5262 4136 5296
rect 4172 5262 4206 5296
rect 4242 5262 4276 5296
rect 4312 5262 4346 5296
rect 4382 5262 4416 5296
rect 4452 5262 4486 5296
rect 4522 5262 4556 5296
rect 4592 5262 4626 5296
rect 4662 5262 4696 5296
rect 4102 5193 4136 5227
rect 4172 5193 4206 5227
rect 4242 5193 4276 5227
rect 4312 5193 4346 5227
rect 4382 5193 4416 5227
rect 4452 5193 4486 5227
rect 4522 5193 4556 5227
rect 4592 5193 4626 5227
rect 4662 5193 4696 5227
rect 4102 5124 4136 5158
rect 4172 5124 4206 5158
rect 4242 5124 4276 5158
rect 4312 5124 4346 5158
rect 4382 5124 4416 5158
rect 4452 5124 4486 5158
rect 4522 5124 4556 5158
rect 4592 5124 4626 5158
rect 4662 5124 4696 5158
rect 4102 5055 4136 5089
rect 4172 5055 4206 5089
rect 4242 5055 4276 5089
rect 4312 5055 4346 5089
rect 4382 5055 4416 5089
rect 4452 5055 4486 5089
rect 4522 5055 4556 5089
rect 4592 5055 4626 5089
rect 4662 5055 4696 5089
rect 4102 4985 4136 5019
rect 4172 4985 4206 5019
rect 4242 4985 4276 5019
rect 4312 4985 4346 5019
rect 4382 4985 4416 5019
rect 4452 4985 4486 5019
rect 4522 4985 4556 5019
rect 4592 4985 4626 5019
rect 4662 4985 4696 5019
rect 4102 4915 4136 4949
rect 4172 4915 4206 4949
rect 4242 4915 4276 4949
rect 4312 4915 4346 4949
rect 4382 4915 4416 4949
rect 4452 4915 4486 4949
rect 4522 4915 4556 4949
rect 4592 4915 4626 4949
rect 4662 4915 4696 4949
rect 4102 4845 4136 4879
rect 4172 4845 4206 4879
rect 4242 4845 4276 4879
rect 4312 4845 4346 4879
rect 4382 4845 4416 4879
rect 4452 4845 4486 4879
rect 4522 4845 4556 4879
rect 4592 4845 4626 4879
rect 4662 4845 4696 4879
rect 4102 4775 4136 4809
rect 4172 4775 4206 4809
rect 4242 4775 4276 4809
rect 4312 4775 4346 4809
rect 4382 4775 4416 4809
rect 4452 4775 4486 4809
rect 4522 4775 4556 4809
rect 4592 4775 4626 4809
rect 4662 4775 4696 4809
rect 4102 4705 4136 4739
rect 4172 4705 4206 4739
rect 4242 4705 4276 4739
rect 4312 4705 4346 4739
rect 4382 4705 4416 4739
rect 4452 4705 4486 4739
rect 4522 4705 4556 4739
rect 4592 4705 4626 4739
rect 4662 4705 4696 4739
rect 4102 4635 4136 4669
rect 4172 4635 4206 4669
rect 4242 4635 4276 4669
rect 4312 4635 4346 4669
rect 4382 4635 4416 4669
rect 4452 4635 4486 4669
rect 4522 4635 4556 4669
rect 4592 4635 4626 4669
rect 4662 4635 4696 4669
rect 4102 4565 4136 4599
rect 4172 4565 4206 4599
rect 4242 4565 4276 4599
rect 4312 4565 4346 4599
rect 4382 4565 4416 4599
rect 4452 4565 4486 4599
rect 4522 4565 4556 4599
rect 4592 4565 4626 4599
rect 4662 4565 4696 4599
rect 4102 4495 4136 4529
rect 4172 4495 4206 4529
rect 4242 4495 4276 4529
rect 4312 4495 4346 4529
rect 4382 4495 4416 4529
rect 4452 4495 4486 4529
rect 4522 4495 4556 4529
rect 4592 4495 4626 4529
rect 4662 4495 4696 4529
rect 4102 4425 4136 4459
rect 4172 4425 4206 4459
rect 4242 4425 4276 4459
rect 4312 4425 4346 4459
rect 4382 4425 4416 4459
rect 4452 4425 4486 4459
rect 4522 4425 4556 4459
rect 4592 4425 4626 4459
rect 4662 4425 4696 4459
rect 4102 4355 4136 4389
rect 4172 4355 4206 4389
rect 4242 4355 4276 4389
rect 4312 4355 4346 4389
rect 4382 4355 4416 4389
rect 4452 4355 4486 4389
rect 4522 4355 4556 4389
rect 4592 4355 4626 4389
rect 4662 4355 4696 4389
rect 4102 4285 4136 4319
rect 4172 4285 4206 4319
rect 4242 4285 4276 4319
rect 4312 4285 4346 4319
rect 4382 4285 4416 4319
rect 4452 4285 4486 4319
rect 4522 4285 4556 4319
rect 4592 4285 4626 4319
rect 4662 4285 4696 4319
rect 4102 4215 4136 4249
rect 4172 4215 4206 4249
rect 4242 4215 4276 4249
rect 4312 4215 4346 4249
rect 4382 4215 4416 4249
rect 4452 4215 4486 4249
rect 4522 4215 4556 4249
rect 4592 4215 4626 4249
rect 4662 4215 4696 4249
rect 4102 4145 4136 4179
rect 4172 4145 4206 4179
rect 4242 4145 4276 4179
rect 4312 4145 4346 4179
rect 4382 4145 4416 4179
rect 4452 4145 4486 4179
rect 4522 4145 4556 4179
rect 4592 4145 4626 4179
rect 4662 4145 4696 4179
rect 4731 4148 4765 4182
rect 4801 4148 4835 4182
rect 4871 4148 4905 4182
rect 4941 4148 4975 4182
rect 5011 4148 5045 4182
rect 5081 4148 5115 4182
rect 5151 4148 5185 4182
rect 5221 4148 5255 4182
rect 5291 4148 5325 4182
rect 5360 4148 5394 4182
rect 5429 4148 5463 4182
rect 5498 4148 5532 4182
rect 5567 4148 5601 4182
rect 5636 4148 5670 4182
rect 5705 4148 5739 4182
rect 5774 4148 5808 4182
rect 5843 4148 5877 4182
rect 5912 4148 5946 4182
rect 5981 4148 6015 4182
rect 6050 4148 6084 4182
rect 6119 4148 6153 4182
rect 6188 4148 6222 4182
rect 6257 4148 6291 4182
rect 6326 4148 6360 4182
rect 6395 4148 6429 4182
rect 6464 4148 6498 4182
rect 6533 4148 6567 4182
rect 6602 4148 6636 4182
rect 6671 4148 6705 4182
rect 6740 4148 6774 4182
rect 6809 4148 6843 4182
rect 6878 4148 6912 4182
rect 6947 4148 6981 4182
rect 7016 4148 7050 4182
rect 7085 4148 7119 4182
rect 7154 4148 7188 4182
rect 7223 4148 7257 4182
rect 7292 4148 7326 4182
rect 7361 4148 7395 4182
rect 7430 4148 7464 4182
rect 7499 4148 7533 4182
rect 7568 4148 7602 4182
rect 7637 4148 7671 4182
rect 7706 4148 7740 4182
rect 7775 4148 7809 4182
rect 7844 4148 7878 4182
rect 7913 4148 7947 4182
rect 7982 4148 8016 4182
rect 8051 4148 8085 4182
rect 8120 4148 8154 4182
rect 8189 4148 8223 4182
rect 8258 4148 8292 4182
rect 4102 4075 4136 4109
rect 4172 4075 4206 4109
rect 4242 4075 4276 4109
rect 4312 4075 4346 4109
rect 4382 4075 4416 4109
rect 4452 4075 4486 4109
rect 4522 4075 4556 4109
rect 4592 4075 4626 4109
rect 4662 4075 4696 4109
rect 4731 4050 4765 4084
rect 4801 4050 4835 4084
rect 4871 4050 4905 4084
rect 4941 4050 4975 4084
rect 5011 4050 5045 4084
rect 5081 4050 5115 4084
rect 5151 4050 5185 4084
rect 5221 4050 5255 4084
rect 5291 4050 5325 4084
rect 5360 4050 5394 4084
rect 5429 4050 5463 4084
rect 5498 4050 5532 4084
rect 5567 4050 5601 4084
rect 5636 4050 5670 4084
rect 5705 4050 5739 4084
rect 5774 4050 5808 4084
rect 5843 4050 5877 4084
rect 5912 4050 5946 4084
rect 5981 4050 6015 4084
rect 6050 4050 6084 4084
rect 6119 4050 6153 4084
rect 6188 4050 6222 4084
rect 6257 4050 6291 4084
rect 6326 4050 6360 4084
rect 6395 4050 6429 4084
rect 6464 4050 6498 4084
rect 6533 4050 6567 4084
rect 6602 4050 6636 4084
rect 6671 4050 6705 4084
rect 6740 4050 6774 4084
rect 6809 4050 6843 4084
rect 6878 4050 6912 4084
rect 6947 4050 6981 4084
rect 7016 4050 7050 4084
rect 7085 4050 7119 4084
rect 7154 4050 7188 4084
rect 7223 4050 7257 4084
rect 7292 4050 7326 4084
rect 7361 4050 7395 4084
rect 7430 4050 7464 4084
rect 7499 4050 7533 4084
rect 7568 4050 7602 4084
rect 7637 4050 7671 4084
rect 7706 4050 7740 4084
rect 7775 4050 7809 4084
rect 7844 4050 7878 4084
rect 7913 4050 7947 4084
rect 7982 4050 8016 4084
rect 8051 4050 8085 4084
rect 8120 4050 8154 4084
rect 8189 4050 8223 4084
rect 8258 4050 8292 4084
rect 4102 4005 4136 4039
rect 4172 4005 4206 4039
rect 4242 4005 4276 4039
rect 4312 4005 4346 4039
rect 4382 4005 4416 4039
rect 4452 4005 4486 4039
rect 4522 4005 4556 4039
rect 4592 4005 4626 4039
rect 4662 4005 4696 4039
rect 4974 3979 5008 4013
rect 5043 3979 5077 4013
rect 5112 3979 5146 4013
rect 5181 3979 5215 4013
rect 5250 3979 5284 4013
rect 5319 3979 5353 4013
rect 5388 3979 5422 4013
rect 5457 3979 5491 4013
rect 5526 3979 5560 4013
rect 5595 3979 5629 4013
rect 5664 3979 5698 4013
rect 5733 3979 5767 4013
rect 5802 3979 5836 4013
rect 5871 3979 5905 4013
rect 5940 3979 5974 4013
rect 6009 3979 6043 4013
rect 6078 3979 6112 4013
rect 6147 3979 6181 4013
rect 6216 3979 6250 4013
rect 6285 3979 6319 4013
rect 6354 3979 6388 4013
rect 6423 3979 6457 4013
rect 6492 3979 6526 4013
rect 6561 3979 6595 4013
rect 6630 3979 6664 4013
rect 6699 3979 6733 4013
rect 6768 3979 6802 4013
rect 6837 3979 6871 4013
rect 6906 3979 6940 4013
rect 6975 3979 7009 4013
rect 7044 3979 7078 4013
rect 7113 3979 7147 4013
rect 7182 3979 7216 4013
rect 7251 3979 7285 4013
rect 7320 3979 7354 4013
rect 7389 3979 7423 4013
rect 7458 3979 7492 4013
rect 7527 3979 7561 4013
rect 7596 3979 7630 4013
rect 7665 3979 7699 4013
rect 7734 3979 7768 4013
rect 7803 3979 7837 4013
rect 7872 3979 7906 4013
rect 7941 3979 7975 4013
rect 8010 3979 8044 4013
rect 8079 3979 8113 4013
rect 8148 3979 8182 4013
rect 8217 3979 8251 4013
rect 8286 3979 8320 4013
rect 8355 3979 8389 4013
rect 8424 3979 8458 4013
rect 8493 3979 8527 4013
rect 8562 3979 8596 4013
rect 8631 3979 8665 4013
rect 8700 3979 8734 4013
rect 8769 3979 8803 4013
rect 8838 3979 8872 4013
rect 8907 3979 8941 4013
rect 8976 3979 9010 4013
rect 9045 3979 9079 4013
rect 9114 3979 9148 4013
rect 9183 3979 9217 4013
rect 9252 3979 9286 4013
rect 9320 3979 9354 4013
rect 9388 3979 9422 4013
rect 4102 3935 4136 3969
rect 4172 3935 4206 3969
rect 4242 3935 4276 3969
rect 4312 3935 4346 3969
rect 4382 3935 4416 3969
rect 4452 3935 4486 3969
rect 4522 3935 4556 3969
rect 4592 3935 4626 3969
rect 4662 3935 4696 3969
rect 4974 3903 5008 3937
rect 5043 3903 5077 3937
rect 5112 3903 5146 3937
rect 5181 3903 5215 3937
rect 5250 3903 5284 3937
rect 5319 3903 5353 3937
rect 5388 3903 5422 3937
rect 5457 3903 5491 3937
rect 5526 3903 5560 3937
rect 5595 3903 5629 3937
rect 5664 3903 5698 3937
rect 5733 3903 5767 3937
rect 5802 3903 5836 3937
rect 5871 3903 5905 3937
rect 5940 3903 5974 3937
rect 6009 3903 6043 3937
rect 6078 3903 6112 3937
rect 6147 3903 6181 3937
rect 6216 3903 6250 3937
rect 6285 3903 6319 3937
rect 6354 3903 6388 3937
rect 6423 3903 6457 3937
rect 6492 3903 6526 3937
rect 6561 3903 6595 3937
rect 6630 3903 6664 3937
rect 6699 3903 6733 3937
rect 6768 3903 6802 3937
rect 6837 3903 6871 3937
rect 6906 3903 6940 3937
rect 6975 3903 7009 3937
rect 7044 3903 7078 3937
rect 7113 3903 7147 3937
rect 7182 3903 7216 3937
rect 7251 3903 7285 3937
rect 7320 3903 7354 3937
rect 7389 3903 7423 3937
rect 7458 3903 7492 3937
rect 7527 3903 7561 3937
rect 7596 3903 7630 3937
rect 7665 3903 7699 3937
rect 7734 3903 7768 3937
rect 7803 3903 7837 3937
rect 7872 3903 7906 3937
rect 7941 3903 7975 3937
rect 8010 3903 8044 3937
rect 8079 3903 8113 3937
rect 8148 3903 8182 3937
rect 8217 3903 8251 3937
rect 8286 3903 8320 3937
rect 8355 3903 8389 3937
rect 8424 3903 8458 3937
rect 8493 3903 8527 3937
rect 8562 3903 8596 3937
rect 8631 3903 8665 3937
rect 8700 3903 8734 3937
rect 8769 3903 8803 3937
rect 8838 3903 8872 3937
rect 8907 3903 8941 3937
rect 8976 3903 9010 3937
rect 9045 3903 9079 3937
rect 9114 3903 9148 3937
rect 9183 3903 9217 3937
rect 9252 3903 9286 3937
rect 9320 3903 9354 3937
rect 9388 3903 9422 3937
rect 3875 2167 4929 3901
rect 4974 3827 5008 3861
rect 5043 3827 5077 3861
rect 5112 3827 5146 3861
rect 5181 3827 5215 3861
rect 5250 3827 5284 3861
rect 5319 3827 5353 3861
rect 5388 3827 5422 3861
rect 5457 3827 5491 3861
rect 5526 3827 5560 3861
rect 5595 3827 5629 3861
rect 5664 3827 5698 3861
rect 5733 3827 5767 3861
rect 5802 3827 5836 3861
rect 5871 3827 5905 3861
rect 5940 3827 5974 3861
rect 6009 3827 6043 3861
rect 6078 3827 6112 3861
rect 6147 3827 6181 3861
rect 6216 3827 6250 3861
rect 6285 3827 6319 3861
rect 6354 3827 6388 3861
rect 6423 3827 6457 3861
rect 6492 3827 6526 3861
rect 6561 3827 6595 3861
rect 6630 3827 6664 3861
rect 6699 3827 6733 3861
rect 6768 3827 6802 3861
rect 6837 3827 6871 3861
rect 6906 3827 6940 3861
rect 6975 3827 7009 3861
rect 7044 3827 7078 3861
rect 7113 3827 7147 3861
rect 7182 3827 7216 3861
rect 7251 3827 7285 3861
rect 7320 3827 7354 3861
rect 7389 3827 7423 3861
rect 7458 3827 7492 3861
rect 7527 3827 7561 3861
rect 7596 3827 7630 3861
rect 7665 3827 7699 3861
rect 7734 3827 7768 3861
rect 7803 3827 7837 3861
rect 7872 3827 7906 3861
rect 7941 3827 7975 3861
rect 8010 3827 8044 3861
rect 8079 3827 8113 3861
rect 8148 3827 8182 3861
rect 8217 3827 8251 3861
rect 8286 3827 8320 3861
rect 8355 3827 8389 3861
rect 8424 3827 8458 3861
rect 8493 3827 8527 3861
rect 8562 3827 8596 3861
rect 8631 3827 8665 3861
rect 8700 3827 8734 3861
rect 8769 3827 8803 3861
rect 8838 3827 8872 3861
rect 8907 3827 8941 3861
rect 8976 3827 9010 3861
rect 9045 3827 9079 3861
rect 9114 3827 9148 3861
rect 9183 3827 9217 3861
rect 9252 3827 9286 3861
rect 9320 3827 9354 3861
rect 9388 3827 9422 3861
rect 4974 3751 5008 3785
rect 5043 3751 5077 3785
rect 5112 3751 5146 3785
rect 5181 3751 5215 3785
rect 5250 3751 5284 3785
rect 5319 3751 5353 3785
rect 5388 3751 5422 3785
rect 5457 3751 5491 3785
rect 5526 3751 5560 3785
rect 5595 3751 5629 3785
rect 5664 3751 5698 3785
rect 5733 3751 5767 3785
rect 5802 3751 5836 3785
rect 5871 3751 5905 3785
rect 5940 3751 5974 3785
rect 6009 3751 6043 3785
rect 6078 3751 6112 3785
rect 6147 3751 6181 3785
rect 6216 3751 6250 3785
rect 6285 3751 6319 3785
rect 6354 3751 6388 3785
rect 6423 3751 6457 3785
rect 6492 3751 6526 3785
rect 6561 3751 6595 3785
rect 6630 3751 6664 3785
rect 6699 3751 6733 3785
rect 6768 3751 6802 3785
rect 6837 3751 6871 3785
rect 6906 3751 6940 3785
rect 6975 3751 7009 3785
rect 7044 3751 7078 3785
rect 7113 3751 7147 3785
rect 7182 3751 7216 3785
rect 7251 3751 7285 3785
rect 7320 3751 7354 3785
rect 7389 3751 7423 3785
rect 7458 3751 7492 3785
rect 7527 3751 7561 3785
rect 7596 3751 7630 3785
rect 7665 3751 7699 3785
rect 7734 3751 7768 3785
rect 7803 3751 7837 3785
rect 7872 3751 7906 3785
rect 7941 3751 7975 3785
rect 8010 3751 8044 3785
rect 8079 3751 8113 3785
rect 8148 3751 8182 3785
rect 8217 3751 8251 3785
rect 8286 3751 8320 3785
rect 8355 3751 8389 3785
rect 8424 3751 8458 3785
rect 8493 3751 8527 3785
rect 8562 3751 8596 3785
rect 8631 3751 8665 3785
rect 8700 3751 8734 3785
rect 8769 3751 8803 3785
rect 8838 3751 8872 3785
rect 8907 3751 8941 3785
rect 8976 3751 9010 3785
rect 9045 3751 9079 3785
rect 9114 3751 9148 3785
rect 9183 3751 9217 3785
rect 9252 3751 9286 3785
rect 9320 3751 9354 3785
rect 9388 3751 9422 3785
rect 4974 3675 5008 3709
rect 5043 3675 5077 3709
rect 5112 3675 5146 3709
rect 5181 3675 5215 3709
rect 5250 3675 5284 3709
rect 5319 3675 5353 3709
rect 5388 3675 5422 3709
rect 5457 3675 5491 3709
rect 5526 3675 5560 3709
rect 5595 3675 5629 3709
rect 5664 3675 5698 3709
rect 5733 3675 5767 3709
rect 5802 3675 5836 3709
rect 5871 3675 5905 3709
rect 5940 3675 5974 3709
rect 6009 3675 6043 3709
rect 6078 3675 6112 3709
rect 6147 3675 6181 3709
rect 6216 3675 6250 3709
rect 6285 3675 6319 3709
rect 6354 3675 6388 3709
rect 6423 3675 6457 3709
rect 6492 3675 6526 3709
rect 6561 3675 6595 3709
rect 6630 3675 6664 3709
rect 6699 3675 6733 3709
rect 6768 3675 6802 3709
rect 6837 3675 6871 3709
rect 6906 3675 6940 3709
rect 6975 3675 7009 3709
rect 7044 3675 7078 3709
rect 7113 3675 7147 3709
rect 7182 3675 7216 3709
rect 7251 3675 7285 3709
rect 7320 3675 7354 3709
rect 7389 3675 7423 3709
rect 7458 3675 7492 3709
rect 7527 3675 7561 3709
rect 7596 3675 7630 3709
rect 7665 3675 7699 3709
rect 7734 3675 7768 3709
rect 7803 3675 7837 3709
rect 7872 3675 7906 3709
rect 7941 3675 7975 3709
rect 8010 3675 8044 3709
rect 8079 3675 8113 3709
rect 8148 3675 8182 3709
rect 8217 3675 8251 3709
rect 8286 3675 8320 3709
rect 8355 3675 8389 3709
rect 8424 3675 8458 3709
rect 8493 3675 8527 3709
rect 8562 3675 8596 3709
rect 8631 3675 8665 3709
rect 8700 3675 8734 3709
rect 8769 3675 8803 3709
rect 8838 3675 8872 3709
rect 8907 3675 8941 3709
rect 8976 3675 9010 3709
rect 9045 3675 9079 3709
rect 9114 3675 9148 3709
rect 9183 3675 9217 3709
rect 9252 3675 9286 3709
rect 9320 3675 9354 3709
rect 9388 3675 9422 3709
rect 13507 4139 13541 4173
rect 13575 4139 13609 4173
rect 13643 4139 13677 4173
rect 13711 4139 13745 4173
rect 13779 4139 13813 4173
rect 13847 4139 13881 4173
rect 13915 4139 13949 4173
rect 13983 4139 14017 4173
rect 14051 4139 14085 4173
rect 14119 4139 14153 4173
rect 14187 4139 14221 4173
rect 14255 4139 14289 4173
rect 14323 4139 14357 4173
rect 14391 4139 14425 4173
rect 14459 4139 14493 4173
rect 14527 4139 14561 4173
rect 13439 4016 13473 4050
rect 13439 3948 13473 3982
rect 13439 3880 13473 3914
rect 13439 3812 13473 3846
rect 13439 3744 13473 3778
rect 13439 3676 13473 3710
rect 13439 3608 13473 3642
rect 13439 3540 13473 3574
rect 13439 3472 13473 3506
rect 13439 3404 13473 3438
rect 13439 3336 13473 3370
rect 13439 3268 13473 3302
rect 11543 3009 11577 3043
rect 11612 3009 11646 3043
rect 11681 3009 11715 3043
rect 11750 3009 11784 3043
rect 11819 3009 11853 3043
rect 11888 3009 11922 3043
rect 11957 3009 11991 3043
rect 12025 3009 12059 3043
rect 12093 3009 12127 3043
rect 12161 3009 12195 3043
rect 12229 3009 12263 3043
rect 12297 3009 12331 3043
rect 11543 2921 11577 2955
rect 11612 2921 11646 2955
rect 11681 2921 11715 2955
rect 11750 2921 11784 2955
rect 11819 2921 11853 2955
rect 11888 2921 11922 2955
rect 11957 2921 11991 2955
rect 12025 2921 12059 2955
rect 12093 2921 12127 2955
rect 12161 2921 12195 2955
rect 12229 2921 12263 2955
rect 12297 2921 12331 2955
rect 11543 2833 11577 2867
rect 11612 2833 11646 2867
rect 11681 2833 11715 2867
rect 11750 2833 11784 2867
rect 11819 2833 11853 2867
rect 11888 2833 11922 2867
rect 11957 2833 11991 2867
rect 12025 2833 12059 2867
rect 12093 2833 12127 2867
rect 12161 2833 12195 2867
rect 12229 2833 12263 2867
rect 12297 2833 12331 2867
rect 11543 2745 11577 2779
rect 11612 2745 11646 2779
rect 11681 2745 11715 2779
rect 11750 2745 11784 2779
rect 11819 2745 11853 2779
rect 11888 2745 11922 2779
rect 11957 2745 11991 2779
rect 12025 2745 12059 2779
rect 12093 2745 12127 2779
rect 12161 2745 12195 2779
rect 12229 2745 12263 2779
rect 12297 2745 12331 2779
rect 11841 2676 11875 2710
rect 11911 2676 11945 2710
rect 11981 2676 12015 2710
rect 12051 2676 12085 2710
rect 12121 2676 12155 2710
rect 12191 2676 12225 2710
rect 12261 2676 12295 2710
rect 12331 2676 12365 2710
rect 11841 2603 11875 2637
rect 11911 2603 11945 2637
rect 11981 2603 12015 2637
rect 12051 2603 12085 2637
rect 12121 2603 12155 2637
rect 12191 2603 12225 2637
rect 12261 2603 12295 2637
rect 12331 2603 12365 2637
rect 11841 2530 11875 2564
rect 11911 2530 11945 2564
rect 11981 2530 12015 2564
rect 12051 2530 12085 2564
rect 12121 2530 12155 2564
rect 12191 2530 12225 2564
rect 12261 2530 12295 2564
rect 12331 2530 12365 2564
rect 11841 2457 11875 2491
rect 11911 2457 11945 2491
rect 11981 2457 12015 2491
rect 12051 2457 12085 2491
rect 12121 2457 12155 2491
rect 12191 2457 12225 2491
rect 12261 2457 12295 2491
rect 12331 2457 12365 2491
rect 11841 2384 11875 2418
rect 11911 2384 11945 2418
rect 11981 2384 12015 2418
rect 12051 2384 12085 2418
rect 12121 2384 12155 2418
rect 12191 2384 12225 2418
rect 12261 2384 12295 2418
rect 12331 2384 12365 2418
rect 11841 2310 11875 2344
rect 11911 2310 11945 2344
rect 11981 2310 12015 2344
rect 12051 2310 12085 2344
rect 12121 2310 12155 2344
rect 12191 2310 12225 2344
rect 12261 2310 12295 2344
rect 12331 2310 12365 2344
rect 11841 2236 11875 2270
rect 11911 2236 11945 2270
rect 11981 2236 12015 2270
rect 12051 2236 12085 2270
rect 12121 2236 12155 2270
rect 12191 2236 12225 2270
rect 12261 2236 12295 2270
rect 12331 2236 12365 2270
rect 3875 2098 3909 2132
rect 3943 2098 3977 2132
rect 4011 2098 4045 2132
rect 4079 2098 4113 2132
rect 4147 2098 4181 2132
rect 4215 2098 4249 2132
rect 4283 2098 4317 2132
rect 4351 2098 4385 2132
rect 4419 2098 4453 2132
rect 4487 2098 4521 2132
rect 4555 2098 4589 2132
rect 4623 2098 4657 2132
rect 4691 2098 4725 2132
rect 4759 2098 4793 2132
rect 4827 2098 4861 2132
rect 4895 2098 4929 2132
rect 3875 2029 3909 2063
rect 3943 2029 3977 2063
rect 4011 2029 4045 2063
rect 4079 2029 4113 2063
rect 4147 2029 4181 2063
rect 4215 2029 4249 2063
rect 4283 2029 4317 2063
rect 4351 2029 4385 2063
rect 4419 2029 4453 2063
rect 4487 2029 4521 2063
rect 4555 2029 4589 2063
rect 4623 2029 4657 2063
rect 4691 2029 4725 2063
rect 4759 2029 4793 2063
rect 4827 2029 4861 2063
rect 4895 2029 4929 2063
rect 3875 1960 3909 1994
rect 3943 1960 3977 1994
rect 4011 1960 4045 1994
rect 4079 1960 4113 1994
rect 4147 1960 4181 1994
rect 4215 1960 4249 1994
rect 4283 1960 4317 1994
rect 4351 1960 4385 1994
rect 4419 1960 4453 1994
rect 4487 1960 4521 1994
rect 4555 1960 4589 1994
rect 4623 1960 4657 1994
rect 4691 1960 4725 1994
rect 4759 1960 4793 1994
rect 4827 1960 4861 1994
rect 4895 1960 4929 1994
rect 3875 1891 3909 1925
rect 3943 1891 3977 1925
rect 4011 1891 4045 1925
rect 4079 1891 4113 1925
rect 4147 1891 4181 1925
rect 4215 1891 4249 1925
rect 4283 1891 4317 1925
rect 4351 1891 4385 1925
rect 4419 1891 4453 1925
rect 4487 1891 4521 1925
rect 4555 1891 4589 1925
rect 4623 1891 4657 1925
rect 4691 1891 4725 1925
rect 4759 1891 4793 1925
rect 4827 1891 4861 1925
rect 4895 1891 4929 1925
rect 3875 1822 3909 1856
rect 3943 1822 3977 1856
rect 4011 1822 4045 1856
rect 4079 1822 4113 1856
rect 4147 1822 4181 1856
rect 4215 1822 4249 1856
rect 4283 1822 4317 1856
rect 4351 1822 4385 1856
rect 4419 1822 4453 1856
rect 4487 1822 4521 1856
rect 4555 1822 4589 1856
rect 4623 1822 4657 1856
rect 4691 1822 4725 1856
rect 4759 1822 4793 1856
rect 4827 1822 4861 1856
rect 4895 1822 4929 1856
rect 3875 1753 3909 1787
rect 3943 1753 3977 1787
rect 4011 1753 4045 1787
rect 4079 1753 4113 1787
rect 4147 1753 4181 1787
rect 4215 1753 4249 1787
rect 4283 1753 4317 1787
rect 4351 1753 4385 1787
rect 4419 1753 4453 1787
rect 4487 1753 4521 1787
rect 4555 1753 4589 1787
rect 4623 1753 4657 1787
rect 4691 1753 4725 1787
rect 4759 1753 4793 1787
rect 4827 1753 4861 1787
rect 4895 1753 4929 1787
rect 3875 1684 3909 1718
rect 3943 1684 3977 1718
rect 4011 1684 4045 1718
rect 4079 1684 4113 1718
rect 4147 1684 4181 1718
rect 4215 1684 4249 1718
rect 4283 1684 4317 1718
rect 4351 1684 4385 1718
rect 4419 1684 4453 1718
rect 4487 1684 4521 1718
rect 4555 1684 4589 1718
rect 4623 1684 4657 1718
rect 4691 1684 4725 1718
rect 4759 1684 4793 1718
rect 4827 1684 4861 1718
rect 4895 1684 4929 1718
rect 3875 1615 3909 1649
rect 3943 1615 3977 1649
rect 4011 1615 4045 1649
rect 4079 1615 4113 1649
rect 4147 1615 4181 1649
rect 4215 1615 4249 1649
rect 4283 1615 4317 1649
rect 4351 1615 4385 1649
rect 4419 1615 4453 1649
rect 4487 1615 4521 1649
rect 4555 1615 4589 1649
rect 4623 1615 4657 1649
rect 4691 1615 4725 1649
rect 4759 1615 4793 1649
rect 4827 1615 4861 1649
rect 4895 1615 4929 1649
rect 3875 1546 3909 1580
rect 3943 1546 3977 1580
rect 4011 1546 4045 1580
rect 4079 1546 4113 1580
rect 4147 1546 4181 1580
rect 4215 1546 4249 1580
rect 4283 1546 4317 1580
rect 4351 1546 4385 1580
rect 4419 1546 4453 1580
rect 4487 1546 4521 1580
rect 4555 1546 4589 1580
rect 4623 1546 4657 1580
rect 4691 1546 4725 1580
rect 4759 1546 4793 1580
rect 4827 1546 4861 1580
rect 4895 1546 4929 1580
rect 3875 1477 3909 1511
rect 3943 1477 3977 1511
rect 4011 1477 4045 1511
rect 4079 1477 4113 1511
rect 4147 1477 4181 1511
rect 4215 1477 4249 1511
rect 4283 1477 4317 1511
rect 4351 1477 4385 1511
rect 4419 1477 4453 1511
rect 4487 1477 4521 1511
rect 4555 1477 4589 1511
rect 4623 1477 4657 1511
rect 4691 1477 4725 1511
rect 4759 1477 4793 1511
rect 4827 1477 4861 1511
rect 4895 1477 4929 1511
rect 3875 1408 3909 1442
rect 3943 1408 3977 1442
rect 4011 1408 4045 1442
rect 4079 1408 4113 1442
rect 4147 1408 4181 1442
rect 4215 1408 4249 1442
rect 4283 1408 4317 1442
rect 4351 1408 4385 1442
rect 4419 1408 4453 1442
rect 4487 1408 4521 1442
rect 4555 1408 4589 1442
rect 4623 1408 4657 1442
rect 4691 1408 4725 1442
rect 4759 1408 4793 1442
rect 4827 1408 4861 1442
rect 4895 1408 4929 1442
rect 3875 1339 3909 1373
rect 3943 1339 3977 1373
rect 4011 1339 4045 1373
rect 4079 1339 4113 1373
rect 4147 1339 4181 1373
rect 4215 1339 4249 1373
rect 4283 1339 4317 1373
rect 4351 1339 4385 1373
rect 4419 1339 4453 1373
rect 4487 1339 4521 1373
rect 4555 1339 4589 1373
rect 4623 1339 4657 1373
rect 4691 1339 4725 1373
rect 4759 1339 4793 1373
rect 4827 1339 4861 1373
rect 4895 1339 4929 1373
rect 3875 1270 3909 1304
rect 3943 1270 3977 1304
rect 4011 1270 4045 1304
rect 4079 1270 4113 1304
rect 4147 1270 4181 1304
rect 4215 1270 4249 1304
rect 4283 1270 4317 1304
rect 4351 1270 4385 1304
rect 4419 1270 4453 1304
rect 4487 1270 4521 1304
rect 4555 1270 4589 1304
rect 4623 1270 4657 1304
rect 4691 1270 4725 1304
rect 4759 1270 4793 1304
rect 4827 1270 4861 1304
rect 4895 1270 4929 1304
rect 3875 1201 3909 1235
rect 3943 1201 3977 1235
rect 4011 1201 4045 1235
rect 4079 1201 4113 1235
rect 4147 1201 4181 1235
rect 4215 1201 4249 1235
rect 4283 1201 4317 1235
rect 4351 1201 4385 1235
rect 4419 1201 4453 1235
rect 4487 1201 4521 1235
rect 4555 1201 4589 1235
rect 4623 1201 4657 1235
rect 4691 1201 4725 1235
rect 4759 1201 4793 1235
rect 4827 1201 4861 1235
rect 4895 1201 4929 1235
rect 3875 1132 3909 1166
rect 3943 1132 3977 1166
rect 4011 1132 4045 1166
rect 4079 1132 4113 1166
rect 4147 1132 4181 1166
rect 4215 1132 4249 1166
rect 4283 1132 4317 1166
rect 4351 1132 4385 1166
rect 4419 1132 4453 1166
rect 4487 1132 4521 1166
rect 4555 1132 4589 1166
rect 4623 1132 4657 1166
rect 4691 1132 4725 1166
rect 4759 1132 4793 1166
rect 4827 1132 4861 1166
rect 4895 1132 4929 1166
rect 3875 1063 3909 1097
rect 3943 1063 3977 1097
rect 4011 1063 4045 1097
rect 4079 1063 4113 1097
rect 4147 1063 4181 1097
rect 4215 1063 4249 1097
rect 4283 1063 4317 1097
rect 4351 1063 4385 1097
rect 4419 1063 4453 1097
rect 4487 1063 4521 1097
rect 4555 1063 4589 1097
rect 4623 1063 4657 1097
rect 4691 1063 4725 1097
rect 4759 1063 4793 1097
rect 4827 1063 4861 1097
rect 4895 1063 4929 1097
rect 3875 994 3909 1028
rect 3943 994 3977 1028
rect 4011 994 4045 1028
rect 4079 994 4113 1028
rect 4147 994 4181 1028
rect 4215 994 4249 1028
rect 4283 994 4317 1028
rect 4351 994 4385 1028
rect 4419 994 4453 1028
rect 4487 994 4521 1028
rect 4555 994 4589 1028
rect 4623 994 4657 1028
rect 4691 994 4725 1028
rect 4759 994 4793 1028
rect 4827 994 4861 1028
rect 4895 994 4929 1028
rect 3875 925 3909 959
rect 3943 925 3977 959
rect 4011 925 4045 959
rect 4079 925 4113 959
rect 4147 925 4181 959
rect 4215 925 4249 959
rect 4283 925 4317 959
rect 4351 925 4385 959
rect 4419 925 4453 959
rect 4487 925 4521 959
rect 4555 925 4589 959
rect 4623 925 4657 959
rect 4691 925 4725 959
rect 4759 925 4793 959
rect 4827 925 4861 959
rect 4895 925 4929 959
rect 3875 856 3909 890
rect 3943 856 3977 890
rect 4011 856 4045 890
rect 4079 856 4113 890
rect 4147 856 4181 890
rect 4215 856 4249 890
rect 4283 856 4317 890
rect 4351 856 4385 890
rect 4419 856 4453 890
rect 4487 856 4521 890
rect 4555 856 4589 890
rect 4623 856 4657 890
rect 4691 856 4725 890
rect 4759 856 4793 890
rect 4827 856 4861 890
rect 4895 856 4929 890
rect 5299 1024 5333 1058
rect 5369 1024 5403 1058
rect 5438 1024 5472 1058
rect 5507 1024 5541 1058
rect 5576 1024 5610 1058
rect 5645 1024 5679 1058
rect 5714 1024 5748 1058
rect 5783 1024 5817 1058
rect 5852 1024 5886 1058
rect 5921 1024 5955 1058
rect 5990 1024 6024 1058
rect 6059 1024 6093 1058
rect 6128 1024 6162 1058
rect 6197 1024 6231 1058
rect 6266 1024 6300 1058
rect 6335 1024 6369 1058
rect 6404 1024 6438 1058
rect 6473 1024 6507 1058
rect 6542 1024 6576 1058
rect 6611 1024 6645 1058
rect 6680 1024 6714 1058
rect 6749 1024 6783 1058
rect 6818 1024 6852 1058
rect 6887 1024 6921 1058
rect 6956 1024 6990 1058
rect 7025 1024 7059 1058
rect 7094 1024 7128 1058
rect 7163 1024 7197 1058
rect 7232 1024 7266 1058
rect 7301 1024 7335 1058
rect 7370 1024 7404 1058
rect 7439 1024 7473 1058
rect 7508 1024 7542 1058
rect 7577 1024 7611 1058
rect 7646 1024 7680 1058
rect 7715 1024 7749 1058
rect 7784 1024 7818 1058
rect 7853 1024 7887 1058
rect 7922 1024 7956 1058
rect 7991 1024 8025 1058
rect 8060 1024 8094 1058
rect 8129 1024 8163 1058
rect 8198 1024 8232 1058
rect 8267 1024 8301 1058
rect 8336 1024 8370 1058
rect 8405 1024 8439 1058
rect 8474 1024 8508 1058
rect 8543 1024 8577 1058
rect 8612 1024 8646 1058
rect 5299 952 5333 986
rect 5369 952 5403 986
rect 5438 952 5472 986
rect 5507 952 5541 986
rect 5576 952 5610 986
rect 5645 952 5679 986
rect 5714 952 5748 986
rect 5783 952 5817 986
rect 5852 952 5886 986
rect 5921 952 5955 986
rect 5990 952 6024 986
rect 6059 952 6093 986
rect 6128 952 6162 986
rect 6197 952 6231 986
rect 6266 952 6300 986
rect 6335 952 6369 986
rect 6404 952 6438 986
rect 6473 952 6507 986
rect 6542 952 6576 986
rect 6611 952 6645 986
rect 6680 952 6714 986
rect 6749 952 6783 986
rect 6818 952 6852 986
rect 6887 952 6921 986
rect 6956 952 6990 986
rect 7025 952 7059 986
rect 7094 952 7128 986
rect 7163 952 7197 986
rect 7232 952 7266 986
rect 7301 952 7335 986
rect 7370 952 7404 986
rect 7439 952 7473 986
rect 7508 952 7542 986
rect 7577 952 7611 986
rect 7646 952 7680 986
rect 7715 952 7749 986
rect 7784 952 7818 986
rect 7853 952 7887 986
rect 7922 952 7956 986
rect 7991 952 8025 986
rect 8060 952 8094 986
rect 8129 952 8163 986
rect 8198 952 8232 986
rect 8267 952 8301 986
rect 8336 952 8370 986
rect 8405 952 8439 986
rect 8474 952 8508 986
rect 8543 952 8577 986
rect 8612 952 8646 986
rect 5299 880 5333 914
rect 5369 880 5403 914
rect 5438 880 5472 914
rect 5507 880 5541 914
rect 5576 880 5610 914
rect 5645 880 5679 914
rect 5714 880 5748 914
rect 5783 880 5817 914
rect 5852 880 5886 914
rect 5921 880 5955 914
rect 5990 880 6024 914
rect 6059 880 6093 914
rect 6128 880 6162 914
rect 6197 880 6231 914
rect 6266 880 6300 914
rect 6335 880 6369 914
rect 6404 880 6438 914
rect 6473 880 6507 914
rect 6542 880 6576 914
rect 6611 880 6645 914
rect 6680 880 6714 914
rect 6749 880 6783 914
rect 6818 880 6852 914
rect 6887 880 6921 914
rect 6956 880 6990 914
rect 7025 880 7059 914
rect 7094 880 7128 914
rect 7163 880 7197 914
rect 7232 880 7266 914
rect 7301 880 7335 914
rect 7370 880 7404 914
rect 7439 880 7473 914
rect 7508 880 7542 914
rect 7577 880 7611 914
rect 7646 880 7680 914
rect 7715 880 7749 914
rect 7784 880 7818 914
rect 7853 880 7887 914
rect 7922 880 7956 914
rect 7991 880 8025 914
rect 8060 880 8094 914
rect 8129 880 8163 914
rect 8198 880 8232 914
rect 8267 880 8301 914
rect 8336 880 8370 914
rect 8405 880 8439 914
rect 8474 880 8508 914
rect 8543 880 8577 914
rect 8612 880 8646 914
rect 3875 787 3909 821
rect 3943 787 3977 821
rect 4011 787 4045 821
rect 4079 787 4113 821
rect 4147 787 4181 821
rect 4215 787 4249 821
rect 4283 787 4317 821
rect 4351 787 4385 821
rect 4419 787 4453 821
rect 4487 787 4521 821
rect 4555 787 4589 821
rect 4623 787 4657 821
rect 4691 787 4725 821
rect 4759 787 4793 821
rect 4827 787 4861 821
rect 4895 787 4929 821
rect 3875 718 3909 752
rect 3943 718 3977 752
rect 4011 718 4045 752
rect 4079 718 4113 752
rect 4147 718 4181 752
rect 4215 718 4249 752
rect 4283 718 4317 752
rect 4351 718 4385 752
rect 4419 718 4453 752
rect 4487 718 4521 752
rect 4555 718 4589 752
rect 4623 718 4657 752
rect 4691 718 4725 752
rect 4759 718 4793 752
rect 4827 718 4861 752
rect 4895 718 4929 752
rect 3875 649 3909 683
rect 3943 649 3977 683
rect 4011 649 4045 683
rect 4079 649 4113 683
rect 4147 649 4181 683
rect 4215 649 4249 683
rect 4283 649 4317 683
rect 4351 649 4385 683
rect 4419 649 4453 683
rect 4487 649 4521 683
rect 4555 649 4589 683
rect 4623 649 4657 683
rect 4691 649 4725 683
rect 4759 649 4793 683
rect 4827 649 4861 683
rect 4895 649 4929 683
rect 3875 580 3909 614
rect 3943 580 3977 614
rect 4011 580 4045 614
rect 4079 580 4113 614
rect 4147 580 4181 614
rect 4215 580 4249 614
rect 4283 580 4317 614
rect 4351 580 4385 614
rect 4419 580 4453 614
rect 4487 580 4521 614
rect 4555 580 4589 614
rect 4623 580 4657 614
rect 4691 580 4725 614
rect 4759 580 4793 614
rect 4827 580 4861 614
rect 4895 580 4929 614
rect 3875 511 3909 545
rect 3943 511 3977 545
rect 4011 511 4045 545
rect 4079 511 4113 545
rect 4147 511 4181 545
rect 4215 511 4249 545
rect 4283 511 4317 545
rect 4351 511 4385 545
rect 4419 511 4453 545
rect 4487 511 4521 545
rect 4555 511 4589 545
rect 4623 511 4657 545
rect 4691 511 4725 545
rect 4759 511 4793 545
rect 4827 511 4861 545
rect 4895 511 4929 545
rect 3875 442 3909 476
rect 3943 442 3977 476
rect 4011 442 4045 476
rect 4079 442 4113 476
rect 4147 442 4181 476
rect 4215 442 4249 476
rect 4283 442 4317 476
rect 4351 442 4385 476
rect 4419 442 4453 476
rect 4487 442 4521 476
rect 4555 442 4589 476
rect 4623 442 4657 476
rect 4691 442 4725 476
rect 4759 442 4793 476
rect 4827 442 4861 476
rect 4895 442 4929 476
rect 3875 373 3909 407
rect 3943 373 3977 407
rect 4011 373 4045 407
rect 4079 373 4113 407
rect 4147 373 4181 407
rect 4215 373 4249 407
rect 4283 373 4317 407
rect 4351 373 4385 407
rect 4419 373 4453 407
rect 4487 373 4521 407
rect 4555 373 4589 407
rect 4623 373 4657 407
rect 4691 373 4725 407
rect 4759 373 4793 407
rect 4827 373 4861 407
rect 4895 373 4929 407
rect 3875 304 3909 338
rect 3943 304 3977 338
rect 4011 304 4045 338
rect 4079 304 4113 338
rect 4147 304 4181 338
rect 4215 304 4249 338
rect 4283 304 4317 338
rect 4351 304 4385 338
rect 4419 304 4453 338
rect 4487 304 4521 338
rect 4555 304 4589 338
rect 4623 304 4657 338
rect 4691 304 4725 338
rect 4759 304 4793 338
rect 4827 304 4861 338
rect 4895 304 4929 338
rect 3875 235 3909 269
rect 3943 235 3977 269
rect 4011 235 4045 269
rect 4079 235 4113 269
rect 4147 235 4181 269
rect 4215 235 4249 269
rect 4283 235 4317 269
rect 4351 235 4385 269
rect 4419 235 4453 269
rect 4487 235 4521 269
rect 4555 235 4589 269
rect 4623 235 4657 269
rect 4691 235 4725 269
rect 4759 235 4793 269
rect 4827 235 4861 269
rect 4895 235 4929 269
rect 3875 166 3909 200
rect 3943 166 3977 200
rect 4011 166 4045 200
rect 4079 166 4113 200
rect 4147 166 4181 200
rect 4215 166 4249 200
rect 4283 166 4317 200
rect 4351 166 4385 200
rect 4419 166 4453 200
rect 4487 166 4521 200
rect 4555 166 4589 200
rect 4623 166 4657 200
rect 4691 166 4725 200
rect 4759 166 4793 200
rect 4827 166 4861 200
rect 4895 166 4929 200
rect 3875 97 3909 131
rect 3943 97 3977 131
rect 4011 97 4045 131
rect 4079 97 4113 131
rect 4147 97 4181 131
rect 4215 97 4249 131
rect 4283 97 4317 131
rect 4351 97 4385 131
rect 4419 97 4453 131
rect 4487 97 4521 131
rect 4555 97 4589 131
rect 4623 97 4657 131
rect 4691 97 4725 131
rect 4759 97 4793 131
rect 4827 97 4861 131
rect 4895 97 4929 131
rect 3875 28 3909 62
rect 3943 28 3977 62
rect 4011 28 4045 62
rect 4079 28 4113 62
rect 4147 28 4181 62
rect 4215 28 4249 62
rect 4283 28 4317 62
rect 4351 28 4385 62
rect 4419 28 4453 62
rect 4487 28 4521 62
rect 4555 28 4589 62
rect 4623 28 4657 62
rect 4691 28 4725 62
rect 4759 28 4793 62
rect 4827 28 4861 62
rect 4895 28 4929 62
rect 11314 805 11348 839
rect 11385 805 11419 839
rect 11456 805 11490 839
rect 11527 805 11561 839
rect 11598 805 11632 839
rect 11669 805 11703 839
rect 11740 805 11774 839
rect 11811 805 11845 839
rect 11882 805 11916 839
rect 11953 805 11987 839
rect 12024 805 12058 839
rect 12095 805 12129 839
rect 12166 805 12200 839
rect 12237 805 12271 839
rect 12308 805 12342 839
rect 12379 805 12413 839
rect 12450 805 12484 839
rect 12521 805 12555 839
rect 12592 805 12626 839
rect 12663 805 12697 839
rect 12734 805 12768 839
rect 12804 805 12838 839
rect 11314 735 11348 769
rect 11385 735 11419 769
rect 11456 735 11490 769
rect 11527 735 11561 769
rect 11598 735 11632 769
rect 11669 735 11703 769
rect 11740 735 11774 769
rect 11811 735 11845 769
rect 11882 735 11916 769
rect 11953 735 11987 769
rect 12024 735 12058 769
rect 12095 735 12129 769
rect 12166 735 12200 769
rect 12237 735 12271 769
rect 12308 735 12342 769
rect 12379 735 12413 769
rect 12450 735 12484 769
rect 12521 735 12555 769
rect 12592 735 12626 769
rect 12663 735 12697 769
rect 12734 735 12768 769
rect 12804 735 12838 769
rect 11314 665 11348 699
rect 11385 665 11419 699
rect 11456 665 11490 699
rect 11527 665 11561 699
rect 11598 665 11632 699
rect 11669 665 11703 699
rect 11740 665 11774 699
rect 11811 665 11845 699
rect 11882 665 11916 699
rect 11953 665 11987 699
rect 12024 665 12058 699
rect 12095 665 12129 699
rect 12166 665 12200 699
rect 12237 665 12271 699
rect 12308 665 12342 699
rect 12379 665 12413 699
rect 12450 665 12484 699
rect 12521 665 12555 699
rect 12592 665 12626 699
rect 12663 665 12697 699
rect 12734 665 12768 699
rect 12804 665 12838 699
rect 11314 595 11348 629
rect 11385 595 11419 629
rect 11456 595 11490 629
rect 11527 595 11561 629
rect 11598 595 11632 629
rect 11669 595 11703 629
rect 11740 595 11774 629
rect 11811 595 11845 629
rect 11882 595 11916 629
rect 11953 595 11987 629
rect 12024 595 12058 629
rect 12095 595 12129 629
rect 12166 595 12200 629
rect 12237 595 12271 629
rect 12308 595 12342 629
rect 12379 595 12413 629
rect 12450 595 12484 629
rect 12521 595 12555 629
rect 12592 595 12626 629
rect 12663 595 12697 629
rect 12734 595 12768 629
rect 12804 595 12838 629
rect 11314 525 11348 559
rect 11385 525 11419 559
rect 11456 525 11490 559
rect 11527 525 11561 559
rect 11598 525 11632 559
rect 11669 525 11703 559
rect 11740 525 11774 559
rect 11811 525 11845 559
rect 11882 525 11916 559
rect 11953 525 11987 559
rect 12024 525 12058 559
rect 12095 525 12129 559
rect 12166 525 12200 559
rect 12237 525 12271 559
rect 12308 525 12342 559
rect 12379 525 12413 559
rect 12450 525 12484 559
rect 12521 525 12555 559
rect 12592 525 12626 559
rect 12663 525 12697 559
rect 12734 525 12768 559
rect 12804 525 12838 559
rect 11314 455 11348 489
rect 11385 455 11419 489
rect 11456 455 11490 489
rect 11527 455 11561 489
rect 11598 455 11632 489
rect 11669 455 11703 489
rect 11740 455 11774 489
rect 11811 455 11845 489
rect 11882 455 11916 489
rect 11953 455 11987 489
rect 12024 455 12058 489
rect 12095 455 12129 489
rect 12166 455 12200 489
rect 12237 455 12271 489
rect 12308 455 12342 489
rect 12379 455 12413 489
rect 12450 455 12484 489
rect 12521 455 12555 489
rect 12592 455 12626 489
rect 12663 455 12697 489
rect 12734 455 12768 489
rect 12804 455 12838 489
rect 11314 385 11348 419
rect 11385 385 11419 419
rect 11456 385 11490 419
rect 11527 385 11561 419
rect 11598 385 11632 419
rect 11669 385 11703 419
rect 11740 385 11774 419
rect 11811 385 11845 419
rect 11882 385 11916 419
rect 11953 385 11987 419
rect 12024 385 12058 419
rect 12095 385 12129 419
rect 12166 385 12200 419
rect 12237 385 12271 419
rect 12308 385 12342 419
rect 12379 385 12413 419
rect 12450 385 12484 419
rect 12521 385 12555 419
rect 12592 385 12626 419
rect 12663 385 12697 419
rect 12734 385 12768 419
rect 12804 385 12838 419
rect 11314 315 11348 349
rect 11385 315 11419 349
rect 11456 315 11490 349
rect 11527 315 11561 349
rect 11598 315 11632 349
rect 11669 315 11703 349
rect 11740 315 11774 349
rect 11811 315 11845 349
rect 11882 315 11916 349
rect 11953 315 11987 349
rect 12024 315 12058 349
rect 12095 315 12129 349
rect 12166 315 12200 349
rect 12237 315 12271 349
rect 12308 315 12342 349
rect 12379 315 12413 349
rect 12450 315 12484 349
rect 12521 315 12555 349
rect 12592 315 12626 349
rect 12663 315 12697 349
rect 12734 315 12768 349
rect 12804 315 12838 349
rect 11314 245 11348 279
rect 11385 245 11419 279
rect 11456 245 11490 279
rect 11527 245 11561 279
rect 11598 245 11632 279
rect 11669 245 11703 279
rect 11740 245 11774 279
rect 11811 245 11845 279
rect 11882 245 11916 279
rect 11953 245 11987 279
rect 12024 245 12058 279
rect 12095 245 12129 279
rect 12166 245 12200 279
rect 12237 245 12271 279
rect 12308 245 12342 279
rect 12379 245 12413 279
rect 12450 245 12484 279
rect 12521 245 12555 279
rect 12592 245 12626 279
rect 12663 245 12697 279
rect 12734 245 12768 279
rect 12804 245 12838 279
rect 11314 175 11348 209
rect 11385 175 11419 209
rect 11456 175 11490 209
rect 11527 175 11561 209
rect 11598 175 11632 209
rect 11669 175 11703 209
rect 11740 175 11774 209
rect 11811 175 11845 209
rect 11882 175 11916 209
rect 11953 175 11987 209
rect 12024 175 12058 209
rect 12095 175 12129 209
rect 12166 175 12200 209
rect 12237 175 12271 209
rect 12308 175 12342 209
rect 12379 175 12413 209
rect 12450 175 12484 209
rect 12521 175 12555 209
rect 12592 175 12626 209
rect 12663 175 12697 209
rect 12734 175 12768 209
rect 12804 175 12838 209
rect 11314 105 11348 139
rect 11385 105 11419 139
rect 11456 105 11490 139
rect 11527 105 11561 139
rect 11598 105 11632 139
rect 11669 105 11703 139
rect 11740 105 11774 139
rect 11811 105 11845 139
rect 11882 105 11916 139
rect 11953 105 11987 139
rect 12024 105 12058 139
rect 12095 105 12129 139
rect 12166 105 12200 139
rect 12237 105 12271 139
rect 12308 105 12342 139
rect 12379 105 12413 139
rect 12450 105 12484 139
rect 12521 105 12555 139
rect 12592 105 12626 139
rect 12663 105 12697 139
rect 12734 105 12768 139
rect 12804 105 12838 139
rect 11314 35 11348 69
rect 11385 35 11419 69
rect 11456 35 11490 69
rect 11527 35 11561 69
rect 11598 35 11632 69
rect 11669 35 11703 69
rect 11740 35 11774 69
rect 11811 35 11845 69
rect 11882 35 11916 69
rect 11953 35 11987 69
rect 12024 35 12058 69
rect 12095 35 12129 69
rect 12166 35 12200 69
rect 12237 35 12271 69
rect 12308 35 12342 69
rect 12379 35 12413 69
rect 12450 35 12484 69
rect 12521 35 12555 69
rect 12592 35 12626 69
rect 12663 35 12697 69
rect 12734 35 12768 69
rect 12804 35 12838 69
rect 11314 -35 11348 -1
rect 11385 -35 11419 -1
rect 11456 -35 11490 -1
rect 11527 -35 11561 -1
rect 11598 -35 11632 -1
rect 11669 -35 11703 -1
rect 11740 -35 11774 -1
rect 11811 -35 11845 -1
rect 11882 -35 11916 -1
rect 11953 -35 11987 -1
rect 12024 -35 12058 -1
rect 12095 -35 12129 -1
rect 12166 -35 12200 -1
rect 12237 -35 12271 -1
rect 12308 -35 12342 -1
rect 12379 -35 12413 -1
rect 12450 -35 12484 -1
rect 12521 -35 12555 -1
rect 12592 -35 12626 -1
rect 12663 -35 12697 -1
rect 12734 -35 12768 -1
rect 12804 -35 12838 -1
rect 13507 2658 13541 2692
rect 13575 2658 13609 2692
rect 13643 2658 13677 2692
rect 13711 2658 13745 2692
rect 13779 2658 13813 2692
rect 13847 2658 13881 2692
rect 13915 2658 13949 2692
rect 13983 2658 14017 2692
rect 14051 2658 14085 2692
rect 14119 2658 14153 2692
rect 14187 2658 14221 2692
rect 14255 2658 14289 2692
rect 14323 2658 14357 2692
rect 14391 2658 14425 2692
rect 14459 2658 14493 2692
rect 14527 2658 14561 2692
rect 14595 2658 14629 2692
rect 13439 2554 13473 2588
rect 14705 2590 14739 2624
rect 13439 2486 13473 2520
rect 13439 2418 13473 2452
rect 13439 2350 13473 2384
rect 13439 2282 13473 2316
rect 13439 2214 13473 2248
rect 13439 2146 13473 2180
rect 13439 2078 13473 2112
rect 13439 2010 13473 2044
rect 13439 1942 13473 1976
rect 13439 1874 13473 1908
rect 13439 1806 13473 1840
rect 13439 1738 13473 1772
rect 13439 1670 13473 1704
rect 13439 1528 13473 1562
rect 13439 1460 13473 1494
rect 13439 1392 13473 1426
rect 13439 1324 13473 1358
rect 13439 1256 13473 1290
rect 13439 1188 13473 1222
rect 13439 1120 13473 1154
rect 13439 1052 13473 1086
rect 13439 984 13473 1018
rect 13439 916 13473 950
rect 13439 848 13473 882
rect 13439 780 13473 814
rect 13439 712 13473 746
rect 13439 644 13473 678
rect 13439 576 13473 610
rect 13439 508 13473 542
rect 13439 440 13473 474
rect 13439 372 13473 406
rect 14705 2522 14739 2556
rect 14705 2454 14739 2488
rect 14705 2386 14739 2420
rect 14705 2318 14739 2352
rect 14705 2250 14739 2284
rect 14705 2182 14739 2216
rect 14705 2114 14739 2148
rect 14705 2046 14739 2080
rect 14705 1978 14739 2012
rect 14705 1910 14739 1944
rect 14705 1842 14739 1876
rect 14705 1774 14739 1808
rect 14705 1706 14739 1740
rect 14705 1638 14739 1672
rect 14705 1570 14739 1604
rect 14705 1502 14739 1536
rect 14705 1434 14739 1468
rect 14705 1366 14739 1400
rect 14705 1298 14739 1332
rect 14705 1230 14739 1264
rect 14705 1162 14739 1196
rect 14705 1094 14739 1128
rect 14705 1026 14739 1060
rect 14705 958 14739 992
rect 14705 890 14739 924
rect 14705 822 14739 856
rect 14705 754 14739 788
rect 14705 686 14739 720
rect 14705 618 14739 652
rect 14705 550 14739 584
rect 14705 482 14739 516
rect 14705 414 14739 448
rect 14705 346 14739 380
rect 13439 304 13473 338
rect 13549 236 13583 270
rect 13617 236 13651 270
rect 13685 236 13719 270
rect 13753 236 13787 270
rect 13821 236 13855 270
rect 13889 236 13923 270
rect 13957 236 13991 270
rect 14025 236 14059 270
rect 14093 236 14127 270
rect 14161 236 14195 270
rect 14229 236 14263 270
rect 14297 236 14331 270
rect 14365 236 14399 270
rect 14433 236 14467 270
rect 14501 236 14535 270
rect 14569 236 14603 270
rect 14637 236 14671 270
rect 8141 -96 8175 -62
rect 8211 -96 8245 -62
rect 8281 -96 8315 -62
rect 8351 -96 8385 -62
rect 8421 -96 8455 -62
rect 8491 -96 8525 -62
rect 8561 -96 8595 -62
rect 8631 -96 8665 -62
rect 8701 -96 8735 -62
rect 8771 -96 8805 -62
rect 8841 -96 8875 -62
rect 8911 -96 8945 -62
rect 8981 -96 9015 -62
rect 9051 -96 9085 -62
rect 9121 -96 9155 -62
rect 9191 -96 9225 -62
rect 9261 -96 9295 -62
rect 9331 -96 9365 -62
rect 9401 -96 9435 -62
rect 9471 -96 9505 -62
rect 9541 -96 9575 -62
rect 9611 -96 9645 -62
rect 9681 -96 9715 -62
rect 9751 -96 9785 -62
rect 9821 -96 9855 -62
rect 9891 -96 9925 -62
rect 9961 -96 9995 -62
rect 10031 -96 10065 -62
rect 10101 -96 10135 -62
rect 10170 -96 10204 -62
rect 10239 -96 10273 -62
rect 10308 -96 10342 -62
rect 10377 -96 10411 -62
rect 10446 -96 10480 -62
rect 11314 -105 11348 -71
rect 11385 -105 11419 -71
rect 11456 -105 11490 -71
rect 11527 -105 11561 -71
rect 11598 -105 11632 -71
rect 11669 -105 11703 -71
rect 11740 -105 11774 -71
rect 11811 -105 11845 -71
rect 11882 -105 11916 -71
rect 11953 -105 11987 -71
rect 12024 -105 12058 -71
rect 12095 -105 12129 -71
rect 12166 -105 12200 -71
rect 12237 -105 12271 -71
rect 12308 -105 12342 -71
rect 12379 -105 12413 -71
rect 12450 -105 12484 -71
rect 12521 -105 12555 -71
rect 12592 -105 12626 -71
rect 12663 -105 12697 -71
rect 12734 -105 12768 -71
rect 12804 -105 12838 -71
rect 8119 -174 8149 -140
rect 8184 -174 8218 -140
rect 8253 -174 8287 -140
rect 8322 -174 8356 -140
rect 8390 -174 8424 -140
rect 8458 -174 8492 -140
rect 8526 -174 8560 -140
rect 8594 -174 8628 -140
rect 8662 -174 8696 -140
rect 8730 -174 8764 -140
rect 8798 -174 8832 -140
rect 8866 -174 8900 -140
rect 8934 -174 8968 -140
rect 9002 -174 9036 -140
rect 9070 -174 9104 -140
rect 9138 -174 9172 -140
rect 9206 -174 9240 -140
rect 9274 -174 9308 -140
rect 9342 -174 9376 -140
rect 9410 -174 9444 -140
rect 9478 -174 9512 -140
rect 9546 -174 9580 -140
rect 9614 -174 9648 -140
rect 9682 -174 9716 -140
rect 9750 -174 9784 -140
rect 9818 -174 9852 -140
rect 9886 -174 9920 -140
rect 9954 -174 9988 -140
rect 10022 -174 10056 -140
rect 10090 -174 10124 -140
rect 10158 -174 10192 -140
rect 10226 -174 10260 -140
rect 10294 -174 10328 -140
rect 10362 -174 10396 -140
rect 10430 -174 10464 -140
rect 10498 -174 10501 -140
rect 11128 -174 11144 -140
rect 11178 -174 11212 -140
rect 11246 -174 11280 -140
rect 11314 -175 11348 -141
rect 11385 -175 11419 -141
rect 11456 -175 11490 -141
rect 11527 -175 11561 -141
rect 11598 -175 11632 -141
rect 11669 -175 11703 -141
rect 11740 -175 11774 -141
rect 11811 -175 11845 -141
rect 11882 -175 11916 -141
rect 11953 -175 11987 -141
rect 12024 -175 12058 -141
rect 12095 -175 12129 -141
rect 12166 -175 12200 -141
rect 12237 -175 12271 -141
rect 12308 -175 12342 -141
rect 12379 -175 12413 -141
rect 12450 -175 12484 -141
rect 12521 -175 12555 -141
rect 12592 -175 12626 -141
rect 12663 -175 12697 -141
rect 12734 -175 12768 -141
rect 12804 -175 12838 -141
<< mvnsubdiffcont >>
rect 1234 8545 1268 8579
rect 1302 8545 1336 8579
rect 1370 8545 1404 8579
rect 1438 8545 1472 8579
rect 1506 8545 1540 8579
rect 1574 8545 1608 8579
rect 1642 8545 1676 8579
rect 1710 8545 1744 8579
rect 1778 8545 1812 8579
rect 1846 8545 1880 8579
rect 1914 8545 1948 8579
rect 1982 8545 2016 8579
rect 2050 8545 2084 8579
rect 2118 8545 2152 8579
rect 2186 8545 2220 8579
rect 2254 8545 2288 8579
rect 2322 8545 2356 8579
rect 2390 8545 2424 8579
rect 2458 8545 2492 8579
rect 2526 8545 2560 8579
rect 2594 8545 2628 8579
rect 2662 8545 2696 8579
rect 2730 8545 2764 8579
rect 2798 8545 2832 8579
rect 2866 8545 2900 8579
rect 2934 8545 2968 8579
rect 3002 8545 3036 8579
rect 3070 8545 3104 8579
rect 3138 8545 3172 8579
rect 3206 8545 3240 8579
rect 3274 8545 3308 8579
rect 3342 8545 3376 8579
rect 3410 8545 3444 8579
rect 3478 8545 3512 8579
rect 3546 8545 3580 8579
rect 3614 8545 3648 8579
rect 3682 8545 3716 8579
rect 3750 8545 3784 8579
rect 3818 8545 3852 8579
rect 3886 8545 3920 8579
rect 3954 8545 3988 8579
rect 4022 8545 4056 8579
rect 4090 8545 4124 8579
rect 4158 8545 4192 8579
rect 4226 8545 4260 8579
rect 4294 8545 4328 8579
rect 1167 8455 1201 8489
rect 4409 8478 4443 8512
rect 1167 8387 1201 8421
rect 1167 8319 1201 8353
rect 1167 8251 1201 8285
rect 1167 8183 1201 8217
rect 1167 8115 1201 8149
rect 1167 8047 1201 8081
rect 1167 7979 1201 8013
rect 1167 7911 1201 7945
rect 1167 7843 1201 7877
rect 1167 7775 1201 7809
rect 1167 7707 1201 7741
rect 1167 7639 1201 7673
rect 1167 7571 1201 7605
rect 1167 7503 1201 7537
rect 1167 7435 1201 7469
rect 1167 7367 1201 7401
rect 4409 8410 4443 8444
rect 4409 8342 4443 8376
rect 4409 8274 4443 8308
rect 4409 8206 4443 8240
rect 4409 8138 4443 8172
rect 4409 8070 4443 8104
rect 4409 8002 4443 8036
rect 4409 7934 4443 7968
rect 4409 7866 4443 7900
rect 4409 7798 4443 7832
rect 4409 7730 4443 7764
rect 4409 7662 4443 7696
rect 4409 7594 4443 7628
rect 4409 7526 4443 7560
rect 4409 7458 4443 7492
rect 4409 7390 4443 7424
rect 1167 7299 1201 7333
rect 4409 7322 4443 7356
rect 1291 7232 1325 7266
rect 1359 7232 1393 7266
rect 1427 7232 1461 7266
rect 1495 7232 1529 7266
rect 1622 7232 1656 7266
rect 1690 7232 1724 7266
rect 1758 7232 1792 7266
rect 1826 7232 1860 7266
rect 1894 7232 1928 7266
rect 1962 7232 1996 7266
rect 2030 7232 2064 7266
rect 2098 7232 2132 7266
rect 2166 7232 2200 7266
rect 2234 7232 2268 7266
rect 2302 7232 2336 7266
rect 2370 7232 2404 7266
rect 2438 7232 2472 7266
rect 2506 7232 2540 7266
rect 2574 7232 2608 7266
rect 2642 7232 2676 7266
rect 2710 7232 2744 7266
rect 2778 7232 2812 7266
rect 2846 7232 2880 7266
rect 2914 7232 2948 7266
rect 2982 7232 3016 7266
rect 3050 7232 3084 7266
rect 3118 7232 3152 7266
rect 3186 7232 3220 7266
rect 3254 7232 3288 7266
rect 3322 7232 3356 7266
rect 3390 7232 3424 7266
rect 3458 7232 3492 7266
rect 3526 7232 3560 7266
rect 3594 7232 3628 7266
rect 3662 7232 3696 7266
rect 3730 7232 3764 7266
rect 3798 7232 3832 7266
rect 3866 7232 3900 7266
rect 3934 7232 3968 7266
rect 4002 7232 4036 7266
rect 4070 7232 4104 7266
rect 4138 7232 4172 7266
rect 4206 7232 4240 7266
rect 4274 7232 4308 7266
rect 4342 7232 4376 7266
rect 13193 4206 13227 4240
rect 14983 4268 15017 4302
rect 14983 4200 15017 4234
rect 13193 4138 13227 4172
rect 13193 4070 13227 4104
rect 13193 4002 13227 4036
rect 13193 3934 13227 3968
rect 13193 3866 13227 3900
rect 13193 3798 13227 3832
rect 13193 3730 13227 3764
rect 13193 3662 13227 3696
rect 13193 3594 13227 3628
rect 13193 3526 13227 3560
rect 13193 3458 13227 3492
rect 13193 3390 13227 3424
rect 13193 3322 13227 3356
rect 13193 3254 13227 3288
rect 14983 4132 15017 4166
rect 14983 4064 15017 4098
rect 14983 3996 15017 4030
rect 14983 3928 15017 3962
rect 14983 3860 15017 3894
rect 14983 3792 15017 3826
rect 14983 3724 15017 3758
rect 14983 3656 15017 3690
rect 14983 3588 15017 3622
rect 14983 3520 15017 3554
rect 14983 3452 15017 3486
rect 14983 3384 15017 3418
rect 14983 3316 15017 3350
rect 14983 3248 15017 3282
rect 13193 3186 13227 3220
rect 13193 3118 13227 3152
rect 14983 3180 15017 3214
rect 13193 3050 13227 3084
rect 14983 3112 15017 3146
rect 14983 3044 15017 3078
rect 13193 2982 13227 3016
rect 13193 2914 13227 2948
rect 14983 2976 15017 3010
rect 14983 2908 15017 2942
rect 13193 2846 13227 2880
rect 13261 2847 13295 2881
rect 13330 2847 13364 2881
rect 13399 2847 13433 2881
rect 13468 2847 13502 2881
rect 13537 2847 13571 2881
rect 13606 2847 13640 2881
rect 13675 2847 13709 2881
rect 13744 2847 13778 2881
rect 13813 2847 13847 2881
rect 13882 2847 13916 2881
rect 13951 2847 13985 2881
rect 14020 2847 14054 2881
rect 14089 2847 14123 2881
rect 14158 2847 14192 2881
rect 14227 2847 14261 2881
rect 14296 2847 14330 2881
rect 14365 2847 14399 2881
rect 14434 2847 14468 2881
rect 14503 2847 14537 2881
rect 14572 2847 14606 2881
rect 14641 2847 14675 2881
rect 14710 2847 14744 2881
rect 14779 2847 14813 2881
rect 14847 2847 14881 2881
rect 14915 2847 14949 2881
rect 13193 2778 13227 2812
rect 13193 2710 13227 2744
rect 14983 2840 15017 2874
rect 14983 2772 15017 2806
rect 14983 2704 15017 2738
rect 13193 2642 13227 2676
rect 13193 2574 13227 2608
rect 13193 2506 13227 2540
rect 13193 2438 13227 2472
rect 13193 2370 13227 2404
rect 13193 2302 13227 2336
rect 13193 2234 13227 2268
rect 13193 2166 13227 2200
rect 13193 2098 13227 2132
rect 13193 2030 13227 2064
rect 13193 1962 13227 1996
rect 13193 1894 13227 1928
rect 13193 1826 13227 1860
rect 13193 1758 13227 1792
rect 13193 1690 13227 1724
rect 13193 1622 13227 1656
rect 13193 1554 13227 1588
rect 13193 1486 13227 1520
rect 13193 1418 13227 1452
rect 13193 1350 13227 1384
rect 13193 1282 13227 1316
rect 13193 1214 13227 1248
rect 13193 1146 13227 1180
rect 13193 1078 13227 1112
rect 13193 1010 13227 1044
rect 13193 942 13227 976
rect 13193 874 13227 908
rect 13193 806 13227 840
rect 13193 738 13227 772
rect 13193 670 13227 704
rect 13193 602 13227 636
rect 13193 534 13227 568
rect 13193 466 13227 500
rect 13193 398 13227 432
rect 13193 330 13227 364
rect 13193 262 13227 296
rect 14983 2636 15017 2670
rect 14983 2568 15017 2602
rect 14983 2500 15017 2534
rect 14983 2432 15017 2466
rect 14983 2364 15017 2398
rect 14983 2296 15017 2330
rect 14983 2228 15017 2262
rect 14983 2160 15017 2194
rect 14983 2092 15017 2126
rect 14983 2024 15017 2058
rect 14983 1956 15017 1990
rect 14983 1888 15017 1922
rect 14983 1820 15017 1854
rect 14983 1752 15017 1786
rect 14983 1684 15017 1718
rect 14983 1616 15017 1650
rect 14983 1548 15017 1582
rect 14983 1480 15017 1514
rect 14983 1412 15017 1446
rect 14983 1344 15017 1378
rect 14983 1276 15017 1310
rect 14983 1208 15017 1242
rect 14983 1140 15017 1174
rect 14983 1072 15017 1106
rect 14983 1004 15017 1038
rect 14983 936 15017 970
rect 14983 868 15017 902
rect 14983 800 15017 834
rect 14983 732 15017 766
rect 14983 664 15017 698
rect 14983 596 15017 630
rect 14983 528 15017 562
rect 14983 460 15017 494
rect 14983 392 15017 426
rect 14983 324 15017 358
rect 14983 256 15017 290
rect 13193 194 13227 228
rect 13193 126 13227 160
rect 13193 58 13227 92
rect 14983 188 15017 222
rect 14983 120 15017 154
rect 14983 52 15017 86
rect 13283 -10 13317 24
rect 13351 -10 13385 24
rect 13419 -10 13453 24
rect 13487 -10 13521 24
rect 13555 -10 13589 24
rect 13623 -10 13657 24
rect 13691 -10 13725 24
rect 13759 -10 13793 24
rect 13827 -10 13861 24
rect 13895 -10 13929 24
rect 13963 -10 13997 24
rect 14031 -10 14065 24
rect 14099 -10 14133 24
rect 14167 -10 14201 24
rect 14235 -10 14269 24
rect 14303 -10 14337 24
rect 14371 -10 14405 24
rect 14439 -10 14473 24
rect 14507 -10 14541 24
rect 14575 -10 14609 24
rect 14643 -10 14677 24
rect 14711 -10 14745 24
rect 14779 -10 14813 24
rect 14847 -10 14881 24
rect 14915 -10 14949 24
<< poly >>
rect 4314 8427 4380 8435
rect 1250 8327 1282 8427
rect 4282 8405 4380 8427
rect 4282 8371 4330 8405
rect 4364 8371 4380 8405
rect 4282 8337 4380 8371
rect 4282 8327 4330 8337
rect 4314 8303 4330 8327
rect 4364 8303 4380 8337
rect 4314 8271 4380 8303
rect 1250 8171 1282 8271
rect 4282 8269 4380 8271
rect 4282 8235 4330 8269
rect 4364 8235 4380 8269
rect 4282 8201 4380 8235
rect 4282 8171 4330 8201
rect 4314 8167 4330 8171
rect 4364 8167 4380 8201
rect 4314 8133 4380 8167
rect 4314 8115 4330 8133
rect 1250 8015 1282 8115
rect 4282 8099 4330 8115
rect 4364 8099 4380 8133
rect 4282 8065 4380 8099
rect 4282 8031 4330 8065
rect 4364 8031 4380 8065
rect 4282 8015 4380 8031
rect 4314 7997 4380 8015
rect 4314 7963 4330 7997
rect 4364 7963 4380 7997
rect 4314 7959 4380 7963
rect 1250 7859 1282 7959
rect 4282 7929 4380 7959
rect 4282 7895 4330 7929
rect 4364 7895 4380 7929
rect 4282 7861 4380 7895
rect 4282 7859 4330 7861
rect 4314 7827 4330 7859
rect 4364 7827 4380 7861
rect 4314 7803 4380 7827
rect 1250 7703 1282 7803
rect 4282 7793 4380 7803
rect 4282 7759 4330 7793
rect 4364 7759 4380 7793
rect 4282 7725 4380 7759
rect 4282 7703 4330 7725
rect 4314 7691 4330 7703
rect 4364 7691 4380 7725
rect 4314 7657 4380 7691
rect 4314 7647 4330 7657
rect 1250 7547 1282 7647
rect 4282 7623 4330 7647
rect 4364 7623 4380 7657
rect 4282 7589 4380 7623
rect 4282 7555 4330 7589
rect 4364 7555 4380 7589
rect 4282 7547 4380 7555
rect 4314 7521 4380 7547
rect 4314 7491 4330 7521
rect 1250 7391 1282 7491
rect 4282 7487 4330 7491
rect 4364 7487 4380 7521
rect 4282 7453 4380 7487
rect 4282 7419 4330 7453
rect 4364 7419 4380 7453
rect 4282 7399 4380 7419
rect 4282 7391 4314 7399
rect 13603 4091 13975 4107
rect 13603 4057 13619 4091
rect 13653 4057 13696 4091
rect 13730 4057 13773 4091
rect 13807 4057 13849 4091
rect 13883 4057 13925 4091
rect 13959 4057 13975 4091
rect 13603 4041 13975 4057
rect 13603 4015 13703 4041
rect 13875 4015 13975 4041
rect 14151 4091 14523 4107
rect 14151 4057 14167 4091
rect 14201 4057 14244 4091
rect 14278 4057 14321 4091
rect 14355 4057 14397 4091
rect 14431 4057 14473 4091
rect 14507 4057 14523 4091
rect 14151 4041 14523 4057
rect 14151 4015 14251 4041
rect 14423 4015 14523 4041
rect 13603 3389 13703 3415
rect 13875 3389 13975 3415
rect 14151 3389 14251 3415
rect 14423 3389 14523 3415
rect 13608 3321 13708 3347
rect 13880 3321 13980 3347
rect 14152 3321 14252 3347
rect 14424 3321 14524 3347
rect 13608 3211 13708 3237
rect 13880 3211 13980 3237
rect 13608 3195 13980 3211
rect 13608 3161 13624 3195
rect 13658 3161 13701 3195
rect 13735 3161 13778 3195
rect 13812 3161 13854 3195
rect 13888 3161 13930 3195
rect 13964 3161 13980 3195
rect 13608 3145 13980 3161
rect 13608 3119 13708 3145
rect 13880 3119 13980 3145
rect 14152 3211 14252 3237
rect 14424 3211 14524 3237
rect 14152 3195 14524 3211
rect 14152 3161 14168 3195
rect 14202 3161 14245 3195
rect 14279 3161 14322 3195
rect 14356 3161 14398 3195
rect 14432 3161 14474 3195
rect 14508 3161 14524 3195
rect 14152 3145 14524 3161
rect 14152 3119 14252 3145
rect 14424 3119 14524 3145
rect 13608 3009 13708 3035
rect 13880 3009 13980 3035
rect 14152 3009 14252 3035
rect 14424 3009 14524 3035
rect 13538 2512 13630 2528
rect 13538 2478 13554 2512
rect 13588 2478 13630 2512
rect 13538 2443 13630 2478
rect 13538 2409 13554 2443
rect 13588 2428 13630 2443
rect 14630 2428 14656 2528
rect 13588 2409 13604 2428
rect 13538 2374 13604 2409
rect 13538 2340 13554 2374
rect 13588 2372 13604 2374
rect 13588 2340 13630 2372
rect 13538 2305 13630 2340
rect 13538 2271 13554 2305
rect 13588 2272 13630 2305
rect 14630 2272 14656 2372
rect 13588 2271 13604 2272
rect 13538 2236 13604 2271
rect 13538 2202 13554 2236
rect 13588 2216 13604 2236
rect 13588 2202 13630 2216
rect 13538 2167 13630 2202
rect 13538 2133 13554 2167
rect 13588 2133 13630 2167
rect 13538 2116 13630 2133
rect 14630 2116 14656 2216
rect 13538 2098 13604 2116
rect 13538 2064 13554 2098
rect 13588 2064 13604 2098
rect 13538 2060 13604 2064
rect 13538 2029 13630 2060
rect 13538 1995 13554 2029
rect 13588 1995 13630 2029
rect 13538 1960 13630 1995
rect 14630 1960 14656 2060
rect 13538 1926 13554 1960
rect 13588 1926 13604 1960
rect 13538 1904 13604 1926
rect 13538 1891 13630 1904
rect 13538 1857 13554 1891
rect 13588 1857 13630 1891
rect 13538 1822 13630 1857
rect 13538 1788 13554 1822
rect 13588 1804 13630 1822
rect 14630 1804 14656 1904
rect 13588 1788 13604 1804
rect 13538 1753 13604 1788
rect 13538 1719 13554 1753
rect 13588 1748 13604 1753
rect 13588 1719 13630 1748
rect 13538 1684 13630 1719
rect 13538 1650 13554 1684
rect 13588 1650 13630 1684
rect 13538 1648 13630 1650
rect 14630 1648 14656 1748
rect 13538 1615 13604 1648
rect 13538 1581 13554 1615
rect 13588 1592 13604 1615
rect 13588 1581 13630 1592
rect 13538 1546 13630 1581
rect 13538 1512 13554 1546
rect 13588 1512 13630 1546
rect 13538 1492 13630 1512
rect 14630 1492 14656 1592
rect 13538 1477 13604 1492
rect 13538 1443 13554 1477
rect 13588 1443 13604 1477
rect 13538 1436 13604 1443
rect 13538 1408 13630 1436
rect 13538 1374 13554 1408
rect 13588 1374 13630 1408
rect 13538 1339 13630 1374
rect 13538 1305 13554 1339
rect 13588 1336 13630 1339
rect 14630 1336 14656 1436
rect 13588 1305 13604 1336
rect 13538 1280 13604 1305
rect 13538 1270 13630 1280
rect 13538 1236 13554 1270
rect 13588 1236 13630 1270
rect 13538 1201 13630 1236
rect 13538 1167 13554 1201
rect 13588 1180 13630 1201
rect 14630 1180 14656 1280
rect 13588 1167 13604 1180
rect 13538 1132 13604 1167
rect 13538 1098 13554 1132
rect 13588 1124 13604 1132
rect 13588 1098 13630 1124
rect 13538 1063 13630 1098
rect 13538 1029 13554 1063
rect 13588 1029 13630 1063
rect 13538 1024 13630 1029
rect 14630 1024 14656 1124
rect 13538 994 13604 1024
rect 13538 960 13554 994
rect 13588 968 13604 994
rect 13588 960 13630 968
rect 13538 926 13630 960
rect 13538 892 13554 926
rect 13588 892 13630 926
rect 13538 868 13630 892
rect 14630 868 14656 968
rect 13538 858 13604 868
rect 13538 824 13554 858
rect 13588 824 13604 858
rect 13538 812 13604 824
rect 13538 790 13630 812
rect 13538 756 13554 790
rect 13588 756 13630 790
rect 13538 722 13630 756
rect 13538 688 13554 722
rect 13588 712 13630 722
rect 14630 712 14656 812
rect 13588 688 13604 712
rect 13538 656 13604 688
rect 13538 654 13630 656
rect 13538 620 13554 654
rect 13588 620 13630 654
rect 13538 586 13630 620
rect 13538 552 13554 586
rect 13588 556 13630 586
rect 14630 556 14656 656
rect 13588 552 13604 556
rect 13538 518 13604 552
rect 13538 484 13554 518
rect 13588 500 13604 518
rect 13588 484 13630 500
rect 13538 450 13630 484
rect 13538 416 13554 450
rect 13588 416 13630 450
rect 13538 400 13630 416
rect 14630 400 14656 500
<< polycont >>
rect 4330 8371 4364 8405
rect 4330 8303 4364 8337
rect 4330 8235 4364 8269
rect 4330 8167 4364 8201
rect 4330 8099 4364 8133
rect 4330 8031 4364 8065
rect 4330 7963 4364 7997
rect 4330 7895 4364 7929
rect 4330 7827 4364 7861
rect 4330 7759 4364 7793
rect 4330 7691 4364 7725
rect 4330 7623 4364 7657
rect 4330 7555 4364 7589
rect 4330 7487 4364 7521
rect 4330 7419 4364 7453
rect 13619 4057 13653 4091
rect 13696 4057 13730 4091
rect 13773 4057 13807 4091
rect 13849 4057 13883 4091
rect 13925 4057 13959 4091
rect 14167 4057 14201 4091
rect 14244 4057 14278 4091
rect 14321 4057 14355 4091
rect 14397 4057 14431 4091
rect 14473 4057 14507 4091
rect 13624 3161 13658 3195
rect 13701 3161 13735 3195
rect 13778 3161 13812 3195
rect 13854 3161 13888 3195
rect 13930 3161 13964 3195
rect 14168 3161 14202 3195
rect 14245 3161 14279 3195
rect 14322 3161 14356 3195
rect 14398 3161 14432 3195
rect 14474 3161 14508 3195
rect 13554 2478 13588 2512
rect 13554 2409 13588 2443
rect 13554 2340 13588 2374
rect 13554 2271 13588 2305
rect 13554 2202 13588 2236
rect 13554 2133 13588 2167
rect 13554 2064 13588 2098
rect 13554 1995 13588 2029
rect 13554 1926 13588 1960
rect 13554 1857 13588 1891
rect 13554 1788 13588 1822
rect 13554 1719 13588 1753
rect 13554 1650 13588 1684
rect 13554 1581 13588 1615
rect 13554 1512 13588 1546
rect 13554 1443 13588 1477
rect 13554 1374 13588 1408
rect 13554 1305 13588 1339
rect 13554 1236 13588 1270
rect 13554 1167 13588 1201
rect 13554 1098 13588 1132
rect 13554 1029 13588 1063
rect 13554 960 13588 994
rect 13554 892 13588 926
rect 13554 824 13588 858
rect 13554 756 13588 790
rect 13554 688 13588 722
rect 13554 620 13588 654
rect 13554 552 13588 586
rect 13554 484 13588 518
rect 13554 416 13588 450
<< locali >>
rect 7860 9779 7942 9813
rect 7826 9739 7976 9779
rect 7860 9705 7942 9739
rect 9391 9779 9473 9813
rect 9357 9739 9507 9779
rect 7826 9665 7976 9705
rect 7860 9631 7942 9665
rect 7826 9591 7976 9631
rect 7860 9557 7942 9591
rect 7826 9517 7976 9557
rect 7860 9483 7942 9517
rect 8640 9507 8736 9716
rect 9391 9705 9473 9739
rect 9357 9665 9507 9705
rect 9391 9631 9473 9665
rect 9357 9591 9507 9631
rect 9391 9557 9473 9591
rect 9357 9517 9507 9557
rect 7826 9443 7976 9483
rect 7860 9409 7942 9443
rect 9391 9483 9473 9517
rect 9357 9443 9507 9483
rect 9391 9409 9473 9443
rect 800 8779 907 8791
rect 834 8757 907 8779
rect 945 8757 975 8791
rect 1017 8757 1043 8791
rect 1089 8757 1111 8791
rect 1161 8757 1179 8791
rect 1233 8757 1247 8791
rect 1305 8757 1315 8791
rect 1377 8757 1383 8791
rect 1449 8757 1451 8791
rect 1485 8757 1487 8791
rect 1553 8757 1559 8791
rect 1621 8757 1631 8791
rect 1689 8757 1703 8791
rect 1757 8757 1775 8791
rect 1825 8757 1847 8791
rect 1893 8757 1919 8791
rect 1961 8757 1991 8791
rect 2029 8757 2063 8791
rect 2097 8757 2131 8791
rect 2169 8757 2199 8791
rect 2241 8757 2267 8791
rect 2313 8757 2335 8791
rect 2385 8757 2403 8791
rect 2457 8757 2471 8791
rect 2529 8757 2539 8791
rect 2601 8757 2607 8791
rect 2673 8757 2675 8791
rect 2709 8757 2711 8791
rect 2777 8757 2783 8791
rect 2845 8757 2855 8791
rect 2913 8757 2927 8791
rect 2981 8757 2999 8791
rect 3049 8757 3071 8791
rect 3117 8757 3143 8791
rect 3185 8757 3215 8791
rect 3253 8757 3287 8791
rect 3321 8757 3355 8791
rect 3393 8757 3423 8791
rect 3465 8757 3491 8791
rect 3537 8757 3559 8791
rect 3609 8757 3627 8791
rect 3681 8757 3695 8791
rect 3753 8757 3763 8791
rect 3825 8757 3831 8791
rect 3897 8757 3899 8791
rect 3933 8757 3935 8791
rect 4001 8757 4007 8791
rect 4069 8757 4079 8791
rect 4137 8757 4151 8791
rect 4205 8757 4223 8791
rect 4273 8757 4295 8791
rect 4341 8757 4367 8791
rect 4409 8757 4439 8791
rect 4477 8757 4511 8791
rect 4545 8757 4579 8791
rect 4617 8757 4647 8791
rect 4689 8757 4715 8791
rect 4761 8757 4773 8791
rect 800 8707 834 8733
rect 800 8635 834 8665
rect 800 8563 834 8597
rect 800 8495 834 8529
rect 800 8427 834 8457
rect 800 8359 834 8385
rect 800 8291 834 8313
rect 800 8223 834 8241
rect 800 8155 834 8169
rect 800 8087 834 8097
rect 800 8019 834 8025
rect 800 7951 834 7953
rect 800 7915 834 7917
rect 800 7843 834 7849
rect 800 7771 834 7781
rect 800 7699 834 7713
rect 800 7627 834 7645
rect 800 7555 834 7577
rect 800 7483 834 7509
rect 800 7411 834 7441
rect 800 7339 834 7373
rect 800 7271 834 7305
rect 800 7203 834 7233
rect 1161 8586 4514 8592
rect 1161 8552 1173 8586
rect 1207 8579 1245 8586
rect 1279 8579 1317 8586
rect 1351 8579 1389 8586
rect 1423 8579 1461 8586
rect 1495 8579 1533 8586
rect 1567 8579 1605 8586
rect 1639 8579 1677 8586
rect 1711 8579 1749 8586
rect 1783 8579 1821 8586
rect 1855 8579 1893 8586
rect 1927 8579 1965 8586
rect 1999 8579 2037 8586
rect 2071 8579 2109 8586
rect 2143 8579 2181 8586
rect 2215 8579 2253 8586
rect 2287 8579 2325 8586
rect 2359 8579 2397 8586
rect 2431 8579 2469 8586
rect 2503 8579 2541 8586
rect 2575 8579 2613 8586
rect 2647 8579 2685 8586
rect 2719 8579 2757 8586
rect 2791 8579 2829 8586
rect 2863 8579 2901 8586
rect 2935 8579 2973 8586
rect 3007 8579 3045 8586
rect 3079 8579 3117 8586
rect 3151 8579 3189 8586
rect 3223 8579 3261 8586
rect 3295 8579 3333 8586
rect 3367 8579 3405 8586
rect 3439 8579 3477 8586
rect 3511 8579 3549 8586
rect 3583 8579 3621 8586
rect 3655 8579 3693 8586
rect 3727 8579 3765 8586
rect 3799 8579 3837 8586
rect 3871 8579 3909 8586
rect 3943 8579 3981 8586
rect 4015 8579 4053 8586
rect 4087 8579 4125 8586
rect 4159 8579 4197 8586
rect 4231 8579 4269 8586
rect 4303 8579 4341 8586
rect 1207 8552 1234 8579
rect 1279 8552 1302 8579
rect 1351 8552 1370 8579
rect 1423 8552 1438 8579
rect 1495 8552 1506 8579
rect 1567 8552 1574 8579
rect 1639 8552 1642 8579
rect 1161 8545 1234 8552
rect 1268 8545 1302 8552
rect 1336 8545 1370 8552
rect 1404 8545 1438 8552
rect 1472 8545 1506 8552
rect 1540 8545 1574 8552
rect 1608 8545 1642 8552
rect 1676 8552 1677 8579
rect 1744 8552 1749 8579
rect 1812 8552 1821 8579
rect 1880 8552 1893 8579
rect 1948 8552 1965 8579
rect 2016 8552 2037 8579
rect 2084 8552 2109 8579
rect 2152 8552 2181 8579
rect 2220 8552 2253 8579
rect 1676 8545 1710 8552
rect 1744 8545 1778 8552
rect 1812 8545 1846 8552
rect 1880 8545 1914 8552
rect 1948 8545 1982 8552
rect 2016 8545 2050 8552
rect 2084 8545 2118 8552
rect 2152 8545 2186 8552
rect 2220 8545 2254 8552
rect 2288 8545 2322 8579
rect 2359 8552 2390 8579
rect 2431 8552 2458 8579
rect 2503 8552 2526 8579
rect 2575 8552 2594 8579
rect 2647 8552 2662 8579
rect 2719 8552 2730 8579
rect 2791 8552 2798 8579
rect 2863 8552 2866 8579
rect 2356 8545 2390 8552
rect 2424 8545 2458 8552
rect 2492 8545 2526 8552
rect 2560 8545 2594 8552
rect 2628 8545 2662 8552
rect 2696 8545 2730 8552
rect 2764 8545 2798 8552
rect 2832 8545 2866 8552
rect 2900 8552 2901 8579
rect 2968 8552 2973 8579
rect 3036 8552 3045 8579
rect 3104 8552 3117 8579
rect 3172 8552 3189 8579
rect 3240 8552 3261 8579
rect 3308 8552 3333 8579
rect 3376 8552 3405 8579
rect 3444 8552 3477 8579
rect 2900 8545 2934 8552
rect 2968 8545 3002 8552
rect 3036 8545 3070 8552
rect 3104 8545 3138 8552
rect 3172 8545 3206 8552
rect 3240 8545 3274 8552
rect 3308 8545 3342 8552
rect 3376 8545 3410 8552
rect 3444 8545 3478 8552
rect 3512 8545 3546 8579
rect 3583 8552 3614 8579
rect 3655 8552 3682 8579
rect 3727 8552 3750 8579
rect 3799 8552 3818 8579
rect 3871 8552 3886 8579
rect 3943 8552 3954 8579
rect 4015 8552 4022 8579
rect 4087 8552 4090 8579
rect 3580 8545 3614 8552
rect 3648 8545 3682 8552
rect 3716 8545 3750 8552
rect 3784 8545 3818 8552
rect 3852 8545 3886 8552
rect 3920 8545 3954 8552
rect 3988 8545 4022 8552
rect 4056 8545 4090 8552
rect 4124 8552 4125 8579
rect 4192 8552 4197 8579
rect 4260 8552 4269 8579
rect 4328 8552 4341 8579
rect 4375 8580 4514 8586
rect 4375 8552 4474 8580
rect 4124 8545 4158 8552
rect 4192 8545 4226 8552
rect 4260 8545 4294 8552
rect 4328 8546 4474 8552
rect 4508 8546 4514 8580
rect 4328 8545 4514 8546
rect 1161 8544 4514 8545
rect 1161 8496 1207 8544
rect 1161 8455 1167 8496
rect 1201 8455 1207 8496
rect 4408 8512 4514 8544
rect 4408 8478 4409 8512
rect 4443 8508 4514 8512
rect 4443 8478 4474 8508
rect 1279 8472 4220 8478
rect 4408 8474 4474 8478
rect 4508 8474 4514 8508
rect 1161 8424 1207 8455
rect 1278 8438 1294 8472
rect 1328 8438 1362 8472
rect 1400 8438 1430 8472
rect 1472 8438 1498 8472
rect 1544 8438 1566 8472
rect 1616 8438 1634 8472
rect 1688 8438 1702 8472
rect 1760 8438 1770 8472
rect 1832 8438 1838 8472
rect 1904 8438 1906 8472
rect 1940 8438 1942 8472
rect 2008 8438 2014 8472
rect 2076 8438 2086 8472
rect 2144 8438 2158 8472
rect 2212 8438 2230 8472
rect 2280 8438 2302 8472
rect 2348 8438 2374 8472
rect 2416 8438 2446 8472
rect 2484 8438 2518 8472
rect 2552 8438 2586 8472
rect 2624 8438 2654 8472
rect 2696 8438 2722 8472
rect 2768 8438 2790 8472
rect 2840 8438 2858 8472
rect 2912 8438 2926 8472
rect 2984 8438 2994 8472
rect 3056 8438 3062 8472
rect 3128 8438 3130 8472
rect 3164 8438 3166 8472
rect 3232 8438 3238 8472
rect 3300 8438 3310 8472
rect 3368 8438 3382 8472
rect 3436 8438 3454 8472
rect 3504 8438 3526 8472
rect 3572 8438 3598 8472
rect 3640 8438 3670 8472
rect 3708 8438 3742 8472
rect 3776 8438 3810 8472
rect 3848 8438 3878 8472
rect 3920 8438 3946 8472
rect 3992 8438 4014 8472
rect 4064 8438 4082 8472
rect 4136 8438 4150 8472
rect 4208 8438 4218 8472
rect 4252 8438 4268 8472
rect 4408 8444 4514 8474
rect 1279 8432 4220 8438
rect 1161 8387 1167 8424
rect 1201 8387 1207 8424
rect 1161 8353 1207 8387
rect 1161 8318 1167 8353
rect 1201 8318 1207 8353
rect 4330 8415 4364 8435
rect 4330 8338 4364 8371
rect 1161 8285 1207 8318
rect 1287 8316 4220 8322
rect 1161 8246 1167 8285
rect 1201 8246 1207 8285
rect 1278 8282 1294 8316
rect 1328 8282 1362 8316
rect 1400 8282 1430 8316
rect 1472 8282 1498 8316
rect 1544 8282 1566 8316
rect 1616 8282 1634 8316
rect 1688 8282 1702 8316
rect 1760 8282 1770 8316
rect 1832 8282 1838 8316
rect 1904 8282 1906 8316
rect 1940 8282 1942 8316
rect 2008 8282 2014 8316
rect 2076 8282 2086 8316
rect 2144 8282 2158 8316
rect 2212 8282 2230 8316
rect 2280 8282 2302 8316
rect 2348 8282 2374 8316
rect 2416 8282 2446 8316
rect 2484 8282 2518 8316
rect 2552 8282 2586 8316
rect 2624 8282 2654 8316
rect 2696 8282 2722 8316
rect 2768 8282 2790 8316
rect 2840 8282 2858 8316
rect 2912 8282 2926 8316
rect 2984 8282 2994 8316
rect 3056 8282 3062 8316
rect 3128 8282 3130 8316
rect 3164 8282 3166 8316
rect 3232 8282 3238 8316
rect 3300 8282 3310 8316
rect 3368 8282 3382 8316
rect 3436 8282 3454 8316
rect 3504 8282 3526 8316
rect 3572 8282 3598 8316
rect 3640 8282 3670 8316
rect 3708 8282 3742 8316
rect 3776 8282 3810 8316
rect 3848 8282 3878 8316
rect 3920 8282 3946 8316
rect 3992 8282 4014 8316
rect 4064 8282 4082 8316
rect 4136 8282 4150 8316
rect 4208 8282 4218 8316
rect 4252 8282 4268 8316
rect 1287 8276 4220 8282
rect 1161 8217 1207 8246
rect 1161 8174 1167 8217
rect 1201 8174 1207 8217
rect 1161 8149 1207 8174
rect 4330 8269 4364 8303
rect 4330 8201 4364 8227
rect 1279 8160 4220 8166
rect 1161 8102 1167 8149
rect 1201 8102 1207 8149
rect 1278 8126 1294 8160
rect 1328 8126 1362 8160
rect 1400 8126 1430 8160
rect 1472 8126 1498 8160
rect 1544 8126 1566 8160
rect 1616 8126 1634 8160
rect 1688 8126 1702 8160
rect 1760 8126 1770 8160
rect 1832 8126 1838 8160
rect 1904 8126 1906 8160
rect 1940 8126 1942 8160
rect 2008 8126 2014 8160
rect 2076 8126 2086 8160
rect 2144 8126 2158 8160
rect 2212 8126 2230 8160
rect 2280 8126 2302 8160
rect 2348 8126 2374 8160
rect 2416 8126 2446 8160
rect 2484 8126 2518 8160
rect 2552 8126 2586 8160
rect 2624 8126 2654 8160
rect 2696 8126 2722 8160
rect 2768 8126 2790 8160
rect 2840 8126 2858 8160
rect 2912 8126 2926 8160
rect 2984 8126 2994 8160
rect 3056 8126 3062 8160
rect 3128 8126 3130 8160
rect 3164 8126 3166 8160
rect 3232 8126 3238 8160
rect 3300 8126 3310 8160
rect 3368 8126 3382 8160
rect 3436 8126 3454 8160
rect 3504 8126 3526 8160
rect 3572 8126 3598 8160
rect 3640 8126 3670 8160
rect 3708 8126 3742 8160
rect 3776 8126 3810 8160
rect 3848 8126 3878 8160
rect 3920 8126 3946 8160
rect 3992 8126 4014 8160
rect 4064 8126 4082 8160
rect 4136 8126 4150 8160
rect 4208 8126 4218 8160
rect 4252 8126 4268 8160
rect 4330 8133 4364 8150
rect 1279 8120 4220 8126
rect 1161 8081 1207 8102
rect 1161 8030 1167 8081
rect 1201 8030 1207 8081
rect 1161 8013 1207 8030
rect 1161 7958 1167 8013
rect 1201 7958 1207 8013
rect 4330 8065 4364 8073
rect 4330 8030 4364 8031
rect 1287 8004 4220 8010
rect 1278 7970 1294 8004
rect 1328 7970 1362 8004
rect 1400 7970 1430 8004
rect 1472 7970 1498 8004
rect 1544 7970 1566 8004
rect 1616 7970 1634 8004
rect 1688 7970 1702 8004
rect 1760 7970 1770 8004
rect 1832 7970 1838 8004
rect 1904 7970 1906 8004
rect 1940 7970 1942 8004
rect 2008 7970 2014 8004
rect 2076 7970 2086 8004
rect 2144 7970 2158 8004
rect 2212 7970 2230 8004
rect 2280 7970 2302 8004
rect 2348 7970 2374 8004
rect 2416 7970 2446 8004
rect 2484 7970 2518 8004
rect 2552 7970 2586 8004
rect 2624 7970 2654 8004
rect 2696 7970 2722 8004
rect 2768 7970 2790 8004
rect 2840 7970 2858 8004
rect 2912 7970 2926 8004
rect 2984 7970 2994 8004
rect 3056 7970 3062 8004
rect 3128 7970 3130 8004
rect 3164 7970 3166 8004
rect 3232 7970 3238 8004
rect 3300 7970 3310 8004
rect 3368 7970 3382 8004
rect 3436 7970 3454 8004
rect 3504 7970 3526 8004
rect 3572 7970 3598 8004
rect 3640 7970 3670 8004
rect 3708 7970 3742 8004
rect 3776 7970 3810 8004
rect 3848 7970 3878 8004
rect 3920 7970 3946 8004
rect 3992 7970 4014 8004
rect 4064 7970 4082 8004
rect 4136 7970 4150 8004
rect 4208 7970 4218 8004
rect 4252 7970 4268 8004
rect 1287 7964 4220 7970
rect 1161 7945 1207 7958
rect 1161 7886 1167 7945
rect 1201 7886 1207 7945
rect 1161 7877 1207 7886
rect 1161 7814 1167 7877
rect 1201 7814 1207 7877
rect 4330 7953 4364 7963
rect 4330 7876 4364 7895
rect 1279 7848 4220 7854
rect 1278 7814 1294 7848
rect 1328 7814 1362 7848
rect 1400 7814 1430 7848
rect 1472 7814 1498 7848
rect 1544 7814 1566 7848
rect 1616 7814 1634 7848
rect 1688 7814 1702 7848
rect 1760 7814 1770 7848
rect 1832 7814 1838 7848
rect 1904 7814 1906 7848
rect 1940 7814 1942 7848
rect 2008 7814 2014 7848
rect 2076 7814 2086 7848
rect 2144 7814 2158 7848
rect 2212 7814 2230 7848
rect 2280 7814 2302 7848
rect 2348 7814 2374 7848
rect 2416 7814 2446 7848
rect 2484 7814 2518 7848
rect 2552 7814 2586 7848
rect 2624 7814 2654 7848
rect 2696 7814 2722 7848
rect 2768 7814 2790 7848
rect 2840 7814 2858 7848
rect 2912 7814 2926 7848
rect 2984 7814 2994 7848
rect 3056 7814 3062 7848
rect 3128 7814 3130 7848
rect 3164 7814 3166 7848
rect 3232 7814 3238 7848
rect 3300 7814 3310 7848
rect 3368 7814 3382 7848
rect 3436 7814 3454 7848
rect 3504 7814 3526 7848
rect 3572 7814 3598 7848
rect 3640 7814 3670 7848
rect 3708 7814 3742 7848
rect 3776 7814 3810 7848
rect 3848 7814 3878 7848
rect 3920 7814 3946 7848
rect 3992 7814 4014 7848
rect 4064 7814 4082 7848
rect 4136 7814 4150 7848
rect 4208 7814 4218 7848
rect 4252 7814 4268 7848
rect 1161 7809 1207 7814
rect 1161 7742 1167 7809
rect 1201 7742 1207 7809
rect 1279 7808 4220 7814
rect 1161 7741 1207 7742
rect 1161 7707 1167 7741
rect 1201 7707 1207 7741
rect 1161 7704 1207 7707
rect 1161 7639 1167 7704
rect 1201 7639 1207 7704
rect 4330 7799 4364 7827
rect 4330 7725 4364 7759
rect 1284 7692 4220 7698
rect 1278 7658 1294 7692
rect 1328 7658 1362 7692
rect 1400 7658 1430 7692
rect 1472 7658 1498 7692
rect 1544 7658 1566 7692
rect 1616 7658 1634 7692
rect 1688 7658 1702 7692
rect 1760 7658 1770 7692
rect 1832 7658 1838 7692
rect 1904 7658 1906 7692
rect 1940 7658 1942 7692
rect 2008 7658 2014 7692
rect 2076 7658 2086 7692
rect 2144 7658 2158 7692
rect 2212 7658 2230 7692
rect 2280 7658 2302 7692
rect 2348 7658 2374 7692
rect 2416 7658 2446 7692
rect 2484 7658 2518 7692
rect 2552 7658 2586 7692
rect 2624 7658 2654 7692
rect 2696 7658 2722 7692
rect 2768 7658 2790 7692
rect 2840 7658 2858 7692
rect 2912 7658 2926 7692
rect 2984 7658 2994 7692
rect 3056 7658 3062 7692
rect 3128 7658 3130 7692
rect 3164 7658 3166 7692
rect 3232 7658 3238 7692
rect 3300 7658 3310 7692
rect 3368 7658 3382 7692
rect 3436 7658 3454 7692
rect 3504 7658 3526 7692
rect 3572 7658 3598 7692
rect 3640 7658 3670 7692
rect 3708 7658 3742 7692
rect 3776 7658 3810 7692
rect 3848 7658 3878 7692
rect 3920 7658 3946 7692
rect 3992 7658 4014 7692
rect 4064 7658 4082 7692
rect 4136 7658 4150 7692
rect 4208 7658 4218 7692
rect 4252 7658 4268 7692
rect 1284 7652 4220 7658
rect 4330 7657 4364 7687
rect 1161 7632 1207 7639
rect 1161 7571 1167 7632
rect 1201 7571 1207 7632
rect 1161 7560 1207 7571
rect 1161 7503 1167 7560
rect 1201 7503 1207 7560
rect 4330 7589 4364 7609
rect 1279 7536 4220 7542
rect 1161 7488 1207 7503
rect 1278 7502 1294 7536
rect 1328 7502 1362 7536
rect 1400 7502 1430 7536
rect 1472 7502 1498 7536
rect 1544 7502 1566 7536
rect 1616 7502 1634 7536
rect 1688 7502 1702 7536
rect 1760 7502 1770 7536
rect 1832 7502 1838 7536
rect 1904 7502 1906 7536
rect 1940 7502 1942 7536
rect 2008 7502 2014 7536
rect 2076 7502 2086 7536
rect 2144 7502 2158 7536
rect 2212 7502 2230 7536
rect 2280 7502 2302 7536
rect 2348 7502 2374 7536
rect 2416 7502 2446 7536
rect 2484 7502 2518 7536
rect 2552 7502 2586 7536
rect 2624 7502 2654 7536
rect 2696 7502 2722 7536
rect 2768 7502 2790 7536
rect 2840 7502 2858 7536
rect 2912 7502 2926 7536
rect 2984 7502 2994 7536
rect 3056 7502 3062 7536
rect 3128 7502 3130 7536
rect 3164 7502 3166 7536
rect 3232 7502 3238 7536
rect 3300 7502 3310 7536
rect 3368 7502 3382 7536
rect 3436 7502 3454 7536
rect 3504 7502 3526 7536
rect 3572 7502 3598 7536
rect 3640 7502 3670 7536
rect 3708 7502 3742 7536
rect 3776 7502 3810 7536
rect 3848 7502 3878 7536
rect 3920 7502 3946 7536
rect 3992 7502 4014 7536
rect 4064 7502 4082 7536
rect 4136 7502 4150 7536
rect 4208 7502 4218 7536
rect 4252 7502 4268 7536
rect 4330 7521 4364 7531
rect 1279 7496 4220 7502
rect 1161 7435 1167 7488
rect 1201 7435 1207 7488
rect 1161 7416 1207 7435
rect 1161 7367 1167 7416
rect 1201 7367 1207 7416
rect 4330 7399 4364 7419
rect 4408 8410 4409 8444
rect 4443 8436 4514 8444
rect 4443 8410 4474 8436
rect 4408 8402 4474 8410
rect 4508 8402 4514 8436
rect 4408 8376 4514 8402
rect 4408 8342 4409 8376
rect 4443 8364 4514 8376
rect 4443 8342 4474 8364
rect 4408 8330 4474 8342
rect 4508 8330 4514 8364
rect 4408 8308 4514 8330
rect 4408 8274 4409 8308
rect 4443 8292 4514 8308
rect 4443 8274 4474 8292
rect 4408 8258 4474 8274
rect 4508 8258 4514 8292
rect 4408 8240 4514 8258
rect 4408 8206 4409 8240
rect 4443 8220 4514 8240
rect 4443 8206 4474 8220
rect 4408 8186 4474 8206
rect 4508 8186 4514 8220
rect 4408 8172 4514 8186
rect 4408 8138 4409 8172
rect 4443 8148 4514 8172
rect 4443 8138 4474 8148
rect 4408 8114 4474 8138
rect 4508 8114 4514 8148
rect 4408 8104 4514 8114
rect 4408 8070 4409 8104
rect 4443 8076 4514 8104
rect 4443 8070 4474 8076
rect 4408 8042 4474 8070
rect 4508 8042 4514 8076
rect 4408 8036 4514 8042
rect 4408 8002 4409 8036
rect 4443 8004 4514 8036
rect 4443 8002 4474 8004
rect 4408 7970 4474 8002
rect 4508 7970 4514 8004
rect 4408 7968 4514 7970
rect 4408 7934 4409 7968
rect 4443 7934 4514 7968
rect 4408 7932 4514 7934
rect 4408 7900 4474 7932
rect 4408 7866 4409 7900
rect 4443 7898 4474 7900
rect 4508 7898 4514 7932
rect 4443 7866 4514 7898
rect 4408 7860 4514 7866
rect 4408 7832 4474 7860
rect 4408 7798 4409 7832
rect 4443 7826 4474 7832
rect 4508 7826 4514 7860
rect 4443 7798 4514 7826
rect 4408 7788 4514 7798
rect 4408 7764 4474 7788
rect 4408 7730 4409 7764
rect 4443 7754 4474 7764
rect 4508 7754 4514 7788
rect 4443 7730 4514 7754
rect 4408 7716 4514 7730
rect 4408 7696 4474 7716
rect 4408 7662 4409 7696
rect 4443 7682 4474 7696
rect 4508 7682 4514 7716
rect 4443 7662 4514 7682
rect 4408 7644 4514 7662
rect 4408 7628 4474 7644
rect 4408 7594 4409 7628
rect 4443 7610 4474 7628
rect 4508 7610 4514 7644
rect 4443 7594 4514 7610
rect 4408 7572 4514 7594
rect 4408 7560 4474 7572
rect 4408 7526 4409 7560
rect 4443 7538 4474 7560
rect 4508 7538 4514 7572
rect 4443 7526 4514 7538
rect 4408 7500 4514 7526
rect 4408 7492 4474 7500
rect 4408 7458 4409 7492
rect 4443 7466 4474 7492
rect 4508 7466 4514 7500
rect 4443 7458 4514 7466
rect 4408 7428 4514 7458
rect 4408 7424 4474 7428
rect 4408 7390 4409 7424
rect 4443 7394 4474 7424
rect 4508 7394 4514 7428
rect 4443 7390 4514 7394
rect 1161 7344 1207 7367
rect 1161 7299 1167 7344
rect 1201 7299 1207 7344
rect 1278 7380 4220 7386
rect 1278 7346 1294 7380
rect 1328 7346 1362 7380
rect 1400 7346 1430 7380
rect 1472 7346 1498 7380
rect 1544 7346 1566 7380
rect 1616 7346 1634 7380
rect 1688 7346 1702 7380
rect 1760 7346 1770 7380
rect 1832 7346 1838 7380
rect 1904 7346 1906 7380
rect 1940 7346 1942 7380
rect 2008 7346 2014 7380
rect 2076 7346 2086 7380
rect 2144 7346 2158 7380
rect 2212 7346 2230 7380
rect 2280 7346 2302 7380
rect 2348 7346 2374 7380
rect 2416 7346 2446 7380
rect 2484 7346 2518 7380
rect 2552 7346 2586 7380
rect 2624 7346 2654 7380
rect 2696 7346 2722 7380
rect 2768 7346 2790 7380
rect 2840 7346 2858 7380
rect 2912 7346 2926 7380
rect 2984 7346 2994 7380
rect 3056 7346 3062 7380
rect 3128 7346 3130 7380
rect 3164 7346 3166 7380
rect 3232 7346 3238 7380
rect 3300 7346 3310 7380
rect 3368 7346 3382 7380
rect 3436 7346 3454 7380
rect 3504 7346 3526 7380
rect 3572 7346 3598 7380
rect 3640 7346 3670 7380
rect 3708 7346 3742 7380
rect 3776 7346 3810 7380
rect 3848 7346 3878 7380
rect 3920 7346 3946 7380
rect 3992 7346 4014 7380
rect 4064 7346 4082 7380
rect 4136 7346 4150 7380
rect 4208 7346 4218 7380
rect 4252 7346 4268 7380
rect 4408 7356 4514 7390
rect 1278 7340 4220 7346
rect 1161 7272 1207 7299
rect 4408 7322 4409 7356
rect 4443 7322 4514 7356
rect 4408 7272 4514 7322
rect 1161 7238 1167 7272
rect 1201 7266 4514 7272
rect 1201 7238 1291 7266
rect 1161 7232 1291 7238
rect 1334 7232 1359 7266
rect 1406 7232 1427 7266
rect 1478 7232 1495 7266
rect 1550 7232 1588 7266
rect 1656 7232 1660 7266
rect 1724 7232 1732 7266
rect 1792 7232 1804 7266
rect 1860 7232 1876 7266
rect 1928 7232 1948 7266
rect 1996 7232 2020 7266
rect 2064 7232 2092 7266
rect 2132 7232 2164 7266
rect 2200 7232 2234 7266
rect 2270 7232 2302 7266
rect 2342 7232 2370 7266
rect 2414 7232 2438 7266
rect 2486 7232 2506 7266
rect 2558 7232 2574 7266
rect 2630 7232 2642 7266
rect 2702 7232 2710 7266
rect 2774 7232 2778 7266
rect 2880 7232 2884 7266
rect 2948 7232 2956 7266
rect 3016 7232 3028 7266
rect 3084 7232 3100 7266
rect 3152 7232 3172 7266
rect 3220 7232 3244 7266
rect 3288 7232 3316 7266
rect 3356 7232 3388 7266
rect 3424 7232 3458 7266
rect 3494 7232 3526 7266
rect 3566 7232 3594 7266
rect 3638 7232 3662 7266
rect 3710 7232 3730 7266
rect 3782 7232 3798 7266
rect 3854 7232 3866 7266
rect 3926 7232 3934 7266
rect 3998 7232 4002 7266
rect 4104 7232 4108 7266
rect 4172 7232 4180 7266
rect 4240 7232 4252 7266
rect 4308 7232 4324 7266
rect 4376 7232 4396 7266
rect 4430 7232 4468 7266
rect 4502 7232 4514 7266
rect 1161 7226 4514 7232
rect 800 7078 834 7161
rect 800 7044 829 7078
rect 875 7044 901 7078
rect 943 7044 973 7078
rect 1011 7044 1045 7078
rect 1079 7044 1113 7078
rect 1151 7044 1181 7078
rect 1223 7044 1249 7078
rect 1295 7044 1317 7078
rect 1367 7044 1385 7078
rect 1439 7044 1453 7078
rect 1511 7044 1521 7078
rect 1583 7044 1589 7078
rect 1655 7044 1657 7078
rect 1691 7044 1693 7078
rect 1759 7044 1765 7078
rect 1827 7044 1837 7078
rect 1895 7044 1909 7078
rect 1963 7044 1981 7078
rect 2031 7044 2053 7078
rect 2099 7044 2125 7078
rect 2167 7044 2197 7078
rect 2235 7044 2269 7078
rect 2303 7044 2337 7078
rect 2375 7044 2405 7078
rect 2447 7044 2473 7078
rect 2519 7044 2541 7078
rect 2591 7044 2609 7078
rect 2663 7044 2677 7078
rect 2735 7044 2745 7078
rect 2807 7044 2813 7078
rect 2879 7044 2881 7078
rect 2915 7044 2917 7078
rect 2983 7044 2989 7078
rect 3051 7044 3061 7078
rect 3119 7044 3133 7078
rect 3187 7044 3205 7078
rect 3255 7044 3277 7078
rect 3323 7044 3349 7078
rect 3391 7044 3421 7078
rect 3459 7044 3493 7078
rect 3527 7044 3561 7078
rect 3599 7044 3629 7078
rect 3671 7044 3697 7078
rect 3743 7044 3765 7078
rect 3815 7044 3833 7078
rect 3887 7044 3901 7078
rect 3959 7044 3969 7078
rect 4031 7044 4037 7078
rect 4103 7044 4105 7078
rect 4139 7044 4141 7078
rect 4207 7044 4213 7078
rect 4275 7044 4285 7078
rect 4343 7044 4357 7078
rect 4411 7044 4429 7078
rect 4479 7044 4501 7078
rect 4547 7044 4573 7078
rect 4615 7044 4645 7078
rect 4683 7044 4731 7078
rect 4411 7007 4731 7044
rect 4411 7006 4446 7007
rect 4480 7006 4518 7007
rect 4411 6972 4424 7006
rect 4480 6973 4507 7006
rect 4552 6973 4590 7007
rect 4624 6973 4662 7007
rect 4696 7006 4731 7007
rect 4458 6972 4507 6973
rect 4541 6972 4590 6973
rect 4624 6972 4672 6973
rect 4706 6972 4731 7006
rect 4411 6939 4731 6972
rect 4411 6934 4446 6939
rect 4480 6934 4518 6939
rect 4411 6900 4424 6934
rect 4480 6905 4507 6934
rect 4552 6905 4590 6939
rect 4624 6905 4662 6939
rect 4696 6934 4731 6939
rect 4458 6900 4507 6905
rect 4541 6900 4590 6905
rect 4624 6900 4672 6905
rect 4706 6900 4731 6934
rect -874 6759 925 6766
rect -874 6725 -850 6759
rect -816 6725 -781 6759
rect -747 6725 -712 6759
rect -678 6725 -643 6759
rect -609 6725 -574 6759
rect -540 6725 -505 6759
rect -471 6725 -436 6759
rect -402 6725 -367 6759
rect -333 6725 -298 6759
rect -264 6725 -229 6759
rect -195 6725 -160 6759
rect -126 6725 -91 6759
rect -57 6725 -22 6759
rect 12 6725 47 6759
rect 81 6725 116 6759
rect 150 6725 185 6759
rect 219 6725 254 6759
rect 288 6725 323 6759
rect 357 6725 391 6759
rect 425 6725 459 6759
rect 493 6725 527 6759
rect 561 6725 595 6759
rect 629 6725 663 6759
rect 697 6725 731 6759
rect 765 6725 799 6759
rect 833 6725 867 6759
rect 901 6725 925 6759
rect -874 6715 925 6725
rect -874 6689 -849 6715
rect -815 6713 925 6715
rect -815 6689 308 6713
rect 342 6689 382 6713
rect 416 6689 456 6713
rect 490 6689 530 6713
rect 564 6689 604 6713
rect 638 6689 678 6713
rect 712 6689 751 6713
rect 785 6689 824 6713
rect 858 6689 925 6713
rect -874 6655 -850 6689
rect -815 6681 -781 6689
rect -816 6655 -781 6681
rect -747 6655 -712 6689
rect -678 6655 -643 6689
rect -609 6655 -574 6689
rect -540 6655 -505 6689
rect -471 6655 -436 6689
rect -402 6655 -367 6689
rect -333 6655 -298 6689
rect -264 6655 -229 6689
rect -195 6655 -160 6689
rect -126 6655 -91 6689
rect -57 6655 -22 6689
rect 12 6655 47 6689
rect 81 6655 116 6689
rect 150 6655 185 6689
rect 219 6655 254 6689
rect 288 6679 308 6689
rect 357 6679 382 6689
rect 425 6679 456 6689
rect 288 6655 323 6679
rect 357 6655 391 6679
rect 425 6655 459 6679
rect 493 6655 527 6689
rect 564 6679 595 6689
rect 638 6679 663 6689
rect 712 6679 731 6689
rect 785 6679 799 6689
rect 858 6679 867 6689
rect 561 6655 595 6679
rect 629 6655 663 6679
rect 697 6655 731 6679
rect 765 6655 799 6679
rect 833 6655 867 6679
rect 901 6655 925 6689
rect -874 6635 925 6655
rect -874 6619 -849 6635
rect -815 6619 925 6635
rect -874 6585 -850 6619
rect -815 6601 -781 6619
rect -816 6585 -781 6601
rect -747 6585 -712 6619
rect -678 6585 -643 6619
rect -609 6585 -574 6619
rect -540 6585 -505 6619
rect -471 6585 -436 6619
rect -402 6585 -367 6619
rect -333 6585 -298 6619
rect -264 6585 -229 6619
rect -195 6585 -160 6619
rect -126 6585 -91 6619
rect -57 6585 -22 6619
rect 12 6585 47 6619
rect 81 6585 116 6619
rect 150 6585 185 6619
rect 219 6585 254 6619
rect 288 6589 323 6619
rect 357 6589 391 6619
rect 425 6589 459 6619
rect 288 6585 308 6589
rect 357 6585 382 6589
rect 425 6585 456 6589
rect 493 6585 527 6619
rect 561 6589 595 6619
rect 629 6589 663 6619
rect 697 6589 731 6619
rect 765 6589 799 6619
rect 833 6589 867 6619
rect 564 6585 595 6589
rect 638 6585 663 6589
rect 712 6585 731 6589
rect 785 6585 799 6589
rect 858 6585 867 6589
rect 901 6585 925 6619
rect -874 6555 308 6585
rect 342 6555 382 6585
rect 416 6555 456 6585
rect 490 6555 530 6585
rect 564 6555 604 6585
rect 638 6555 678 6585
rect 712 6555 751 6585
rect 785 6555 824 6585
rect 858 6555 925 6585
rect -874 6549 -849 6555
rect -815 6549 925 6555
rect -874 6515 -850 6549
rect -815 6521 -781 6549
rect -816 6515 -781 6521
rect -747 6515 -712 6549
rect -678 6515 -643 6549
rect -609 6515 -574 6549
rect -540 6515 -505 6549
rect -471 6515 -436 6549
rect -402 6515 -367 6549
rect -333 6515 -298 6549
rect -264 6515 -229 6549
rect -195 6515 -160 6549
rect -126 6515 -91 6549
rect -57 6515 -22 6549
rect 12 6515 47 6549
rect 81 6515 116 6549
rect 150 6515 185 6549
rect 219 6515 254 6549
rect 288 6515 323 6549
rect 357 6515 391 6549
rect 425 6515 459 6549
rect 493 6515 527 6549
rect 561 6515 595 6549
rect 629 6515 663 6549
rect 697 6515 731 6549
rect 765 6515 799 6549
rect 833 6515 867 6549
rect 901 6515 925 6549
rect -874 6479 925 6515
rect -874 6445 -850 6479
rect -816 6475 -781 6479
rect -815 6445 -781 6475
rect -747 6445 -712 6479
rect -678 6445 -643 6479
rect -609 6445 -574 6479
rect -540 6445 -505 6479
rect -471 6445 -436 6479
rect -402 6445 -367 6479
rect -333 6445 -298 6479
rect -264 6445 -229 6479
rect -195 6445 -160 6479
rect -126 6445 -91 6479
rect -57 6445 -22 6479
rect 12 6445 47 6479
rect 81 6445 116 6479
rect 150 6445 185 6479
rect 219 6445 254 6479
rect 288 6445 323 6479
rect 357 6445 391 6479
rect 425 6445 459 6479
rect 493 6445 527 6479
rect 561 6445 595 6479
rect 629 6445 663 6479
rect 697 6445 731 6479
rect 765 6445 799 6479
rect 833 6445 867 6479
rect 901 6445 925 6479
rect 1053 6548 1135 6582
rect 1019 6498 1169 6548
rect 1053 6464 1135 6498
rect 2549 6546 3353 6879
rect 4411 6871 4731 6900
rect 4411 6837 4446 6871
rect 4480 6861 4518 6871
rect 4552 6861 4590 6871
rect 4624 6861 4662 6871
rect 4480 6837 4502 6861
rect 4552 6837 4576 6861
rect 4624 6837 4649 6861
rect 4696 6837 4731 6871
rect 4411 6827 4502 6837
rect 4536 6827 4576 6837
rect 4610 6827 4649 6837
rect 4683 6827 4731 6837
rect 4411 6803 4731 6827
rect 4411 6769 4446 6803
rect 4480 6769 4518 6803
rect 4552 6769 4590 6803
rect 4624 6769 4662 6803
rect 4696 6769 4731 6803
rect 4411 6735 4596 6769
rect 4630 6735 4668 6769
rect 4702 6735 4731 6769
rect 4411 6701 4446 6735
rect 4480 6701 4518 6735
rect 4552 6701 4590 6735
rect 4624 6701 4662 6735
rect 4696 6701 4731 6735
rect 4411 6667 4731 6701
rect 4411 6633 4446 6667
rect 4480 6633 4518 6667
rect 4552 6633 4590 6667
rect 4624 6633 4662 6667
rect 4696 6633 4731 6667
rect 4411 6599 4731 6633
rect 2549 6512 2551 6546
rect 2585 6512 2627 6546
rect 2661 6512 2703 6546
rect 2737 6512 2779 6546
rect 2813 6512 2854 6546
rect 2888 6512 2929 6546
rect 2963 6512 3004 6546
rect 3038 6512 3079 6546
rect 3113 6512 3154 6546
rect 3188 6512 3229 6546
rect 3263 6512 3353 6546
rect 2549 6475 3353 6512
rect 4092 6560 4174 6594
rect 4058 6510 4208 6560
rect 4092 6476 4174 6510
rect 4411 6565 4446 6599
rect 4480 6565 4518 6599
rect 4552 6565 4590 6599
rect 4624 6565 4662 6599
rect 4696 6565 4731 6599
rect 4411 6531 4731 6565
rect 4411 6497 4446 6531
rect 4480 6497 4518 6531
rect 4552 6497 4590 6531
rect 4624 6497 4662 6531
rect 4696 6497 4731 6531
rect 2549 6472 3270 6475
rect -874 6441 -849 6445
rect -815 6441 925 6445
rect -874 6409 925 6441
rect -874 6375 -850 6409
rect -816 6395 -781 6409
rect -815 6375 -781 6395
rect -747 6375 -712 6409
rect -678 6375 -643 6409
rect -609 6375 -574 6409
rect -540 6375 -505 6409
rect -471 6375 -436 6409
rect -402 6375 -367 6409
rect -333 6375 -298 6409
rect -264 6375 -229 6409
rect -195 6375 -160 6409
rect -126 6375 -91 6409
rect -57 6375 -22 6409
rect 12 6375 47 6409
rect 81 6375 116 6409
rect 150 6375 185 6409
rect 219 6375 254 6409
rect 288 6375 323 6409
rect 357 6375 391 6409
rect 425 6375 459 6409
rect 493 6375 527 6409
rect 561 6375 595 6409
rect 629 6375 663 6409
rect 697 6375 731 6409
rect 765 6375 799 6409
rect 833 6375 867 6409
rect 901 6375 925 6409
rect 2549 6438 2551 6472
rect 2585 6438 2627 6472
rect 2661 6438 2703 6472
rect 2737 6438 2779 6472
rect 2813 6438 2854 6472
rect 2888 6438 2929 6472
rect 2963 6438 3004 6472
rect 3038 6438 3079 6472
rect 3113 6438 3154 6472
rect 3188 6438 3229 6472
rect 3263 6438 3270 6472
rect 2549 6398 3270 6438
rect 2549 6379 2551 6398
rect -874 6361 -849 6375
rect -815 6361 925 6375
rect -874 6339 925 6361
rect -874 6305 -850 6339
rect -816 6315 -781 6339
rect -815 6305 -781 6315
rect -747 6305 -712 6339
rect -678 6305 -643 6339
rect -609 6305 -574 6339
rect -540 6305 -505 6339
rect -471 6305 -436 6339
rect -402 6305 -367 6339
rect -333 6305 -298 6339
rect -264 6305 -229 6339
rect -195 6305 -160 6339
rect -126 6305 -91 6339
rect -57 6305 -22 6339
rect 12 6305 47 6339
rect 81 6305 116 6339
rect 150 6305 185 6339
rect 219 6305 254 6339
rect 288 6305 323 6339
rect 357 6305 391 6339
rect 425 6305 459 6339
rect 493 6305 527 6339
rect 561 6305 595 6339
rect 629 6305 663 6339
rect 697 6305 731 6339
rect 765 6305 799 6339
rect 833 6305 867 6339
rect 901 6305 925 6339
rect -874 6281 -849 6305
rect -815 6281 925 6305
rect -874 6269 925 6281
rect -874 6235 -850 6269
rect -816 6235 -781 6269
rect -747 6235 -712 6269
rect -678 6235 -643 6269
rect -609 6235 -574 6269
rect -540 6235 -505 6269
rect -471 6235 -436 6269
rect -402 6235 -367 6269
rect -333 6235 -298 6269
rect -264 6235 -229 6269
rect -195 6235 -160 6269
rect -126 6235 -91 6269
rect -57 6235 -22 6269
rect 12 6235 47 6269
rect 81 6235 116 6269
rect 150 6235 185 6269
rect 219 6235 254 6269
rect 288 6235 323 6269
rect 357 6235 391 6269
rect 425 6235 459 6269
rect 493 6235 527 6269
rect 561 6235 595 6269
rect 629 6235 663 6269
rect 697 6235 731 6269
rect 765 6235 799 6269
rect 833 6235 867 6269
rect 901 6235 925 6269
rect 1053 6345 1135 6379
rect 1019 6295 1169 6345
rect 1053 6261 1135 6295
rect 1969 6364 2551 6379
rect 2585 6364 2627 6398
rect 2661 6364 2703 6398
rect 2737 6364 2779 6398
rect 2813 6364 2854 6398
rect 2888 6364 2929 6398
rect 2963 6364 3004 6398
rect 3038 6364 3079 6398
rect 3113 6364 3154 6398
rect 3188 6364 3229 6398
rect 3263 6364 3270 6398
rect 1969 6324 3270 6364
rect 1969 6290 2551 6324
rect 2585 6290 2627 6324
rect 2661 6290 2703 6324
rect 2737 6290 2779 6324
rect 2813 6290 2854 6324
rect 2888 6290 2929 6324
rect 2963 6290 3004 6324
rect 3038 6290 3079 6324
rect 3113 6290 3154 6324
rect 3188 6290 3229 6324
rect 3263 6290 3270 6324
rect -874 6234 925 6235
rect -874 6200 -849 6234
rect -815 6200 925 6234
rect -874 6199 925 6200
rect -874 6165 -850 6199
rect -816 6165 -781 6199
rect -747 6165 -712 6199
rect -678 6165 -643 6199
rect -609 6165 -574 6199
rect -540 6165 -505 6199
rect -471 6165 -436 6199
rect -402 6165 -367 6199
rect -333 6165 -298 6199
rect -264 6165 -229 6199
rect -195 6165 -160 6199
rect -126 6165 -91 6199
rect -57 6165 -22 6199
rect 12 6165 47 6199
rect 81 6165 116 6199
rect 150 6165 185 6199
rect 219 6165 254 6199
rect 288 6165 323 6199
rect 357 6165 391 6199
rect 425 6165 459 6199
rect 493 6165 527 6199
rect 561 6165 595 6199
rect 629 6165 663 6199
rect 697 6165 731 6199
rect 765 6165 799 6199
rect 833 6165 867 6199
rect 901 6165 925 6199
rect -874 6153 925 6165
rect -874 6129 -849 6153
rect -815 6129 925 6153
rect -874 6095 -850 6129
rect -815 6119 -781 6129
rect -816 6095 -781 6119
rect -747 6095 -712 6129
rect -678 6095 -643 6129
rect -609 6095 -574 6129
rect -540 6095 -505 6129
rect -471 6095 -436 6129
rect -402 6095 -367 6129
rect -333 6095 -298 6129
rect -264 6095 -229 6129
rect -195 6095 -160 6129
rect -126 6095 -91 6129
rect -57 6095 -22 6129
rect 12 6095 47 6129
rect 81 6095 116 6129
rect 150 6095 185 6129
rect 219 6095 254 6129
rect 288 6095 323 6129
rect 357 6095 391 6129
rect 425 6095 459 6129
rect 493 6095 527 6129
rect 561 6095 595 6129
rect 629 6095 663 6129
rect 697 6095 731 6129
rect 765 6095 799 6129
rect 833 6095 867 6129
rect 901 6095 925 6129
rect -874 6088 925 6095
rect 1969 6250 3270 6290
rect 1969 6216 2551 6250
rect 2585 6216 2627 6250
rect 2661 6216 2703 6250
rect 2737 6216 2779 6250
rect 2813 6216 2854 6250
rect 2888 6216 2929 6250
rect 2963 6216 3004 6250
rect 3038 6216 3079 6250
rect 3113 6216 3154 6250
rect 3188 6216 3229 6250
rect 3263 6216 3270 6250
rect 1969 5975 3270 6216
rect 4411 6463 4731 6497
rect 4411 6429 4446 6463
rect 4480 6429 4518 6463
rect 4552 6429 4590 6463
rect 4624 6429 4662 6463
rect 4696 6429 4731 6463
rect 4411 6395 4731 6429
rect 4411 6361 4446 6395
rect 4480 6361 4518 6395
rect 4552 6361 4590 6395
rect 4624 6361 4662 6395
rect 4696 6361 4731 6395
rect 4411 6327 4731 6361
rect 4411 6293 4446 6327
rect 4480 6293 4518 6327
rect 4552 6293 4590 6327
rect 4624 6293 4662 6327
rect 4696 6293 4731 6327
rect 4411 6259 4731 6293
rect 4411 6225 4446 6259
rect 4480 6225 4518 6259
rect 4552 6225 4590 6259
rect 4624 6225 4662 6259
rect 4696 6225 4731 6259
rect 4411 6191 4731 6225
rect 4092 6127 4174 6161
rect 4058 6077 4208 6127
rect 4092 6043 4174 6077
rect 4411 6157 4446 6191
rect 4480 6157 4518 6191
rect 4552 6157 4590 6191
rect 4624 6157 4662 6191
rect 4696 6157 4731 6191
rect 4411 6123 4731 6157
rect 4411 6089 4446 6123
rect 4480 6089 4518 6123
rect 4552 6089 4590 6123
rect 4624 6089 4662 6123
rect 4696 6089 4731 6123
rect 4411 6055 4731 6089
rect 4411 6021 4446 6055
rect 4480 6021 4518 6055
rect 4552 6021 4590 6055
rect 4624 6021 4662 6055
rect 4696 6021 4731 6055
rect 4411 5987 4731 6021
rect 4411 5953 4446 5987
rect 4480 5953 4518 5987
rect 4552 5953 4590 5987
rect 4624 5953 4662 5987
rect 4696 5953 4731 5987
rect 4411 5919 4731 5953
rect 2845 5844 3988 5915
rect 3821 4203 3988 5844
rect 4411 5885 4446 5919
rect 4480 5885 4518 5919
rect 4552 5885 4590 5919
rect 4624 5885 4662 5919
rect 4696 5885 4731 5919
rect 4411 5850 4731 5885
rect 4411 5816 4446 5850
rect 4480 5816 4518 5850
rect 4552 5816 4590 5850
rect 4624 5816 4662 5850
rect 4696 5816 4731 5850
rect 4411 5779 4731 5816
rect 4067 5745 4102 5779
rect 4136 5745 4172 5779
rect 4206 5745 4242 5779
rect 4276 5745 4312 5779
rect 4346 5745 4382 5779
rect 4416 5745 4452 5779
rect 4486 5745 4522 5779
rect 4556 5745 4592 5779
rect 4626 5745 4662 5779
rect 4696 5745 4731 5779
rect 4067 5710 4731 5745
rect 4067 5676 4102 5710
rect 4136 5676 4172 5710
rect 4206 5676 4242 5710
rect 4276 5676 4312 5710
rect 4346 5676 4382 5710
rect 4416 5676 4452 5710
rect 4486 5676 4522 5710
rect 4556 5676 4592 5710
rect 4626 5676 4662 5710
rect 4696 5676 4731 5710
rect 4067 5641 4731 5676
rect 4067 5607 4102 5641
rect 4136 5607 4172 5641
rect 4206 5607 4242 5641
rect 4276 5607 4312 5641
rect 4346 5607 4382 5641
rect 4416 5607 4452 5641
rect 4486 5607 4522 5641
rect 4556 5607 4592 5641
rect 4626 5607 4662 5641
rect 4696 5607 4731 5641
rect 4067 5572 4731 5607
rect 4067 5538 4102 5572
rect 4136 5538 4172 5572
rect 4206 5538 4242 5572
rect 4276 5538 4312 5572
rect 4346 5538 4382 5572
rect 4416 5538 4452 5572
rect 4486 5538 4522 5572
rect 4556 5538 4592 5572
rect 4626 5538 4662 5572
rect 4696 5538 4731 5572
rect 4067 5503 4731 5538
rect 4067 5469 4102 5503
rect 4136 5469 4172 5503
rect 4206 5469 4242 5503
rect 4276 5469 4312 5503
rect 4346 5469 4382 5503
rect 4416 5469 4452 5503
rect 4486 5469 4522 5503
rect 4556 5469 4592 5503
rect 4626 5469 4662 5503
rect 4696 5469 4731 5503
rect 4067 5434 4731 5469
rect 4067 5400 4102 5434
rect 4136 5400 4172 5434
rect 4206 5400 4242 5434
rect 4276 5400 4312 5434
rect 4346 5400 4382 5434
rect 4416 5400 4452 5434
rect 4486 5400 4522 5434
rect 4556 5400 4592 5434
rect 4626 5400 4662 5434
rect 4696 5400 4731 5434
rect 4067 5365 4731 5400
rect 4067 5331 4102 5365
rect 4136 5331 4172 5365
rect 4206 5331 4242 5365
rect 4276 5331 4312 5365
rect 4346 5331 4382 5365
rect 4416 5331 4452 5365
rect 4486 5331 4522 5365
rect 4556 5335 4592 5365
rect 4626 5335 4662 5365
rect 4556 5331 4579 5335
rect 4626 5331 4651 5335
rect 4696 5331 4731 5365
rect 4067 5301 4579 5331
rect 4613 5301 4651 5331
rect 4685 5301 4731 5331
rect 4067 5296 4731 5301
rect 4067 5262 4102 5296
rect 4136 5262 4172 5296
rect 4206 5262 4242 5296
rect 4276 5262 4312 5296
rect 4346 5262 4382 5296
rect 4416 5262 4452 5296
rect 4486 5262 4522 5296
rect 4556 5262 4592 5296
rect 4626 5262 4662 5296
rect 4696 5262 4731 5296
rect 4067 5245 4731 5262
rect 4067 5227 4466 5245
rect 4500 5227 4556 5245
rect 4067 5193 4102 5227
rect 4136 5193 4172 5227
rect 4206 5193 4242 5227
rect 4276 5193 4312 5227
rect 4346 5193 4382 5227
rect 4416 5193 4452 5227
rect 4500 5211 4522 5227
rect 4486 5193 4522 5211
rect 4590 5227 4646 5245
rect 4680 5227 4731 5245
rect 4590 5211 4592 5227
rect 4556 5193 4592 5211
rect 4626 5211 4646 5227
rect 4626 5193 4662 5211
rect 4696 5193 4731 5227
rect 4067 5171 4731 5193
rect 4067 5158 4466 5171
rect 4500 5158 4556 5171
rect 4067 5124 4102 5158
rect 4136 5124 4172 5158
rect 4206 5124 4242 5158
rect 4276 5124 4312 5158
rect 4346 5124 4382 5158
rect 4416 5124 4452 5158
rect 4500 5137 4522 5158
rect 4486 5124 4522 5137
rect 4590 5158 4646 5171
rect 4680 5158 4731 5171
rect 4590 5137 4592 5158
rect 4556 5124 4592 5137
rect 4626 5137 4646 5158
rect 4626 5124 4662 5137
rect 4696 5124 4731 5158
rect 4067 5097 4731 5124
rect 4067 5089 4466 5097
rect 4500 5089 4556 5097
rect 4067 5055 4102 5089
rect 4136 5055 4172 5089
rect 4206 5055 4242 5089
rect 4276 5055 4312 5089
rect 4346 5055 4382 5089
rect 4416 5055 4452 5089
rect 4500 5063 4522 5089
rect 4486 5055 4522 5063
rect 4590 5089 4646 5097
rect 4680 5089 4731 5097
rect 4590 5063 4592 5089
rect 4556 5055 4592 5063
rect 4626 5063 4646 5089
rect 4626 5055 4662 5063
rect 4696 5055 4731 5089
rect 4067 5023 4731 5055
rect 4067 5019 4466 5023
rect 4500 5019 4556 5023
rect 4067 4985 4102 5019
rect 4136 4985 4172 5019
rect 4206 4985 4242 5019
rect 4276 4985 4312 5019
rect 4346 4985 4382 5019
rect 4416 4985 4452 5019
rect 4500 4989 4522 5019
rect 4486 4985 4522 4989
rect 4590 5019 4646 5023
rect 4680 5019 4731 5023
rect 4590 4989 4592 5019
rect 4556 4985 4592 4989
rect 4626 4989 4646 5019
rect 4626 4985 4662 4989
rect 4696 4985 4731 5019
rect 4067 4949 4731 4985
rect 4067 4915 4102 4949
rect 4136 4915 4172 4949
rect 4206 4915 4242 4949
rect 4276 4915 4312 4949
rect 4346 4915 4382 4949
rect 4416 4915 4452 4949
rect 4500 4915 4522 4949
rect 4590 4915 4592 4949
rect 4626 4915 4646 4949
rect 4696 4915 4731 4949
rect 4067 4879 4731 4915
rect 4067 4845 4102 4879
rect 4136 4845 4172 4879
rect 4206 4845 4242 4879
rect 4276 4845 4312 4879
rect 4346 4845 4382 4879
rect 4416 4845 4452 4879
rect 4486 4875 4522 4879
rect 4500 4845 4522 4875
rect 4556 4875 4592 4879
rect 4067 4841 4466 4845
rect 4500 4841 4556 4845
rect 4590 4845 4592 4875
rect 4626 4875 4662 4879
rect 4626 4845 4646 4875
rect 4696 4845 4731 4879
rect 4590 4841 4646 4845
rect 4680 4841 4731 4845
rect 4067 4809 4731 4841
rect 4067 4775 4102 4809
rect 4136 4775 4172 4809
rect 4206 4775 4242 4809
rect 4276 4775 4312 4809
rect 4346 4775 4382 4809
rect 4416 4775 4452 4809
rect 4486 4801 4522 4809
rect 4500 4775 4522 4801
rect 4556 4801 4592 4809
rect 4067 4767 4466 4775
rect 4500 4767 4556 4775
rect 4590 4775 4592 4801
rect 4626 4801 4662 4809
rect 4626 4775 4646 4801
rect 4696 4775 4731 4809
rect 4590 4767 4646 4775
rect 4680 4767 4731 4775
rect 4067 4739 4731 4767
rect 4067 4705 4102 4739
rect 4136 4705 4172 4739
rect 4206 4705 4242 4739
rect 4276 4705 4312 4739
rect 4346 4705 4382 4739
rect 4416 4705 4452 4739
rect 4486 4727 4522 4739
rect 4500 4705 4522 4727
rect 4556 4727 4592 4739
rect 4067 4693 4466 4705
rect 4500 4693 4556 4705
rect 4590 4705 4592 4727
rect 4626 4727 4662 4739
rect 4626 4705 4646 4727
rect 4696 4705 4731 4739
rect 4590 4693 4646 4705
rect 4680 4693 4731 4705
rect 4067 4669 4731 4693
rect 4067 4635 4102 4669
rect 4136 4635 4172 4669
rect 4206 4635 4242 4669
rect 4276 4635 4312 4669
rect 4346 4635 4382 4669
rect 4416 4635 4452 4669
rect 4486 4635 4522 4669
rect 4556 4635 4592 4669
rect 4626 4635 4662 4669
rect 4696 4635 4731 4669
rect 4067 4626 4731 4635
rect 4067 4599 4579 4626
rect 4613 4599 4651 4626
rect 4685 4599 4731 4626
rect 4067 4565 4102 4599
rect 4136 4565 4172 4599
rect 4206 4565 4242 4599
rect 4276 4565 4312 4599
rect 4346 4565 4382 4599
rect 4416 4565 4452 4599
rect 4486 4565 4522 4599
rect 4556 4592 4579 4599
rect 4626 4592 4651 4599
rect 4556 4565 4592 4592
rect 4626 4565 4662 4592
rect 4696 4565 4731 4599
rect 4067 4529 4731 4565
rect 4067 4495 4102 4529
rect 4136 4495 4172 4529
rect 4206 4495 4242 4529
rect 4276 4495 4312 4529
rect 4346 4495 4382 4529
rect 4416 4495 4452 4529
rect 4486 4495 4522 4529
rect 4556 4495 4592 4529
rect 4626 4495 4662 4529
rect 4696 4495 4731 4529
rect 4067 4459 4731 4495
rect 4067 4425 4102 4459
rect 4136 4425 4172 4459
rect 4206 4425 4242 4459
rect 4276 4425 4312 4459
rect 4346 4425 4382 4459
rect 4416 4425 4452 4459
rect 4486 4425 4522 4459
rect 4556 4425 4592 4459
rect 4626 4425 4662 4459
rect 4696 4425 4731 4459
rect 4067 4389 4731 4425
rect 4067 4355 4102 4389
rect 4136 4355 4172 4389
rect 4206 4355 4242 4389
rect 4276 4355 4312 4389
rect 4346 4355 4382 4389
rect 4416 4355 4452 4389
rect 4486 4355 4522 4389
rect 4556 4355 4592 4389
rect 4626 4355 4662 4389
rect 4696 4355 4731 4389
rect 4067 4319 4731 4355
rect 4067 4285 4102 4319
rect 4136 4285 4172 4319
rect 4206 4285 4242 4319
rect 4276 4285 4312 4319
rect 4346 4285 4382 4319
rect 4416 4285 4452 4319
rect 4486 4285 4522 4319
rect 4556 4285 4592 4319
rect 4626 4285 4662 4319
rect 4696 4285 4731 4319
rect 4067 4249 4731 4285
rect 4067 4215 4102 4249
rect 4136 4215 4172 4249
rect 4206 4215 4242 4249
rect 4276 4215 4312 4249
rect 4346 4215 4382 4249
rect 4416 4215 4452 4249
rect 4486 4215 4522 4249
rect 4556 4215 4592 4249
rect 4626 4215 4662 4249
rect 4696 4216 4731 4249
rect 13193 4314 13239 4326
rect 13193 4280 13205 4314
rect 13193 4242 13239 4280
rect 13193 4240 13205 4242
rect 4696 4215 8292 4216
rect 4067 4182 8292 4215
rect 4067 4179 4731 4182
rect 4067 4145 4102 4179
rect 4136 4145 4172 4179
rect 4206 4145 4242 4179
rect 4276 4145 4312 4179
rect 4346 4145 4382 4179
rect 4416 4145 4452 4179
rect 4486 4145 4522 4179
rect 4556 4145 4592 4179
rect 4626 4145 4662 4179
rect 4696 4148 4731 4179
rect 4765 4148 4801 4182
rect 4835 4148 4871 4182
rect 4905 4148 4941 4182
rect 4975 4148 5011 4182
rect 5045 4148 5081 4182
rect 5115 4148 5151 4182
rect 5185 4148 5221 4182
rect 5255 4148 5291 4182
rect 5325 4148 5360 4182
rect 5394 4148 5429 4182
rect 5463 4148 5498 4182
rect 5532 4148 5567 4182
rect 5601 4148 5636 4182
rect 5670 4148 5705 4182
rect 5739 4148 5774 4182
rect 5808 4148 5843 4182
rect 5877 4148 5912 4182
rect 5946 4148 5981 4182
rect 6015 4148 6050 4182
rect 6084 4148 6119 4182
rect 6153 4148 6188 4182
rect 6222 4148 6257 4182
rect 6291 4148 6326 4182
rect 6360 4148 6395 4182
rect 6429 4148 6464 4182
rect 6498 4148 6533 4182
rect 6567 4148 6602 4182
rect 6636 4148 6671 4182
rect 6705 4148 6740 4182
rect 6774 4148 6809 4182
rect 6843 4148 6878 4182
rect 6912 4148 6947 4182
rect 6981 4148 7016 4182
rect 7050 4148 7085 4182
rect 7119 4148 7154 4182
rect 7188 4148 7223 4182
rect 7257 4148 7292 4182
rect 7326 4148 7361 4182
rect 7395 4148 7430 4182
rect 7464 4148 7499 4182
rect 7533 4148 7568 4182
rect 7602 4148 7637 4182
rect 7671 4148 7706 4182
rect 7740 4148 7775 4182
rect 7809 4148 7844 4182
rect 7878 4148 7913 4182
rect 7947 4148 7982 4182
rect 8016 4148 8051 4182
rect 8085 4148 8120 4182
rect 8154 4148 8189 4182
rect 8223 4148 8258 4182
rect 4696 4145 8292 4148
rect 4067 4109 8292 4145
rect 4067 4075 4102 4109
rect 4136 4075 4172 4109
rect 4206 4075 4242 4109
rect 4276 4075 4312 4109
rect 4346 4075 4382 4109
rect 4416 4075 4452 4109
rect 4486 4075 4522 4109
rect 4556 4075 4592 4109
rect 4626 4075 4662 4109
rect 4696 4084 8292 4109
rect 4696 4075 4731 4084
rect 4067 4050 4731 4075
rect 4765 4050 4801 4084
rect 4835 4050 4871 4084
rect 4905 4050 4941 4084
rect 4975 4050 5011 4084
rect 5045 4050 5081 4084
rect 5115 4050 5151 4084
rect 5185 4050 5221 4084
rect 5255 4050 5291 4084
rect 5325 4050 5360 4084
rect 5394 4050 5429 4084
rect 5463 4050 5498 4084
rect 5532 4050 5567 4084
rect 5601 4050 5636 4084
rect 5670 4050 5705 4084
rect 5739 4050 5774 4084
rect 5808 4050 5843 4084
rect 5877 4050 5912 4084
rect 5946 4050 5981 4084
rect 6015 4050 6050 4084
rect 6084 4050 6119 4084
rect 6153 4050 6188 4084
rect 6222 4050 6257 4084
rect 6291 4050 6326 4084
rect 6360 4050 6395 4084
rect 6429 4050 6464 4084
rect 6498 4050 6533 4084
rect 6567 4050 6602 4084
rect 6636 4050 6671 4084
rect 6705 4050 6740 4084
rect 6774 4050 6809 4084
rect 6843 4050 6878 4084
rect 6912 4050 6947 4084
rect 6981 4050 7016 4084
rect 7050 4050 7085 4084
rect 7119 4050 7154 4084
rect 7188 4050 7223 4084
rect 7257 4050 7292 4084
rect 7326 4050 7361 4084
rect 7395 4050 7430 4084
rect 7464 4050 7499 4084
rect 7533 4050 7568 4084
rect 7602 4050 7637 4084
rect 7671 4050 7706 4084
rect 7740 4050 7775 4084
rect 7809 4050 7844 4084
rect 7878 4050 7913 4084
rect 7947 4050 7982 4084
rect 8016 4050 8051 4084
rect 8085 4050 8120 4084
rect 8154 4050 8189 4084
rect 8223 4050 8258 4084
rect 4067 4039 8292 4050
rect 4067 4005 4102 4039
rect 4136 4005 4172 4039
rect 4206 4005 4242 4039
rect 4276 4005 4312 4039
rect 4346 4005 4382 4039
rect 4416 4005 4452 4039
rect 4486 4005 4522 4039
rect 4556 4005 4592 4039
rect 4626 4005 4662 4039
rect 4696 4016 8292 4039
rect 13227 4206 13239 4208
rect 13193 4172 13239 4206
rect 14983 4314 15017 4326
rect 14983 4241 15017 4268
rect 13227 4170 13239 4172
rect 13193 4136 13205 4138
rect 13193 4104 13239 4136
rect 13227 4098 13239 4104
rect 13193 4064 13205 4070
rect 13193 4036 13239 4064
rect 13227 4026 13239 4036
rect 4696 4013 9456 4016
rect 4696 4005 4974 4013
rect 4067 3979 4974 4005
rect 5008 3979 5043 4013
rect 5077 3979 5112 4013
rect 5146 3979 5181 4013
rect 5215 3979 5250 4013
rect 5284 3979 5319 4013
rect 5353 3979 5388 4013
rect 5422 3979 5457 4013
rect 5491 3979 5526 4013
rect 5560 3979 5595 4013
rect 5629 3979 5664 4013
rect 5698 3979 5733 4013
rect 5767 3979 5802 4013
rect 5836 3979 5871 4013
rect 5905 3979 5940 4013
rect 5974 3979 6009 4013
rect 6043 3979 6078 4013
rect 6112 3979 6147 4013
rect 6181 3979 6216 4013
rect 6250 3979 6285 4013
rect 6319 3979 6354 4013
rect 6388 3979 6423 4013
rect 6457 3979 6492 4013
rect 6526 3979 6561 4013
rect 6595 3979 6630 4013
rect 6664 3979 6699 4013
rect 6733 3979 6768 4013
rect 6802 3979 6837 4013
rect 6871 3979 6906 4013
rect 6940 3979 6975 4013
rect 7009 3979 7044 4013
rect 7078 3979 7113 4013
rect 7147 3979 7182 4013
rect 7216 3979 7251 4013
rect 7285 3979 7320 4013
rect 7354 3979 7389 4013
rect 7423 3979 7458 4013
rect 7492 3979 7527 4013
rect 7561 3979 7596 4013
rect 7630 3979 7665 4013
rect 7699 3979 7734 4013
rect 7768 3979 7803 4013
rect 7837 3979 7872 4013
rect 7906 3979 7941 4013
rect 7975 3979 8010 4013
rect 8044 3979 8079 4013
rect 8113 3979 8148 4013
rect 8182 3979 8217 4013
rect 8251 3979 8286 4013
rect 8320 3979 8355 4013
rect 8389 3979 8424 4013
rect 8458 3979 8493 4013
rect 8527 3979 8562 4013
rect 8596 3979 8631 4013
rect 8665 3979 8700 4013
rect 8734 3979 8769 4013
rect 8803 3979 8838 4013
rect 8872 3979 8907 4013
rect 8941 3979 8976 4013
rect 9010 3979 9045 4013
rect 9079 3979 9114 4013
rect 9148 3979 9183 4013
rect 9217 3979 9252 4013
rect 9286 3979 9320 4013
rect 9354 3979 9388 4013
rect 9422 3979 9456 4013
rect 4067 3969 9456 3979
rect 4067 3935 4102 3969
rect 4136 3935 4172 3969
rect 4206 3935 4242 3969
rect 4276 3935 4312 3969
rect 4346 3935 4382 3969
rect 4416 3935 4452 3969
rect 4486 3935 4522 3969
rect 4556 3935 4592 3969
rect 4626 3935 4662 3969
rect 4696 3937 9456 3969
rect 4696 3935 4974 3937
rect 4067 3925 4974 3935
rect 3864 3903 4974 3925
rect 5008 3903 5043 3937
rect 5077 3903 5112 3937
rect 5146 3903 5181 3937
rect 5215 3903 5250 3937
rect 5284 3903 5319 3937
rect 5353 3903 5388 3937
rect 5422 3903 5457 3937
rect 5491 3903 5526 3937
rect 5560 3903 5595 3937
rect 5629 3903 5664 3937
rect 5698 3903 5733 3937
rect 5767 3903 5802 3937
rect 5836 3903 5871 3937
rect 5905 3903 5940 3937
rect 5974 3903 6009 3937
rect 6043 3903 6078 3937
rect 6112 3903 6147 3937
rect 6181 3903 6216 3937
rect 6250 3903 6285 3937
rect 6319 3903 6354 3937
rect 6388 3903 6423 3937
rect 6457 3903 6492 3937
rect 6526 3903 6561 3937
rect 6595 3903 6630 3937
rect 6664 3903 6699 3937
rect 6733 3903 6768 3937
rect 6802 3903 6837 3937
rect 6871 3903 6906 3937
rect 6940 3903 6975 3937
rect 7009 3903 7044 3937
rect 7078 3903 7113 3937
rect 7147 3903 7182 3937
rect 7216 3903 7251 3937
rect 7285 3903 7320 3937
rect 7354 3903 7389 3937
rect 7423 3903 7458 3937
rect 7492 3903 7527 3937
rect 7561 3903 7596 3937
rect 7630 3903 7665 3937
rect 7699 3903 7734 3937
rect 7768 3903 7803 3937
rect 7837 3903 7872 3937
rect 7906 3903 7941 3937
rect 7975 3903 8010 3937
rect 8044 3903 8079 3937
rect 8113 3903 8148 3937
rect 8182 3903 8217 3937
rect 8251 3903 8286 3937
rect 8320 3903 8355 3937
rect 8389 3903 8424 3937
rect 8458 3903 8493 3937
rect 8527 3903 8562 3937
rect 8596 3903 8631 3937
rect 8665 3903 8700 3937
rect 8734 3903 8769 3937
rect 8803 3903 8838 3937
rect 8872 3903 8907 3937
rect 8941 3903 8976 3937
rect 9010 3903 9045 3937
rect 9079 3903 9114 3937
rect 9148 3903 9183 3937
rect 9217 3903 9252 3937
rect 9286 3903 9320 3937
rect 9354 3903 9388 3937
rect 9422 3903 9456 3937
rect 3864 3901 9456 3903
rect 3864 2167 3875 3901
rect 4929 3861 9456 3901
rect 11498 3984 11538 4018
rect 11572 3984 11612 4018
rect 11646 3984 11686 4018
rect 11720 3984 11760 4018
rect 11794 3984 11834 4018
rect 11464 3902 11868 3984
rect 11498 3868 11538 3902
rect 11572 3868 11612 3902
rect 11646 3868 11686 3902
rect 11720 3868 11760 3902
rect 11794 3868 11834 3902
rect 11998 3984 12038 4018
rect 12072 3984 12112 4018
rect 12146 3984 12186 4018
rect 12220 3984 12260 4018
rect 12294 3984 12334 4018
rect 11964 3902 12368 3984
rect 11998 3868 12038 3902
rect 12072 3868 12112 3902
rect 12146 3868 12186 3902
rect 12220 3868 12260 3902
rect 12294 3868 12334 3902
rect 12499 3984 12539 4018
rect 12573 3984 12613 4018
rect 12647 3984 12687 4018
rect 12721 3984 12761 4018
rect 12795 3984 12835 4018
rect 12465 3902 12869 3984
rect 12499 3868 12539 3902
rect 12573 3868 12613 3902
rect 12647 3868 12687 3902
rect 12721 3868 12761 3902
rect 12795 3868 12835 3902
rect 13193 3992 13205 4002
rect 13193 3968 13239 3992
rect 13227 3954 13239 3968
rect 13193 3920 13205 3934
rect 13193 3900 13239 3920
rect 13227 3882 13239 3900
rect 4929 3827 4974 3861
rect 5008 3827 5043 3861
rect 5077 3827 5112 3861
rect 5146 3827 5181 3861
rect 5215 3827 5250 3861
rect 5284 3827 5319 3861
rect 5353 3827 5388 3861
rect 5422 3827 5457 3861
rect 5491 3827 5526 3861
rect 5560 3827 5595 3861
rect 5629 3827 5664 3861
rect 5698 3827 5733 3861
rect 5767 3827 5802 3861
rect 5836 3827 5871 3861
rect 5905 3827 5940 3861
rect 5974 3827 6009 3861
rect 6043 3827 6078 3861
rect 6112 3827 6147 3861
rect 6181 3827 6216 3861
rect 6250 3827 6285 3861
rect 6319 3827 6354 3861
rect 6388 3827 6423 3861
rect 6457 3827 6492 3861
rect 6526 3827 6561 3861
rect 6595 3827 6630 3861
rect 6664 3827 6699 3861
rect 6733 3827 6768 3861
rect 6802 3827 6837 3861
rect 6871 3827 6906 3861
rect 6940 3827 6975 3861
rect 7009 3827 7044 3861
rect 7078 3827 7113 3861
rect 7147 3827 7182 3861
rect 7216 3827 7251 3861
rect 7285 3827 7320 3861
rect 7354 3827 7389 3861
rect 7423 3827 7458 3861
rect 7492 3827 7527 3861
rect 7561 3827 7596 3861
rect 7630 3827 7665 3861
rect 7699 3827 7734 3861
rect 7768 3827 7803 3861
rect 7837 3827 7872 3861
rect 7906 3827 7941 3861
rect 7975 3827 8010 3861
rect 8044 3827 8079 3861
rect 8113 3827 8148 3861
rect 8182 3827 8217 3861
rect 8251 3827 8286 3861
rect 8320 3827 8355 3861
rect 8389 3827 8424 3861
rect 8458 3827 8493 3861
rect 8527 3827 8562 3861
rect 8596 3827 8631 3861
rect 8665 3827 8700 3861
rect 8734 3827 8769 3861
rect 8803 3827 8838 3861
rect 8872 3827 8907 3861
rect 8941 3827 8976 3861
rect 9010 3827 9045 3861
rect 9079 3827 9114 3861
rect 9148 3827 9183 3861
rect 9217 3827 9252 3861
rect 9286 3827 9320 3861
rect 9354 3827 9388 3861
rect 9422 3827 9456 3861
rect 4929 3785 9456 3827
rect 4929 3751 4974 3785
rect 5008 3751 5043 3785
rect 5077 3751 5112 3785
rect 5146 3751 5181 3785
rect 5215 3751 5250 3785
rect 5284 3751 5319 3785
rect 5353 3751 5388 3785
rect 5422 3751 5457 3785
rect 5491 3751 5526 3785
rect 5560 3751 5595 3785
rect 5629 3751 5664 3785
rect 5698 3751 5733 3785
rect 5767 3751 5802 3785
rect 5836 3751 5871 3785
rect 5905 3751 5940 3785
rect 5974 3751 6009 3785
rect 6043 3751 6078 3785
rect 6112 3751 6147 3785
rect 6181 3751 6216 3785
rect 6250 3751 6285 3785
rect 6319 3751 6354 3785
rect 6388 3751 6423 3785
rect 6457 3751 6492 3785
rect 6526 3751 6561 3785
rect 6595 3751 6630 3785
rect 6664 3751 6699 3785
rect 6733 3751 6768 3785
rect 6802 3751 6837 3785
rect 6871 3751 6906 3785
rect 6940 3751 6975 3785
rect 7009 3751 7044 3785
rect 7078 3751 7113 3785
rect 7147 3751 7182 3785
rect 7216 3751 7251 3785
rect 7285 3751 7320 3785
rect 7354 3751 7389 3785
rect 7423 3751 7458 3785
rect 7492 3751 7527 3785
rect 7561 3751 7596 3785
rect 7630 3751 7665 3785
rect 7699 3751 7734 3785
rect 7768 3751 7803 3785
rect 7837 3751 7872 3785
rect 7906 3751 7941 3785
rect 7975 3751 8010 3785
rect 8044 3751 8079 3785
rect 8113 3751 8148 3785
rect 8182 3751 8217 3785
rect 8251 3751 8286 3785
rect 8320 3751 8355 3785
rect 8389 3751 8424 3785
rect 8458 3758 8493 3785
rect 8527 3758 8562 3785
rect 8596 3758 8631 3785
rect 8665 3758 8700 3785
rect 8734 3758 8769 3785
rect 8458 3751 8474 3758
rect 8527 3751 8547 3758
rect 8596 3751 8620 3758
rect 8665 3751 8693 3758
rect 8734 3751 8766 3758
rect 8803 3751 8838 3785
rect 8872 3758 8907 3785
rect 8941 3758 8976 3785
rect 9010 3758 9045 3785
rect 9079 3758 9114 3785
rect 9148 3758 9183 3785
rect 9217 3758 9252 3785
rect 9286 3758 9320 3785
rect 9354 3758 9388 3785
rect 8873 3751 8907 3758
rect 8946 3751 8976 3758
rect 9018 3751 9045 3758
rect 9090 3751 9114 3758
rect 9162 3751 9183 3758
rect 9234 3751 9252 3758
rect 9306 3751 9320 3758
rect 9378 3751 9388 3758
rect 9422 3751 9456 3785
rect 4929 3724 8474 3751
rect 8508 3724 8547 3751
rect 8581 3724 8620 3751
rect 8654 3724 8693 3751
rect 8727 3724 8766 3751
rect 8800 3724 8839 3751
rect 8873 3724 8912 3751
rect 8946 3724 8984 3751
rect 9018 3724 9056 3751
rect 9090 3724 9128 3751
rect 9162 3724 9200 3751
rect 9234 3724 9272 3751
rect 9306 3724 9344 3751
rect 9378 3724 9456 3751
rect 4929 3709 9456 3724
rect 4929 3675 4974 3709
rect 5008 3675 5043 3709
rect 5077 3675 5112 3709
rect 5146 3675 5181 3709
rect 5215 3675 5250 3709
rect 5284 3675 5319 3709
rect 5353 3675 5388 3709
rect 5422 3675 5457 3709
rect 5491 3675 5526 3709
rect 5560 3675 5595 3709
rect 5629 3675 5664 3709
rect 5698 3675 5733 3709
rect 5767 3675 5802 3709
rect 5836 3675 5871 3709
rect 5905 3675 5940 3709
rect 5974 3675 6009 3709
rect 6043 3675 6078 3709
rect 6112 3675 6147 3709
rect 6181 3675 6216 3709
rect 6250 3675 6285 3709
rect 6319 3675 6354 3709
rect 6388 3675 6423 3709
rect 6457 3675 6492 3709
rect 6526 3675 6561 3709
rect 6595 3675 6630 3709
rect 6664 3675 6699 3709
rect 6733 3675 6768 3709
rect 6802 3675 6837 3709
rect 6871 3675 6906 3709
rect 6940 3675 6975 3709
rect 7009 3675 7044 3709
rect 7078 3675 7113 3709
rect 7147 3675 7182 3709
rect 7216 3675 7251 3709
rect 7285 3675 7320 3709
rect 7354 3675 7389 3709
rect 7423 3675 7458 3709
rect 7492 3675 7527 3709
rect 7561 3675 7596 3709
rect 7630 3675 7665 3709
rect 7699 3675 7734 3709
rect 7768 3675 7803 3709
rect 7837 3675 7872 3709
rect 7906 3675 7941 3709
rect 7975 3675 8010 3709
rect 8044 3675 8079 3709
rect 8113 3675 8148 3709
rect 8182 3675 8217 3709
rect 8251 3675 8286 3709
rect 8320 3675 8355 3709
rect 8389 3675 8424 3709
rect 8458 3675 8493 3709
rect 8527 3675 8562 3709
rect 8596 3675 8631 3709
rect 8665 3675 8700 3709
rect 8734 3675 8769 3709
rect 8803 3675 8838 3709
rect 8872 3675 8907 3709
rect 8941 3675 8976 3709
rect 9010 3675 9045 3709
rect 9079 3675 9114 3709
rect 9148 3675 9183 3709
rect 9217 3675 9252 3709
rect 9286 3675 9320 3709
rect 9354 3675 9388 3709
rect 9422 3675 9456 3709
rect 4929 3672 9456 3675
rect 13193 3848 13205 3866
rect 13193 3832 13239 3848
rect 13227 3810 13239 3832
rect 13193 3776 13205 3798
rect 13193 3764 13239 3776
rect 13227 3738 13239 3764
rect 13193 3704 13205 3730
rect 13193 3696 13239 3704
rect 4929 3623 9400 3672
rect 13227 3666 13239 3696
rect 13193 3632 13205 3662
rect 13193 3628 13239 3632
rect 4929 3589 5176 3623
rect 13227 3594 13239 3628
rect 4929 2167 4940 3589
rect 13193 3560 13205 3594
rect 13227 3526 13239 3560
rect 13193 3522 13239 3526
rect 13193 3492 13205 3522
rect 13227 3458 13239 3488
rect 13193 3450 13239 3458
rect 13193 3424 13205 3450
rect 13227 3390 13239 3416
rect 13193 3378 13239 3390
rect 13193 3356 13205 3378
rect 13227 3322 13239 3344
rect 13193 3306 13239 3322
rect 13193 3288 13205 3306
rect 11498 3252 11537 3286
rect 11571 3252 11610 3286
rect 11644 3252 11683 3286
rect 11717 3252 11756 3286
rect 11790 3252 11828 3286
rect 11862 3252 11900 3286
rect 11934 3252 11972 3286
rect 12006 3252 12044 3286
rect 12078 3252 12116 3286
rect 12150 3252 12188 3286
rect 12222 3252 12260 3286
rect 12294 3252 12332 3286
rect 12366 3252 12404 3286
rect 12438 3252 12464 3286
rect 11464 3170 12464 3252
rect 11498 3136 11537 3170
rect 11571 3136 11610 3170
rect 11644 3136 11683 3170
rect 11717 3136 11756 3170
rect 11790 3136 11828 3170
rect 11862 3136 11900 3170
rect 11934 3136 11972 3170
rect 12006 3136 12044 3170
rect 12078 3136 12116 3170
rect 12150 3136 12188 3170
rect 12222 3136 12260 3170
rect 12294 3136 12332 3170
rect 12366 3136 12404 3170
rect 12438 3136 12464 3170
rect 12514 3252 12558 3286
rect 12592 3252 12635 3286
rect 12669 3252 12712 3286
rect 12746 3252 12789 3286
rect 12823 3252 12866 3286
rect 12480 3194 12900 3252
rect 12514 3160 12558 3194
rect 12592 3160 12635 3194
rect 12669 3160 12712 3194
rect 12746 3160 12789 3194
rect 12823 3160 12866 3194
rect 12480 3102 12900 3160
rect 12514 3068 12558 3102
rect 12592 3068 12635 3102
rect 12669 3068 12712 3102
rect 12746 3068 12789 3102
rect 12823 3068 12866 3102
rect 13227 3254 13239 3272
rect 13193 3234 13239 3254
rect 13193 3220 13205 3234
rect 13431 4180 14615 4186
rect 13431 4173 13509 4180
rect 13543 4173 13583 4180
rect 13617 4173 13657 4180
rect 13691 4173 13731 4180
rect 13765 4173 13805 4180
rect 13839 4173 13879 4180
rect 13913 4173 13953 4180
rect 13987 4173 14027 4180
rect 14061 4173 14101 4180
rect 14135 4173 14175 4180
rect 14209 4173 14249 4180
rect 14283 4173 14323 4180
rect 14357 4173 14397 4180
rect 14431 4173 14470 4180
rect 14504 4173 14543 4180
rect 13431 4139 13507 4173
rect 13543 4146 13575 4173
rect 13617 4146 13643 4173
rect 13691 4146 13711 4173
rect 13765 4146 13779 4173
rect 13839 4146 13847 4173
rect 13913 4146 13915 4173
rect 13541 4139 13575 4146
rect 13609 4139 13643 4146
rect 13677 4139 13711 4146
rect 13745 4139 13779 4146
rect 13813 4139 13847 4146
rect 13881 4139 13915 4146
rect 13949 4146 13953 4173
rect 14017 4146 14027 4173
rect 14085 4146 14101 4173
rect 14153 4146 14175 4173
rect 14221 4146 14249 4173
rect 13949 4139 13983 4146
rect 14017 4139 14051 4146
rect 14085 4139 14119 4146
rect 14153 4139 14187 4146
rect 14221 4139 14255 4146
rect 14289 4139 14323 4173
rect 14357 4139 14391 4173
rect 14431 4146 14459 4173
rect 14504 4146 14527 4173
rect 14577 4146 14615 4180
rect 14425 4139 14459 4146
rect 14493 4139 14527 4146
rect 14561 4139 14615 4146
rect 14983 4168 15017 4200
rect 13431 4107 13477 4139
rect 13431 4073 13437 4107
rect 13471 4073 13477 4107
rect 14983 4098 15017 4132
rect 13431 4050 13477 4073
rect 13603 4057 13619 4091
rect 13653 4057 13686 4091
rect 13730 4057 13768 4091
rect 13807 4057 13849 4091
rect 13884 4057 13925 4091
rect 13966 4057 13975 4091
rect 14151 4057 14167 4091
rect 14202 4057 14244 4091
rect 14283 4057 14321 4091
rect 14364 4057 14397 4091
rect 14445 4057 14473 4091
rect 13431 4034 13439 4050
rect 13431 4000 13437 4034
rect 13473 4016 13477 4050
rect 13471 4000 13477 4016
rect 13431 3982 13477 4000
rect 13431 3961 13439 3982
rect 13431 3927 13437 3961
rect 13473 3948 13477 3982
rect 14983 4030 15017 4061
rect 14983 3962 15017 3988
rect 13471 3927 13477 3948
rect 13431 3914 13477 3927
rect 13431 3888 13439 3914
rect 13431 3854 13437 3888
rect 13473 3880 13477 3914
rect 13471 3854 13477 3880
rect 13431 3846 13477 3854
rect 13431 3815 13439 3846
rect 13431 3781 13437 3815
rect 13473 3812 13477 3846
rect 13471 3781 13477 3812
rect 13431 3778 13477 3781
rect 13431 3744 13439 3778
rect 13473 3744 13477 3778
rect 13431 3742 13477 3744
rect 13431 3708 13437 3742
rect 13471 3710 13477 3742
rect 13431 3676 13439 3708
rect 13473 3676 13477 3710
rect 13431 3669 13477 3676
rect 13431 3635 13437 3669
rect 13471 3642 13477 3669
rect 13431 3608 13439 3635
rect 13473 3608 13477 3642
rect 13431 3596 13477 3608
rect 13431 3562 13437 3596
rect 13471 3574 13477 3596
rect 13431 3540 13439 3562
rect 13473 3540 13477 3574
rect 13431 3523 13477 3540
rect 13431 3489 13437 3523
rect 13471 3506 13477 3523
rect 13431 3472 13439 3489
rect 13473 3472 13477 3506
rect 13431 3450 13477 3472
rect 13431 3416 13437 3450
rect 13471 3438 13477 3450
rect 13431 3404 13439 3416
rect 13473 3404 13477 3438
rect 13558 3937 13592 3953
rect 13558 3869 13592 3882
rect 13558 3801 13592 3808
rect 13558 3665 13592 3699
rect 13558 3597 13592 3631
rect 13558 3529 13592 3563
rect 13558 3461 13592 3495
rect 13558 3411 13592 3427
rect 13714 3937 13748 3953
rect 13714 3869 13748 3882
rect 13714 3801 13748 3808
rect 13714 3665 13748 3699
rect 13714 3597 13748 3631
rect 13714 3529 13748 3563
rect 13714 3461 13748 3495
rect 13714 3411 13748 3427
rect 13830 3937 13864 3953
rect 13830 3869 13864 3903
rect 13830 3801 13864 3835
rect 13830 3733 13864 3767
rect 13830 3672 13864 3699
rect 13830 3597 13864 3631
rect 13830 3529 13864 3563
rect 13830 3461 13864 3487
rect 13986 3938 14020 3953
rect 14106 3938 14140 3953
rect 13986 3869 14020 3903
rect 13986 3804 14020 3835
rect 13986 3733 14020 3767
rect 13986 3665 14020 3699
rect 13986 3597 14020 3631
rect 13986 3529 14020 3563
rect 13986 3461 14020 3495
rect 13986 3411 14020 3427
rect 14109 3937 14140 3938
rect 14075 3903 14106 3904
rect 14075 3869 14140 3903
rect 14075 3846 14106 3869
rect 14109 3812 14140 3835
rect 14075 3801 14140 3812
rect 14075 3767 14106 3801
rect 14075 3753 14140 3767
rect 14109 3733 14140 3753
rect 14075 3699 14106 3719
rect 14075 3665 14140 3699
rect 14075 3631 14106 3665
rect 14075 3597 14140 3631
rect 14075 3563 14106 3597
rect 14075 3529 14140 3563
rect 14075 3495 14106 3529
rect 14075 3461 14140 3495
rect 14075 3427 14106 3461
rect 14075 3411 14140 3427
rect 14262 3937 14296 3953
rect 14262 3869 14296 3903
rect 14262 3801 14296 3835
rect 14262 3733 14296 3767
rect 14262 3678 14296 3699
rect 14262 3597 14296 3631
rect 14262 3529 14296 3548
rect 14262 3486 14296 3495
rect 14262 3411 14296 3427
rect 14378 3937 14412 3953
rect 14378 3869 14412 3903
rect 14378 3801 14412 3835
rect 14378 3733 14412 3767
rect 14378 3678 14412 3699
rect 14378 3597 14412 3631
rect 14378 3529 14412 3548
rect 14378 3486 14412 3495
rect 14378 3411 14412 3427
rect 14534 3940 14568 3953
rect 14534 3869 14568 3903
rect 14534 3801 14568 3827
rect 14534 3733 14568 3747
rect 14534 3665 14568 3667
rect 14534 3621 14568 3631
rect 14534 3541 14568 3563
rect 14534 3461 14568 3495
rect 14534 3411 14568 3427
rect 14983 3894 15017 3915
rect 14983 3826 15017 3842
rect 14983 3758 15017 3769
rect 14983 3690 15017 3696
rect 14983 3622 15017 3623
rect 14983 3584 15017 3588
rect 14983 3511 15017 3520
rect 14983 3438 15017 3452
rect 13431 3376 13477 3404
rect 13431 3342 13437 3376
rect 13471 3370 13477 3376
rect 13431 3336 13439 3342
rect 13473 3336 13477 3370
rect 13431 3302 13477 3336
rect 13431 3268 13437 3302
rect 13473 3268 13477 3302
rect 13431 3230 13477 3268
rect 13955 3336 13993 3370
rect 14027 3336 14209 3368
rect 13563 3309 13597 3330
rect 13719 3309 13869 3336
rect 13753 3250 13835 3309
rect 13922 3309 14209 3336
rect 14983 3365 15017 3384
rect 13922 3275 13991 3309
rect 14025 3275 14107 3309
rect 14141 3275 14209 3309
rect 13922 3261 14209 3275
rect 13959 3259 14209 3261
rect 14263 3309 14413 3329
rect 13719 3238 13869 3250
rect 14297 3250 14379 3309
rect 14505 3324 14611 3335
rect 14505 3309 14556 3324
rect 14505 3275 14535 3309
rect 14590 3290 14611 3324
rect 14569 3275 14611 3290
rect 14505 3259 14611 3275
rect 14983 3292 15017 3316
rect 14263 3238 14413 3250
rect 14556 3252 14590 3259
rect 14983 3219 15017 3248
rect 13227 3186 13239 3200
rect 14025 3195 14412 3198
rect 13193 3162 13239 3186
rect 13193 3152 13205 3162
rect 13608 3161 13617 3195
rect 13658 3161 13701 3195
rect 13735 3161 13751 3195
rect 13812 3161 13854 3195
rect 13888 3161 13930 3195
rect 13964 3161 13980 3195
rect 14059 3161 14114 3195
rect 14148 3161 14168 3195
rect 14236 3161 14245 3195
rect 14279 3161 14290 3195
rect 14356 3161 14378 3195
rect 14432 3161 14474 3195
rect 14508 3161 14524 3195
rect 14025 3158 14412 3161
rect 13227 3118 13239 3128
rect 14983 3146 15017 3180
rect 13193 3089 13239 3118
rect 13719 3106 13869 3118
rect 13193 3084 13205 3089
rect 13227 3050 13239 3055
rect 11509 3043 12365 3044
rect 11509 3009 11543 3043
rect 11577 3009 11612 3043
rect 11646 3009 11681 3043
rect 11715 3009 11750 3043
rect 11784 3009 11819 3043
rect 11853 3009 11888 3043
rect 11922 3009 11957 3043
rect 11991 3009 12025 3043
rect 12059 3009 12093 3043
rect 12127 3009 12161 3043
rect 12195 3009 12229 3043
rect 12263 3009 12297 3043
rect 12331 3009 12365 3043
rect 11509 2956 12365 3009
rect 11509 2955 11564 2956
rect 11598 2955 11640 2956
rect 11674 2955 11716 2956
rect 11509 2921 11543 2955
rect 11598 2922 11612 2955
rect 11674 2922 11681 2955
rect 11577 2921 11612 2922
rect 11646 2921 11681 2922
rect 11715 2922 11716 2955
rect 11750 2955 11792 2956
rect 11826 2955 11868 2956
rect 11902 2955 11943 2956
rect 11977 2955 12018 2956
rect 12052 2955 12093 2956
rect 12127 2955 12168 2956
rect 12202 2955 12243 2956
rect 12277 2955 12318 2956
rect 11715 2921 11750 2922
rect 11784 2922 11792 2955
rect 11853 2922 11868 2955
rect 11922 2922 11943 2955
rect 11991 2922 12018 2955
rect 11784 2921 11819 2922
rect 11853 2921 11888 2922
rect 11922 2921 11957 2922
rect 11991 2921 12025 2922
rect 12059 2921 12093 2955
rect 12127 2921 12161 2955
rect 12202 2922 12229 2955
rect 12277 2922 12297 2955
rect 12352 2922 12365 2956
rect 12195 2921 12229 2922
rect 12263 2921 12297 2922
rect 12331 2921 12365 2922
rect 11509 2880 12365 2921
rect 11509 2867 11564 2880
rect 11598 2867 11640 2880
rect 11674 2867 11716 2880
rect 11509 2833 11543 2867
rect 11598 2846 11612 2867
rect 11674 2846 11681 2867
rect 11577 2833 11612 2846
rect 11646 2833 11681 2846
rect 11715 2846 11716 2867
rect 11750 2867 11792 2880
rect 11826 2867 11868 2880
rect 11902 2867 11943 2880
rect 11977 2867 12018 2880
rect 12052 2867 12093 2880
rect 12127 2867 12168 2880
rect 12202 2867 12243 2880
rect 12277 2867 12318 2880
rect 11715 2833 11750 2846
rect 11784 2846 11792 2867
rect 11853 2846 11868 2867
rect 11922 2846 11943 2867
rect 11991 2846 12018 2867
rect 11784 2833 11819 2846
rect 11853 2833 11888 2846
rect 11922 2833 11957 2846
rect 11991 2833 12025 2846
rect 12059 2833 12093 2867
rect 12127 2833 12161 2867
rect 12202 2846 12229 2867
rect 12277 2846 12297 2867
rect 12352 2846 12365 2880
rect 12195 2833 12229 2846
rect 12263 2833 12297 2846
rect 12331 2833 12365 2846
rect 11509 2804 12365 2833
rect 11509 2779 11564 2804
rect 11598 2779 11640 2804
rect 11674 2779 11716 2804
rect 11509 2745 11543 2779
rect 11598 2770 11612 2779
rect 11674 2770 11681 2779
rect 11577 2745 11612 2770
rect 11646 2745 11681 2770
rect 11715 2770 11716 2779
rect 11750 2779 11792 2804
rect 11826 2779 11868 2804
rect 11902 2779 11943 2804
rect 11977 2779 12018 2804
rect 12052 2779 12093 2804
rect 12127 2779 12168 2804
rect 12202 2779 12243 2804
rect 12277 2779 12318 2804
rect 11715 2745 11750 2770
rect 11784 2770 11792 2779
rect 11853 2770 11868 2779
rect 11922 2770 11943 2779
rect 11991 2770 12018 2779
rect 11784 2745 11819 2770
rect 11853 2745 11888 2770
rect 11922 2745 11957 2770
rect 11991 2745 12025 2770
rect 12059 2745 12093 2779
rect 12127 2745 12161 2779
rect 12202 2770 12229 2779
rect 12277 2770 12297 2779
rect 12352 2770 12365 2804
rect 12195 2745 12229 2770
rect 12263 2745 12297 2770
rect 12331 2745 12365 2770
rect 11509 2744 12365 2745
rect 11564 2728 12365 2744
rect 11598 2694 11640 2728
rect 11674 2694 11716 2728
rect 11750 2694 11792 2728
rect 11826 2710 11868 2728
rect 11902 2710 11943 2728
rect 11977 2710 12018 2728
rect 12052 2710 12093 2728
rect 12127 2710 12168 2728
rect 12202 2710 12243 2728
rect 12277 2710 12318 2728
rect 12352 2710 12365 2728
rect 11826 2694 11841 2710
rect 11902 2694 11911 2710
rect 11977 2694 11981 2710
rect 11564 2676 11841 2694
rect 11875 2676 11911 2694
rect 11945 2676 11981 2694
rect 12015 2694 12018 2710
rect 12085 2694 12093 2710
rect 12155 2694 12168 2710
rect 12225 2694 12243 2710
rect 12295 2694 12318 2710
rect 12015 2676 12051 2694
rect 12085 2676 12121 2694
rect 12155 2676 12191 2694
rect 12225 2676 12261 2694
rect 12295 2676 12331 2694
rect 11564 2652 12365 2676
rect 11598 2618 11640 2652
rect 11674 2618 11716 2652
rect 11750 2618 11792 2652
rect 11826 2637 11868 2652
rect 11902 2637 11943 2652
rect 11977 2637 12018 2652
rect 12052 2637 12093 2652
rect 12127 2637 12168 2652
rect 12202 2637 12243 2652
rect 12277 2637 12318 2652
rect 12352 2637 12365 2652
rect 11826 2618 11841 2637
rect 11902 2618 11911 2637
rect 11977 2618 11981 2637
rect 11564 2603 11841 2618
rect 11875 2603 11911 2618
rect 11945 2603 11981 2618
rect 12015 2618 12018 2637
rect 12085 2618 12093 2637
rect 12155 2618 12168 2637
rect 12225 2618 12243 2637
rect 12295 2618 12318 2637
rect 12015 2603 12051 2618
rect 12085 2603 12121 2618
rect 12155 2603 12191 2618
rect 12225 2603 12261 2618
rect 12295 2603 12331 2618
rect 11564 2576 12365 2603
rect 11598 2542 11640 2576
rect 11674 2542 11716 2576
rect 11750 2542 11792 2576
rect 11826 2564 11868 2576
rect 11902 2564 11943 2576
rect 11977 2564 12018 2576
rect 12052 2564 12093 2576
rect 12127 2564 12168 2576
rect 12202 2564 12243 2576
rect 12277 2564 12318 2576
rect 12352 2564 12365 2576
rect 11826 2542 11841 2564
rect 11902 2542 11911 2564
rect 11977 2542 11981 2564
rect 11564 2530 11841 2542
rect 11875 2530 11911 2542
rect 11945 2530 11981 2542
rect 12015 2542 12018 2564
rect 12085 2542 12093 2564
rect 12155 2542 12168 2564
rect 12225 2542 12243 2564
rect 12295 2542 12318 2564
rect 12015 2530 12051 2542
rect 12085 2530 12121 2542
rect 12155 2530 12191 2542
rect 12225 2530 12261 2542
rect 12295 2530 12331 2542
rect 11564 2500 12365 2530
rect 11598 2466 11640 2500
rect 11674 2466 11716 2500
rect 11750 2466 11792 2500
rect 11826 2491 11868 2500
rect 11902 2491 11943 2500
rect 11977 2491 12018 2500
rect 12052 2491 12093 2500
rect 12127 2491 12168 2500
rect 12202 2491 12243 2500
rect 12277 2491 12318 2500
rect 12352 2491 12365 2500
rect 11826 2466 11841 2491
rect 11902 2466 11911 2491
rect 11977 2466 11981 2491
rect 11564 2457 11841 2466
rect 11875 2457 11911 2466
rect 11945 2457 11981 2466
rect 12015 2466 12018 2491
rect 12085 2466 12093 2491
rect 12155 2466 12168 2491
rect 12225 2466 12243 2491
rect 12295 2466 12318 2491
rect 13193 3016 13239 3050
rect 13563 3025 13597 3047
rect 13753 3047 13835 3106
rect 14263 3106 14413 3118
rect 13719 3031 13869 3047
rect 13991 3081 14141 3097
rect 14025 3047 14107 3081
rect 13991 3016 14141 3047
rect 14297 3047 14379 3106
rect 14263 3031 14413 3047
rect 14474 3094 14569 3097
rect 14508 3081 14569 3094
rect 14508 3060 14535 3081
rect 14474 3047 14535 3060
rect 13193 2948 13239 2982
rect 14025 2982 14107 3016
rect 14474 3022 14569 3047
rect 14508 2988 14569 3022
rect 14983 3078 15017 3112
rect 14983 3010 15017 3039
rect 13991 2979 14141 2982
rect 13227 2943 13239 2948
rect 13193 2909 13205 2914
rect 13193 2883 13239 2909
rect 14983 2942 15017 2966
rect 14983 2883 15017 2893
rect 13193 2881 15017 2883
rect 13193 2880 13261 2881
rect 13227 2870 13261 2880
rect 13295 2877 13330 2881
rect 13364 2877 13399 2881
rect 13433 2877 13468 2881
rect 13239 2847 13261 2870
rect 13311 2847 13330 2877
rect 13386 2847 13399 2877
rect 13461 2847 13468 2877
rect 13502 2877 13537 2881
rect 13193 2836 13205 2846
rect 13239 2843 13277 2847
rect 13311 2843 13352 2847
rect 13386 2843 13427 2847
rect 13461 2843 13502 2847
rect 13536 2847 13537 2877
rect 13571 2877 13606 2881
rect 13640 2877 13675 2881
rect 13709 2877 13744 2881
rect 13778 2877 13813 2881
rect 13847 2877 13882 2881
rect 13916 2877 13951 2881
rect 13571 2847 13577 2877
rect 13640 2847 13652 2877
rect 13709 2847 13727 2877
rect 13778 2847 13801 2877
rect 13847 2847 13875 2877
rect 13916 2847 13949 2877
rect 13985 2847 14020 2881
rect 14054 2877 14089 2881
rect 14123 2877 14158 2881
rect 14192 2877 14227 2881
rect 14261 2877 14296 2881
rect 14330 2877 14365 2881
rect 14399 2877 14434 2881
rect 14468 2877 14503 2881
rect 14057 2847 14089 2877
rect 14131 2847 14158 2877
rect 14205 2847 14227 2877
rect 14279 2847 14296 2877
rect 14353 2847 14365 2877
rect 14427 2847 14434 2877
rect 14501 2847 14503 2877
rect 14537 2877 14572 2881
rect 14606 2877 14641 2881
rect 14675 2877 14710 2881
rect 14744 2877 14779 2881
rect 14813 2877 14847 2881
rect 14881 2877 14915 2881
rect 14537 2847 14541 2877
rect 14606 2847 14615 2877
rect 14675 2847 14689 2877
rect 14744 2847 14763 2877
rect 14813 2847 14837 2877
rect 14881 2847 14911 2877
rect 14949 2874 15017 2881
rect 14949 2847 14983 2874
rect 13536 2843 13577 2847
rect 13611 2843 13652 2847
rect 13686 2843 13727 2847
rect 13761 2843 13801 2847
rect 13835 2843 13875 2847
rect 13909 2843 13949 2847
rect 13983 2843 14023 2847
rect 14057 2843 14097 2847
rect 14131 2843 14171 2847
rect 14205 2843 14245 2847
rect 14279 2843 14319 2847
rect 14353 2843 14393 2847
rect 14427 2843 14467 2847
rect 14501 2843 14541 2847
rect 14575 2843 14615 2847
rect 14649 2843 14689 2847
rect 14723 2843 14763 2847
rect 14797 2843 14837 2847
rect 14871 2843 14911 2847
rect 14945 2843 14983 2847
rect 13239 2837 14983 2843
rect 13193 2812 13239 2836
rect 13227 2797 13239 2812
rect 13193 2763 13205 2778
rect 13193 2744 13239 2763
rect 13227 2724 13239 2744
rect 13193 2690 13205 2710
rect 14983 2806 15017 2820
rect 14983 2738 15017 2747
rect 13193 2676 13239 2690
rect 13227 2651 13239 2676
rect 13193 2617 13205 2642
rect 13193 2608 13239 2617
rect 13227 2578 13239 2608
rect 13193 2544 13205 2574
rect 13193 2540 13239 2544
rect 13227 2506 13239 2540
rect 13193 2505 13239 2506
rect 12015 2457 12051 2466
rect 12085 2457 12121 2466
rect 12155 2457 12191 2466
rect 12225 2457 12261 2466
rect 12295 2457 12331 2466
rect 11564 2424 12365 2457
rect 11598 2390 11640 2424
rect 11674 2390 11716 2424
rect 11750 2390 11792 2424
rect 11826 2418 11868 2424
rect 11902 2418 11943 2424
rect 11977 2418 12018 2424
rect 12052 2418 12093 2424
rect 12127 2418 12168 2424
rect 12202 2418 12243 2424
rect 12277 2418 12318 2424
rect 12352 2418 12365 2424
rect 11826 2390 11841 2418
rect 11902 2390 11911 2418
rect 11977 2390 11981 2418
rect 11564 2384 11841 2390
rect 11875 2384 11911 2390
rect 11945 2384 11981 2390
rect 12015 2390 12018 2418
rect 12085 2390 12093 2418
rect 12155 2390 12168 2418
rect 12225 2390 12243 2418
rect 12295 2390 12318 2418
rect 12015 2384 12051 2390
rect 12085 2384 12121 2390
rect 12155 2384 12191 2390
rect 12225 2384 12261 2390
rect 12295 2384 12331 2390
rect 11564 2348 12365 2384
rect 11598 2314 11640 2348
rect 11674 2314 11716 2348
rect 11750 2314 11792 2348
rect 11826 2344 11868 2348
rect 11902 2344 11943 2348
rect 11977 2344 12018 2348
rect 12052 2344 12093 2348
rect 12127 2344 12168 2348
rect 12202 2344 12243 2348
rect 12277 2344 12318 2348
rect 12352 2344 12365 2348
rect 11826 2314 11841 2344
rect 11902 2314 11911 2344
rect 11977 2314 11981 2344
rect 11564 2310 11841 2314
rect 11875 2310 11911 2314
rect 11945 2310 11981 2314
rect 12015 2314 12018 2344
rect 12085 2314 12093 2344
rect 12155 2314 12168 2344
rect 12225 2314 12243 2344
rect 12295 2314 12318 2344
rect 12499 2452 12539 2486
rect 12573 2452 12613 2486
rect 12647 2452 12687 2486
rect 12721 2452 12761 2486
rect 12795 2452 12835 2486
rect 12465 2370 12869 2452
rect 12499 2336 12539 2370
rect 12573 2336 12613 2370
rect 12647 2336 12687 2370
rect 12721 2336 12761 2370
rect 12795 2336 12835 2370
rect 13193 2472 13205 2505
rect 13227 2438 13239 2471
rect 13193 2432 13239 2438
rect 13193 2404 13205 2432
rect 13227 2370 13239 2398
rect 13193 2359 13239 2370
rect 13193 2336 13205 2359
rect 12015 2310 12051 2314
rect 12085 2310 12121 2314
rect 12155 2310 12191 2314
rect 12225 2310 12261 2314
rect 12295 2310 12331 2314
rect 11564 2272 12365 2310
rect 11598 2238 11640 2272
rect 11674 2238 11716 2272
rect 11750 2238 11792 2272
rect 11826 2270 11868 2272
rect 11902 2270 11943 2272
rect 11977 2270 12018 2272
rect 12052 2270 12093 2272
rect 12127 2270 12168 2272
rect 12202 2270 12243 2272
rect 12277 2270 12318 2272
rect 12352 2270 12365 2272
rect 11826 2238 11841 2270
rect 11902 2238 11911 2270
rect 11977 2238 11981 2270
rect 11875 2236 11911 2238
rect 11945 2236 11981 2238
rect 12015 2238 12018 2270
rect 12085 2238 12093 2270
rect 12155 2238 12168 2270
rect 12225 2238 12243 2270
rect 12295 2238 12318 2270
rect 12015 2236 12051 2238
rect 12085 2236 12121 2238
rect 12155 2236 12191 2238
rect 12225 2236 12261 2238
rect 12295 2236 12331 2238
rect 11841 2202 12365 2236
rect 13227 2302 13239 2325
rect 13193 2286 13239 2302
rect 13193 2268 13205 2286
rect 13227 2234 13239 2252
rect 13193 2213 13239 2234
rect 3864 2132 4940 2167
rect 3864 2098 3875 2132
rect 3909 2098 3943 2132
rect 3977 2098 4011 2132
rect 4045 2098 4079 2132
rect 4113 2098 4147 2132
rect 4181 2098 4215 2132
rect 4249 2098 4283 2132
rect 4317 2098 4351 2132
rect 4385 2098 4419 2132
rect 4453 2098 4487 2132
rect 4521 2098 4555 2132
rect 4589 2098 4623 2132
rect 4657 2098 4691 2132
rect 4725 2098 4759 2132
rect 4793 2098 4827 2132
rect 4861 2098 4895 2132
rect 4929 2098 4940 2132
rect 3864 2063 4940 2098
rect 3864 2029 3875 2063
rect 3909 2029 3943 2063
rect 3977 2029 4011 2063
rect 4045 2029 4079 2063
rect 4113 2029 4147 2063
rect 4181 2029 4215 2063
rect 4249 2029 4283 2063
rect 4317 2029 4351 2063
rect 4385 2029 4419 2063
rect 4453 2029 4487 2063
rect 4521 2029 4555 2063
rect 4589 2029 4623 2063
rect 4657 2029 4691 2063
rect 4725 2029 4759 2063
rect 4793 2029 4827 2063
rect 4861 2029 4895 2063
rect 4929 2029 4940 2063
rect 3864 1994 4940 2029
rect 3864 1960 3875 1994
rect 3909 1960 3943 1994
rect 3977 1960 4011 1994
rect 4045 1960 4079 1994
rect 4113 1960 4147 1994
rect 4181 1960 4215 1994
rect 4249 1960 4283 1994
rect 4317 1960 4351 1994
rect 4385 1960 4419 1994
rect 4453 1960 4487 1994
rect 4521 1960 4555 1994
rect 4589 1960 4623 1994
rect 4657 1960 4691 1994
rect 4725 1960 4759 1994
rect 4793 1960 4827 1994
rect 4861 1960 4895 1994
rect 4929 1960 4940 1994
rect 3864 1925 4940 1960
rect 3864 1891 3875 1925
rect 3909 1891 3943 1925
rect 3977 1891 4011 1925
rect 4045 1891 4079 1925
rect 4113 1891 4147 1925
rect 4181 1891 4215 1925
rect 4249 1891 4283 1925
rect 4317 1891 4351 1925
rect 4385 1891 4419 1925
rect 4453 1891 4487 1925
rect 4521 1891 4555 1925
rect 4589 1891 4623 1925
rect 4657 1891 4691 1925
rect 4725 1891 4759 1925
rect 4793 1891 4827 1925
rect 4861 1891 4895 1925
rect 4929 1891 4940 1925
rect 3864 1856 4940 1891
rect 3864 1822 3875 1856
rect 3909 1822 3943 1856
rect 3977 1822 4011 1856
rect 4045 1822 4079 1856
rect 4113 1822 4147 1856
rect 4181 1822 4215 1856
rect 4249 1822 4283 1856
rect 4317 1822 4351 1856
rect 4385 1822 4419 1856
rect 4453 1822 4487 1856
rect 4521 1822 4555 1856
rect 4589 1822 4623 1856
rect 4657 1822 4691 1856
rect 4725 1822 4759 1856
rect 4793 1822 4827 1856
rect 4861 1822 4895 1856
rect 4929 1822 4940 1856
rect 3864 1787 4940 1822
rect 3864 1753 3875 1787
rect 3909 1753 3943 1787
rect 3977 1753 4011 1787
rect 4045 1753 4079 1787
rect 4113 1753 4147 1787
rect 4181 1753 4215 1787
rect 4249 1753 4283 1787
rect 4317 1753 4351 1787
rect 4385 1753 4419 1787
rect 4453 1753 4487 1787
rect 4521 1753 4555 1787
rect 4589 1753 4623 1787
rect 4657 1753 4691 1787
rect 4725 1753 4759 1787
rect 4793 1753 4827 1787
rect 4861 1753 4895 1787
rect 4929 1753 4940 1787
rect 3864 1718 4940 1753
rect 3864 1684 3875 1718
rect 3909 1684 3943 1718
rect 3977 1684 4011 1718
rect 4045 1684 4079 1718
rect 4113 1684 4147 1718
rect 4181 1684 4215 1718
rect 4249 1684 4283 1718
rect 4317 1684 4351 1718
rect 4385 1684 4419 1718
rect 4453 1684 4487 1718
rect 4521 1684 4555 1718
rect 4589 1684 4623 1718
rect 4657 1684 4691 1718
rect 4725 1684 4759 1718
rect 4793 1684 4827 1718
rect 4861 1684 4895 1718
rect 4929 1684 4940 1718
rect 3864 1649 4940 1684
rect 3864 1615 3875 1649
rect 3909 1615 3943 1649
rect 3977 1615 4011 1649
rect 4045 1615 4079 1649
rect 4113 1615 4147 1649
rect 4181 1615 4215 1649
rect 4249 1615 4283 1649
rect 4317 1615 4351 1649
rect 4385 1615 4419 1649
rect 4453 1615 4487 1649
rect 4521 1615 4555 1649
rect 4589 1615 4623 1649
rect 4657 1615 4691 1649
rect 4725 1615 4759 1649
rect 4793 1615 4827 1649
rect 4861 1615 4895 1649
rect 4929 1615 4940 1649
rect 3864 1580 4940 1615
rect 3864 1546 3875 1580
rect 3909 1546 3943 1580
rect 3977 1546 4011 1580
rect 4045 1546 4079 1580
rect 4113 1546 4147 1580
rect 4181 1546 4215 1580
rect 4249 1546 4283 1580
rect 4317 1546 4351 1580
rect 4385 1546 4419 1580
rect 4453 1546 4487 1580
rect 4521 1546 4555 1580
rect 4589 1546 4623 1580
rect 4657 1546 4691 1580
rect 4725 1546 4759 1580
rect 4793 1546 4827 1580
rect 4861 1546 4895 1580
rect 4929 1546 4940 1580
rect 3864 1511 4940 1546
rect 3864 1477 3875 1511
rect 3909 1477 3943 1511
rect 3977 1477 4011 1511
rect 4045 1477 4079 1511
rect 4113 1477 4147 1511
rect 4181 1477 4215 1511
rect 4249 1477 4283 1511
rect 4317 1477 4351 1511
rect 4385 1477 4419 1511
rect 4453 1477 4487 1511
rect 4521 1477 4555 1511
rect 4589 1477 4623 1511
rect 4657 1477 4691 1511
rect 4725 1477 4759 1511
rect 4793 1477 4827 1511
rect 4861 1477 4895 1511
rect 4929 1477 4940 1511
rect 3864 1442 4940 1477
rect 3864 1408 3875 1442
rect 3909 1408 3943 1442
rect 3977 1408 4011 1442
rect 4045 1408 4079 1442
rect 4113 1408 4147 1442
rect 4181 1408 4215 1442
rect 4249 1408 4283 1442
rect 4317 1408 4351 1442
rect 4385 1408 4419 1442
rect 4453 1408 4487 1442
rect 4521 1408 4555 1442
rect 4589 1408 4623 1442
rect 4657 1408 4691 1442
rect 4725 1408 4759 1442
rect 4793 1408 4827 1442
rect 4861 1408 4895 1442
rect 4929 1408 4940 1442
rect 3864 1373 4940 1408
rect 3864 1339 3875 1373
rect 3909 1339 3943 1373
rect 3977 1339 4011 1373
rect 4045 1339 4079 1373
rect 4113 1339 4147 1373
rect 4181 1339 4215 1373
rect 4249 1339 4283 1373
rect 4317 1339 4351 1373
rect 4385 1339 4419 1373
rect 4453 1339 4487 1373
rect 4521 1339 4555 1373
rect 4589 1339 4623 1373
rect 4657 1339 4691 1373
rect 4725 1339 4759 1373
rect 4793 1339 4827 1373
rect 4861 1339 4895 1373
rect 4929 1339 4940 1373
rect 3864 1304 4940 1339
rect 3864 1270 3875 1304
rect 3909 1270 3943 1304
rect 3977 1270 4011 1304
rect 4045 1270 4079 1304
rect 4113 1270 4147 1304
rect 4181 1270 4215 1304
rect 4249 1270 4283 1304
rect 4317 1270 4351 1304
rect 4385 1270 4419 1304
rect 4453 1270 4487 1304
rect 4521 1270 4555 1304
rect 4589 1270 4623 1304
rect 4657 1270 4691 1304
rect 4725 1270 4759 1304
rect 4793 1270 4827 1304
rect 4861 1270 4895 1304
rect 4929 1270 4940 1304
rect 3864 1235 4940 1270
rect 3864 1201 3875 1235
rect 3909 1201 3943 1235
rect 3977 1201 4011 1235
rect 4045 1201 4079 1235
rect 4113 1201 4147 1235
rect 4181 1201 4215 1235
rect 4249 1201 4283 1235
rect 4317 1201 4351 1235
rect 4385 1201 4419 1235
rect 4453 1201 4487 1235
rect 4521 1201 4555 1235
rect 4589 1201 4623 1235
rect 4657 1201 4691 1235
rect 4725 1201 4759 1235
rect 4793 1201 4827 1235
rect 4861 1201 4895 1235
rect 4929 1201 4940 1235
rect 3864 1166 4940 1201
rect 3864 1132 3875 1166
rect 3909 1132 3943 1166
rect 3977 1132 4011 1166
rect 4045 1132 4079 1166
rect 4113 1132 4147 1166
rect 4181 1132 4215 1166
rect 4249 1132 4283 1166
rect 4317 1132 4351 1166
rect 4385 1132 4419 1166
rect 4453 1132 4487 1166
rect 4521 1132 4555 1166
rect 4589 1132 4623 1166
rect 4657 1132 4691 1166
rect 4725 1132 4759 1166
rect 4793 1132 4827 1166
rect 4861 1132 4895 1166
rect 4929 1132 4940 1166
rect 3864 1097 4940 1132
rect 3864 1063 3875 1097
rect 3909 1063 3943 1097
rect 3977 1063 4011 1097
rect 4045 1063 4079 1097
rect 4113 1063 4147 1097
rect 4181 1063 4215 1097
rect 4249 1063 4283 1097
rect 4317 1063 4351 1097
rect 4385 1063 4419 1097
rect 4453 1063 4487 1097
rect 4521 1063 4555 1097
rect 4589 1063 4623 1097
rect 4657 1063 4691 1097
rect 4725 1063 4759 1097
rect 4793 1063 4827 1097
rect 4861 1063 4895 1097
rect 4929 1063 4940 1097
rect 13193 2200 13205 2213
rect 13227 2166 13239 2179
rect 13193 2140 13239 2166
rect 13193 2132 13205 2140
rect 13227 2098 13239 2106
rect 13193 2067 13239 2098
rect 13193 2064 13205 2067
rect 13227 2030 13239 2033
rect 13193 1996 13239 2030
rect 13227 1994 13239 1996
rect 13193 1960 13205 1962
rect 13193 1928 13239 1960
rect 13227 1921 13239 1928
rect 13193 1887 13205 1894
rect 13193 1860 13239 1887
rect 13227 1848 13239 1860
rect 13193 1814 13205 1826
rect 13193 1792 13239 1814
rect 13227 1775 13239 1792
rect 13193 1741 13205 1758
rect 13193 1724 13239 1741
rect 13227 1702 13239 1724
rect 13193 1668 13205 1690
rect 13193 1656 13239 1668
rect 13227 1629 13239 1656
rect 13193 1595 13205 1622
rect 13193 1588 13239 1595
rect 13227 1556 13239 1588
rect 13193 1522 13205 1554
rect 13193 1520 13239 1522
rect 13227 1486 13239 1520
rect 13193 1483 13239 1486
rect 13193 1452 13205 1483
rect 13227 1418 13239 1449
rect 13193 1410 13239 1418
rect 13193 1384 13205 1410
rect 13227 1350 13239 1376
rect 13193 1337 13239 1350
rect 13193 1316 13205 1337
rect 13227 1282 13239 1303
rect 13193 1264 13239 1282
rect 13193 1248 13205 1264
rect 13227 1214 13239 1230
rect 13193 1191 13239 1214
rect 13193 1180 13205 1191
rect 13227 1146 13239 1157
rect 13193 1118 13239 1146
rect 13193 1112 13205 1118
rect 3864 1028 4940 1063
rect 3864 994 3875 1028
rect 3909 994 3943 1028
rect 3977 994 4011 1028
rect 4045 994 4079 1028
rect 4113 994 4147 1028
rect 4181 994 4215 1028
rect 4249 994 4283 1028
rect 4317 994 4351 1028
rect 4385 994 4419 1028
rect 4453 994 4487 1028
rect 4521 994 4555 1028
rect 4589 994 4623 1028
rect 4657 994 4691 1028
rect 4725 994 4759 1028
rect 4793 994 4827 1028
rect 4861 994 4895 1028
rect 4929 994 4940 1028
rect 3864 959 4940 994
rect 3864 925 3875 959
rect 3909 925 3943 959
rect 3977 925 4011 959
rect 4045 925 4079 959
rect 4113 925 4147 959
rect 4181 925 4215 959
rect 4249 925 4283 959
rect 4317 925 4351 959
rect 4385 925 4419 959
rect 4453 925 4487 959
rect 4521 925 4555 959
rect 4589 925 4623 959
rect 4657 925 4691 959
rect 4725 925 4759 959
rect 4793 925 4827 959
rect 4861 925 4895 959
rect 4929 925 4940 959
rect 3864 890 4940 925
rect 3864 856 3875 890
rect 3909 856 3943 890
rect 3977 856 4011 890
rect 4045 856 4079 890
rect 4113 856 4147 890
rect 4181 856 4215 890
rect 4249 856 4283 890
rect 4317 856 4351 890
rect 4385 856 4419 890
rect 4453 856 4487 890
rect 4521 856 4555 890
rect 4589 856 4623 890
rect 4657 856 4691 890
rect 4725 856 4759 890
rect 4793 856 4827 890
rect 4861 856 4895 890
rect 4929 856 4940 890
rect 3864 821 4940 856
rect 5299 1058 8646 1093
rect 5333 1024 5369 1058
rect 5403 1024 5438 1058
rect 5472 1024 5507 1058
rect 5541 1024 5576 1058
rect 5610 1024 5645 1058
rect 5679 1024 5714 1058
rect 5748 1024 5783 1058
rect 5817 1024 5852 1058
rect 5886 1024 5921 1058
rect 5955 1024 5990 1058
rect 6024 1024 6059 1058
rect 6093 1024 6128 1058
rect 6162 1024 6197 1058
rect 6231 1024 6266 1058
rect 6300 1024 6335 1058
rect 6369 1024 6404 1058
rect 6438 1024 6473 1058
rect 6507 1024 6542 1058
rect 6576 1024 6611 1058
rect 6645 1024 6680 1058
rect 6714 1024 6749 1058
rect 6783 1024 6818 1058
rect 6852 1024 6887 1058
rect 6921 1024 6956 1058
rect 6990 1024 7025 1058
rect 7059 1024 7094 1058
rect 7128 1024 7163 1058
rect 7197 1024 7232 1058
rect 7266 1024 7301 1058
rect 7335 1024 7370 1058
rect 7404 1024 7439 1058
rect 7473 1024 7508 1058
rect 7542 1024 7577 1058
rect 7611 1024 7646 1058
rect 7680 1024 7715 1058
rect 7749 1024 7784 1058
rect 7818 1024 7853 1058
rect 7887 1024 7922 1058
rect 7956 1024 7991 1058
rect 8025 1024 8060 1058
rect 8094 1024 8129 1058
rect 8163 1024 8198 1058
rect 8232 1024 8267 1058
rect 8301 1024 8336 1058
rect 8370 1024 8405 1058
rect 8439 1024 8474 1058
rect 8508 1024 8543 1058
rect 8577 1024 8612 1058
rect 5299 986 8646 1024
rect 5333 952 5369 986
rect 5403 952 5438 986
rect 5472 952 5507 986
rect 5541 952 5576 986
rect 5610 952 5645 986
rect 5679 952 5714 986
rect 5748 952 5783 986
rect 5817 952 5852 986
rect 5886 952 5921 986
rect 5955 952 5990 986
rect 6024 952 6059 986
rect 6093 952 6128 986
rect 6162 952 6197 986
rect 6231 952 6266 986
rect 6300 952 6335 986
rect 6369 952 6404 986
rect 6438 952 6473 986
rect 6507 952 6542 986
rect 6576 952 6611 986
rect 6645 952 6680 986
rect 6714 952 6749 986
rect 6783 952 6818 986
rect 6852 952 6887 986
rect 6921 952 6956 986
rect 6990 952 7025 986
rect 7059 952 7094 986
rect 7128 952 7163 986
rect 7197 952 7232 986
rect 7266 952 7301 986
rect 7335 952 7370 986
rect 7404 952 7439 986
rect 7473 952 7508 986
rect 7542 952 7577 986
rect 7611 952 7646 986
rect 7680 952 7715 986
rect 7749 952 7784 986
rect 7818 952 7853 986
rect 7887 952 7922 986
rect 7956 952 7991 986
rect 8025 952 8060 986
rect 8094 952 8129 986
rect 8163 952 8198 986
rect 8232 952 8267 986
rect 8301 952 8336 986
rect 8370 952 8405 986
rect 8439 952 8474 986
rect 8508 952 8543 986
rect 8577 952 8612 986
rect 5299 914 8646 952
rect 5333 880 5369 914
rect 5403 880 5438 914
rect 5472 880 5507 914
rect 5541 880 5576 914
rect 5610 880 5645 914
rect 5679 880 5714 914
rect 5748 880 5783 914
rect 5817 880 5852 914
rect 5886 880 5921 914
rect 5955 880 5990 914
rect 6024 880 6059 914
rect 6093 880 6128 914
rect 6162 880 6197 914
rect 6231 880 6266 914
rect 6300 880 6335 914
rect 6369 880 6404 914
rect 6438 880 6473 914
rect 6507 880 6542 914
rect 6576 880 6611 914
rect 6645 880 6680 914
rect 6714 880 6749 914
rect 6783 880 6818 914
rect 6852 880 6887 914
rect 6921 880 6956 914
rect 6990 880 7025 914
rect 7059 880 7094 914
rect 7128 880 7163 914
rect 7197 880 7232 914
rect 7266 880 7301 914
rect 7335 880 7370 914
rect 7404 880 7439 914
rect 7473 880 7508 914
rect 7542 880 7577 914
rect 7611 880 7646 914
rect 7680 880 7715 914
rect 7749 880 7784 914
rect 7818 880 7853 914
rect 7887 880 7922 914
rect 7956 880 7991 914
rect 8025 880 8060 914
rect 8094 880 8129 914
rect 8163 880 8198 914
rect 8232 880 8267 914
rect 8301 880 8336 914
rect 8370 880 8405 914
rect 8439 880 8474 914
rect 8508 880 8543 914
rect 8577 880 8612 914
rect 5299 845 8646 880
rect 13227 1078 13239 1084
rect 13193 1045 13239 1078
rect 13193 1044 13205 1045
rect 13227 1010 13239 1011
rect 13193 976 13239 1010
rect 13227 972 13239 976
rect 13193 938 13205 942
rect 13193 908 13239 938
rect 13227 899 13239 908
rect 3864 787 3875 821
rect 3909 787 3943 821
rect 3977 787 4011 821
rect 4045 787 4079 821
rect 4113 787 4147 821
rect 4181 787 4215 821
rect 4249 787 4283 821
rect 4317 787 4351 821
rect 4385 787 4419 821
rect 4453 787 4487 821
rect 4521 787 4555 821
rect 4589 787 4623 821
rect 4657 787 4691 821
rect 4725 787 4759 821
rect 4793 787 4827 821
rect 4861 787 4895 821
rect 4929 787 4940 821
rect 3864 752 4940 787
rect 3864 718 3875 752
rect 3909 718 3943 752
rect 3977 718 4011 752
rect 4045 718 4079 752
rect 4113 718 4147 752
rect 4181 718 4215 752
rect 4249 718 4283 752
rect 4317 718 4351 752
rect 4385 718 4419 752
rect 4453 718 4487 752
rect 4521 718 4555 752
rect 4589 718 4623 752
rect 4657 718 4691 752
rect 4725 718 4759 752
rect 4793 718 4827 752
rect 4861 718 4895 752
rect 4929 718 4940 752
rect 3864 683 4940 718
rect 3864 649 3875 683
rect 3909 649 3943 683
rect 3977 649 4011 683
rect 4045 649 4079 683
rect 4113 649 4147 683
rect 4181 649 4215 683
rect 4249 649 4283 683
rect 4317 649 4351 683
rect 4385 649 4419 683
rect 4453 649 4487 683
rect 4521 649 4555 683
rect 4589 649 4623 683
rect 4657 649 4691 683
rect 4725 649 4759 683
rect 4793 649 4827 683
rect 4861 649 4895 683
rect 4929 649 4940 683
rect 3864 614 4940 649
rect 3864 580 3875 614
rect 3909 580 3943 614
rect 3977 580 4011 614
rect 4045 580 4079 614
rect 4113 580 4147 614
rect 4181 580 4215 614
rect 4249 580 4283 614
rect 4317 580 4351 614
rect 4385 580 4419 614
rect 4453 580 4487 614
rect 4521 580 4555 614
rect 4589 580 4623 614
rect 4657 580 4691 614
rect 4725 580 4759 614
rect 4793 580 4827 614
rect 4861 580 4895 614
rect 4929 580 4940 614
rect 3864 545 4940 580
rect 3864 511 3875 545
rect 3909 511 3943 545
rect 3977 511 4011 545
rect 4045 511 4079 545
rect 4113 511 4147 545
rect 4181 511 4215 545
rect 4249 511 4283 545
rect 4317 511 4351 545
rect 4385 511 4419 545
rect 4453 511 4487 545
rect 4521 511 4555 545
rect 4589 511 4623 545
rect 4657 511 4691 545
rect 4725 511 4759 545
rect 4793 511 4827 545
rect 4861 511 4895 545
rect 4929 511 4940 545
rect 3864 476 4940 511
rect 3864 442 3875 476
rect 3909 442 3943 476
rect 3977 442 4011 476
rect 4045 442 4079 476
rect 4113 442 4147 476
rect 4181 442 4215 476
rect 4249 442 4283 476
rect 4317 442 4351 476
rect 4385 442 4419 476
rect 4453 442 4487 476
rect 4521 442 4555 476
rect 4589 442 4623 476
rect 4657 442 4691 476
rect 4725 442 4759 476
rect 4793 442 4827 476
rect 4861 442 4895 476
rect 4929 442 4940 476
rect 3864 407 4940 442
rect 3864 373 3875 407
rect 3909 373 3943 407
rect 3977 373 4011 407
rect 4045 373 4079 407
rect 4113 373 4147 407
rect 4181 373 4215 407
rect 4249 373 4283 407
rect 4317 373 4351 407
rect 4385 373 4419 407
rect 4453 373 4487 407
rect 4521 373 4555 407
rect 4589 373 4623 407
rect 4657 373 4691 407
rect 4725 373 4759 407
rect 4793 373 4827 407
rect 4861 373 4895 407
rect 4929 373 4940 407
rect 3864 338 4940 373
rect 3864 304 3875 338
rect 3909 304 3943 338
rect 3977 304 4011 338
rect 4045 304 4079 338
rect 4113 304 4147 338
rect 4181 304 4215 338
rect 4249 304 4283 338
rect 4317 304 4351 338
rect 4385 304 4419 338
rect 4453 304 4487 338
rect 4521 304 4555 338
rect 4589 304 4623 338
rect 4657 304 4691 338
rect 4725 304 4759 338
rect 4793 304 4827 338
rect 4861 304 4895 338
rect 4929 304 4940 338
rect 3864 269 4940 304
rect 3864 235 3875 269
rect 3909 235 3943 269
rect 3977 235 4011 269
rect 4045 235 4079 269
rect 4113 235 4147 269
rect 4181 235 4215 269
rect 4249 235 4283 269
rect 4317 235 4351 269
rect 4385 235 4419 269
rect 4453 235 4487 269
rect 4521 235 4555 269
rect 4589 235 4623 269
rect 4657 235 4691 269
rect 4725 235 4759 269
rect 4793 235 4827 269
rect 4861 235 4895 269
rect 4929 235 4940 269
rect 3864 200 4940 235
rect 3864 166 3875 200
rect 3909 166 3943 200
rect 3977 166 4011 200
rect 4045 166 4079 200
rect 4113 166 4147 200
rect 4181 166 4215 200
rect 4249 166 4283 200
rect 4317 166 4351 200
rect 4385 166 4419 200
rect 4453 166 4487 200
rect 4521 166 4555 200
rect 4589 166 4623 200
rect 4657 166 4691 200
rect 4725 166 4759 200
rect 4793 166 4827 200
rect 4861 166 4895 200
rect 4929 166 4940 200
rect 3864 131 4940 166
rect 3864 97 3875 131
rect 3909 97 3943 131
rect 3977 97 4011 131
rect 4045 97 4079 131
rect 4113 97 4147 131
rect 4181 97 4215 131
rect 4249 97 4283 131
rect 4317 97 4351 131
rect 4385 97 4419 131
rect 4453 97 4487 131
rect 4521 97 4555 131
rect 4589 97 4623 131
rect 4657 97 4691 131
rect 4725 97 4759 131
rect 4793 97 4827 131
rect 4861 97 4895 131
rect 4929 97 4940 131
rect 3864 62 4940 97
rect 3864 28 3875 62
rect 3909 28 3943 62
rect 3977 28 4011 62
rect 4045 28 4079 62
rect 4113 28 4147 62
rect 4181 28 4215 62
rect 4249 28 4283 62
rect 4317 28 4351 62
rect 4385 28 4419 62
rect 4453 28 4487 62
rect 4521 28 4555 62
rect 4589 28 4623 62
rect 4657 28 4691 62
rect 4725 28 4759 62
rect 4793 28 4827 62
rect 4861 28 4895 62
rect 4929 28 4940 62
rect 3864 4 4940 28
rect 11314 839 12838 879
rect 11348 805 11385 839
rect 11419 805 11456 839
rect 11490 837 11527 839
rect 11561 837 11598 839
rect 11632 837 11669 839
rect 11703 837 11740 839
rect 11774 837 11811 839
rect 11845 837 11882 839
rect 11916 837 11953 839
rect 11987 837 12024 839
rect 12058 837 12095 839
rect 11490 805 11502 837
rect 11561 805 11576 837
rect 11632 805 11650 837
rect 11703 805 11724 837
rect 11774 805 11798 837
rect 11845 805 11872 837
rect 11916 805 11946 837
rect 11987 805 12020 837
rect 12058 805 12094 837
rect 12129 805 12166 839
rect 12200 837 12237 839
rect 12271 837 12308 839
rect 12342 837 12379 839
rect 12413 837 12450 839
rect 12484 837 12521 839
rect 12555 837 12592 839
rect 12626 837 12663 839
rect 12697 837 12734 839
rect 12768 837 12804 839
rect 12202 805 12237 837
rect 12276 805 12308 837
rect 12350 805 12379 837
rect 12424 805 12450 837
rect 12498 805 12521 837
rect 12572 805 12592 837
rect 12645 805 12663 837
rect 12718 805 12734 837
rect 12791 805 12804 837
rect 11314 803 11502 805
rect 11536 803 11576 805
rect 11610 803 11650 805
rect 11684 803 11724 805
rect 11758 803 11798 805
rect 11832 803 11872 805
rect 11906 803 11946 805
rect 11980 803 12020 805
rect 12054 803 12094 805
rect 12128 803 12168 805
rect 12202 803 12242 805
rect 12276 803 12316 805
rect 12350 803 12390 805
rect 12424 803 12464 805
rect 12498 803 12538 805
rect 12572 803 12611 805
rect 12645 803 12684 805
rect 12718 803 12757 805
rect 12791 803 12838 805
rect 11314 769 12838 803
rect 11348 735 11385 769
rect 11419 735 11456 769
rect 11490 765 11527 769
rect 11561 765 11598 769
rect 11632 765 11669 769
rect 11703 765 11740 769
rect 11774 765 11811 769
rect 11845 765 11882 769
rect 11916 765 11953 769
rect 11987 765 12024 769
rect 12058 765 12095 769
rect 11490 735 11502 765
rect 11561 735 11576 765
rect 11632 735 11650 765
rect 11703 735 11724 765
rect 11774 735 11798 765
rect 11845 735 11872 765
rect 11916 735 11946 765
rect 11987 735 12020 765
rect 12058 735 12094 765
rect 12129 735 12166 769
rect 12200 765 12237 769
rect 12271 765 12308 769
rect 12342 765 12379 769
rect 12413 765 12450 769
rect 12484 765 12521 769
rect 12555 765 12592 769
rect 12626 765 12663 769
rect 12697 765 12734 769
rect 12768 765 12804 769
rect 12202 735 12237 765
rect 12276 735 12308 765
rect 12350 735 12379 765
rect 12424 735 12450 765
rect 12498 735 12521 765
rect 12572 735 12592 765
rect 12645 735 12663 765
rect 12718 735 12734 765
rect 12791 735 12804 765
rect 11314 731 11502 735
rect 11536 731 11576 735
rect 11610 731 11650 735
rect 11684 731 11724 735
rect 11758 731 11798 735
rect 11832 731 11872 735
rect 11906 731 11946 735
rect 11980 731 12020 735
rect 12054 731 12094 735
rect 12128 731 12168 735
rect 12202 731 12242 735
rect 12276 731 12316 735
rect 12350 731 12390 735
rect 12424 731 12464 735
rect 12498 731 12538 735
rect 12572 731 12611 735
rect 12645 731 12684 735
rect 12718 731 12757 735
rect 12791 731 12838 735
rect 11314 699 12838 731
rect 11348 665 11385 699
rect 11419 665 11456 699
rect 11490 693 11527 699
rect 11561 693 11598 699
rect 11632 693 11669 699
rect 11703 693 11740 699
rect 11774 693 11811 699
rect 11845 693 11882 699
rect 11916 693 11953 699
rect 11987 693 12024 699
rect 12058 693 12095 699
rect 11490 665 11502 693
rect 11561 665 11576 693
rect 11632 665 11650 693
rect 11703 665 11724 693
rect 11774 665 11798 693
rect 11845 665 11872 693
rect 11916 665 11946 693
rect 11987 665 12020 693
rect 12058 665 12094 693
rect 12129 665 12166 699
rect 12200 693 12237 699
rect 12271 693 12308 699
rect 12342 693 12379 699
rect 12413 693 12450 699
rect 12484 693 12521 699
rect 12555 693 12592 699
rect 12626 693 12663 699
rect 12697 693 12734 699
rect 12768 693 12804 699
rect 12202 665 12237 693
rect 12276 665 12308 693
rect 12350 665 12379 693
rect 12424 665 12450 693
rect 12498 665 12521 693
rect 12572 665 12592 693
rect 12645 665 12663 693
rect 12718 665 12734 693
rect 12791 665 12804 693
rect 11314 659 11502 665
rect 11536 659 11576 665
rect 11610 659 11650 665
rect 11684 659 11724 665
rect 11758 659 11798 665
rect 11832 659 11872 665
rect 11906 659 11946 665
rect 11980 659 12020 665
rect 12054 659 12094 665
rect 12128 659 12168 665
rect 12202 659 12242 665
rect 12276 659 12316 665
rect 12350 659 12390 665
rect 12424 659 12464 665
rect 12498 659 12538 665
rect 12572 659 12611 665
rect 12645 659 12684 665
rect 12718 659 12757 665
rect 12791 659 12838 665
rect 11314 629 12838 659
rect 11348 595 11385 629
rect 11419 595 11456 629
rect 11490 621 11527 629
rect 11561 621 11598 629
rect 11632 621 11669 629
rect 11703 621 11740 629
rect 11774 621 11811 629
rect 11845 621 11882 629
rect 11916 621 11953 629
rect 11987 621 12024 629
rect 12058 621 12095 629
rect 11490 595 11502 621
rect 11561 595 11576 621
rect 11632 595 11650 621
rect 11703 595 11724 621
rect 11774 595 11798 621
rect 11845 595 11872 621
rect 11916 595 11946 621
rect 11987 595 12020 621
rect 12058 595 12094 621
rect 12129 595 12166 629
rect 12200 621 12237 629
rect 12271 621 12308 629
rect 12342 621 12379 629
rect 12413 621 12450 629
rect 12484 621 12521 629
rect 12555 621 12592 629
rect 12626 621 12663 629
rect 12697 621 12734 629
rect 12768 621 12804 629
rect 12202 595 12237 621
rect 12276 595 12308 621
rect 12350 595 12379 621
rect 12424 595 12450 621
rect 12498 595 12521 621
rect 12572 595 12592 621
rect 12645 595 12663 621
rect 12718 595 12734 621
rect 12791 595 12804 621
rect 11314 587 11502 595
rect 11536 587 11576 595
rect 11610 587 11650 595
rect 11684 587 11724 595
rect 11758 587 11798 595
rect 11832 587 11872 595
rect 11906 587 11946 595
rect 11980 587 12020 595
rect 12054 587 12094 595
rect 12128 587 12168 595
rect 12202 587 12242 595
rect 12276 587 12316 595
rect 12350 587 12390 595
rect 12424 587 12464 595
rect 12498 587 12538 595
rect 12572 587 12611 595
rect 12645 587 12684 595
rect 12718 587 12757 595
rect 12791 587 12838 595
rect 11314 559 12838 587
rect 11348 525 11385 559
rect 11419 525 11456 559
rect 11490 549 11527 559
rect 11561 549 11598 559
rect 11632 549 11669 559
rect 11703 549 11740 559
rect 11774 549 11811 559
rect 11845 549 11882 559
rect 11916 549 11953 559
rect 11987 549 12024 559
rect 12058 549 12095 559
rect 11490 525 11502 549
rect 11561 525 11576 549
rect 11632 525 11650 549
rect 11703 525 11724 549
rect 11774 525 11798 549
rect 11845 525 11872 549
rect 11916 525 11946 549
rect 11987 525 12020 549
rect 12058 525 12094 549
rect 12129 525 12166 559
rect 12200 549 12237 559
rect 12271 549 12308 559
rect 12342 549 12379 559
rect 12413 549 12450 559
rect 12484 549 12521 559
rect 12555 549 12592 559
rect 12626 549 12663 559
rect 12697 549 12734 559
rect 12768 549 12804 559
rect 12202 525 12237 549
rect 12276 525 12308 549
rect 12350 525 12379 549
rect 12424 525 12450 549
rect 12498 525 12521 549
rect 12572 525 12592 549
rect 12645 525 12663 549
rect 12718 525 12734 549
rect 12791 525 12804 549
rect 11314 515 11502 525
rect 11536 515 11576 525
rect 11610 515 11650 525
rect 11684 515 11724 525
rect 11758 515 11798 525
rect 11832 515 11872 525
rect 11906 515 11946 525
rect 11980 515 12020 525
rect 12054 515 12094 525
rect 12128 515 12168 525
rect 12202 515 12242 525
rect 12276 515 12316 525
rect 12350 515 12390 525
rect 12424 515 12464 525
rect 12498 515 12538 525
rect 12572 515 12611 525
rect 12645 515 12684 525
rect 12718 515 12757 525
rect 12791 515 12838 525
rect 11314 489 12838 515
rect 11348 455 11385 489
rect 11419 455 11456 489
rect 11490 477 11527 489
rect 11561 477 11598 489
rect 11632 477 11669 489
rect 11703 477 11740 489
rect 11774 477 11811 489
rect 11845 477 11882 489
rect 11916 477 11953 489
rect 11987 477 12024 489
rect 12058 477 12095 489
rect 11490 455 11502 477
rect 11561 455 11576 477
rect 11632 455 11650 477
rect 11703 455 11724 477
rect 11774 455 11798 477
rect 11845 455 11872 477
rect 11916 455 11946 477
rect 11987 455 12020 477
rect 12058 455 12094 477
rect 12129 455 12166 489
rect 12200 477 12237 489
rect 12271 477 12308 489
rect 12342 477 12379 489
rect 12413 477 12450 489
rect 12484 477 12521 489
rect 12555 477 12592 489
rect 12626 477 12663 489
rect 12697 477 12734 489
rect 12768 477 12804 489
rect 12202 455 12237 477
rect 12276 455 12308 477
rect 12350 455 12379 477
rect 12424 455 12450 477
rect 12498 455 12521 477
rect 12572 455 12592 477
rect 12645 455 12663 477
rect 12718 455 12734 477
rect 12791 455 12804 477
rect 11314 443 11502 455
rect 11536 443 11576 455
rect 11610 443 11650 455
rect 11684 443 11724 455
rect 11758 443 11798 455
rect 11832 443 11872 455
rect 11906 443 11946 455
rect 11980 443 12020 455
rect 12054 443 12094 455
rect 12128 443 12168 455
rect 12202 443 12242 455
rect 12276 443 12316 455
rect 12350 443 12390 455
rect 12424 443 12464 455
rect 12498 443 12538 455
rect 12572 443 12611 455
rect 12645 443 12684 455
rect 12718 443 12757 455
rect 12791 443 12838 455
rect 11314 419 12838 443
rect 11348 385 11385 419
rect 11419 385 11456 419
rect 11490 405 11527 419
rect 11561 405 11598 419
rect 11632 405 11669 419
rect 11703 405 11740 419
rect 11774 405 11811 419
rect 11845 405 11882 419
rect 11916 405 11953 419
rect 11987 405 12024 419
rect 12058 405 12095 419
rect 11490 385 11502 405
rect 11561 385 11576 405
rect 11632 385 11650 405
rect 11703 385 11724 405
rect 11774 385 11798 405
rect 11845 385 11872 405
rect 11916 385 11946 405
rect 11987 385 12020 405
rect 12058 385 12094 405
rect 12129 385 12166 419
rect 12200 405 12237 419
rect 12271 405 12308 419
rect 12342 405 12379 419
rect 12413 405 12450 419
rect 12484 405 12521 419
rect 12555 405 12592 419
rect 12626 405 12663 419
rect 12697 405 12734 419
rect 12768 405 12804 419
rect 12202 385 12237 405
rect 12276 385 12308 405
rect 12350 385 12379 405
rect 12424 385 12450 405
rect 12498 385 12521 405
rect 12572 385 12592 405
rect 12645 385 12663 405
rect 12718 385 12734 405
rect 12791 385 12804 405
rect 11314 371 11502 385
rect 11536 371 11576 385
rect 11610 371 11650 385
rect 11684 371 11724 385
rect 11758 371 11798 385
rect 11832 371 11872 385
rect 11906 371 11946 385
rect 11980 371 12020 385
rect 12054 371 12094 385
rect 12128 371 12168 385
rect 12202 371 12242 385
rect 12276 371 12316 385
rect 12350 371 12390 385
rect 12424 371 12464 385
rect 12498 371 12538 385
rect 12572 371 12611 385
rect 12645 371 12684 385
rect 12718 371 12757 385
rect 12791 371 12838 385
rect 11314 349 12838 371
rect 11348 315 11385 349
rect 11419 315 11456 349
rect 11490 333 11527 349
rect 11561 333 11598 349
rect 11632 333 11669 349
rect 11703 333 11740 349
rect 11774 333 11811 349
rect 11845 333 11882 349
rect 11916 333 11953 349
rect 11987 333 12024 349
rect 12058 333 12095 349
rect 11490 315 11502 333
rect 11561 315 11576 333
rect 11632 315 11650 333
rect 11703 315 11724 333
rect 11774 315 11798 333
rect 11845 315 11872 333
rect 11916 315 11946 333
rect 11987 315 12020 333
rect 12058 315 12094 333
rect 12129 315 12166 349
rect 12200 333 12237 349
rect 12271 333 12308 349
rect 12342 333 12379 349
rect 12413 333 12450 349
rect 12484 333 12521 349
rect 12555 333 12592 349
rect 12626 333 12663 349
rect 12697 333 12734 349
rect 12768 333 12804 349
rect 12202 315 12237 333
rect 12276 315 12308 333
rect 12350 315 12379 333
rect 12424 315 12450 333
rect 12498 315 12521 333
rect 12572 315 12592 333
rect 12645 315 12663 333
rect 12718 315 12734 333
rect 12791 315 12804 333
rect 11314 299 11502 315
rect 11536 299 11576 315
rect 11610 299 11650 315
rect 11684 299 11724 315
rect 11758 299 11798 315
rect 11832 299 11872 315
rect 11906 299 11946 315
rect 11980 299 12020 315
rect 12054 299 12094 315
rect 12128 299 12168 315
rect 12202 299 12242 315
rect 12276 299 12316 315
rect 12350 299 12390 315
rect 12424 299 12464 315
rect 12498 299 12538 315
rect 12572 299 12611 315
rect 12645 299 12684 315
rect 12718 299 12757 315
rect 12791 299 12838 315
rect 11314 279 12838 299
rect 11348 245 11385 279
rect 11419 245 11456 279
rect 11490 261 11527 279
rect 11561 261 11598 279
rect 11632 261 11669 279
rect 11703 261 11740 279
rect 11774 261 11811 279
rect 11845 261 11882 279
rect 11916 261 11953 279
rect 11987 261 12024 279
rect 12058 261 12095 279
rect 11490 245 11502 261
rect 11561 245 11576 261
rect 11632 245 11650 261
rect 11703 245 11724 261
rect 11774 245 11798 261
rect 11845 245 11872 261
rect 11916 245 11946 261
rect 11987 245 12020 261
rect 12058 245 12094 261
rect 12129 245 12166 279
rect 12200 261 12237 279
rect 12271 261 12308 279
rect 12342 261 12379 279
rect 12413 261 12450 279
rect 12484 261 12521 279
rect 12555 261 12592 279
rect 12626 261 12663 279
rect 12697 261 12734 279
rect 12768 261 12804 279
rect 12202 245 12237 261
rect 12276 245 12308 261
rect 12350 245 12379 261
rect 12424 245 12450 261
rect 12498 245 12521 261
rect 12572 245 12592 261
rect 12645 245 12663 261
rect 12718 245 12734 261
rect 12791 245 12804 261
rect 11314 227 11502 245
rect 11536 227 11576 245
rect 11610 227 11650 245
rect 11684 227 11724 245
rect 11758 227 11798 245
rect 11832 227 11872 245
rect 11906 227 11946 245
rect 11980 227 12020 245
rect 12054 227 12094 245
rect 12128 227 12168 245
rect 12202 227 12242 245
rect 12276 227 12316 245
rect 12350 227 12390 245
rect 12424 227 12464 245
rect 12498 227 12538 245
rect 12572 227 12611 245
rect 12645 227 12684 245
rect 12718 227 12757 245
rect 12791 227 12838 245
rect 11314 209 12838 227
rect 11348 175 11385 209
rect 11419 175 11456 209
rect 11490 189 11527 209
rect 11561 189 11598 209
rect 11632 189 11669 209
rect 11703 189 11740 209
rect 11774 189 11811 209
rect 11845 189 11882 209
rect 11916 189 11953 209
rect 11987 189 12024 209
rect 12058 189 12095 209
rect 11490 175 11502 189
rect 11561 175 11576 189
rect 11632 175 11650 189
rect 11703 175 11724 189
rect 11774 175 11798 189
rect 11845 175 11872 189
rect 11916 175 11946 189
rect 11987 175 12020 189
rect 12058 175 12094 189
rect 12129 175 12166 209
rect 12200 189 12237 209
rect 12271 189 12308 209
rect 12342 189 12379 209
rect 12413 189 12450 209
rect 12484 189 12521 209
rect 12555 189 12592 209
rect 12626 189 12663 209
rect 12697 189 12734 209
rect 12768 189 12804 209
rect 12202 175 12237 189
rect 12276 175 12308 189
rect 12350 175 12379 189
rect 12424 175 12450 189
rect 12498 175 12521 189
rect 12572 175 12592 189
rect 12645 175 12663 189
rect 12718 175 12734 189
rect 12791 175 12804 189
rect 11314 155 11502 175
rect 11536 155 11576 175
rect 11610 155 11650 175
rect 11684 155 11724 175
rect 11758 155 11798 175
rect 11832 155 11872 175
rect 11906 155 11946 175
rect 11980 155 12020 175
rect 12054 155 12094 175
rect 12128 155 12168 175
rect 12202 155 12242 175
rect 12276 155 12316 175
rect 12350 155 12390 175
rect 12424 155 12464 175
rect 12498 155 12538 175
rect 12572 155 12611 175
rect 12645 155 12684 175
rect 12718 155 12757 175
rect 12791 155 12838 175
rect 11314 139 12838 155
rect 11348 105 11385 139
rect 11419 105 11456 139
rect 11490 117 11527 139
rect 11561 117 11598 139
rect 11632 117 11669 139
rect 11703 117 11740 139
rect 11774 117 11811 139
rect 11845 117 11882 139
rect 11916 117 11953 139
rect 11987 117 12024 139
rect 12058 117 12095 139
rect 11490 105 11502 117
rect 11561 105 11576 117
rect 11632 105 11650 117
rect 11703 105 11724 117
rect 11774 105 11798 117
rect 11845 105 11872 117
rect 11916 105 11946 117
rect 11987 105 12020 117
rect 12058 105 12094 117
rect 12129 105 12166 139
rect 12200 117 12237 139
rect 12271 117 12308 139
rect 12342 117 12379 139
rect 12413 117 12450 139
rect 12484 117 12521 139
rect 12555 117 12592 139
rect 12626 117 12663 139
rect 12697 117 12734 139
rect 12768 117 12804 139
rect 12202 105 12237 117
rect 12276 105 12308 117
rect 12350 105 12379 117
rect 12424 105 12450 117
rect 12498 105 12521 117
rect 12572 105 12592 117
rect 12645 105 12663 117
rect 12718 105 12734 117
rect 12791 105 12804 117
rect 11314 83 11502 105
rect 11536 83 11576 105
rect 11610 83 11650 105
rect 11684 83 11724 105
rect 11758 83 11798 105
rect 11832 83 11872 105
rect 11906 83 11946 105
rect 11980 83 12020 105
rect 12054 83 12094 105
rect 12128 83 12168 105
rect 12202 83 12242 105
rect 12276 83 12316 105
rect 12350 83 12390 105
rect 12424 83 12464 105
rect 12498 83 12538 105
rect 12572 83 12611 105
rect 12645 83 12684 105
rect 12718 83 12757 105
rect 12791 83 12838 105
rect 11314 69 12838 83
rect 11348 35 11385 69
rect 11419 35 11456 69
rect 11490 35 11527 69
rect 11561 35 11598 69
rect 11632 35 11669 69
rect 11703 35 11740 69
rect 11774 35 11811 69
rect 11845 35 11882 69
rect 11916 35 11953 69
rect 11987 35 12024 69
rect 12058 35 12095 69
rect 12129 35 12166 69
rect 12200 35 12237 69
rect 12271 35 12308 69
rect 12342 35 12379 69
rect 12413 35 12450 69
rect 12484 35 12521 69
rect 12555 35 12592 69
rect 12626 35 12663 69
rect 12697 35 12734 69
rect 12768 35 12804 69
rect 11314 15 12838 35
rect 11314 -1 11346 15
rect 11380 -1 11420 15
rect 11380 -19 11385 -1
rect 11348 -35 11385 -19
rect 11419 -19 11420 -1
rect 11454 -1 11494 15
rect 11528 -1 11567 15
rect 11601 -1 11640 15
rect 11674 -1 12838 15
rect 11454 -19 11456 -1
rect 11419 -35 11456 -19
rect 11490 -19 11494 -1
rect 11561 -19 11567 -1
rect 11632 -19 11640 -1
rect 11490 -35 11527 -19
rect 11561 -35 11598 -19
rect 11632 -35 11669 -19
rect 11703 -35 11740 -1
rect 11774 -35 11811 -1
rect 11845 -35 11882 -1
rect 11916 -35 11953 -1
rect 11987 -35 12024 -1
rect 12058 -35 12095 -1
rect 12129 -35 12166 -1
rect 12200 -35 12237 -1
rect 12271 -35 12308 -1
rect 12342 -35 12379 -1
rect 12413 -35 12450 -1
rect 12484 -35 12521 -1
rect 12555 -35 12592 -1
rect 12626 -35 12663 -1
rect 12697 -35 12734 -1
rect 12768 -35 12804 -1
rect 13193 865 13205 874
rect 13193 840 13239 865
rect 13227 826 13239 840
rect 13193 792 13205 806
rect 13193 772 13239 792
rect 13227 753 13239 772
rect 13193 719 13205 738
rect 13193 704 13239 719
rect 13227 680 13239 704
rect 13193 646 13205 670
rect 13193 636 13239 646
rect 13227 607 13239 636
rect 13193 573 13205 602
rect 13193 568 13239 573
rect 13227 534 13239 568
rect 13193 500 13205 534
rect 13227 466 13239 500
rect 13193 461 13239 466
rect 13193 432 13205 461
rect 13227 398 13239 427
rect 13193 388 13239 398
rect 13193 364 13205 388
rect 13227 330 13239 354
rect 13193 315 13239 330
rect 13193 296 13205 315
rect 13227 262 13239 281
rect 13193 242 13239 262
rect 13193 228 13205 242
rect 13433 2692 14745 2698
rect 13433 2658 13507 2692
rect 13545 2658 13575 2692
rect 13620 2658 13643 2692
rect 13695 2658 13711 2692
rect 13770 2658 13779 2692
rect 13845 2658 13847 2692
rect 13881 2658 13886 2692
rect 13949 2658 13961 2692
rect 14017 2658 14036 2692
rect 14085 2658 14111 2692
rect 14153 2658 14186 2692
rect 14221 2658 14255 2692
rect 14295 2658 14323 2692
rect 14369 2658 14391 2692
rect 14443 2658 14459 2692
rect 14517 2658 14527 2692
rect 14591 2658 14595 2692
rect 14629 2658 14631 2692
rect 14665 2658 14745 2692
rect 13433 2652 14745 2658
rect 13433 2592 13479 2652
rect 13433 2554 13439 2592
rect 13473 2554 13479 2592
rect 14699 2624 14745 2652
rect 14699 2586 14705 2624
rect 14739 2586 14745 2624
rect 13433 2520 13479 2554
rect 13684 2539 13700 2573
rect 13734 2539 13768 2573
rect 13802 2539 13836 2573
rect 13870 2539 13904 2573
rect 13938 2539 13972 2573
rect 14006 2539 14040 2573
rect 14074 2539 14108 2573
rect 14142 2539 14167 2573
rect 14210 2539 14240 2573
rect 14278 2539 14312 2573
rect 14346 2539 14380 2573
rect 14418 2539 14448 2573
rect 14490 2539 14516 2573
rect 14562 2539 14584 2573
rect 14699 2556 14745 2586
rect 13433 2458 13439 2520
rect 13473 2458 13479 2520
rect 13433 2452 13479 2458
rect 13433 2418 13439 2452
rect 13473 2418 13479 2452
rect 13433 2384 13479 2418
rect 13433 2348 13439 2384
rect 13473 2348 13479 2384
rect 13433 2316 13479 2348
rect 13433 2276 13439 2316
rect 13473 2276 13479 2316
rect 13433 2248 13479 2276
rect 13433 2204 13439 2248
rect 13473 2204 13479 2248
rect 13433 2180 13479 2204
rect 13433 2132 13439 2180
rect 13473 2132 13479 2180
rect 13433 2112 13479 2132
rect 13433 2060 13439 2112
rect 13473 2060 13479 2112
rect 13433 2044 13479 2060
rect 13433 1987 13439 2044
rect 13473 1987 13479 2044
rect 13433 1976 13479 1987
rect 13433 1914 13439 1976
rect 13473 1914 13479 1976
rect 13433 1908 13479 1914
rect 13433 1841 13439 1908
rect 13473 1841 13479 1908
rect 13433 1840 13479 1841
rect 13433 1806 13439 1840
rect 13473 1806 13479 1840
rect 13433 1802 13479 1806
rect 13433 1738 13439 1802
rect 13473 1738 13479 1802
rect 13433 1729 13479 1738
rect 13433 1670 13439 1729
rect 13473 1670 13479 1729
rect 13433 1656 13479 1670
rect 13433 1622 13439 1656
rect 13473 1622 13479 1656
rect 13433 1583 13479 1622
rect 13433 1528 13439 1583
rect 13473 1528 13479 1583
rect 13433 1510 13479 1528
rect 13433 1460 13439 1510
rect 13473 1460 13479 1510
rect 13433 1437 13479 1460
rect 13433 1392 13439 1437
rect 13473 1392 13479 1437
rect 13433 1364 13479 1392
rect 13433 1324 13439 1364
rect 13473 1324 13479 1364
rect 13433 1291 13479 1324
rect 13433 1256 13439 1291
rect 13473 1256 13479 1291
rect 13433 1222 13479 1256
rect 13433 1184 13439 1222
rect 13473 1184 13479 1222
rect 13433 1154 13479 1184
rect 13433 1111 13439 1154
rect 13473 1111 13479 1154
rect 13433 1086 13479 1111
rect 13433 1038 13439 1086
rect 13473 1038 13479 1086
rect 13433 1018 13479 1038
rect 13433 965 13439 1018
rect 13473 965 13479 1018
rect 13433 950 13479 965
rect 13433 892 13439 950
rect 13473 892 13479 950
rect 13433 882 13479 892
rect 13433 819 13439 882
rect 13473 819 13479 882
rect 13433 814 13479 819
rect 13433 712 13439 814
rect 13473 712 13479 814
rect 13433 707 13479 712
rect 13433 644 13439 707
rect 13473 644 13479 707
rect 13433 634 13479 644
rect 13433 576 13439 634
rect 13473 576 13479 634
rect 13433 561 13479 576
rect 13433 508 13439 561
rect 13473 508 13479 561
rect 13433 488 13479 508
rect 13433 440 13439 488
rect 13473 440 13479 488
rect 13433 415 13479 440
rect 13433 372 13439 415
rect 13473 372 13479 415
rect 13554 2516 13588 2528
rect 13554 2443 13588 2478
rect 14699 2512 14705 2556
rect 14739 2512 14745 2556
rect 14699 2488 14745 2512
rect 14699 2438 14705 2488
rect 14739 2438 14745 2488
rect 14699 2420 14745 2438
rect 13554 2374 13588 2409
rect 13734 2383 13757 2417
rect 13802 2383 13830 2417
rect 13870 2383 13903 2417
rect 13938 2383 13972 2417
rect 14009 2383 14040 2417
rect 14081 2383 14108 2417
rect 14142 2383 14176 2417
rect 14210 2383 14244 2417
rect 14278 2383 14312 2417
rect 14346 2383 14380 2417
rect 14414 2383 14448 2417
rect 14482 2383 14516 2417
rect 14550 2383 14584 2417
rect 14618 2383 14634 2417
rect 13554 2305 13588 2336
rect 13554 2236 13588 2263
rect 14699 2364 14705 2420
rect 14739 2364 14745 2420
rect 14699 2352 14745 2364
rect 14699 2290 14705 2352
rect 14739 2290 14745 2352
rect 14699 2284 14745 2290
rect 13684 2227 13700 2261
rect 13734 2227 13768 2261
rect 13802 2227 13836 2261
rect 13870 2227 13904 2261
rect 13938 2227 13972 2261
rect 14006 2227 14040 2261
rect 14074 2227 14108 2261
rect 14142 2227 14167 2261
rect 14210 2227 14240 2261
rect 14278 2227 14312 2261
rect 14346 2227 14380 2261
rect 14418 2227 14448 2261
rect 14490 2227 14516 2261
rect 14562 2227 14584 2261
rect 13554 2167 13588 2190
rect 13554 2098 13588 2116
rect 14699 2182 14705 2284
rect 14739 2182 14745 2284
rect 14699 2176 14745 2182
rect 14699 2114 14705 2176
rect 14739 2114 14745 2176
rect 13734 2071 13757 2105
rect 13802 2071 13830 2105
rect 13870 2071 13903 2105
rect 13938 2071 13972 2105
rect 14009 2071 14040 2105
rect 14081 2071 14108 2105
rect 14142 2071 14176 2105
rect 14210 2071 14244 2105
rect 14278 2071 14312 2105
rect 14346 2071 14380 2105
rect 14414 2071 14448 2105
rect 14482 2071 14516 2105
rect 14550 2071 14584 2105
rect 14618 2071 14634 2105
rect 14699 2102 14745 2114
rect 13554 2029 13588 2042
rect 13554 1960 13588 1968
rect 14699 2046 14705 2102
rect 14739 2046 14745 2102
rect 14699 2028 14745 2046
rect 14699 1978 14705 2028
rect 14739 1978 14745 2028
rect 14699 1954 14745 1978
rect 13684 1915 13700 1949
rect 13734 1915 13768 1949
rect 13802 1915 13836 1949
rect 13870 1915 13904 1949
rect 13938 1915 13972 1949
rect 14006 1915 14040 1949
rect 14074 1915 14108 1949
rect 14142 1915 14167 1949
rect 14210 1915 14240 1949
rect 14278 1915 14312 1949
rect 14346 1915 14380 1949
rect 14418 1915 14448 1949
rect 14490 1915 14516 1949
rect 14562 1915 14584 1949
rect 13554 1891 13588 1894
rect 13554 1854 13588 1857
rect 14699 1910 14705 1954
rect 14739 1910 14745 1954
rect 14699 1880 14745 1910
rect 14699 1842 14705 1880
rect 14739 1842 14745 1880
rect 14699 1808 14745 1842
rect 13554 1780 13588 1788
rect 13734 1759 13757 1793
rect 13802 1759 13830 1793
rect 13870 1759 13903 1793
rect 13938 1759 13972 1793
rect 14009 1759 14040 1793
rect 14081 1759 14108 1793
rect 14142 1759 14176 1793
rect 14210 1759 14244 1793
rect 14278 1759 14312 1793
rect 14346 1759 14380 1793
rect 14414 1759 14448 1793
rect 14482 1759 14516 1793
rect 14550 1759 14584 1793
rect 14618 1759 14634 1793
rect 14699 1772 14705 1808
rect 14739 1772 14745 1808
rect 13554 1706 13588 1719
rect 13554 1632 13588 1650
rect 14699 1740 14745 1772
rect 14699 1698 14705 1740
rect 14739 1698 14745 1740
rect 14699 1672 14745 1698
rect 13684 1603 13700 1637
rect 13734 1603 13768 1637
rect 13802 1603 13836 1637
rect 13870 1603 13904 1637
rect 13938 1603 13972 1637
rect 14006 1603 14040 1637
rect 14074 1603 14108 1637
rect 14142 1603 14167 1637
rect 14210 1603 14240 1637
rect 14278 1603 14312 1637
rect 14346 1603 14380 1637
rect 14418 1603 14448 1637
rect 14490 1603 14516 1637
rect 14562 1603 14584 1637
rect 14699 1624 14705 1672
rect 14739 1624 14745 1672
rect 14699 1604 14745 1624
rect 13554 1558 13588 1581
rect 13554 1484 13588 1512
rect 14699 1550 14705 1604
rect 14739 1550 14745 1604
rect 14699 1536 14745 1550
rect 13734 1447 13757 1481
rect 13802 1447 13830 1481
rect 13870 1447 13903 1481
rect 13938 1447 13972 1481
rect 14009 1447 14040 1481
rect 14081 1447 14108 1481
rect 14142 1447 14176 1481
rect 14210 1447 14244 1481
rect 14278 1447 14312 1481
rect 14346 1447 14380 1481
rect 14414 1447 14448 1481
rect 14482 1447 14516 1481
rect 14550 1447 14584 1481
rect 14618 1447 14634 1481
rect 14699 1477 14705 1536
rect 14739 1477 14745 1536
rect 14699 1468 14745 1477
rect 13554 1410 13588 1443
rect 13554 1339 13588 1374
rect 14699 1404 14705 1468
rect 14739 1404 14745 1468
rect 14699 1400 14745 1404
rect 14699 1366 14705 1400
rect 14739 1366 14745 1400
rect 14699 1365 14745 1366
rect 13554 1270 13588 1302
rect 13684 1291 13700 1325
rect 13734 1291 13768 1325
rect 13802 1291 13836 1325
rect 13870 1291 13904 1325
rect 13938 1291 13972 1325
rect 14006 1291 14040 1325
rect 14074 1291 14108 1325
rect 14142 1291 14167 1325
rect 14210 1291 14240 1325
rect 14278 1291 14312 1325
rect 14346 1291 14380 1325
rect 14418 1291 14448 1325
rect 14490 1291 14516 1325
rect 14562 1291 14584 1325
rect 14699 1298 14705 1365
rect 14739 1298 14745 1365
rect 14699 1292 14745 1298
rect 13554 1201 13588 1228
rect 14699 1230 14705 1292
rect 14739 1230 14745 1292
rect 14699 1219 14745 1230
rect 13554 1132 13588 1154
rect 13734 1135 13757 1169
rect 13802 1135 13830 1169
rect 13870 1135 13903 1169
rect 13938 1135 13972 1169
rect 14009 1135 14040 1169
rect 14081 1135 14108 1169
rect 14142 1135 14176 1169
rect 14210 1135 14244 1169
rect 14278 1135 14312 1169
rect 14346 1135 14380 1169
rect 14414 1135 14448 1169
rect 14482 1135 14516 1169
rect 14550 1135 14584 1169
rect 14618 1135 14634 1169
rect 14699 1162 14705 1219
rect 14739 1162 14745 1219
rect 14699 1146 14745 1162
rect 13554 1063 13588 1080
rect 14699 1094 14705 1146
rect 14739 1094 14745 1146
rect 14699 1073 14745 1094
rect 14699 1026 14705 1073
rect 14739 1026 14745 1073
rect 13554 994 13588 1006
rect 13684 979 13700 1013
rect 13734 979 13768 1013
rect 13802 979 13836 1013
rect 13870 979 13904 1013
rect 13938 979 13972 1013
rect 14006 979 14040 1013
rect 14074 979 14108 1013
rect 14142 979 14167 1013
rect 14210 979 14240 1013
rect 14278 979 14312 1013
rect 14346 979 14380 1013
rect 14418 979 14448 1013
rect 14490 979 14516 1013
rect 14562 979 14584 1013
rect 14699 1000 14745 1026
rect 13554 926 13588 932
rect 14699 958 14705 1000
rect 14739 958 14745 1000
rect 14699 927 14745 958
rect 14699 890 14705 927
rect 14739 890 14745 927
rect 13554 818 13588 824
rect 13734 823 13757 857
rect 13802 823 13830 857
rect 13870 823 13903 857
rect 13938 823 13972 857
rect 14009 823 14040 857
rect 14081 823 14108 857
rect 14142 823 14176 857
rect 14210 823 14244 857
rect 14278 823 14312 857
rect 14346 823 14380 857
rect 14414 823 14448 857
rect 14482 823 14516 857
rect 14550 823 14584 857
rect 14618 823 14634 857
rect 14699 856 14745 890
rect 13554 744 13588 756
rect 14699 820 14705 856
rect 14739 820 14745 856
rect 14699 788 14745 820
rect 14699 747 14705 788
rect 14739 747 14745 788
rect 14699 720 14745 747
rect 13554 670 13588 688
rect 13684 667 13700 701
rect 13734 667 13768 701
rect 13802 667 13836 701
rect 13870 667 13904 701
rect 13938 667 13972 701
rect 14006 667 14040 701
rect 14074 667 14108 701
rect 14142 667 14167 701
rect 14210 667 14240 701
rect 14278 667 14312 701
rect 14346 667 14380 701
rect 14418 667 14448 701
rect 14490 667 14516 701
rect 14562 667 14584 701
rect 14699 674 14705 720
rect 14739 674 14745 720
rect 13554 596 13588 620
rect 13554 522 13588 552
rect 14699 652 14745 674
rect 14699 601 14705 652
rect 14739 601 14745 652
rect 14699 584 14745 601
rect 13734 511 13757 545
rect 13802 511 13830 545
rect 13870 511 13903 545
rect 13938 511 13972 545
rect 14009 511 14040 545
rect 14081 511 14108 545
rect 14142 511 14176 545
rect 14210 511 14244 545
rect 14278 511 14312 545
rect 14346 511 14380 545
rect 14414 511 14448 545
rect 14482 511 14516 545
rect 14550 511 14584 545
rect 14618 511 14634 545
rect 14699 528 14705 584
rect 14739 528 14745 584
rect 14699 516 14745 528
rect 13554 450 13588 484
rect 13554 400 13588 416
rect 14699 455 14705 516
rect 14739 455 14745 516
rect 14699 448 14745 455
rect 13433 342 13479 372
rect 13684 355 13700 389
rect 13734 355 13768 389
rect 13802 355 13836 389
rect 13870 355 13904 389
rect 13938 355 13972 389
rect 14006 355 14040 389
rect 14074 355 14108 389
rect 14142 355 14167 389
rect 14210 355 14240 389
rect 14278 355 14312 389
rect 14346 355 14380 389
rect 14418 355 14448 389
rect 14490 355 14516 389
rect 14562 355 14584 389
rect 14699 382 14705 448
rect 14739 382 14745 448
rect 14699 380 14745 382
rect 13433 304 13439 342
rect 13473 304 13479 342
rect 13433 276 13479 304
rect 14699 346 14705 380
rect 14739 346 14745 380
rect 14699 343 14745 346
rect 14699 309 14705 343
rect 14739 309 14745 343
rect 14699 276 14745 309
rect 13433 270 14745 276
rect 13433 236 13513 270
rect 13547 236 13549 270
rect 13583 236 13587 270
rect 13651 236 13661 270
rect 13719 236 13735 270
rect 13787 236 13809 270
rect 13855 236 13883 270
rect 13923 236 13957 270
rect 13992 236 14025 270
rect 14067 236 14093 270
rect 14142 236 14161 270
rect 14217 236 14229 270
rect 14292 236 14297 270
rect 14331 236 14333 270
rect 14399 236 14408 270
rect 14467 236 14483 270
rect 14535 236 14558 270
rect 14603 236 14633 270
rect 14671 236 14745 270
rect 13433 230 14745 236
rect 14983 2670 15017 2674
rect 14983 2635 15017 2636
rect 14983 2562 15017 2568
rect 14983 2489 15017 2500
rect 14983 2416 15017 2432
rect 14983 2343 15017 2364
rect 14983 2270 15017 2296
rect 14983 2197 15017 2228
rect 14983 2126 15017 2160
rect 14983 2058 15017 2090
rect 14983 1990 15017 2017
rect 14983 1922 15017 1944
rect 14983 1854 15017 1871
rect 14983 1786 15017 1798
rect 14983 1718 15017 1725
rect 14983 1650 15017 1652
rect 14983 1613 15017 1616
rect 14983 1540 15017 1548
rect 14983 1467 15017 1480
rect 14983 1394 15017 1412
rect 14983 1321 15017 1344
rect 14983 1248 15017 1276
rect 14983 1176 15017 1208
rect 14983 1106 15017 1140
rect 14983 1038 15017 1070
rect 14983 970 15017 998
rect 14983 902 15017 926
rect 14983 834 15017 854
rect 14983 766 15017 782
rect 14983 698 15017 710
rect 14983 630 15017 638
rect 14983 562 15017 566
rect 14983 456 15017 460
rect 14983 384 15017 392
rect 14983 312 15017 324
rect 14983 240 15017 256
rect 13227 194 13239 208
rect 13193 169 13239 194
rect 13193 160 13205 169
rect 13227 126 13239 135
rect 13193 96 13239 126
rect 13193 92 13205 96
rect 13227 58 13239 62
rect 13193 45 13239 58
rect 14983 168 15017 188
rect 14983 96 15017 120
rect 14983 45 15017 52
rect 13193 24 15017 45
rect 13193 -10 13279 24
rect 13317 -10 13351 24
rect 13387 -10 13419 24
rect 13461 -10 13487 24
rect 13535 -10 13555 24
rect 13609 -10 13623 24
rect 13683 -10 13691 24
rect 13757 -10 13759 24
rect 13793 -10 13797 24
rect 13861 -10 13871 24
rect 13929 -10 13945 24
rect 13997 -10 14019 24
rect 14065 -10 14093 24
rect 14133 -10 14167 24
rect 14201 -10 14235 24
rect 14275 -10 14303 24
rect 14349 -10 14371 24
rect 14423 -10 14439 24
rect 14497 -10 14507 24
rect 14571 -10 14575 24
rect 14609 -10 14611 24
rect 14677 -10 14686 24
rect 14745 -10 14761 24
rect 14813 -10 14836 24
rect 14881 -10 14911 24
rect 14949 -10 15017 24
rect 11314 -57 12838 -35
rect 11314 -62 11346 -57
rect 5776 -128 5810 -65
rect 6128 -128 6162 -65
rect 8037 -96 8071 -62
rect 8105 -96 8141 -62
rect 8175 -96 8211 -62
rect 8245 -96 8281 -62
rect 8315 -96 8351 -62
rect 8385 -96 8421 -62
rect 8455 -96 8491 -62
rect 8525 -96 8561 -62
rect 8595 -96 8631 -62
rect 8665 -96 8701 -62
rect 8735 -96 8771 -62
rect 8805 -96 8841 -62
rect 8875 -96 8911 -62
rect 8945 -96 8981 -62
rect 9015 -96 9051 -62
rect 9085 -96 9121 -62
rect 9155 -96 9191 -62
rect 9225 -96 9261 -62
rect 9295 -96 9331 -62
rect 9365 -96 9401 -62
rect 9435 -96 9471 -62
rect 9505 -96 9541 -62
rect 9575 -96 9611 -62
rect 9645 -96 9681 -62
rect 9715 -96 9751 -62
rect 9785 -96 9821 -62
rect 9855 -96 9891 -62
rect 9925 -96 9961 -62
rect 9995 -96 10031 -62
rect 10065 -96 10101 -62
rect 10135 -96 10170 -62
rect 10204 -96 10239 -62
rect 10273 -96 10308 -62
rect 10342 -96 10377 -62
rect 10411 -96 10446 -62
rect 10480 -96 10515 -62
rect 10549 -96 10583 -62
rect 11072 -71 11346 -62
rect 11380 -71 11420 -57
rect 11072 -96 11314 -71
rect 11380 -91 11385 -71
rect 7548 -105 11314 -96
rect 11348 -105 11385 -91
rect 11419 -91 11420 -71
rect 11454 -71 11494 -57
rect 11528 -71 11567 -57
rect 11601 -71 11640 -57
rect 11674 -71 12838 -57
rect 11454 -91 11456 -71
rect 11419 -105 11456 -91
rect 11490 -91 11494 -71
rect 11561 -91 11567 -71
rect 11632 -91 11640 -71
rect 11490 -105 11527 -91
rect 11561 -105 11598 -91
rect 11632 -105 11669 -91
rect 11703 -105 11740 -71
rect 11774 -105 11811 -71
rect 11845 -105 11882 -71
rect 11916 -105 11953 -71
rect 11987 -105 12024 -71
rect 12058 -105 12095 -71
rect 12129 -105 12166 -71
rect 12200 -105 12237 -71
rect 12271 -105 12308 -71
rect 12342 -105 12379 -71
rect 12413 -105 12450 -71
rect 12484 -105 12521 -71
rect 12555 -105 12592 -71
rect 12626 -105 12663 -71
rect 12697 -105 12734 -71
rect 12768 -105 12804 -71
rect 7548 -128 12838 -105
rect 5735 -140 12838 -128
rect 5735 -174 5769 -140
rect 5803 -174 5838 -140
rect 5872 -174 5907 -140
rect 5941 -174 5976 -140
rect 6010 -174 6045 -140
rect 6079 -174 6114 -140
rect 6148 -174 6183 -140
rect 6217 -174 6252 -140
rect 6286 -174 6321 -140
rect 6355 -174 6390 -140
rect 6424 -174 6459 -140
rect 6493 -174 6528 -140
rect 6562 -174 6597 -140
rect 6631 -174 6666 -140
rect 6700 -174 6735 -140
rect 6769 -174 6804 -140
rect 6838 -174 6873 -140
rect 6907 -174 6942 -140
rect 6976 -174 7011 -140
rect 7045 -174 7080 -140
rect 7114 -174 7149 -140
rect 7183 -174 7218 -140
rect 7252 -174 7287 -140
rect 7321 -174 7356 -140
rect 7390 -174 7425 -140
rect 7459 -174 7494 -140
rect 7528 -174 7563 -140
rect 7597 -174 7632 -140
rect 7666 -174 7701 -140
rect 7735 -174 7770 -140
rect 7804 -174 7839 -140
rect 7873 -174 7908 -140
rect 7942 -174 7977 -140
rect 8011 -174 8046 -140
rect 8080 -174 8115 -140
rect 8149 -174 8184 -140
rect 8218 -174 8253 -140
rect 8287 -174 8322 -140
rect 8356 -174 8390 -140
rect 8424 -174 8458 -140
rect 8492 -174 8526 -140
rect 8560 -174 8594 -140
rect 8628 -174 8662 -140
rect 8696 -174 8730 -140
rect 8764 -174 8798 -140
rect 8832 -174 8866 -140
rect 8900 -174 8934 -140
rect 8968 -174 9002 -140
rect 9036 -174 9070 -140
rect 9104 -174 9138 -140
rect 9172 -174 9206 -140
rect 9240 -174 9274 -140
rect 9308 -174 9342 -140
rect 9376 -174 9410 -140
rect 9444 -174 9478 -140
rect 9512 -174 9546 -140
rect 9580 -174 9614 -140
rect 9648 -174 9682 -140
rect 9716 -174 9750 -140
rect 9784 -174 9818 -140
rect 9852 -174 9886 -140
rect 9920 -174 9954 -140
rect 9988 -174 10022 -140
rect 10056 -174 10090 -140
rect 10124 -174 10158 -140
rect 10192 -174 10226 -140
rect 10260 -174 10294 -140
rect 10328 -174 10362 -140
rect 10396 -174 10430 -140
rect 10464 -174 10498 -140
rect 10532 -174 10566 -140
rect 10600 -174 10634 -140
rect 10668 -174 10702 -140
rect 10736 -174 10770 -140
rect 10804 -174 10838 -140
rect 10872 -174 10906 -140
rect 10940 -174 10974 -140
rect 11008 -174 11042 -140
rect 11076 -174 11110 -140
rect 11144 -174 11178 -140
rect 11212 -174 11246 -140
rect 11280 -141 12838 -140
rect 11280 -174 11314 -141
rect 5735 -175 11314 -174
rect 11348 -175 11385 -141
rect 11419 -175 11456 -141
rect 11490 -175 11527 -141
rect 11561 -175 11598 -141
rect 11632 -175 11669 -141
rect 11703 -175 11740 -141
rect 11774 -175 11811 -141
rect 11845 -175 11882 -141
rect 11916 -175 11953 -141
rect 11987 -175 12024 -141
rect 12058 -175 12095 -141
rect 12129 -175 12166 -141
rect 12200 -175 12237 -141
rect 12271 -175 12308 -141
rect 12342 -175 12379 -141
rect 12413 -175 12450 -141
rect 12484 -175 12521 -141
rect 12555 -175 12592 -141
rect 12626 -175 12663 -141
rect 12697 -175 12734 -141
rect 12768 -175 12804 -141
rect 5735 -215 12838 -175
rect 5735 -249 11332 -215
rect 12277 -255 12831 -215
rect 12277 -289 12316 -255
rect 12350 -289 12384 -255
rect 12418 -289 12452 -255
rect 12486 -289 12520 -255
rect 12554 -289 12588 -255
rect 12622 -289 12656 -255
rect 12690 -289 12724 -255
rect 12758 -289 12831 -255
rect 12277 -325 12831 -289
rect 12277 -359 12316 -325
rect 12350 -359 12384 -325
rect 12418 -359 12452 -325
rect 12486 -359 12520 -325
rect 12554 -359 12588 -325
rect 12622 -359 12656 -325
rect 12690 -359 12724 -325
rect 12758 -359 12831 -325
rect 12277 -395 12831 -359
rect 12277 -429 12316 -395
rect 12350 -429 12384 -395
rect 12418 -429 12452 -395
rect 12486 -429 12520 -395
rect 12554 -429 12588 -395
rect 12622 -429 12656 -395
rect 12690 -429 12724 -395
rect 12758 -429 12831 -395
rect 12277 -465 12831 -429
rect 12277 -499 12316 -465
rect 12350 -499 12384 -465
rect 12418 -499 12452 -465
rect 12486 -499 12520 -465
rect 12554 -499 12588 -465
rect 12622 -499 12656 -465
rect 12690 -499 12724 -465
rect 12758 -499 12831 -465
rect 12277 -507 12831 -499
rect 12277 -535 12797 -507
rect 12277 -569 12316 -535
rect 12350 -569 12384 -535
rect 12418 -569 12452 -535
rect 12486 -569 12520 -535
rect 12554 -569 12588 -535
rect 12622 -569 12656 -535
rect 12690 -569 12724 -535
rect 12758 -569 12797 -535
rect 12277 -606 12797 -569
rect 12277 -640 12316 -606
rect 12350 -640 12384 -606
rect 12418 -640 12452 -606
rect 12486 -640 12520 -606
rect 12554 -640 12588 -606
rect 12622 -640 12656 -606
rect 12690 -640 12724 -606
rect 12758 -640 12797 -606
rect 12277 -677 12797 -640
rect 12277 -711 12316 -677
rect 12350 -711 12384 -677
rect 12418 -711 12452 -677
rect 12486 -711 12520 -677
rect 12554 -711 12588 -677
rect 12622 -711 12656 -677
rect 12690 -711 12724 -677
rect 12758 -711 12797 -677
rect 12277 -748 12797 -711
rect 12277 -782 12316 -748
rect 12350 -768 12384 -748
rect 12418 -768 12452 -748
rect 12486 -768 12520 -748
rect 12554 -768 12588 -748
rect 12356 -782 12384 -768
rect 12433 -782 12452 -768
rect 12509 -782 12520 -768
rect 12585 -782 12588 -768
rect 12622 -768 12656 -748
rect 12690 -768 12724 -748
rect 12622 -782 12627 -768
rect 12690 -782 12703 -768
rect 12758 -782 12797 -748
rect 12277 -802 12322 -782
rect 12356 -802 12399 -782
rect 12433 -802 12475 -782
rect 12509 -802 12551 -782
rect 12585 -802 12627 -782
rect 12661 -802 12703 -782
rect 12737 -802 12797 -782
rect 12277 -819 12797 -802
rect 12277 -853 12316 -819
rect 12350 -840 12384 -819
rect 12418 -840 12452 -819
rect 12486 -840 12520 -819
rect 12554 -840 12588 -819
rect 12356 -853 12384 -840
rect 12433 -853 12452 -840
rect 12509 -853 12520 -840
rect 12585 -853 12588 -840
rect 12622 -840 12656 -819
rect 12690 -840 12724 -819
rect 12622 -853 12627 -840
rect 12690 -853 12703 -840
rect 12758 -853 12797 -819
rect 12277 -874 12322 -853
rect 12356 -874 12399 -853
rect 12433 -874 12475 -853
rect 12509 -874 12551 -853
rect 12585 -874 12627 -853
rect 12661 -874 12703 -853
rect 12737 -874 12797 -853
rect 12277 -890 12797 -874
rect 12277 -924 12316 -890
rect 12350 -912 12384 -890
rect 12418 -912 12452 -890
rect 12486 -912 12520 -890
rect 12554 -912 12588 -890
rect 12356 -924 12384 -912
rect 12433 -924 12452 -912
rect 12509 -924 12520 -912
rect 12585 -924 12588 -912
rect 12622 -912 12656 -890
rect 12690 -912 12724 -890
rect 12622 -924 12627 -912
rect 12690 -924 12703 -912
rect 12758 -924 12797 -890
rect 12277 -946 12322 -924
rect 12356 -946 12399 -924
rect 12433 -946 12475 -924
rect 12509 -946 12551 -924
rect 12585 -946 12627 -924
rect 12661 -946 12703 -924
rect 12737 -946 12797 -924
rect 12277 -961 12797 -946
rect 12277 -995 12316 -961
rect 12350 -995 12384 -961
rect 12418 -995 12452 -961
rect 12486 -995 12520 -961
rect 12554 -995 12588 -961
rect 12622 -995 12656 -961
rect 12690 -995 12724 -961
rect 12758 -995 12797 -961
<< viali >>
rect 7826 9779 7860 9813
rect 7942 9779 7976 9813
rect 7826 9705 7860 9739
rect 7942 9705 7976 9739
rect 9357 9779 9391 9813
rect 9473 9779 9507 9813
rect 7826 9631 7860 9665
rect 7942 9631 7976 9665
rect 7826 9557 7860 9591
rect 7942 9557 7976 9591
rect 7826 9483 7860 9517
rect 7942 9483 7976 9517
rect 9357 9705 9391 9739
rect 9473 9705 9507 9739
rect 9357 9631 9391 9665
rect 9473 9631 9507 9665
rect 9357 9557 9391 9591
rect 9473 9557 9507 9591
rect 7826 9409 7860 9443
rect 7942 9409 7976 9443
rect 9357 9483 9391 9517
rect 9473 9483 9507 9517
rect 9357 9409 9391 9443
rect 9473 9409 9507 9443
rect 800 8767 834 8779
rect 800 8745 834 8767
rect 911 8757 941 8791
rect 941 8757 945 8791
rect 983 8757 1009 8791
rect 1009 8757 1017 8791
rect 1055 8757 1077 8791
rect 1077 8757 1089 8791
rect 1127 8757 1145 8791
rect 1145 8757 1161 8791
rect 1199 8757 1213 8791
rect 1213 8757 1233 8791
rect 1271 8757 1281 8791
rect 1281 8757 1305 8791
rect 1343 8757 1349 8791
rect 1349 8757 1377 8791
rect 1415 8757 1417 8791
rect 1417 8757 1449 8791
rect 1487 8757 1519 8791
rect 1519 8757 1521 8791
rect 1559 8757 1587 8791
rect 1587 8757 1593 8791
rect 1631 8757 1655 8791
rect 1655 8757 1665 8791
rect 1703 8757 1723 8791
rect 1723 8757 1737 8791
rect 1775 8757 1791 8791
rect 1791 8757 1809 8791
rect 1847 8757 1859 8791
rect 1859 8757 1881 8791
rect 1919 8757 1927 8791
rect 1927 8757 1953 8791
rect 1991 8757 1995 8791
rect 1995 8757 2025 8791
rect 2063 8757 2097 8791
rect 2135 8757 2165 8791
rect 2165 8757 2169 8791
rect 2207 8757 2233 8791
rect 2233 8757 2241 8791
rect 2279 8757 2301 8791
rect 2301 8757 2313 8791
rect 2351 8757 2369 8791
rect 2369 8757 2385 8791
rect 2423 8757 2437 8791
rect 2437 8757 2457 8791
rect 2495 8757 2505 8791
rect 2505 8757 2529 8791
rect 2567 8757 2573 8791
rect 2573 8757 2601 8791
rect 2639 8757 2641 8791
rect 2641 8757 2673 8791
rect 2711 8757 2743 8791
rect 2743 8757 2745 8791
rect 2783 8757 2811 8791
rect 2811 8757 2817 8791
rect 2855 8757 2879 8791
rect 2879 8757 2889 8791
rect 2927 8757 2947 8791
rect 2947 8757 2961 8791
rect 2999 8757 3015 8791
rect 3015 8757 3033 8791
rect 3071 8757 3083 8791
rect 3083 8757 3105 8791
rect 3143 8757 3151 8791
rect 3151 8757 3177 8791
rect 3215 8757 3219 8791
rect 3219 8757 3249 8791
rect 3287 8757 3321 8791
rect 3359 8757 3389 8791
rect 3389 8757 3393 8791
rect 3431 8757 3457 8791
rect 3457 8757 3465 8791
rect 3503 8757 3525 8791
rect 3525 8757 3537 8791
rect 3575 8757 3593 8791
rect 3593 8757 3609 8791
rect 3647 8757 3661 8791
rect 3661 8757 3681 8791
rect 3719 8757 3729 8791
rect 3729 8757 3753 8791
rect 3791 8757 3797 8791
rect 3797 8757 3825 8791
rect 3863 8757 3865 8791
rect 3865 8757 3897 8791
rect 3935 8757 3967 8791
rect 3967 8757 3969 8791
rect 4007 8757 4035 8791
rect 4035 8757 4041 8791
rect 4079 8757 4103 8791
rect 4103 8757 4113 8791
rect 4151 8757 4171 8791
rect 4171 8757 4185 8791
rect 4223 8757 4239 8791
rect 4239 8757 4257 8791
rect 4295 8757 4307 8791
rect 4307 8757 4329 8791
rect 4367 8757 4375 8791
rect 4375 8757 4401 8791
rect 4439 8757 4443 8791
rect 4443 8757 4473 8791
rect 4511 8757 4545 8791
rect 4583 8757 4613 8791
rect 4613 8757 4617 8791
rect 4655 8757 4681 8791
rect 4681 8757 4689 8791
rect 4727 8766 4749 8791
rect 4749 8766 4761 8791
rect 4727 8757 4731 8766
rect 4731 8757 4761 8766
rect 800 8699 834 8707
rect 800 8673 834 8699
rect 800 8631 834 8635
rect 800 8601 834 8631
rect 800 8529 834 8563
rect 800 8461 834 8491
rect 800 8457 834 8461
rect 800 8393 834 8419
rect 800 8385 834 8393
rect 800 8325 834 8347
rect 800 8313 834 8325
rect 800 8257 834 8275
rect 800 8241 834 8257
rect 800 8189 834 8203
rect 800 8169 834 8189
rect 800 8121 834 8131
rect 800 8097 834 8121
rect 800 8053 834 8059
rect 800 8025 834 8053
rect 800 7985 834 7987
rect 800 7953 834 7985
rect 800 7883 834 7915
rect 800 7881 834 7883
rect 800 7815 834 7843
rect 800 7809 834 7815
rect 800 7747 834 7771
rect 800 7737 834 7747
rect 800 7679 834 7699
rect 800 7665 834 7679
rect 800 7611 834 7627
rect 800 7593 834 7611
rect 800 7543 834 7555
rect 800 7521 834 7543
rect 800 7475 834 7483
rect 800 7449 834 7475
rect 800 7407 834 7411
rect 800 7377 834 7407
rect 800 7305 834 7339
rect 800 7237 834 7267
rect 800 7233 834 7237
rect 1173 8552 1207 8586
rect 1245 8579 1279 8586
rect 1317 8579 1351 8586
rect 1389 8579 1423 8586
rect 1461 8579 1495 8586
rect 1533 8579 1567 8586
rect 1605 8579 1639 8586
rect 1677 8579 1711 8586
rect 1749 8579 1783 8586
rect 1821 8579 1855 8586
rect 1893 8579 1927 8586
rect 1965 8579 1999 8586
rect 2037 8579 2071 8586
rect 2109 8579 2143 8586
rect 2181 8579 2215 8586
rect 2253 8579 2287 8586
rect 2325 8579 2359 8586
rect 2397 8579 2431 8586
rect 2469 8579 2503 8586
rect 2541 8579 2575 8586
rect 2613 8579 2647 8586
rect 2685 8579 2719 8586
rect 2757 8579 2791 8586
rect 2829 8579 2863 8586
rect 2901 8579 2935 8586
rect 2973 8579 3007 8586
rect 3045 8579 3079 8586
rect 3117 8579 3151 8586
rect 3189 8579 3223 8586
rect 3261 8579 3295 8586
rect 3333 8579 3367 8586
rect 3405 8579 3439 8586
rect 3477 8579 3511 8586
rect 3549 8579 3583 8586
rect 3621 8579 3655 8586
rect 3693 8579 3727 8586
rect 3765 8579 3799 8586
rect 3837 8579 3871 8586
rect 3909 8579 3943 8586
rect 3981 8579 4015 8586
rect 4053 8579 4087 8586
rect 4125 8579 4159 8586
rect 4197 8579 4231 8586
rect 4269 8579 4303 8586
rect 1245 8552 1268 8579
rect 1268 8552 1279 8579
rect 1317 8552 1336 8579
rect 1336 8552 1351 8579
rect 1389 8552 1404 8579
rect 1404 8552 1423 8579
rect 1461 8552 1472 8579
rect 1472 8552 1495 8579
rect 1533 8552 1540 8579
rect 1540 8552 1567 8579
rect 1605 8552 1608 8579
rect 1608 8552 1639 8579
rect 1677 8552 1710 8579
rect 1710 8552 1711 8579
rect 1749 8552 1778 8579
rect 1778 8552 1783 8579
rect 1821 8552 1846 8579
rect 1846 8552 1855 8579
rect 1893 8552 1914 8579
rect 1914 8552 1927 8579
rect 1965 8552 1982 8579
rect 1982 8552 1999 8579
rect 2037 8552 2050 8579
rect 2050 8552 2071 8579
rect 2109 8552 2118 8579
rect 2118 8552 2143 8579
rect 2181 8552 2186 8579
rect 2186 8552 2215 8579
rect 2253 8552 2254 8579
rect 2254 8552 2287 8579
rect 2325 8552 2356 8579
rect 2356 8552 2359 8579
rect 2397 8552 2424 8579
rect 2424 8552 2431 8579
rect 2469 8552 2492 8579
rect 2492 8552 2503 8579
rect 2541 8552 2560 8579
rect 2560 8552 2575 8579
rect 2613 8552 2628 8579
rect 2628 8552 2647 8579
rect 2685 8552 2696 8579
rect 2696 8552 2719 8579
rect 2757 8552 2764 8579
rect 2764 8552 2791 8579
rect 2829 8552 2832 8579
rect 2832 8552 2863 8579
rect 2901 8552 2934 8579
rect 2934 8552 2935 8579
rect 2973 8552 3002 8579
rect 3002 8552 3007 8579
rect 3045 8552 3070 8579
rect 3070 8552 3079 8579
rect 3117 8552 3138 8579
rect 3138 8552 3151 8579
rect 3189 8552 3206 8579
rect 3206 8552 3223 8579
rect 3261 8552 3274 8579
rect 3274 8552 3295 8579
rect 3333 8552 3342 8579
rect 3342 8552 3367 8579
rect 3405 8552 3410 8579
rect 3410 8552 3439 8579
rect 3477 8552 3478 8579
rect 3478 8552 3511 8579
rect 3549 8552 3580 8579
rect 3580 8552 3583 8579
rect 3621 8552 3648 8579
rect 3648 8552 3655 8579
rect 3693 8552 3716 8579
rect 3716 8552 3727 8579
rect 3765 8552 3784 8579
rect 3784 8552 3799 8579
rect 3837 8552 3852 8579
rect 3852 8552 3871 8579
rect 3909 8552 3920 8579
rect 3920 8552 3943 8579
rect 3981 8552 3988 8579
rect 3988 8552 4015 8579
rect 4053 8552 4056 8579
rect 4056 8552 4087 8579
rect 4125 8552 4158 8579
rect 4158 8552 4159 8579
rect 4197 8552 4226 8579
rect 4226 8552 4231 8579
rect 4269 8552 4294 8579
rect 4294 8552 4303 8579
rect 4341 8552 4375 8586
rect 4474 8546 4508 8580
rect 1167 8489 1201 8496
rect 1167 8462 1201 8489
rect 4474 8474 4508 8508
rect 1294 8438 1328 8472
rect 1366 8438 1396 8472
rect 1396 8438 1400 8472
rect 1438 8438 1464 8472
rect 1464 8438 1472 8472
rect 1510 8438 1532 8472
rect 1532 8438 1544 8472
rect 1582 8438 1600 8472
rect 1600 8438 1616 8472
rect 1654 8438 1668 8472
rect 1668 8438 1688 8472
rect 1726 8438 1736 8472
rect 1736 8438 1760 8472
rect 1798 8438 1804 8472
rect 1804 8438 1832 8472
rect 1870 8438 1872 8472
rect 1872 8438 1904 8472
rect 1942 8438 1974 8472
rect 1974 8438 1976 8472
rect 2014 8438 2042 8472
rect 2042 8438 2048 8472
rect 2086 8438 2110 8472
rect 2110 8438 2120 8472
rect 2158 8438 2178 8472
rect 2178 8438 2192 8472
rect 2230 8438 2246 8472
rect 2246 8438 2264 8472
rect 2302 8438 2314 8472
rect 2314 8438 2336 8472
rect 2374 8438 2382 8472
rect 2382 8438 2408 8472
rect 2446 8438 2450 8472
rect 2450 8438 2480 8472
rect 2518 8438 2552 8472
rect 2590 8438 2620 8472
rect 2620 8438 2624 8472
rect 2662 8438 2688 8472
rect 2688 8438 2696 8472
rect 2734 8438 2756 8472
rect 2756 8438 2768 8472
rect 2806 8438 2824 8472
rect 2824 8438 2840 8472
rect 2878 8438 2892 8472
rect 2892 8438 2912 8472
rect 2950 8438 2960 8472
rect 2960 8438 2984 8472
rect 3022 8438 3028 8472
rect 3028 8438 3056 8472
rect 3094 8438 3096 8472
rect 3096 8438 3128 8472
rect 3166 8438 3198 8472
rect 3198 8438 3200 8472
rect 3238 8438 3266 8472
rect 3266 8438 3272 8472
rect 3310 8438 3334 8472
rect 3334 8438 3344 8472
rect 3382 8438 3402 8472
rect 3402 8438 3416 8472
rect 3454 8438 3470 8472
rect 3470 8438 3488 8472
rect 3526 8438 3538 8472
rect 3538 8438 3560 8472
rect 3598 8438 3606 8472
rect 3606 8438 3632 8472
rect 3670 8438 3674 8472
rect 3674 8438 3704 8472
rect 3742 8438 3776 8472
rect 3814 8438 3844 8472
rect 3844 8438 3848 8472
rect 3886 8438 3912 8472
rect 3912 8438 3920 8472
rect 3958 8438 3980 8472
rect 3980 8438 3992 8472
rect 4030 8438 4048 8472
rect 4048 8438 4064 8472
rect 4102 8438 4116 8472
rect 4116 8438 4136 8472
rect 4174 8438 4184 8472
rect 4184 8438 4208 8472
rect 1167 8421 1201 8424
rect 1167 8390 1201 8421
rect 1167 8319 1201 8352
rect 1167 8318 1201 8319
rect 4330 8405 4364 8415
rect 4330 8381 4364 8405
rect 4330 8337 4364 8338
rect 1167 8251 1201 8280
rect 1167 8246 1201 8251
rect 1366 8282 1396 8316
rect 1396 8282 1400 8316
rect 1438 8282 1464 8316
rect 1464 8282 1472 8316
rect 1510 8282 1532 8316
rect 1532 8282 1544 8316
rect 1582 8282 1600 8316
rect 1600 8282 1616 8316
rect 1654 8282 1668 8316
rect 1668 8282 1688 8316
rect 1726 8282 1736 8316
rect 1736 8282 1760 8316
rect 1798 8282 1804 8316
rect 1804 8282 1832 8316
rect 1870 8282 1872 8316
rect 1872 8282 1904 8316
rect 1942 8282 1974 8316
rect 1974 8282 1976 8316
rect 2014 8282 2042 8316
rect 2042 8282 2048 8316
rect 2086 8282 2110 8316
rect 2110 8282 2120 8316
rect 2158 8282 2178 8316
rect 2178 8282 2192 8316
rect 2230 8282 2246 8316
rect 2246 8282 2264 8316
rect 2302 8282 2314 8316
rect 2314 8282 2336 8316
rect 2374 8282 2382 8316
rect 2382 8282 2408 8316
rect 2446 8282 2450 8316
rect 2450 8282 2480 8316
rect 2518 8282 2552 8316
rect 2590 8282 2620 8316
rect 2620 8282 2624 8316
rect 2662 8282 2688 8316
rect 2688 8282 2696 8316
rect 2734 8282 2756 8316
rect 2756 8282 2768 8316
rect 2806 8282 2824 8316
rect 2824 8282 2840 8316
rect 2878 8282 2892 8316
rect 2892 8282 2912 8316
rect 2950 8282 2960 8316
rect 2960 8282 2984 8316
rect 3022 8282 3028 8316
rect 3028 8282 3056 8316
rect 3094 8282 3096 8316
rect 3096 8282 3128 8316
rect 3166 8282 3198 8316
rect 3198 8282 3200 8316
rect 3238 8282 3266 8316
rect 3266 8282 3272 8316
rect 3310 8282 3334 8316
rect 3334 8282 3344 8316
rect 3382 8282 3402 8316
rect 3402 8282 3416 8316
rect 3454 8282 3470 8316
rect 3470 8282 3488 8316
rect 3526 8282 3538 8316
rect 3538 8282 3560 8316
rect 3598 8282 3606 8316
rect 3606 8282 3632 8316
rect 3670 8282 3674 8316
rect 3674 8282 3704 8316
rect 3742 8282 3776 8316
rect 3814 8282 3844 8316
rect 3844 8282 3848 8316
rect 3886 8282 3912 8316
rect 3912 8282 3920 8316
rect 3958 8282 3980 8316
rect 3980 8282 3992 8316
rect 4030 8282 4048 8316
rect 4048 8282 4064 8316
rect 4102 8282 4116 8316
rect 4116 8282 4136 8316
rect 4174 8282 4184 8316
rect 4184 8282 4208 8316
rect 4330 8304 4364 8337
rect 1167 8183 1201 8208
rect 1167 8174 1201 8183
rect 4330 8235 4364 8261
rect 4330 8227 4364 8235
rect 4330 8167 4364 8184
rect 1167 8115 1201 8136
rect 1167 8102 1201 8115
rect 1294 8126 1328 8160
rect 1366 8126 1396 8160
rect 1396 8126 1400 8160
rect 1438 8126 1464 8160
rect 1464 8126 1472 8160
rect 1510 8126 1532 8160
rect 1532 8126 1544 8160
rect 1582 8126 1600 8160
rect 1600 8126 1616 8160
rect 1654 8126 1668 8160
rect 1668 8126 1688 8160
rect 1726 8126 1736 8160
rect 1736 8126 1760 8160
rect 1798 8126 1804 8160
rect 1804 8126 1832 8160
rect 1870 8126 1872 8160
rect 1872 8126 1904 8160
rect 1942 8126 1974 8160
rect 1974 8126 1976 8160
rect 2014 8126 2042 8160
rect 2042 8126 2048 8160
rect 2086 8126 2110 8160
rect 2110 8126 2120 8160
rect 2158 8126 2178 8160
rect 2178 8126 2192 8160
rect 2230 8126 2246 8160
rect 2246 8126 2264 8160
rect 2302 8126 2314 8160
rect 2314 8126 2336 8160
rect 2374 8126 2382 8160
rect 2382 8126 2408 8160
rect 2446 8126 2450 8160
rect 2450 8126 2480 8160
rect 2518 8126 2552 8160
rect 2590 8126 2620 8160
rect 2620 8126 2624 8160
rect 2662 8126 2688 8160
rect 2688 8126 2696 8160
rect 2734 8126 2756 8160
rect 2756 8126 2768 8160
rect 2806 8126 2824 8160
rect 2824 8126 2840 8160
rect 2878 8126 2892 8160
rect 2892 8126 2912 8160
rect 2950 8126 2960 8160
rect 2960 8126 2984 8160
rect 3022 8126 3028 8160
rect 3028 8126 3056 8160
rect 3094 8126 3096 8160
rect 3096 8126 3128 8160
rect 3166 8126 3198 8160
rect 3198 8126 3200 8160
rect 3238 8126 3266 8160
rect 3266 8126 3272 8160
rect 3310 8126 3334 8160
rect 3334 8126 3344 8160
rect 3382 8126 3402 8160
rect 3402 8126 3416 8160
rect 3454 8126 3470 8160
rect 3470 8126 3488 8160
rect 3526 8126 3538 8160
rect 3538 8126 3560 8160
rect 3598 8126 3606 8160
rect 3606 8126 3632 8160
rect 3670 8126 3674 8160
rect 3674 8126 3704 8160
rect 3742 8126 3776 8160
rect 3814 8126 3844 8160
rect 3844 8126 3848 8160
rect 3886 8126 3912 8160
rect 3912 8126 3920 8160
rect 3958 8126 3980 8160
rect 3980 8126 3992 8160
rect 4030 8126 4048 8160
rect 4048 8126 4064 8160
rect 4102 8126 4116 8160
rect 4116 8126 4136 8160
rect 4174 8126 4184 8160
rect 4184 8126 4208 8160
rect 4330 8150 4364 8167
rect 1167 8047 1201 8064
rect 1167 8030 1201 8047
rect 1167 7979 1201 7992
rect 1167 7958 1201 7979
rect 4330 8099 4364 8107
rect 4330 8073 4364 8099
rect 1366 7970 1396 8004
rect 1396 7970 1400 8004
rect 1438 7970 1464 8004
rect 1464 7970 1472 8004
rect 1510 7970 1532 8004
rect 1532 7970 1544 8004
rect 1582 7970 1600 8004
rect 1600 7970 1616 8004
rect 1654 7970 1668 8004
rect 1668 7970 1688 8004
rect 1726 7970 1736 8004
rect 1736 7970 1760 8004
rect 1798 7970 1804 8004
rect 1804 7970 1832 8004
rect 1870 7970 1872 8004
rect 1872 7970 1904 8004
rect 1942 7970 1974 8004
rect 1974 7970 1976 8004
rect 2014 7970 2042 8004
rect 2042 7970 2048 8004
rect 2086 7970 2110 8004
rect 2110 7970 2120 8004
rect 2158 7970 2178 8004
rect 2178 7970 2192 8004
rect 2230 7970 2246 8004
rect 2246 7970 2264 8004
rect 2302 7970 2314 8004
rect 2314 7970 2336 8004
rect 2374 7970 2382 8004
rect 2382 7970 2408 8004
rect 2446 7970 2450 8004
rect 2450 7970 2480 8004
rect 2518 7970 2552 8004
rect 2590 7970 2620 8004
rect 2620 7970 2624 8004
rect 2662 7970 2688 8004
rect 2688 7970 2696 8004
rect 2734 7970 2756 8004
rect 2756 7970 2768 8004
rect 2806 7970 2824 8004
rect 2824 7970 2840 8004
rect 2878 7970 2892 8004
rect 2892 7970 2912 8004
rect 2950 7970 2960 8004
rect 2960 7970 2984 8004
rect 3022 7970 3028 8004
rect 3028 7970 3056 8004
rect 3094 7970 3096 8004
rect 3096 7970 3128 8004
rect 3166 7970 3198 8004
rect 3198 7970 3200 8004
rect 3238 7970 3266 8004
rect 3266 7970 3272 8004
rect 3310 7970 3334 8004
rect 3334 7970 3344 8004
rect 3382 7970 3402 8004
rect 3402 7970 3416 8004
rect 3454 7970 3470 8004
rect 3470 7970 3488 8004
rect 3526 7970 3538 8004
rect 3538 7970 3560 8004
rect 3598 7970 3606 8004
rect 3606 7970 3632 8004
rect 3670 7970 3674 8004
rect 3674 7970 3704 8004
rect 3742 7970 3776 8004
rect 3814 7970 3844 8004
rect 3844 7970 3848 8004
rect 3886 7970 3912 8004
rect 3912 7970 3920 8004
rect 3958 7970 3980 8004
rect 3980 7970 3992 8004
rect 4030 7970 4048 8004
rect 4048 7970 4064 8004
rect 4102 7970 4116 8004
rect 4116 7970 4136 8004
rect 4174 7970 4184 8004
rect 4184 7970 4208 8004
rect 4330 7997 4364 8030
rect 4330 7996 4364 7997
rect 1167 7911 1201 7920
rect 1167 7886 1201 7911
rect 1167 7843 1201 7848
rect 1167 7814 1201 7843
rect 4330 7929 4364 7953
rect 4330 7919 4364 7929
rect 4330 7861 4364 7876
rect 1294 7814 1328 7848
rect 1366 7814 1396 7848
rect 1396 7814 1400 7848
rect 1438 7814 1464 7848
rect 1464 7814 1472 7848
rect 1510 7814 1532 7848
rect 1532 7814 1544 7848
rect 1582 7814 1600 7848
rect 1600 7814 1616 7848
rect 1654 7814 1668 7848
rect 1668 7814 1688 7848
rect 1726 7814 1736 7848
rect 1736 7814 1760 7848
rect 1798 7814 1804 7848
rect 1804 7814 1832 7848
rect 1870 7814 1872 7848
rect 1872 7814 1904 7848
rect 1942 7814 1974 7848
rect 1974 7814 1976 7848
rect 2014 7814 2042 7848
rect 2042 7814 2048 7848
rect 2086 7814 2110 7848
rect 2110 7814 2120 7848
rect 2158 7814 2178 7848
rect 2178 7814 2192 7848
rect 2230 7814 2246 7848
rect 2246 7814 2264 7848
rect 2302 7814 2314 7848
rect 2314 7814 2336 7848
rect 2374 7814 2382 7848
rect 2382 7814 2408 7848
rect 2446 7814 2450 7848
rect 2450 7814 2480 7848
rect 2518 7814 2552 7848
rect 2590 7814 2620 7848
rect 2620 7814 2624 7848
rect 2662 7814 2688 7848
rect 2688 7814 2696 7848
rect 2734 7814 2756 7848
rect 2756 7814 2768 7848
rect 2806 7814 2824 7848
rect 2824 7814 2840 7848
rect 2878 7814 2892 7848
rect 2892 7814 2912 7848
rect 2950 7814 2960 7848
rect 2960 7814 2984 7848
rect 3022 7814 3028 7848
rect 3028 7814 3056 7848
rect 3094 7814 3096 7848
rect 3096 7814 3128 7848
rect 3166 7814 3198 7848
rect 3198 7814 3200 7848
rect 3238 7814 3266 7848
rect 3266 7814 3272 7848
rect 3310 7814 3334 7848
rect 3334 7814 3344 7848
rect 3382 7814 3402 7848
rect 3402 7814 3416 7848
rect 3454 7814 3470 7848
rect 3470 7814 3488 7848
rect 3526 7814 3538 7848
rect 3538 7814 3560 7848
rect 3598 7814 3606 7848
rect 3606 7814 3632 7848
rect 3670 7814 3674 7848
rect 3674 7814 3704 7848
rect 3742 7814 3776 7848
rect 3814 7814 3844 7848
rect 3844 7814 3848 7848
rect 3886 7814 3912 7848
rect 3912 7814 3920 7848
rect 3958 7814 3980 7848
rect 3980 7814 3992 7848
rect 4030 7814 4048 7848
rect 4048 7814 4064 7848
rect 4102 7814 4116 7848
rect 4116 7814 4136 7848
rect 4174 7814 4184 7848
rect 4184 7814 4208 7848
rect 4330 7842 4364 7861
rect 1167 7775 1201 7776
rect 1167 7742 1201 7775
rect 1167 7673 1201 7704
rect 1167 7670 1201 7673
rect 4330 7793 4364 7799
rect 4330 7765 4364 7793
rect 1366 7658 1396 7692
rect 1396 7658 1400 7692
rect 1438 7658 1464 7692
rect 1464 7658 1472 7692
rect 1510 7658 1532 7692
rect 1532 7658 1544 7692
rect 1582 7658 1600 7692
rect 1600 7658 1616 7692
rect 1654 7658 1668 7692
rect 1668 7658 1688 7692
rect 1726 7658 1736 7692
rect 1736 7658 1760 7692
rect 1798 7658 1804 7692
rect 1804 7658 1832 7692
rect 1870 7658 1872 7692
rect 1872 7658 1904 7692
rect 1942 7658 1974 7692
rect 1974 7658 1976 7692
rect 2014 7658 2042 7692
rect 2042 7658 2048 7692
rect 2086 7658 2110 7692
rect 2110 7658 2120 7692
rect 2158 7658 2178 7692
rect 2178 7658 2192 7692
rect 2230 7658 2246 7692
rect 2246 7658 2264 7692
rect 2302 7658 2314 7692
rect 2314 7658 2336 7692
rect 2374 7658 2382 7692
rect 2382 7658 2408 7692
rect 2446 7658 2450 7692
rect 2450 7658 2480 7692
rect 2518 7658 2552 7692
rect 2590 7658 2620 7692
rect 2620 7658 2624 7692
rect 2662 7658 2688 7692
rect 2688 7658 2696 7692
rect 2734 7658 2756 7692
rect 2756 7658 2768 7692
rect 2806 7658 2824 7692
rect 2824 7658 2840 7692
rect 2878 7658 2892 7692
rect 2892 7658 2912 7692
rect 2950 7658 2960 7692
rect 2960 7658 2984 7692
rect 3022 7658 3028 7692
rect 3028 7658 3056 7692
rect 3094 7658 3096 7692
rect 3096 7658 3128 7692
rect 3166 7658 3198 7692
rect 3198 7658 3200 7692
rect 3238 7658 3266 7692
rect 3266 7658 3272 7692
rect 3310 7658 3334 7692
rect 3334 7658 3344 7692
rect 3382 7658 3402 7692
rect 3402 7658 3416 7692
rect 3454 7658 3470 7692
rect 3470 7658 3488 7692
rect 3526 7658 3538 7692
rect 3538 7658 3560 7692
rect 3598 7658 3606 7692
rect 3606 7658 3632 7692
rect 3670 7658 3674 7692
rect 3674 7658 3704 7692
rect 3742 7658 3776 7692
rect 3814 7658 3844 7692
rect 3844 7658 3848 7692
rect 3886 7658 3912 7692
rect 3912 7658 3920 7692
rect 3958 7658 3980 7692
rect 3980 7658 3992 7692
rect 4030 7658 4048 7692
rect 4048 7658 4064 7692
rect 4102 7658 4116 7692
rect 4116 7658 4136 7692
rect 4174 7658 4184 7692
rect 4184 7658 4208 7692
rect 4330 7691 4364 7721
rect 4330 7687 4364 7691
rect 1167 7605 1201 7632
rect 1167 7598 1201 7605
rect 1167 7537 1201 7560
rect 1167 7526 1201 7537
rect 4330 7623 4364 7643
rect 4330 7609 4364 7623
rect 4330 7555 4364 7565
rect 1294 7502 1328 7536
rect 1366 7502 1396 7536
rect 1396 7502 1400 7536
rect 1438 7502 1464 7536
rect 1464 7502 1472 7536
rect 1510 7502 1532 7536
rect 1532 7502 1544 7536
rect 1582 7502 1600 7536
rect 1600 7502 1616 7536
rect 1654 7502 1668 7536
rect 1668 7502 1688 7536
rect 1726 7502 1736 7536
rect 1736 7502 1760 7536
rect 1798 7502 1804 7536
rect 1804 7502 1832 7536
rect 1870 7502 1872 7536
rect 1872 7502 1904 7536
rect 1942 7502 1974 7536
rect 1974 7502 1976 7536
rect 2014 7502 2042 7536
rect 2042 7502 2048 7536
rect 2086 7502 2110 7536
rect 2110 7502 2120 7536
rect 2158 7502 2178 7536
rect 2178 7502 2192 7536
rect 2230 7502 2246 7536
rect 2246 7502 2264 7536
rect 2302 7502 2314 7536
rect 2314 7502 2336 7536
rect 2374 7502 2382 7536
rect 2382 7502 2408 7536
rect 2446 7502 2450 7536
rect 2450 7502 2480 7536
rect 2518 7502 2552 7536
rect 2590 7502 2620 7536
rect 2620 7502 2624 7536
rect 2662 7502 2688 7536
rect 2688 7502 2696 7536
rect 2734 7502 2756 7536
rect 2756 7502 2768 7536
rect 2806 7502 2824 7536
rect 2824 7502 2840 7536
rect 2878 7502 2892 7536
rect 2892 7502 2912 7536
rect 2950 7502 2960 7536
rect 2960 7502 2984 7536
rect 3022 7502 3028 7536
rect 3028 7502 3056 7536
rect 3094 7502 3096 7536
rect 3096 7502 3128 7536
rect 3166 7502 3198 7536
rect 3198 7502 3200 7536
rect 3238 7502 3266 7536
rect 3266 7502 3272 7536
rect 3310 7502 3334 7536
rect 3334 7502 3344 7536
rect 3382 7502 3402 7536
rect 3402 7502 3416 7536
rect 3454 7502 3470 7536
rect 3470 7502 3488 7536
rect 3526 7502 3538 7536
rect 3538 7502 3560 7536
rect 3598 7502 3606 7536
rect 3606 7502 3632 7536
rect 3670 7502 3674 7536
rect 3674 7502 3704 7536
rect 3742 7502 3776 7536
rect 3814 7502 3844 7536
rect 3844 7502 3848 7536
rect 3886 7502 3912 7536
rect 3912 7502 3920 7536
rect 3958 7502 3980 7536
rect 3980 7502 3992 7536
rect 4030 7502 4048 7536
rect 4048 7502 4064 7536
rect 4102 7502 4116 7536
rect 4116 7502 4136 7536
rect 4174 7502 4184 7536
rect 4184 7502 4208 7536
rect 4330 7531 4364 7555
rect 1167 7469 1201 7488
rect 1167 7454 1201 7469
rect 1167 7401 1201 7416
rect 1167 7382 1201 7401
rect 4330 7453 4364 7487
rect 4474 8402 4508 8436
rect 4474 8330 4508 8364
rect 4474 8258 4508 8292
rect 4474 8186 4508 8220
rect 4474 8114 4508 8148
rect 4474 8042 4508 8076
rect 4474 7970 4508 8004
rect 4474 7898 4508 7932
rect 4474 7826 4508 7860
rect 4474 7754 4508 7788
rect 4474 7682 4508 7716
rect 4474 7610 4508 7644
rect 4474 7538 4508 7572
rect 4474 7466 4508 7500
rect 4474 7394 4508 7428
rect 1167 7333 1201 7344
rect 1167 7310 1201 7333
rect 1294 7346 1328 7380
rect 1366 7346 1396 7380
rect 1396 7346 1400 7380
rect 1438 7346 1464 7380
rect 1464 7346 1472 7380
rect 1510 7346 1532 7380
rect 1532 7346 1544 7380
rect 1582 7346 1600 7380
rect 1600 7346 1616 7380
rect 1654 7346 1668 7380
rect 1668 7346 1688 7380
rect 1726 7346 1736 7380
rect 1736 7346 1760 7380
rect 1798 7346 1804 7380
rect 1804 7346 1832 7380
rect 1870 7346 1872 7380
rect 1872 7346 1904 7380
rect 1942 7346 1974 7380
rect 1974 7346 1976 7380
rect 2014 7346 2042 7380
rect 2042 7346 2048 7380
rect 2086 7346 2110 7380
rect 2110 7346 2120 7380
rect 2158 7346 2178 7380
rect 2178 7346 2192 7380
rect 2230 7346 2246 7380
rect 2246 7346 2264 7380
rect 2302 7346 2314 7380
rect 2314 7346 2336 7380
rect 2374 7346 2382 7380
rect 2382 7346 2408 7380
rect 2446 7346 2450 7380
rect 2450 7346 2480 7380
rect 2518 7346 2552 7380
rect 2590 7346 2620 7380
rect 2620 7346 2624 7380
rect 2662 7346 2688 7380
rect 2688 7346 2696 7380
rect 2734 7346 2756 7380
rect 2756 7346 2768 7380
rect 2806 7346 2824 7380
rect 2824 7346 2840 7380
rect 2878 7346 2892 7380
rect 2892 7346 2912 7380
rect 2950 7346 2960 7380
rect 2960 7346 2984 7380
rect 3022 7346 3028 7380
rect 3028 7346 3056 7380
rect 3094 7346 3096 7380
rect 3096 7346 3128 7380
rect 3166 7346 3198 7380
rect 3198 7346 3200 7380
rect 3238 7346 3266 7380
rect 3266 7346 3272 7380
rect 3310 7346 3334 7380
rect 3334 7346 3344 7380
rect 3382 7346 3402 7380
rect 3402 7346 3416 7380
rect 3454 7346 3470 7380
rect 3470 7346 3488 7380
rect 3526 7346 3538 7380
rect 3538 7346 3560 7380
rect 3598 7346 3606 7380
rect 3606 7346 3632 7380
rect 3670 7346 3674 7380
rect 3674 7346 3704 7380
rect 3742 7346 3776 7380
rect 3814 7346 3844 7380
rect 3844 7346 3848 7380
rect 3886 7346 3912 7380
rect 3912 7346 3920 7380
rect 3958 7346 3980 7380
rect 3980 7346 3992 7380
rect 4030 7346 4048 7380
rect 4048 7346 4064 7380
rect 4102 7346 4116 7380
rect 4116 7346 4136 7380
rect 4174 7346 4184 7380
rect 4184 7346 4208 7380
rect 1167 7238 1201 7272
rect 1300 7232 1325 7266
rect 1325 7232 1334 7266
rect 1372 7232 1393 7266
rect 1393 7232 1406 7266
rect 1444 7232 1461 7266
rect 1461 7232 1478 7266
rect 1516 7232 1529 7266
rect 1529 7232 1550 7266
rect 1588 7232 1622 7266
rect 1660 7232 1690 7266
rect 1690 7232 1694 7266
rect 1732 7232 1758 7266
rect 1758 7232 1766 7266
rect 1804 7232 1826 7266
rect 1826 7232 1838 7266
rect 1876 7232 1894 7266
rect 1894 7232 1910 7266
rect 1948 7232 1962 7266
rect 1962 7232 1982 7266
rect 2020 7232 2030 7266
rect 2030 7232 2054 7266
rect 2092 7232 2098 7266
rect 2098 7232 2126 7266
rect 2164 7232 2166 7266
rect 2166 7232 2198 7266
rect 2236 7232 2268 7266
rect 2268 7232 2270 7266
rect 2308 7232 2336 7266
rect 2336 7232 2342 7266
rect 2380 7232 2404 7266
rect 2404 7232 2414 7266
rect 2452 7232 2472 7266
rect 2472 7232 2486 7266
rect 2524 7232 2540 7266
rect 2540 7232 2558 7266
rect 2596 7232 2608 7266
rect 2608 7232 2630 7266
rect 2668 7232 2676 7266
rect 2676 7232 2702 7266
rect 2740 7232 2744 7266
rect 2744 7232 2774 7266
rect 2812 7232 2846 7266
rect 2884 7232 2914 7266
rect 2914 7232 2918 7266
rect 2956 7232 2982 7266
rect 2982 7232 2990 7266
rect 3028 7232 3050 7266
rect 3050 7232 3062 7266
rect 3100 7232 3118 7266
rect 3118 7232 3134 7266
rect 3172 7232 3186 7266
rect 3186 7232 3206 7266
rect 3244 7232 3254 7266
rect 3254 7232 3278 7266
rect 3316 7232 3322 7266
rect 3322 7232 3350 7266
rect 3388 7232 3390 7266
rect 3390 7232 3422 7266
rect 3460 7232 3492 7266
rect 3492 7232 3494 7266
rect 3532 7232 3560 7266
rect 3560 7232 3566 7266
rect 3604 7232 3628 7266
rect 3628 7232 3638 7266
rect 3676 7232 3696 7266
rect 3696 7232 3710 7266
rect 3748 7232 3764 7266
rect 3764 7232 3782 7266
rect 3820 7232 3832 7266
rect 3832 7232 3854 7266
rect 3892 7232 3900 7266
rect 3900 7232 3926 7266
rect 3964 7232 3968 7266
rect 3968 7232 3998 7266
rect 4036 7232 4070 7266
rect 4108 7232 4138 7266
rect 4138 7232 4142 7266
rect 4180 7232 4206 7266
rect 4206 7232 4214 7266
rect 4252 7232 4274 7266
rect 4274 7232 4286 7266
rect 4324 7232 4342 7266
rect 4342 7232 4358 7266
rect 4396 7232 4430 7266
rect 4468 7232 4502 7266
rect 800 7169 834 7195
rect 800 7161 834 7169
rect 829 7044 841 7078
rect 841 7044 863 7078
rect 901 7044 909 7078
rect 909 7044 935 7078
rect 973 7044 977 7078
rect 977 7044 1007 7078
rect 1045 7044 1079 7078
rect 1117 7044 1147 7078
rect 1147 7044 1151 7078
rect 1189 7044 1215 7078
rect 1215 7044 1223 7078
rect 1261 7044 1283 7078
rect 1283 7044 1295 7078
rect 1333 7044 1351 7078
rect 1351 7044 1367 7078
rect 1405 7044 1419 7078
rect 1419 7044 1439 7078
rect 1477 7044 1487 7078
rect 1487 7044 1511 7078
rect 1549 7044 1555 7078
rect 1555 7044 1583 7078
rect 1621 7044 1623 7078
rect 1623 7044 1655 7078
rect 1693 7044 1725 7078
rect 1725 7044 1727 7078
rect 1765 7044 1793 7078
rect 1793 7044 1799 7078
rect 1837 7044 1861 7078
rect 1861 7044 1871 7078
rect 1909 7044 1929 7078
rect 1929 7044 1943 7078
rect 1981 7044 1997 7078
rect 1997 7044 2015 7078
rect 2053 7044 2065 7078
rect 2065 7044 2087 7078
rect 2125 7044 2133 7078
rect 2133 7044 2159 7078
rect 2197 7044 2201 7078
rect 2201 7044 2231 7078
rect 2269 7044 2303 7078
rect 2341 7044 2371 7078
rect 2371 7044 2375 7078
rect 2413 7044 2439 7078
rect 2439 7044 2447 7078
rect 2485 7044 2507 7078
rect 2507 7044 2519 7078
rect 2557 7044 2575 7078
rect 2575 7044 2591 7078
rect 2629 7044 2643 7078
rect 2643 7044 2663 7078
rect 2701 7044 2711 7078
rect 2711 7044 2735 7078
rect 2773 7044 2779 7078
rect 2779 7044 2807 7078
rect 2845 7044 2847 7078
rect 2847 7044 2879 7078
rect 2917 7044 2949 7078
rect 2949 7044 2951 7078
rect 2989 7044 3017 7078
rect 3017 7044 3023 7078
rect 3061 7044 3085 7078
rect 3085 7044 3095 7078
rect 3133 7044 3153 7078
rect 3153 7044 3167 7078
rect 3205 7044 3221 7078
rect 3221 7044 3239 7078
rect 3277 7044 3289 7078
rect 3289 7044 3311 7078
rect 3349 7044 3357 7078
rect 3357 7044 3383 7078
rect 3421 7044 3425 7078
rect 3425 7044 3455 7078
rect 3493 7044 3527 7078
rect 3565 7044 3595 7078
rect 3595 7044 3599 7078
rect 3637 7044 3663 7078
rect 3663 7044 3671 7078
rect 3709 7044 3731 7078
rect 3731 7044 3743 7078
rect 3781 7044 3799 7078
rect 3799 7044 3815 7078
rect 3853 7044 3867 7078
rect 3867 7044 3887 7078
rect 3925 7044 3935 7078
rect 3935 7044 3959 7078
rect 3997 7044 4003 7078
rect 4003 7044 4031 7078
rect 4069 7044 4071 7078
rect 4071 7044 4103 7078
rect 4141 7044 4173 7078
rect 4173 7044 4175 7078
rect 4213 7044 4241 7078
rect 4241 7044 4247 7078
rect 4285 7044 4309 7078
rect 4309 7044 4319 7078
rect 4357 7044 4377 7078
rect 4377 7044 4391 7078
rect 4429 7044 4445 7078
rect 4445 7044 4463 7078
rect 4501 7044 4513 7078
rect 4513 7044 4535 7078
rect 4573 7044 4581 7078
rect 4581 7044 4607 7078
rect 4645 7044 4649 7078
rect 4649 7044 4679 7078
rect 4424 6973 4446 7006
rect 4446 6973 4458 7006
rect 4507 6973 4518 7006
rect 4518 6973 4541 7006
rect 4590 6973 4624 7006
rect 4672 6973 4696 7006
rect 4696 6973 4706 7006
rect 4424 6972 4458 6973
rect 4507 6972 4541 6973
rect 4590 6972 4624 6973
rect 4672 6972 4706 6973
rect 4424 6905 4446 6934
rect 4446 6905 4458 6934
rect 4507 6905 4518 6934
rect 4518 6905 4541 6934
rect 4590 6905 4624 6934
rect 4672 6905 4696 6934
rect 4696 6905 4706 6934
rect 4424 6900 4458 6905
rect 4507 6900 4541 6905
rect 4590 6900 4624 6905
rect 4672 6900 4706 6905
rect -849 6689 -815 6715
rect 308 6689 342 6713
rect 382 6689 416 6713
rect 456 6689 490 6713
rect 530 6689 564 6713
rect 604 6689 638 6713
rect 678 6689 712 6713
rect 751 6689 785 6713
rect 824 6689 858 6713
rect -849 6681 -816 6689
rect -816 6681 -815 6689
rect 308 6679 323 6689
rect 323 6679 342 6689
rect 382 6679 391 6689
rect 391 6679 416 6689
rect 456 6679 459 6689
rect 459 6679 490 6689
rect 530 6679 561 6689
rect 561 6679 564 6689
rect 604 6679 629 6689
rect 629 6679 638 6689
rect 678 6679 697 6689
rect 697 6679 712 6689
rect 751 6679 765 6689
rect 765 6679 785 6689
rect 824 6679 833 6689
rect 833 6679 858 6689
rect -849 6619 -815 6635
rect -849 6601 -816 6619
rect -816 6601 -815 6619
rect 308 6585 323 6589
rect 323 6585 342 6589
rect 382 6585 391 6589
rect 391 6585 416 6589
rect 456 6585 459 6589
rect 459 6585 490 6589
rect 530 6585 561 6589
rect 561 6585 564 6589
rect 604 6585 629 6589
rect 629 6585 638 6589
rect 678 6585 697 6589
rect 697 6585 712 6589
rect 751 6585 765 6589
rect 765 6585 785 6589
rect 824 6585 833 6589
rect 833 6585 858 6589
rect 308 6555 342 6585
rect 382 6555 416 6585
rect 456 6555 490 6585
rect 530 6555 564 6585
rect 604 6555 638 6585
rect 678 6555 712 6585
rect 751 6555 785 6585
rect 824 6555 858 6585
rect -849 6549 -815 6555
rect -849 6521 -816 6549
rect -816 6521 -815 6549
rect -849 6445 -816 6475
rect -816 6445 -815 6475
rect 1019 6548 1053 6582
rect 1135 6548 1169 6582
rect 1019 6464 1053 6498
rect 1135 6464 1169 6498
rect 4502 6837 4518 6861
rect 4518 6837 4536 6861
rect 4576 6837 4590 6861
rect 4590 6837 4610 6861
rect 4649 6837 4662 6861
rect 4662 6837 4683 6861
rect 4502 6827 4536 6837
rect 4576 6827 4610 6837
rect 4649 6827 4683 6837
rect 4596 6735 4630 6769
rect 4668 6735 4702 6769
rect 2551 6512 2585 6546
rect 2627 6512 2661 6546
rect 2703 6512 2737 6546
rect 2779 6512 2813 6546
rect 2854 6512 2888 6546
rect 2929 6512 2963 6546
rect 3004 6512 3038 6546
rect 3079 6512 3113 6546
rect 3154 6512 3188 6546
rect 3229 6512 3263 6546
rect 4058 6560 4092 6594
rect 4174 6560 4208 6594
rect 4058 6476 4092 6510
rect 4174 6476 4208 6510
rect -849 6441 -815 6445
rect -849 6375 -816 6395
rect -816 6375 -815 6395
rect 2551 6438 2585 6472
rect 2627 6438 2661 6472
rect 2703 6438 2737 6472
rect 2779 6438 2813 6472
rect 2854 6438 2888 6472
rect 2929 6438 2963 6472
rect 3004 6438 3038 6472
rect 3079 6438 3113 6472
rect 3154 6438 3188 6472
rect 3229 6438 3263 6472
rect -849 6361 -815 6375
rect -849 6305 -816 6315
rect -816 6305 -815 6315
rect -849 6281 -815 6305
rect 1019 6345 1053 6379
rect 1135 6345 1169 6379
rect 1019 6261 1053 6295
rect 1135 6261 1169 6295
rect 2551 6364 2585 6398
rect 2627 6364 2661 6398
rect 2703 6364 2737 6398
rect 2779 6364 2813 6398
rect 2854 6364 2888 6398
rect 2929 6364 2963 6398
rect 3004 6364 3038 6398
rect 3079 6364 3113 6398
rect 3154 6364 3188 6398
rect 3229 6364 3263 6398
rect 2551 6290 2585 6324
rect 2627 6290 2661 6324
rect 2703 6290 2737 6324
rect 2779 6290 2813 6324
rect 2854 6290 2888 6324
rect 2929 6290 2963 6324
rect 3004 6290 3038 6324
rect 3079 6290 3113 6324
rect 3154 6290 3188 6324
rect 3229 6290 3263 6324
rect -849 6200 -815 6234
rect -849 6129 -815 6153
rect -849 6119 -816 6129
rect -816 6119 -815 6129
rect 2551 6216 2585 6250
rect 2627 6216 2661 6250
rect 2703 6216 2737 6250
rect 2779 6216 2813 6250
rect 2854 6216 2888 6250
rect 2929 6216 2963 6250
rect 3004 6216 3038 6250
rect 3079 6216 3113 6250
rect 3154 6216 3188 6250
rect 3229 6216 3263 6250
rect 4058 6127 4092 6161
rect 4174 6127 4208 6161
rect 4058 6043 4092 6077
rect 4174 6043 4208 6077
rect 4579 5331 4592 5335
rect 4592 5331 4613 5335
rect 4651 5331 4662 5335
rect 4662 5331 4685 5335
rect 4579 5301 4613 5331
rect 4651 5301 4685 5331
rect 4466 5227 4500 5245
rect 4466 5211 4486 5227
rect 4486 5211 4500 5227
rect 4556 5211 4590 5245
rect 4646 5227 4680 5245
rect 4646 5211 4662 5227
rect 4662 5211 4680 5227
rect 4466 5158 4500 5171
rect 4466 5137 4486 5158
rect 4486 5137 4500 5158
rect 4556 5137 4590 5171
rect 4646 5158 4680 5171
rect 4646 5137 4662 5158
rect 4662 5137 4680 5158
rect 4466 5089 4500 5097
rect 4466 5063 4486 5089
rect 4486 5063 4500 5089
rect 4556 5063 4590 5097
rect 4646 5089 4680 5097
rect 4646 5063 4662 5089
rect 4662 5063 4680 5089
rect 4466 5019 4500 5023
rect 4466 4989 4486 5019
rect 4486 4989 4500 5019
rect 4556 4989 4590 5023
rect 4646 5019 4680 5023
rect 4646 4989 4662 5019
rect 4662 4989 4680 5019
rect 4466 4915 4486 4949
rect 4486 4915 4500 4949
rect 4556 4915 4590 4949
rect 4646 4915 4662 4949
rect 4662 4915 4680 4949
rect 4466 4845 4486 4875
rect 4486 4845 4500 4875
rect 4466 4841 4500 4845
rect 4556 4841 4590 4875
rect 4646 4845 4662 4875
rect 4662 4845 4680 4875
rect 4646 4841 4680 4845
rect 4466 4775 4486 4801
rect 4486 4775 4500 4801
rect 4466 4767 4500 4775
rect 4556 4767 4590 4801
rect 4646 4775 4662 4801
rect 4662 4775 4680 4801
rect 4646 4767 4680 4775
rect 4466 4705 4486 4727
rect 4486 4705 4500 4727
rect 4466 4693 4500 4705
rect 4556 4693 4590 4727
rect 4646 4705 4662 4727
rect 4662 4705 4680 4727
rect 4646 4693 4680 4705
rect 4579 4599 4613 4626
rect 4651 4599 4685 4626
rect 4579 4592 4592 4599
rect 4592 4592 4613 4599
rect 4651 4592 4662 4599
rect 4662 4592 4685 4599
rect 13205 4280 13239 4314
rect 13205 4240 13239 4242
rect 13205 4208 13227 4240
rect 13227 4208 13239 4240
rect 14983 4302 15017 4314
rect 14983 4280 15017 4302
rect 14983 4234 15017 4241
rect 14983 4207 15017 4234
rect 13205 4138 13227 4170
rect 13227 4138 13239 4170
rect 13205 4136 13239 4138
rect 13205 4070 13227 4098
rect 13227 4070 13239 4098
rect 13205 4064 13239 4070
rect 11464 3984 11498 4018
rect 11538 3984 11572 4018
rect 11612 3984 11646 4018
rect 11686 3984 11720 4018
rect 11760 3984 11794 4018
rect 11834 3984 11868 4018
rect 11464 3868 11498 3902
rect 11538 3868 11572 3902
rect 11612 3868 11646 3902
rect 11686 3868 11720 3902
rect 11760 3868 11794 3902
rect 11834 3868 11868 3902
rect 11964 3984 11998 4018
rect 12038 3984 12072 4018
rect 12112 3984 12146 4018
rect 12186 3984 12220 4018
rect 12260 3984 12294 4018
rect 12334 3984 12368 4018
rect 11964 3868 11998 3902
rect 12038 3868 12072 3902
rect 12112 3868 12146 3902
rect 12186 3868 12220 3902
rect 12260 3868 12294 3902
rect 12334 3868 12368 3902
rect 12465 3984 12499 4018
rect 12539 3984 12573 4018
rect 12613 3984 12647 4018
rect 12687 3984 12721 4018
rect 12761 3984 12795 4018
rect 12835 3984 12869 4018
rect 12465 3868 12499 3902
rect 12539 3868 12573 3902
rect 12613 3868 12647 3902
rect 12687 3868 12721 3902
rect 12761 3868 12795 3902
rect 12835 3868 12869 3902
rect 13205 4002 13227 4026
rect 13227 4002 13239 4026
rect 13205 3992 13239 4002
rect 13205 3934 13227 3954
rect 13227 3934 13239 3954
rect 13205 3920 13239 3934
rect 8474 3751 8493 3758
rect 8493 3751 8508 3758
rect 8547 3751 8562 3758
rect 8562 3751 8581 3758
rect 8620 3751 8631 3758
rect 8631 3751 8654 3758
rect 8693 3751 8700 3758
rect 8700 3751 8727 3758
rect 8766 3751 8769 3758
rect 8769 3751 8800 3758
rect 8839 3751 8872 3758
rect 8872 3751 8873 3758
rect 8912 3751 8941 3758
rect 8941 3751 8946 3758
rect 8984 3751 9010 3758
rect 9010 3751 9018 3758
rect 9056 3751 9079 3758
rect 9079 3751 9090 3758
rect 9128 3751 9148 3758
rect 9148 3751 9162 3758
rect 9200 3751 9217 3758
rect 9217 3751 9234 3758
rect 9272 3751 9286 3758
rect 9286 3751 9306 3758
rect 9344 3751 9354 3758
rect 9354 3751 9378 3758
rect 8474 3724 8508 3751
rect 8547 3724 8581 3751
rect 8620 3724 8654 3751
rect 8693 3724 8727 3751
rect 8766 3724 8800 3751
rect 8839 3724 8873 3751
rect 8912 3724 8946 3751
rect 8984 3724 9018 3751
rect 9056 3724 9090 3751
rect 9128 3724 9162 3751
rect 9200 3724 9234 3751
rect 9272 3724 9306 3751
rect 9344 3724 9378 3751
rect 13205 3866 13227 3882
rect 13227 3866 13239 3882
rect 13205 3848 13239 3866
rect 13205 3798 13227 3810
rect 13227 3798 13239 3810
rect 13205 3776 13239 3798
rect 13205 3730 13227 3738
rect 13227 3730 13239 3738
rect 13205 3704 13239 3730
rect 13205 3662 13227 3666
rect 13227 3662 13239 3666
rect 13205 3632 13239 3662
rect 13205 3560 13239 3594
rect 13205 3492 13239 3522
rect 13205 3488 13227 3492
rect 13227 3488 13239 3492
rect 13205 3424 13239 3450
rect 13205 3416 13227 3424
rect 13227 3416 13239 3424
rect 13205 3356 13239 3378
rect 13205 3344 13227 3356
rect 13227 3344 13239 3356
rect 13205 3288 13239 3306
rect 11464 3252 11498 3286
rect 11537 3252 11571 3286
rect 11610 3252 11644 3286
rect 11683 3252 11717 3286
rect 11756 3252 11790 3286
rect 11828 3252 11862 3286
rect 11900 3252 11934 3286
rect 11972 3252 12006 3286
rect 12044 3252 12078 3286
rect 12116 3252 12150 3286
rect 12188 3252 12222 3286
rect 12260 3252 12294 3286
rect 12332 3252 12366 3286
rect 12404 3252 12438 3286
rect 11464 3136 11498 3170
rect 11537 3136 11571 3170
rect 11610 3136 11644 3170
rect 11683 3136 11717 3170
rect 11756 3136 11790 3170
rect 11828 3136 11862 3170
rect 11900 3136 11934 3170
rect 11972 3136 12006 3170
rect 12044 3136 12078 3170
rect 12116 3136 12150 3170
rect 12188 3136 12222 3170
rect 12260 3136 12294 3170
rect 12332 3136 12366 3170
rect 12404 3136 12438 3170
rect 12480 3252 12514 3286
rect 12558 3252 12592 3286
rect 12635 3252 12669 3286
rect 12712 3252 12746 3286
rect 12789 3252 12823 3286
rect 12866 3252 12900 3286
rect 12480 3160 12514 3194
rect 12558 3160 12592 3194
rect 12635 3160 12669 3194
rect 12712 3160 12746 3194
rect 12789 3160 12823 3194
rect 12866 3160 12900 3194
rect 12480 3068 12514 3102
rect 12558 3068 12592 3102
rect 12635 3068 12669 3102
rect 12712 3068 12746 3102
rect 12789 3068 12823 3102
rect 12866 3068 12900 3102
rect 13205 3272 13227 3288
rect 13227 3272 13239 3288
rect 13205 3220 13239 3234
rect 13509 4173 13543 4180
rect 13583 4173 13617 4180
rect 13657 4173 13691 4180
rect 13731 4173 13765 4180
rect 13805 4173 13839 4180
rect 13879 4173 13913 4180
rect 13953 4173 13987 4180
rect 14027 4173 14061 4180
rect 14101 4173 14135 4180
rect 14175 4173 14209 4180
rect 14249 4173 14283 4180
rect 14323 4173 14357 4180
rect 14397 4173 14431 4180
rect 14470 4173 14504 4180
rect 14543 4173 14577 4180
rect 13509 4146 13541 4173
rect 13541 4146 13543 4173
rect 13583 4146 13609 4173
rect 13609 4146 13617 4173
rect 13657 4146 13677 4173
rect 13677 4146 13691 4173
rect 13731 4146 13745 4173
rect 13745 4146 13765 4173
rect 13805 4146 13813 4173
rect 13813 4146 13839 4173
rect 13879 4146 13881 4173
rect 13881 4146 13913 4173
rect 13953 4146 13983 4173
rect 13983 4146 13987 4173
rect 14027 4146 14051 4173
rect 14051 4146 14061 4173
rect 14101 4146 14119 4173
rect 14119 4146 14135 4173
rect 14175 4146 14187 4173
rect 14187 4146 14209 4173
rect 14249 4146 14255 4173
rect 14255 4146 14283 4173
rect 14323 4146 14357 4173
rect 14397 4146 14425 4173
rect 14425 4146 14431 4173
rect 14470 4146 14493 4173
rect 14493 4146 14504 4173
rect 14543 4146 14561 4173
rect 14561 4146 14577 4173
rect 14983 4166 15017 4168
rect 13437 4073 13471 4107
rect 14983 4134 15017 4166
rect 13686 4057 13696 4091
rect 13696 4057 13720 4091
rect 13768 4057 13773 4091
rect 13773 4057 13802 4091
rect 13850 4057 13883 4091
rect 13883 4057 13884 4091
rect 13932 4057 13959 4091
rect 13959 4057 13966 4091
rect 14168 4057 14201 4091
rect 14201 4057 14202 4091
rect 14249 4057 14278 4091
rect 14278 4057 14283 4091
rect 14330 4057 14355 4091
rect 14355 4057 14364 4091
rect 14411 4057 14431 4091
rect 14431 4057 14445 4091
rect 14492 4057 14507 4091
rect 14507 4057 14526 4091
rect 14983 4064 15017 4095
rect 14983 4061 15017 4064
rect 13437 4016 13439 4034
rect 13439 4016 13471 4034
rect 13437 4000 13471 4016
rect 13437 3948 13439 3961
rect 13439 3948 13471 3961
rect 14983 3996 15017 4022
rect 14983 3988 15017 3996
rect 13437 3927 13471 3948
rect 13437 3880 13439 3888
rect 13439 3880 13471 3888
rect 13437 3854 13471 3880
rect 13437 3812 13439 3815
rect 13439 3812 13471 3815
rect 13437 3781 13471 3812
rect 13437 3710 13471 3742
rect 13437 3708 13439 3710
rect 13439 3708 13471 3710
rect 13437 3642 13471 3669
rect 13437 3635 13439 3642
rect 13439 3635 13471 3642
rect 13437 3574 13471 3596
rect 13437 3562 13439 3574
rect 13439 3562 13471 3574
rect 13437 3506 13471 3523
rect 13437 3489 13439 3506
rect 13439 3489 13471 3506
rect 13437 3438 13471 3450
rect 13437 3416 13439 3438
rect 13439 3416 13471 3438
rect 13558 3903 13592 3916
rect 13558 3882 13592 3903
rect 13558 3835 13592 3842
rect 13558 3808 13592 3835
rect 13558 3733 13592 3767
rect 13714 3903 13748 3916
rect 13714 3882 13748 3903
rect 13714 3835 13748 3842
rect 13714 3808 13748 3835
rect 13714 3733 13748 3767
rect 13830 3665 13864 3672
rect 13830 3638 13864 3665
rect 13830 3563 13864 3597
rect 13830 3495 13864 3521
rect 13830 3487 13864 3495
rect 13830 3427 13864 3445
rect 13830 3411 13864 3427
rect 13986 3937 14020 3938
rect 13986 3904 14020 3937
rect 13986 3801 14020 3804
rect 13986 3770 14020 3801
rect 14075 3937 14109 3938
rect 14075 3904 14106 3937
rect 14106 3904 14109 3937
rect 14075 3835 14106 3846
rect 14106 3835 14109 3846
rect 14075 3812 14109 3835
rect 14075 3733 14109 3753
rect 14075 3719 14106 3733
rect 14106 3719 14109 3733
rect 14262 3665 14296 3678
rect 14262 3644 14296 3665
rect 14262 3563 14296 3582
rect 14262 3548 14296 3563
rect 14262 3461 14296 3486
rect 14262 3452 14296 3461
rect 14378 3665 14412 3678
rect 14378 3644 14412 3665
rect 14378 3563 14412 3582
rect 14378 3548 14412 3563
rect 14378 3461 14412 3486
rect 14378 3452 14412 3461
rect 14534 3937 14568 3940
rect 14534 3906 14568 3937
rect 14534 3835 14568 3861
rect 14534 3827 14568 3835
rect 14534 3767 14568 3781
rect 14534 3747 14568 3767
rect 14534 3699 14568 3701
rect 14534 3667 14568 3699
rect 14534 3597 14568 3621
rect 14534 3587 14568 3597
rect 14534 3529 14568 3541
rect 14534 3507 14568 3529
rect 14983 3928 15017 3949
rect 14983 3915 15017 3928
rect 14983 3860 15017 3876
rect 14983 3842 15017 3860
rect 14983 3792 15017 3803
rect 14983 3769 15017 3792
rect 14983 3724 15017 3730
rect 14983 3696 15017 3724
rect 14983 3656 15017 3657
rect 14983 3623 15017 3656
rect 14983 3554 15017 3584
rect 14983 3550 15017 3554
rect 14983 3486 15017 3511
rect 14983 3477 15017 3486
rect 14983 3418 15017 3438
rect 13437 3370 13471 3376
rect 14983 3404 15017 3418
rect 13437 3342 13439 3370
rect 13439 3342 13471 3370
rect 13437 3268 13439 3302
rect 13439 3268 13471 3302
rect 13563 3330 13597 3364
rect 13921 3336 13955 3370
rect 13993 3336 14027 3370
rect 13563 3275 13597 3292
rect 13563 3258 13597 3275
rect 13719 3275 13753 3284
rect 13719 3250 13753 3275
rect 13835 3275 13869 3284
rect 13835 3250 13869 3275
rect 14983 3350 15017 3365
rect 14263 3275 14297 3284
rect 14263 3250 14297 3275
rect 14379 3275 14413 3284
rect 14379 3250 14413 3275
rect 14556 3309 14590 3324
rect 14556 3290 14569 3309
rect 14569 3290 14590 3309
rect 14983 3331 15017 3350
rect 14983 3282 15017 3292
rect 13205 3200 13227 3220
rect 13227 3200 13239 3220
rect 14556 3218 14590 3252
rect 14983 3258 15017 3282
rect 14983 3214 15017 3219
rect 13205 3152 13239 3162
rect 13617 3161 13624 3195
rect 13624 3161 13651 3195
rect 13751 3161 13778 3195
rect 13778 3161 13785 3195
rect 14025 3161 14059 3195
rect 14114 3161 14148 3195
rect 14202 3161 14236 3195
rect 14290 3161 14322 3195
rect 14322 3161 14324 3195
rect 14378 3161 14398 3195
rect 14398 3161 14412 3195
rect 14983 3185 15017 3214
rect 13205 3128 13227 3152
rect 13227 3128 13239 3152
rect 13205 3084 13239 3089
rect 13205 3055 13227 3084
rect 13227 3055 13239 3084
rect 11564 2955 11598 2956
rect 11640 2955 11674 2956
rect 11564 2922 11577 2955
rect 11577 2922 11598 2955
rect 11640 2922 11646 2955
rect 11646 2922 11674 2955
rect 11716 2922 11750 2956
rect 11792 2955 11826 2956
rect 11868 2955 11902 2956
rect 11943 2955 11977 2956
rect 12018 2955 12052 2956
rect 12093 2955 12127 2956
rect 12168 2955 12202 2956
rect 12243 2955 12277 2956
rect 12318 2955 12352 2956
rect 11792 2922 11819 2955
rect 11819 2922 11826 2955
rect 11868 2922 11888 2955
rect 11888 2922 11902 2955
rect 11943 2922 11957 2955
rect 11957 2922 11977 2955
rect 12018 2922 12025 2955
rect 12025 2922 12052 2955
rect 12093 2922 12127 2955
rect 12168 2922 12195 2955
rect 12195 2922 12202 2955
rect 12243 2922 12263 2955
rect 12263 2922 12277 2955
rect 12318 2922 12331 2955
rect 12331 2922 12352 2955
rect 11564 2867 11598 2880
rect 11640 2867 11674 2880
rect 11564 2846 11577 2867
rect 11577 2846 11598 2867
rect 11640 2846 11646 2867
rect 11646 2846 11674 2867
rect 11716 2846 11750 2880
rect 11792 2867 11826 2880
rect 11868 2867 11902 2880
rect 11943 2867 11977 2880
rect 12018 2867 12052 2880
rect 12093 2867 12127 2880
rect 12168 2867 12202 2880
rect 12243 2867 12277 2880
rect 12318 2867 12352 2880
rect 11792 2846 11819 2867
rect 11819 2846 11826 2867
rect 11868 2846 11888 2867
rect 11888 2846 11902 2867
rect 11943 2846 11957 2867
rect 11957 2846 11977 2867
rect 12018 2846 12025 2867
rect 12025 2846 12052 2867
rect 12093 2846 12127 2867
rect 12168 2846 12195 2867
rect 12195 2846 12202 2867
rect 12243 2846 12263 2867
rect 12263 2846 12277 2867
rect 12318 2846 12331 2867
rect 12331 2846 12352 2867
rect 11564 2779 11598 2804
rect 11640 2779 11674 2804
rect 11564 2770 11577 2779
rect 11577 2770 11598 2779
rect 11640 2770 11646 2779
rect 11646 2770 11674 2779
rect 11716 2770 11750 2804
rect 11792 2779 11826 2804
rect 11868 2779 11902 2804
rect 11943 2779 11977 2804
rect 12018 2779 12052 2804
rect 12093 2779 12127 2804
rect 12168 2779 12202 2804
rect 12243 2779 12277 2804
rect 12318 2779 12352 2804
rect 11792 2770 11819 2779
rect 11819 2770 11826 2779
rect 11868 2770 11888 2779
rect 11888 2770 11902 2779
rect 11943 2770 11957 2779
rect 11957 2770 11977 2779
rect 12018 2770 12025 2779
rect 12025 2770 12052 2779
rect 12093 2770 12127 2779
rect 12168 2770 12195 2779
rect 12195 2770 12202 2779
rect 12243 2770 12263 2779
rect 12263 2770 12277 2779
rect 12318 2770 12331 2779
rect 12331 2770 12352 2779
rect 11564 2694 11598 2728
rect 11640 2694 11674 2728
rect 11716 2694 11750 2728
rect 11792 2694 11826 2728
rect 11868 2710 11902 2728
rect 11943 2710 11977 2728
rect 12018 2710 12052 2728
rect 12093 2710 12127 2728
rect 12168 2710 12202 2728
rect 12243 2710 12277 2728
rect 12318 2710 12352 2728
rect 11868 2694 11875 2710
rect 11875 2694 11902 2710
rect 11943 2694 11945 2710
rect 11945 2694 11977 2710
rect 12018 2694 12051 2710
rect 12051 2694 12052 2710
rect 12093 2694 12121 2710
rect 12121 2694 12127 2710
rect 12168 2694 12191 2710
rect 12191 2694 12202 2710
rect 12243 2694 12261 2710
rect 12261 2694 12277 2710
rect 12318 2694 12331 2710
rect 12331 2694 12352 2710
rect 11564 2618 11598 2652
rect 11640 2618 11674 2652
rect 11716 2618 11750 2652
rect 11792 2618 11826 2652
rect 11868 2637 11902 2652
rect 11943 2637 11977 2652
rect 12018 2637 12052 2652
rect 12093 2637 12127 2652
rect 12168 2637 12202 2652
rect 12243 2637 12277 2652
rect 12318 2637 12352 2652
rect 11868 2618 11875 2637
rect 11875 2618 11902 2637
rect 11943 2618 11945 2637
rect 11945 2618 11977 2637
rect 12018 2618 12051 2637
rect 12051 2618 12052 2637
rect 12093 2618 12121 2637
rect 12121 2618 12127 2637
rect 12168 2618 12191 2637
rect 12191 2618 12202 2637
rect 12243 2618 12261 2637
rect 12261 2618 12277 2637
rect 12318 2618 12331 2637
rect 12331 2618 12352 2637
rect 11564 2542 11598 2576
rect 11640 2542 11674 2576
rect 11716 2542 11750 2576
rect 11792 2542 11826 2576
rect 11868 2564 11902 2576
rect 11943 2564 11977 2576
rect 12018 2564 12052 2576
rect 12093 2564 12127 2576
rect 12168 2564 12202 2576
rect 12243 2564 12277 2576
rect 12318 2564 12352 2576
rect 11868 2542 11875 2564
rect 11875 2542 11902 2564
rect 11943 2542 11945 2564
rect 11945 2542 11977 2564
rect 12018 2542 12051 2564
rect 12051 2542 12052 2564
rect 12093 2542 12121 2564
rect 12121 2542 12127 2564
rect 12168 2542 12191 2564
rect 12191 2542 12202 2564
rect 12243 2542 12261 2564
rect 12261 2542 12277 2564
rect 12318 2542 12331 2564
rect 12331 2542 12352 2564
rect 11564 2466 11598 2500
rect 11640 2466 11674 2500
rect 11716 2466 11750 2500
rect 11792 2466 11826 2500
rect 11868 2491 11902 2500
rect 11943 2491 11977 2500
rect 12018 2491 12052 2500
rect 12093 2491 12127 2500
rect 12168 2491 12202 2500
rect 12243 2491 12277 2500
rect 12318 2491 12352 2500
rect 11868 2466 11875 2491
rect 11875 2466 11902 2491
rect 11943 2466 11945 2491
rect 11945 2466 11977 2491
rect 12018 2466 12051 2491
rect 12051 2466 12052 2491
rect 12093 2466 12121 2491
rect 12121 2466 12127 2491
rect 12168 2466 12191 2491
rect 12191 2466 12202 2491
rect 12243 2466 12261 2491
rect 12261 2466 12277 2491
rect 12318 2466 12331 2491
rect 12331 2466 12352 2491
rect 13205 2982 13227 3016
rect 13227 2982 13239 3016
rect 13563 3081 13597 3097
rect 13563 3063 13597 3081
rect 13719 3081 13753 3106
rect 13719 3072 13753 3081
rect 13835 3081 13869 3106
rect 13835 3072 13869 3081
rect 13563 2991 13597 3025
rect 14263 3081 14297 3106
rect 14263 3072 14297 3081
rect 14379 3081 14413 3106
rect 14983 3112 15017 3146
rect 14379 3072 14413 3081
rect 14474 3060 14508 3094
rect 13991 2982 14025 3016
rect 14107 2982 14141 3016
rect 14474 2988 14508 3022
rect 14983 3044 15017 3073
rect 14983 3039 15017 3044
rect 13205 2914 13227 2943
rect 13227 2914 13239 2943
rect 13205 2909 13239 2914
rect 14983 2976 15017 3000
rect 14983 2966 15017 2976
rect 14983 2908 15017 2927
rect 14983 2893 15017 2908
rect 13205 2846 13227 2870
rect 13227 2846 13239 2870
rect 13277 2847 13295 2877
rect 13295 2847 13311 2877
rect 13352 2847 13364 2877
rect 13364 2847 13386 2877
rect 13427 2847 13433 2877
rect 13433 2847 13461 2877
rect 13205 2836 13239 2846
rect 13277 2843 13311 2847
rect 13352 2843 13386 2847
rect 13427 2843 13461 2847
rect 13502 2843 13536 2877
rect 13577 2847 13606 2877
rect 13606 2847 13611 2877
rect 13652 2847 13675 2877
rect 13675 2847 13686 2877
rect 13727 2847 13744 2877
rect 13744 2847 13761 2877
rect 13801 2847 13813 2877
rect 13813 2847 13835 2877
rect 13875 2847 13882 2877
rect 13882 2847 13909 2877
rect 13949 2847 13951 2877
rect 13951 2847 13983 2877
rect 14023 2847 14054 2877
rect 14054 2847 14057 2877
rect 14097 2847 14123 2877
rect 14123 2847 14131 2877
rect 14171 2847 14192 2877
rect 14192 2847 14205 2877
rect 14245 2847 14261 2877
rect 14261 2847 14279 2877
rect 14319 2847 14330 2877
rect 14330 2847 14353 2877
rect 14393 2847 14399 2877
rect 14399 2847 14427 2877
rect 14467 2847 14468 2877
rect 14468 2847 14501 2877
rect 14541 2847 14572 2877
rect 14572 2847 14575 2877
rect 14615 2847 14641 2877
rect 14641 2847 14649 2877
rect 14689 2847 14710 2877
rect 14710 2847 14723 2877
rect 14763 2847 14779 2877
rect 14779 2847 14797 2877
rect 14837 2847 14847 2877
rect 14847 2847 14871 2877
rect 14911 2847 14915 2877
rect 14915 2847 14945 2877
rect 13577 2843 13611 2847
rect 13652 2843 13686 2847
rect 13727 2843 13761 2847
rect 13801 2843 13835 2847
rect 13875 2843 13909 2847
rect 13949 2843 13983 2847
rect 14023 2843 14057 2847
rect 14097 2843 14131 2847
rect 14171 2843 14205 2847
rect 14245 2843 14279 2847
rect 14319 2843 14353 2847
rect 14393 2843 14427 2847
rect 14467 2843 14501 2847
rect 14541 2843 14575 2847
rect 14615 2843 14649 2847
rect 14689 2843 14723 2847
rect 14763 2843 14797 2847
rect 14837 2843 14871 2847
rect 14911 2843 14945 2847
rect 14983 2840 15017 2854
rect 13205 2778 13227 2797
rect 13227 2778 13239 2797
rect 13205 2763 13239 2778
rect 13205 2710 13227 2724
rect 13227 2710 13239 2724
rect 13205 2690 13239 2710
rect 14983 2820 15017 2840
rect 14983 2772 15017 2781
rect 14983 2747 15017 2772
rect 14983 2704 15017 2708
rect 13205 2642 13227 2651
rect 13227 2642 13239 2651
rect 13205 2617 13239 2642
rect 13205 2574 13227 2578
rect 13227 2574 13239 2578
rect 13205 2544 13239 2574
rect 11564 2390 11598 2424
rect 11640 2390 11674 2424
rect 11716 2390 11750 2424
rect 11792 2390 11826 2424
rect 11868 2418 11902 2424
rect 11943 2418 11977 2424
rect 12018 2418 12052 2424
rect 12093 2418 12127 2424
rect 12168 2418 12202 2424
rect 12243 2418 12277 2424
rect 12318 2418 12352 2424
rect 11868 2390 11875 2418
rect 11875 2390 11902 2418
rect 11943 2390 11945 2418
rect 11945 2390 11977 2418
rect 12018 2390 12051 2418
rect 12051 2390 12052 2418
rect 12093 2390 12121 2418
rect 12121 2390 12127 2418
rect 12168 2390 12191 2418
rect 12191 2390 12202 2418
rect 12243 2390 12261 2418
rect 12261 2390 12277 2418
rect 12318 2390 12331 2418
rect 12331 2390 12352 2418
rect 11564 2314 11598 2348
rect 11640 2314 11674 2348
rect 11716 2314 11750 2348
rect 11792 2314 11826 2348
rect 11868 2344 11902 2348
rect 11943 2344 11977 2348
rect 12018 2344 12052 2348
rect 12093 2344 12127 2348
rect 12168 2344 12202 2348
rect 12243 2344 12277 2348
rect 12318 2344 12352 2348
rect 11868 2314 11875 2344
rect 11875 2314 11902 2344
rect 11943 2314 11945 2344
rect 11945 2314 11977 2344
rect 12018 2314 12051 2344
rect 12051 2314 12052 2344
rect 12093 2314 12121 2344
rect 12121 2314 12127 2344
rect 12168 2314 12191 2344
rect 12191 2314 12202 2344
rect 12243 2314 12261 2344
rect 12261 2314 12277 2344
rect 12318 2314 12331 2344
rect 12331 2314 12352 2344
rect 12465 2452 12499 2486
rect 12539 2452 12573 2486
rect 12613 2452 12647 2486
rect 12687 2452 12721 2486
rect 12761 2452 12795 2486
rect 12835 2452 12869 2486
rect 12465 2336 12499 2370
rect 12539 2336 12573 2370
rect 12613 2336 12647 2370
rect 12687 2336 12721 2370
rect 12761 2336 12795 2370
rect 12835 2336 12869 2370
rect 13205 2472 13239 2505
rect 13205 2471 13227 2472
rect 13227 2471 13239 2472
rect 13205 2404 13239 2432
rect 13205 2398 13227 2404
rect 13227 2398 13239 2404
rect 13205 2336 13239 2359
rect 11564 2238 11598 2272
rect 11640 2238 11674 2272
rect 11716 2238 11750 2272
rect 11792 2238 11826 2272
rect 11868 2270 11902 2272
rect 11943 2270 11977 2272
rect 12018 2270 12052 2272
rect 12093 2270 12127 2272
rect 12168 2270 12202 2272
rect 12243 2270 12277 2272
rect 12318 2270 12352 2272
rect 11868 2238 11875 2270
rect 11875 2238 11902 2270
rect 11943 2238 11945 2270
rect 11945 2238 11977 2270
rect 12018 2238 12051 2270
rect 12051 2238 12052 2270
rect 12093 2238 12121 2270
rect 12121 2238 12127 2270
rect 12168 2238 12191 2270
rect 12191 2238 12202 2270
rect 12243 2238 12261 2270
rect 12261 2238 12277 2270
rect 12318 2238 12331 2270
rect 12331 2238 12352 2270
rect 13205 2325 13227 2336
rect 13227 2325 13239 2336
rect 13205 2268 13239 2286
rect 13205 2252 13227 2268
rect 13227 2252 13239 2268
rect 13205 2200 13239 2213
rect 13205 2179 13227 2200
rect 13227 2179 13239 2200
rect 13205 2132 13239 2140
rect 13205 2106 13227 2132
rect 13227 2106 13239 2132
rect 13205 2064 13239 2067
rect 13205 2033 13227 2064
rect 13227 2033 13239 2064
rect 13205 1962 13227 1994
rect 13227 1962 13239 1994
rect 13205 1960 13239 1962
rect 13205 1894 13227 1921
rect 13227 1894 13239 1921
rect 13205 1887 13239 1894
rect 13205 1826 13227 1848
rect 13227 1826 13239 1848
rect 13205 1814 13239 1826
rect 13205 1758 13227 1775
rect 13227 1758 13239 1775
rect 13205 1741 13239 1758
rect 13205 1690 13227 1702
rect 13227 1690 13239 1702
rect 13205 1668 13239 1690
rect 13205 1622 13227 1629
rect 13227 1622 13239 1629
rect 13205 1595 13239 1622
rect 13205 1554 13227 1556
rect 13227 1554 13239 1556
rect 13205 1522 13239 1554
rect 13205 1452 13239 1483
rect 13205 1449 13227 1452
rect 13227 1449 13239 1452
rect 13205 1384 13239 1410
rect 13205 1376 13227 1384
rect 13227 1376 13239 1384
rect 13205 1316 13239 1337
rect 13205 1303 13227 1316
rect 13227 1303 13239 1316
rect 13205 1248 13239 1264
rect 13205 1230 13227 1248
rect 13227 1230 13239 1248
rect 13205 1180 13239 1191
rect 13205 1157 13227 1180
rect 13227 1157 13239 1180
rect 13205 1112 13239 1118
rect 13205 1084 13227 1112
rect 13227 1084 13239 1112
rect 13205 1044 13239 1045
rect 13205 1011 13227 1044
rect 13227 1011 13239 1044
rect 13205 942 13227 972
rect 13227 942 13239 972
rect 13205 938 13239 942
rect 11502 805 11527 837
rect 11527 805 11536 837
rect 11576 805 11598 837
rect 11598 805 11610 837
rect 11650 805 11669 837
rect 11669 805 11684 837
rect 11724 805 11740 837
rect 11740 805 11758 837
rect 11798 805 11811 837
rect 11811 805 11832 837
rect 11872 805 11882 837
rect 11882 805 11906 837
rect 11946 805 11953 837
rect 11953 805 11980 837
rect 12020 805 12024 837
rect 12024 805 12054 837
rect 12094 805 12095 837
rect 12095 805 12128 837
rect 12168 805 12200 837
rect 12200 805 12202 837
rect 12242 805 12271 837
rect 12271 805 12276 837
rect 12316 805 12342 837
rect 12342 805 12350 837
rect 12390 805 12413 837
rect 12413 805 12424 837
rect 12464 805 12484 837
rect 12484 805 12498 837
rect 12538 805 12555 837
rect 12555 805 12572 837
rect 12611 805 12626 837
rect 12626 805 12645 837
rect 12684 805 12697 837
rect 12697 805 12718 837
rect 12757 805 12768 837
rect 12768 805 12791 837
rect 11502 803 11536 805
rect 11576 803 11610 805
rect 11650 803 11684 805
rect 11724 803 11758 805
rect 11798 803 11832 805
rect 11872 803 11906 805
rect 11946 803 11980 805
rect 12020 803 12054 805
rect 12094 803 12128 805
rect 12168 803 12202 805
rect 12242 803 12276 805
rect 12316 803 12350 805
rect 12390 803 12424 805
rect 12464 803 12498 805
rect 12538 803 12572 805
rect 12611 803 12645 805
rect 12684 803 12718 805
rect 12757 803 12791 805
rect 11502 735 11527 765
rect 11527 735 11536 765
rect 11576 735 11598 765
rect 11598 735 11610 765
rect 11650 735 11669 765
rect 11669 735 11684 765
rect 11724 735 11740 765
rect 11740 735 11758 765
rect 11798 735 11811 765
rect 11811 735 11832 765
rect 11872 735 11882 765
rect 11882 735 11906 765
rect 11946 735 11953 765
rect 11953 735 11980 765
rect 12020 735 12024 765
rect 12024 735 12054 765
rect 12094 735 12095 765
rect 12095 735 12128 765
rect 12168 735 12200 765
rect 12200 735 12202 765
rect 12242 735 12271 765
rect 12271 735 12276 765
rect 12316 735 12342 765
rect 12342 735 12350 765
rect 12390 735 12413 765
rect 12413 735 12424 765
rect 12464 735 12484 765
rect 12484 735 12498 765
rect 12538 735 12555 765
rect 12555 735 12572 765
rect 12611 735 12626 765
rect 12626 735 12645 765
rect 12684 735 12697 765
rect 12697 735 12718 765
rect 12757 735 12768 765
rect 12768 735 12791 765
rect 11502 731 11536 735
rect 11576 731 11610 735
rect 11650 731 11684 735
rect 11724 731 11758 735
rect 11798 731 11832 735
rect 11872 731 11906 735
rect 11946 731 11980 735
rect 12020 731 12054 735
rect 12094 731 12128 735
rect 12168 731 12202 735
rect 12242 731 12276 735
rect 12316 731 12350 735
rect 12390 731 12424 735
rect 12464 731 12498 735
rect 12538 731 12572 735
rect 12611 731 12645 735
rect 12684 731 12718 735
rect 12757 731 12791 735
rect 11502 665 11527 693
rect 11527 665 11536 693
rect 11576 665 11598 693
rect 11598 665 11610 693
rect 11650 665 11669 693
rect 11669 665 11684 693
rect 11724 665 11740 693
rect 11740 665 11758 693
rect 11798 665 11811 693
rect 11811 665 11832 693
rect 11872 665 11882 693
rect 11882 665 11906 693
rect 11946 665 11953 693
rect 11953 665 11980 693
rect 12020 665 12024 693
rect 12024 665 12054 693
rect 12094 665 12095 693
rect 12095 665 12128 693
rect 12168 665 12200 693
rect 12200 665 12202 693
rect 12242 665 12271 693
rect 12271 665 12276 693
rect 12316 665 12342 693
rect 12342 665 12350 693
rect 12390 665 12413 693
rect 12413 665 12424 693
rect 12464 665 12484 693
rect 12484 665 12498 693
rect 12538 665 12555 693
rect 12555 665 12572 693
rect 12611 665 12626 693
rect 12626 665 12645 693
rect 12684 665 12697 693
rect 12697 665 12718 693
rect 12757 665 12768 693
rect 12768 665 12791 693
rect 11502 659 11536 665
rect 11576 659 11610 665
rect 11650 659 11684 665
rect 11724 659 11758 665
rect 11798 659 11832 665
rect 11872 659 11906 665
rect 11946 659 11980 665
rect 12020 659 12054 665
rect 12094 659 12128 665
rect 12168 659 12202 665
rect 12242 659 12276 665
rect 12316 659 12350 665
rect 12390 659 12424 665
rect 12464 659 12498 665
rect 12538 659 12572 665
rect 12611 659 12645 665
rect 12684 659 12718 665
rect 12757 659 12791 665
rect 11502 595 11527 621
rect 11527 595 11536 621
rect 11576 595 11598 621
rect 11598 595 11610 621
rect 11650 595 11669 621
rect 11669 595 11684 621
rect 11724 595 11740 621
rect 11740 595 11758 621
rect 11798 595 11811 621
rect 11811 595 11832 621
rect 11872 595 11882 621
rect 11882 595 11906 621
rect 11946 595 11953 621
rect 11953 595 11980 621
rect 12020 595 12024 621
rect 12024 595 12054 621
rect 12094 595 12095 621
rect 12095 595 12128 621
rect 12168 595 12200 621
rect 12200 595 12202 621
rect 12242 595 12271 621
rect 12271 595 12276 621
rect 12316 595 12342 621
rect 12342 595 12350 621
rect 12390 595 12413 621
rect 12413 595 12424 621
rect 12464 595 12484 621
rect 12484 595 12498 621
rect 12538 595 12555 621
rect 12555 595 12572 621
rect 12611 595 12626 621
rect 12626 595 12645 621
rect 12684 595 12697 621
rect 12697 595 12718 621
rect 12757 595 12768 621
rect 12768 595 12791 621
rect 11502 587 11536 595
rect 11576 587 11610 595
rect 11650 587 11684 595
rect 11724 587 11758 595
rect 11798 587 11832 595
rect 11872 587 11906 595
rect 11946 587 11980 595
rect 12020 587 12054 595
rect 12094 587 12128 595
rect 12168 587 12202 595
rect 12242 587 12276 595
rect 12316 587 12350 595
rect 12390 587 12424 595
rect 12464 587 12498 595
rect 12538 587 12572 595
rect 12611 587 12645 595
rect 12684 587 12718 595
rect 12757 587 12791 595
rect 11502 525 11527 549
rect 11527 525 11536 549
rect 11576 525 11598 549
rect 11598 525 11610 549
rect 11650 525 11669 549
rect 11669 525 11684 549
rect 11724 525 11740 549
rect 11740 525 11758 549
rect 11798 525 11811 549
rect 11811 525 11832 549
rect 11872 525 11882 549
rect 11882 525 11906 549
rect 11946 525 11953 549
rect 11953 525 11980 549
rect 12020 525 12024 549
rect 12024 525 12054 549
rect 12094 525 12095 549
rect 12095 525 12128 549
rect 12168 525 12200 549
rect 12200 525 12202 549
rect 12242 525 12271 549
rect 12271 525 12276 549
rect 12316 525 12342 549
rect 12342 525 12350 549
rect 12390 525 12413 549
rect 12413 525 12424 549
rect 12464 525 12484 549
rect 12484 525 12498 549
rect 12538 525 12555 549
rect 12555 525 12572 549
rect 12611 525 12626 549
rect 12626 525 12645 549
rect 12684 525 12697 549
rect 12697 525 12718 549
rect 12757 525 12768 549
rect 12768 525 12791 549
rect 11502 515 11536 525
rect 11576 515 11610 525
rect 11650 515 11684 525
rect 11724 515 11758 525
rect 11798 515 11832 525
rect 11872 515 11906 525
rect 11946 515 11980 525
rect 12020 515 12054 525
rect 12094 515 12128 525
rect 12168 515 12202 525
rect 12242 515 12276 525
rect 12316 515 12350 525
rect 12390 515 12424 525
rect 12464 515 12498 525
rect 12538 515 12572 525
rect 12611 515 12645 525
rect 12684 515 12718 525
rect 12757 515 12791 525
rect 11502 455 11527 477
rect 11527 455 11536 477
rect 11576 455 11598 477
rect 11598 455 11610 477
rect 11650 455 11669 477
rect 11669 455 11684 477
rect 11724 455 11740 477
rect 11740 455 11758 477
rect 11798 455 11811 477
rect 11811 455 11832 477
rect 11872 455 11882 477
rect 11882 455 11906 477
rect 11946 455 11953 477
rect 11953 455 11980 477
rect 12020 455 12024 477
rect 12024 455 12054 477
rect 12094 455 12095 477
rect 12095 455 12128 477
rect 12168 455 12200 477
rect 12200 455 12202 477
rect 12242 455 12271 477
rect 12271 455 12276 477
rect 12316 455 12342 477
rect 12342 455 12350 477
rect 12390 455 12413 477
rect 12413 455 12424 477
rect 12464 455 12484 477
rect 12484 455 12498 477
rect 12538 455 12555 477
rect 12555 455 12572 477
rect 12611 455 12626 477
rect 12626 455 12645 477
rect 12684 455 12697 477
rect 12697 455 12718 477
rect 12757 455 12768 477
rect 12768 455 12791 477
rect 11502 443 11536 455
rect 11576 443 11610 455
rect 11650 443 11684 455
rect 11724 443 11758 455
rect 11798 443 11832 455
rect 11872 443 11906 455
rect 11946 443 11980 455
rect 12020 443 12054 455
rect 12094 443 12128 455
rect 12168 443 12202 455
rect 12242 443 12276 455
rect 12316 443 12350 455
rect 12390 443 12424 455
rect 12464 443 12498 455
rect 12538 443 12572 455
rect 12611 443 12645 455
rect 12684 443 12718 455
rect 12757 443 12791 455
rect 11502 385 11527 405
rect 11527 385 11536 405
rect 11576 385 11598 405
rect 11598 385 11610 405
rect 11650 385 11669 405
rect 11669 385 11684 405
rect 11724 385 11740 405
rect 11740 385 11758 405
rect 11798 385 11811 405
rect 11811 385 11832 405
rect 11872 385 11882 405
rect 11882 385 11906 405
rect 11946 385 11953 405
rect 11953 385 11980 405
rect 12020 385 12024 405
rect 12024 385 12054 405
rect 12094 385 12095 405
rect 12095 385 12128 405
rect 12168 385 12200 405
rect 12200 385 12202 405
rect 12242 385 12271 405
rect 12271 385 12276 405
rect 12316 385 12342 405
rect 12342 385 12350 405
rect 12390 385 12413 405
rect 12413 385 12424 405
rect 12464 385 12484 405
rect 12484 385 12498 405
rect 12538 385 12555 405
rect 12555 385 12572 405
rect 12611 385 12626 405
rect 12626 385 12645 405
rect 12684 385 12697 405
rect 12697 385 12718 405
rect 12757 385 12768 405
rect 12768 385 12791 405
rect 11502 371 11536 385
rect 11576 371 11610 385
rect 11650 371 11684 385
rect 11724 371 11758 385
rect 11798 371 11832 385
rect 11872 371 11906 385
rect 11946 371 11980 385
rect 12020 371 12054 385
rect 12094 371 12128 385
rect 12168 371 12202 385
rect 12242 371 12276 385
rect 12316 371 12350 385
rect 12390 371 12424 385
rect 12464 371 12498 385
rect 12538 371 12572 385
rect 12611 371 12645 385
rect 12684 371 12718 385
rect 12757 371 12791 385
rect 11502 315 11527 333
rect 11527 315 11536 333
rect 11576 315 11598 333
rect 11598 315 11610 333
rect 11650 315 11669 333
rect 11669 315 11684 333
rect 11724 315 11740 333
rect 11740 315 11758 333
rect 11798 315 11811 333
rect 11811 315 11832 333
rect 11872 315 11882 333
rect 11882 315 11906 333
rect 11946 315 11953 333
rect 11953 315 11980 333
rect 12020 315 12024 333
rect 12024 315 12054 333
rect 12094 315 12095 333
rect 12095 315 12128 333
rect 12168 315 12200 333
rect 12200 315 12202 333
rect 12242 315 12271 333
rect 12271 315 12276 333
rect 12316 315 12342 333
rect 12342 315 12350 333
rect 12390 315 12413 333
rect 12413 315 12424 333
rect 12464 315 12484 333
rect 12484 315 12498 333
rect 12538 315 12555 333
rect 12555 315 12572 333
rect 12611 315 12626 333
rect 12626 315 12645 333
rect 12684 315 12697 333
rect 12697 315 12718 333
rect 12757 315 12768 333
rect 12768 315 12791 333
rect 11502 299 11536 315
rect 11576 299 11610 315
rect 11650 299 11684 315
rect 11724 299 11758 315
rect 11798 299 11832 315
rect 11872 299 11906 315
rect 11946 299 11980 315
rect 12020 299 12054 315
rect 12094 299 12128 315
rect 12168 299 12202 315
rect 12242 299 12276 315
rect 12316 299 12350 315
rect 12390 299 12424 315
rect 12464 299 12498 315
rect 12538 299 12572 315
rect 12611 299 12645 315
rect 12684 299 12718 315
rect 12757 299 12791 315
rect 11502 245 11527 261
rect 11527 245 11536 261
rect 11576 245 11598 261
rect 11598 245 11610 261
rect 11650 245 11669 261
rect 11669 245 11684 261
rect 11724 245 11740 261
rect 11740 245 11758 261
rect 11798 245 11811 261
rect 11811 245 11832 261
rect 11872 245 11882 261
rect 11882 245 11906 261
rect 11946 245 11953 261
rect 11953 245 11980 261
rect 12020 245 12024 261
rect 12024 245 12054 261
rect 12094 245 12095 261
rect 12095 245 12128 261
rect 12168 245 12200 261
rect 12200 245 12202 261
rect 12242 245 12271 261
rect 12271 245 12276 261
rect 12316 245 12342 261
rect 12342 245 12350 261
rect 12390 245 12413 261
rect 12413 245 12424 261
rect 12464 245 12484 261
rect 12484 245 12498 261
rect 12538 245 12555 261
rect 12555 245 12572 261
rect 12611 245 12626 261
rect 12626 245 12645 261
rect 12684 245 12697 261
rect 12697 245 12718 261
rect 12757 245 12768 261
rect 12768 245 12791 261
rect 11502 227 11536 245
rect 11576 227 11610 245
rect 11650 227 11684 245
rect 11724 227 11758 245
rect 11798 227 11832 245
rect 11872 227 11906 245
rect 11946 227 11980 245
rect 12020 227 12054 245
rect 12094 227 12128 245
rect 12168 227 12202 245
rect 12242 227 12276 245
rect 12316 227 12350 245
rect 12390 227 12424 245
rect 12464 227 12498 245
rect 12538 227 12572 245
rect 12611 227 12645 245
rect 12684 227 12718 245
rect 12757 227 12791 245
rect 11502 175 11527 189
rect 11527 175 11536 189
rect 11576 175 11598 189
rect 11598 175 11610 189
rect 11650 175 11669 189
rect 11669 175 11684 189
rect 11724 175 11740 189
rect 11740 175 11758 189
rect 11798 175 11811 189
rect 11811 175 11832 189
rect 11872 175 11882 189
rect 11882 175 11906 189
rect 11946 175 11953 189
rect 11953 175 11980 189
rect 12020 175 12024 189
rect 12024 175 12054 189
rect 12094 175 12095 189
rect 12095 175 12128 189
rect 12168 175 12200 189
rect 12200 175 12202 189
rect 12242 175 12271 189
rect 12271 175 12276 189
rect 12316 175 12342 189
rect 12342 175 12350 189
rect 12390 175 12413 189
rect 12413 175 12424 189
rect 12464 175 12484 189
rect 12484 175 12498 189
rect 12538 175 12555 189
rect 12555 175 12572 189
rect 12611 175 12626 189
rect 12626 175 12645 189
rect 12684 175 12697 189
rect 12697 175 12718 189
rect 12757 175 12768 189
rect 12768 175 12791 189
rect 11502 155 11536 175
rect 11576 155 11610 175
rect 11650 155 11684 175
rect 11724 155 11758 175
rect 11798 155 11832 175
rect 11872 155 11906 175
rect 11946 155 11980 175
rect 12020 155 12054 175
rect 12094 155 12128 175
rect 12168 155 12202 175
rect 12242 155 12276 175
rect 12316 155 12350 175
rect 12390 155 12424 175
rect 12464 155 12498 175
rect 12538 155 12572 175
rect 12611 155 12645 175
rect 12684 155 12718 175
rect 12757 155 12791 175
rect 11502 105 11527 117
rect 11527 105 11536 117
rect 11576 105 11598 117
rect 11598 105 11610 117
rect 11650 105 11669 117
rect 11669 105 11684 117
rect 11724 105 11740 117
rect 11740 105 11758 117
rect 11798 105 11811 117
rect 11811 105 11832 117
rect 11872 105 11882 117
rect 11882 105 11906 117
rect 11946 105 11953 117
rect 11953 105 11980 117
rect 12020 105 12024 117
rect 12024 105 12054 117
rect 12094 105 12095 117
rect 12095 105 12128 117
rect 12168 105 12200 117
rect 12200 105 12202 117
rect 12242 105 12271 117
rect 12271 105 12276 117
rect 12316 105 12342 117
rect 12342 105 12350 117
rect 12390 105 12413 117
rect 12413 105 12424 117
rect 12464 105 12484 117
rect 12484 105 12498 117
rect 12538 105 12555 117
rect 12555 105 12572 117
rect 12611 105 12626 117
rect 12626 105 12645 117
rect 12684 105 12697 117
rect 12697 105 12718 117
rect 12757 105 12768 117
rect 12768 105 12791 117
rect 11502 83 11536 105
rect 11576 83 11610 105
rect 11650 83 11684 105
rect 11724 83 11758 105
rect 11798 83 11832 105
rect 11872 83 11906 105
rect 11946 83 11980 105
rect 12020 83 12054 105
rect 12094 83 12128 105
rect 12168 83 12202 105
rect 12242 83 12276 105
rect 12316 83 12350 105
rect 12390 83 12424 105
rect 12464 83 12498 105
rect 12538 83 12572 105
rect 12611 83 12645 105
rect 12684 83 12718 105
rect 12757 83 12791 105
rect 11346 -1 11380 15
rect 11346 -19 11348 -1
rect 11348 -19 11380 -1
rect 11420 -19 11454 15
rect 11494 -1 11528 15
rect 11567 -1 11601 15
rect 11640 -1 11674 15
rect 11494 -19 11527 -1
rect 11527 -19 11528 -1
rect 11567 -19 11598 -1
rect 11598 -19 11601 -1
rect 11640 -19 11669 -1
rect 11669 -19 11674 -1
rect 13205 874 13227 899
rect 13227 874 13239 899
rect 13205 865 13239 874
rect 13205 806 13227 826
rect 13227 806 13239 826
rect 13205 792 13239 806
rect 13205 738 13227 753
rect 13227 738 13239 753
rect 13205 719 13239 738
rect 13205 670 13227 680
rect 13227 670 13239 680
rect 13205 646 13239 670
rect 13205 602 13227 607
rect 13227 602 13239 607
rect 13205 573 13239 602
rect 13205 500 13239 534
rect 13205 432 13239 461
rect 13205 427 13227 432
rect 13227 427 13239 432
rect 13205 364 13239 388
rect 13205 354 13227 364
rect 13227 354 13239 364
rect 13205 296 13239 315
rect 13205 281 13227 296
rect 13227 281 13239 296
rect 13205 228 13239 242
rect 13511 2658 13541 2692
rect 13541 2658 13545 2692
rect 13586 2658 13609 2692
rect 13609 2658 13620 2692
rect 13661 2658 13677 2692
rect 13677 2658 13695 2692
rect 13736 2658 13745 2692
rect 13745 2658 13770 2692
rect 13811 2658 13813 2692
rect 13813 2658 13845 2692
rect 13886 2658 13915 2692
rect 13915 2658 13920 2692
rect 13961 2658 13983 2692
rect 13983 2658 13995 2692
rect 14036 2658 14051 2692
rect 14051 2658 14070 2692
rect 14111 2658 14119 2692
rect 14119 2658 14145 2692
rect 14186 2658 14187 2692
rect 14187 2658 14220 2692
rect 14261 2658 14289 2692
rect 14289 2658 14295 2692
rect 14335 2658 14357 2692
rect 14357 2658 14369 2692
rect 14409 2658 14425 2692
rect 14425 2658 14443 2692
rect 14483 2658 14493 2692
rect 14493 2658 14517 2692
rect 14557 2658 14561 2692
rect 14561 2658 14591 2692
rect 14631 2658 14665 2692
rect 13439 2588 13473 2592
rect 13439 2558 13473 2588
rect 14705 2590 14739 2620
rect 14705 2586 14739 2590
rect 14167 2539 14176 2573
rect 14176 2539 14201 2573
rect 14240 2539 14244 2573
rect 14244 2539 14274 2573
rect 14312 2539 14346 2573
rect 14384 2539 14414 2573
rect 14414 2539 14418 2573
rect 14456 2539 14482 2573
rect 14482 2539 14490 2573
rect 14528 2539 14550 2573
rect 14550 2539 14562 2573
rect 14600 2539 14618 2573
rect 14618 2539 14634 2573
rect 13439 2486 13473 2492
rect 13439 2458 13473 2486
rect 13439 2350 13473 2382
rect 13439 2348 13473 2350
rect 13439 2282 13473 2310
rect 13439 2276 13473 2282
rect 13439 2214 13473 2238
rect 13439 2204 13473 2214
rect 13439 2146 13473 2166
rect 13439 2132 13473 2146
rect 13439 2078 13473 2094
rect 13439 2060 13473 2078
rect 13439 2010 13473 2021
rect 13439 1987 13473 2010
rect 13439 1942 13473 1948
rect 13439 1914 13473 1942
rect 13439 1874 13473 1875
rect 13439 1841 13473 1874
rect 13439 1772 13473 1802
rect 13439 1768 13473 1772
rect 13439 1704 13473 1729
rect 13439 1695 13473 1704
rect 13439 1622 13473 1656
rect 13439 1562 13473 1583
rect 13439 1549 13473 1562
rect 13439 1494 13473 1510
rect 13439 1476 13473 1494
rect 13439 1426 13473 1437
rect 13439 1403 13473 1426
rect 13439 1358 13473 1364
rect 13439 1330 13473 1358
rect 13439 1290 13473 1291
rect 13439 1257 13473 1290
rect 13439 1188 13473 1218
rect 13439 1184 13473 1188
rect 13439 1120 13473 1145
rect 13439 1111 13473 1120
rect 13439 1052 13473 1072
rect 13439 1038 13473 1052
rect 13439 984 13473 999
rect 13439 965 13473 984
rect 13439 916 13473 926
rect 13439 892 13473 916
rect 13439 848 13473 853
rect 13439 819 13473 848
rect 13439 746 13473 780
rect 13439 678 13473 707
rect 13439 673 13473 678
rect 13439 610 13473 634
rect 13439 600 13473 610
rect 13439 542 13473 561
rect 13439 527 13473 542
rect 13439 474 13473 488
rect 13439 454 13473 474
rect 13439 406 13473 415
rect 13439 381 13473 406
rect 13554 2512 13588 2516
rect 13554 2482 13588 2512
rect 13554 2409 13588 2443
rect 14705 2522 14739 2546
rect 14705 2512 14739 2522
rect 14705 2454 14739 2472
rect 14705 2438 14739 2454
rect 13684 2383 13700 2417
rect 13700 2383 13718 2417
rect 13757 2383 13768 2417
rect 13768 2383 13791 2417
rect 13830 2383 13836 2417
rect 13836 2383 13864 2417
rect 13903 2383 13904 2417
rect 13904 2383 13937 2417
rect 13975 2383 14006 2417
rect 14006 2383 14009 2417
rect 14047 2383 14074 2417
rect 14074 2383 14081 2417
rect 13554 2340 13588 2370
rect 13554 2336 13588 2340
rect 13554 2271 13588 2297
rect 13554 2263 13588 2271
rect 14705 2386 14739 2398
rect 14705 2364 14739 2386
rect 14705 2318 14739 2324
rect 14705 2290 14739 2318
rect 14167 2227 14176 2261
rect 14176 2227 14201 2261
rect 14240 2227 14244 2261
rect 14244 2227 14274 2261
rect 14312 2227 14346 2261
rect 14384 2227 14414 2261
rect 14414 2227 14418 2261
rect 14456 2227 14482 2261
rect 14482 2227 14490 2261
rect 14528 2227 14550 2261
rect 14550 2227 14562 2261
rect 14600 2227 14618 2261
rect 14618 2227 14634 2261
rect 13554 2202 13588 2224
rect 13554 2190 13588 2202
rect 13554 2133 13588 2150
rect 13554 2116 13588 2133
rect 14705 2216 14739 2250
rect 14705 2148 14739 2176
rect 14705 2142 14739 2148
rect 13554 2064 13588 2076
rect 13684 2071 13700 2105
rect 13700 2071 13718 2105
rect 13757 2071 13768 2105
rect 13768 2071 13791 2105
rect 13830 2071 13836 2105
rect 13836 2071 13864 2105
rect 13903 2071 13904 2105
rect 13904 2071 13937 2105
rect 13975 2071 14006 2105
rect 14006 2071 14009 2105
rect 14047 2071 14074 2105
rect 14074 2071 14081 2105
rect 13554 2042 13588 2064
rect 13554 1995 13588 2002
rect 13554 1968 13588 1995
rect 14705 2080 14739 2102
rect 14705 2068 14739 2080
rect 14705 2012 14739 2028
rect 14705 1994 14739 2012
rect 13554 1926 13588 1928
rect 13554 1894 13588 1926
rect 14167 1915 14176 1949
rect 14176 1915 14201 1949
rect 14240 1915 14244 1949
rect 14244 1915 14274 1949
rect 14312 1915 14346 1949
rect 14384 1915 14414 1949
rect 14414 1915 14418 1949
rect 14456 1915 14482 1949
rect 14482 1915 14490 1949
rect 14528 1915 14550 1949
rect 14550 1915 14562 1949
rect 14600 1915 14618 1949
rect 14618 1915 14634 1949
rect 13554 1822 13588 1854
rect 13554 1820 13588 1822
rect 14705 1944 14739 1954
rect 14705 1920 14739 1944
rect 14705 1876 14739 1880
rect 14705 1846 14739 1876
rect 13554 1753 13588 1780
rect 13684 1759 13700 1793
rect 13700 1759 13718 1793
rect 13757 1759 13768 1793
rect 13768 1759 13791 1793
rect 13830 1759 13836 1793
rect 13836 1759 13864 1793
rect 13903 1759 13904 1793
rect 13904 1759 13937 1793
rect 13975 1759 14006 1793
rect 14006 1759 14009 1793
rect 14047 1759 14074 1793
rect 14074 1759 14081 1793
rect 14705 1774 14739 1806
rect 14705 1772 14739 1774
rect 13554 1746 13588 1753
rect 13554 1684 13588 1706
rect 13554 1672 13588 1684
rect 14705 1706 14739 1732
rect 14705 1698 14739 1706
rect 13554 1615 13588 1632
rect 13554 1598 13588 1615
rect 14167 1603 14176 1637
rect 14176 1603 14201 1637
rect 14240 1603 14244 1637
rect 14244 1603 14274 1637
rect 14312 1603 14346 1637
rect 14384 1603 14414 1637
rect 14414 1603 14418 1637
rect 14456 1603 14482 1637
rect 14482 1603 14490 1637
rect 14528 1603 14550 1637
rect 14550 1603 14562 1637
rect 14600 1603 14618 1637
rect 14618 1603 14634 1637
rect 14705 1638 14739 1658
rect 14705 1624 14739 1638
rect 13554 1546 13588 1558
rect 13554 1524 13588 1546
rect 13554 1477 13588 1484
rect 14705 1570 14739 1584
rect 14705 1550 14739 1570
rect 13554 1450 13588 1477
rect 13684 1447 13700 1481
rect 13700 1447 13718 1481
rect 13757 1447 13768 1481
rect 13768 1447 13791 1481
rect 13830 1447 13836 1481
rect 13836 1447 13864 1481
rect 13903 1447 13904 1481
rect 13904 1447 13937 1481
rect 13975 1447 14006 1481
rect 14006 1447 14009 1481
rect 14047 1447 14074 1481
rect 14074 1447 14081 1481
rect 14705 1502 14739 1511
rect 14705 1477 14739 1502
rect 13554 1408 13588 1410
rect 13554 1376 13588 1408
rect 13554 1305 13588 1336
rect 14705 1434 14739 1438
rect 14705 1404 14739 1434
rect 13554 1302 13588 1305
rect 14167 1291 14176 1325
rect 14176 1291 14201 1325
rect 14240 1291 14244 1325
rect 14244 1291 14274 1325
rect 14312 1291 14346 1325
rect 14384 1291 14414 1325
rect 14414 1291 14418 1325
rect 14456 1291 14482 1325
rect 14482 1291 14490 1325
rect 14528 1291 14550 1325
rect 14550 1291 14562 1325
rect 14600 1291 14618 1325
rect 14618 1291 14634 1325
rect 14705 1332 14739 1365
rect 14705 1331 14739 1332
rect 13554 1236 13588 1262
rect 13554 1228 13588 1236
rect 13554 1167 13588 1188
rect 14705 1264 14739 1292
rect 14705 1258 14739 1264
rect 13554 1154 13588 1167
rect 13684 1135 13700 1169
rect 13700 1135 13718 1169
rect 13757 1135 13768 1169
rect 13768 1135 13791 1169
rect 13830 1135 13836 1169
rect 13836 1135 13864 1169
rect 13903 1135 13904 1169
rect 13904 1135 13937 1169
rect 13975 1135 14006 1169
rect 14006 1135 14009 1169
rect 14047 1135 14074 1169
rect 14074 1135 14081 1169
rect 14705 1196 14739 1219
rect 14705 1185 14739 1196
rect 13554 1098 13588 1114
rect 13554 1080 13588 1098
rect 13554 1029 13588 1040
rect 13554 1006 13588 1029
rect 14705 1128 14739 1146
rect 14705 1112 14739 1128
rect 14705 1060 14739 1073
rect 14705 1039 14739 1060
rect 14167 979 14176 1013
rect 14176 979 14201 1013
rect 14240 979 14244 1013
rect 14244 979 14274 1013
rect 14312 979 14346 1013
rect 14384 979 14414 1013
rect 14414 979 14418 1013
rect 14456 979 14482 1013
rect 14482 979 14490 1013
rect 14528 979 14550 1013
rect 14550 979 14562 1013
rect 14600 979 14618 1013
rect 14618 979 14634 1013
rect 13554 960 13588 966
rect 13554 932 13588 960
rect 13554 858 13588 892
rect 14705 992 14739 1000
rect 14705 966 14739 992
rect 14705 924 14739 927
rect 14705 893 14739 924
rect 13684 823 13700 857
rect 13700 823 13718 857
rect 13757 823 13768 857
rect 13768 823 13791 857
rect 13830 823 13836 857
rect 13836 823 13864 857
rect 13903 823 13904 857
rect 13904 823 13937 857
rect 13975 823 14006 857
rect 14006 823 14009 857
rect 14047 823 14074 857
rect 14074 823 14081 857
rect 13554 790 13588 818
rect 13554 784 13588 790
rect 13554 722 13588 744
rect 13554 710 13588 722
rect 14705 822 14739 854
rect 14705 820 14739 822
rect 14705 754 14739 781
rect 14705 747 14739 754
rect 13554 654 13588 670
rect 14167 667 14176 701
rect 14176 667 14201 701
rect 14240 667 14244 701
rect 14244 667 14274 701
rect 14312 667 14346 701
rect 14384 667 14414 701
rect 14414 667 14418 701
rect 14456 667 14482 701
rect 14482 667 14490 701
rect 14528 667 14550 701
rect 14550 667 14562 701
rect 14600 667 14618 701
rect 14618 667 14634 701
rect 14705 686 14739 708
rect 14705 674 14739 686
rect 13554 636 13588 654
rect 13554 586 13588 596
rect 13554 562 13588 586
rect 14705 618 14739 635
rect 14705 601 14739 618
rect 13554 518 13588 522
rect 13554 488 13588 518
rect 13684 511 13700 545
rect 13700 511 13718 545
rect 13757 511 13768 545
rect 13768 511 13791 545
rect 13830 511 13836 545
rect 13836 511 13864 545
rect 13903 511 13904 545
rect 13904 511 13937 545
rect 13975 511 14006 545
rect 14006 511 14009 545
rect 14047 511 14074 545
rect 14074 511 14081 545
rect 14705 550 14739 562
rect 14705 528 14739 550
rect 14705 482 14739 489
rect 14705 455 14739 482
rect 14167 355 14176 389
rect 14176 355 14201 389
rect 14240 355 14244 389
rect 14244 355 14274 389
rect 14312 355 14346 389
rect 14384 355 14414 389
rect 14414 355 14418 389
rect 14456 355 14482 389
rect 14482 355 14490 389
rect 14528 355 14550 389
rect 14550 355 14562 389
rect 14600 355 14618 389
rect 14618 355 14634 389
rect 14705 414 14739 416
rect 14705 382 14739 414
rect 13439 338 13473 342
rect 13439 308 13473 338
rect 14705 309 14739 343
rect 13513 236 13547 270
rect 13587 236 13617 270
rect 13617 236 13621 270
rect 13661 236 13685 270
rect 13685 236 13695 270
rect 13735 236 13753 270
rect 13753 236 13769 270
rect 13809 236 13821 270
rect 13821 236 13843 270
rect 13883 236 13889 270
rect 13889 236 13917 270
rect 13958 236 13991 270
rect 13991 236 13992 270
rect 14033 236 14059 270
rect 14059 236 14067 270
rect 14108 236 14127 270
rect 14127 236 14142 270
rect 14183 236 14195 270
rect 14195 236 14217 270
rect 14258 236 14263 270
rect 14263 236 14292 270
rect 14333 236 14365 270
rect 14365 236 14367 270
rect 14408 236 14433 270
rect 14433 236 14442 270
rect 14483 236 14501 270
rect 14501 236 14517 270
rect 14558 236 14569 270
rect 14569 236 14592 270
rect 14633 236 14637 270
rect 14637 236 14667 270
rect 14983 2674 15017 2704
rect 14983 2602 15017 2635
rect 14983 2601 15017 2602
rect 14983 2534 15017 2562
rect 14983 2528 15017 2534
rect 14983 2466 15017 2489
rect 14983 2455 15017 2466
rect 14983 2398 15017 2416
rect 14983 2382 15017 2398
rect 14983 2330 15017 2343
rect 14983 2309 15017 2330
rect 14983 2262 15017 2270
rect 14983 2236 15017 2262
rect 14983 2194 15017 2197
rect 14983 2163 15017 2194
rect 14983 2092 15017 2124
rect 14983 2090 15017 2092
rect 14983 2024 15017 2051
rect 14983 2017 15017 2024
rect 14983 1956 15017 1978
rect 14983 1944 15017 1956
rect 14983 1888 15017 1905
rect 14983 1871 15017 1888
rect 14983 1820 15017 1832
rect 14983 1798 15017 1820
rect 14983 1752 15017 1759
rect 14983 1725 15017 1752
rect 14983 1684 15017 1686
rect 14983 1652 15017 1684
rect 14983 1582 15017 1613
rect 14983 1579 15017 1582
rect 14983 1514 15017 1540
rect 14983 1506 15017 1514
rect 14983 1446 15017 1467
rect 14983 1433 15017 1446
rect 14983 1378 15017 1394
rect 14983 1360 15017 1378
rect 14983 1310 15017 1321
rect 14983 1287 15017 1310
rect 14983 1242 15017 1248
rect 14983 1214 15017 1242
rect 14983 1174 15017 1176
rect 14983 1142 15017 1174
rect 14983 1072 15017 1104
rect 14983 1070 15017 1072
rect 14983 1004 15017 1032
rect 14983 998 15017 1004
rect 14983 936 15017 960
rect 14983 926 15017 936
rect 14983 868 15017 888
rect 14983 854 15017 868
rect 14983 800 15017 816
rect 14983 782 15017 800
rect 14983 732 15017 744
rect 14983 710 15017 732
rect 14983 664 15017 672
rect 14983 638 15017 664
rect 14983 596 15017 600
rect 14983 566 15017 596
rect 14983 494 15017 528
rect 14983 426 15017 456
rect 14983 422 15017 426
rect 14983 358 15017 384
rect 14983 350 15017 358
rect 14983 290 15017 312
rect 14983 278 15017 290
rect 13205 208 13227 228
rect 13227 208 13239 228
rect 13205 160 13239 169
rect 13205 135 13227 160
rect 13227 135 13239 160
rect 13205 92 13239 96
rect 13205 62 13227 92
rect 13227 62 13239 92
rect 14983 222 15017 240
rect 14983 206 15017 222
rect 14983 154 15017 168
rect 14983 134 15017 154
rect 14983 86 15017 96
rect 14983 62 15017 86
rect 13279 -10 13283 24
rect 13283 -10 13313 24
rect 13353 -10 13385 24
rect 13385 -10 13387 24
rect 13427 -10 13453 24
rect 13453 -10 13461 24
rect 13501 -10 13521 24
rect 13521 -10 13535 24
rect 13575 -10 13589 24
rect 13589 -10 13609 24
rect 13649 -10 13657 24
rect 13657 -10 13683 24
rect 13723 -10 13725 24
rect 13725 -10 13757 24
rect 13797 -10 13827 24
rect 13827 -10 13831 24
rect 13871 -10 13895 24
rect 13895 -10 13905 24
rect 13945 -10 13963 24
rect 13963 -10 13979 24
rect 14019 -10 14031 24
rect 14031 -10 14053 24
rect 14093 -10 14099 24
rect 14099 -10 14127 24
rect 14167 -10 14201 24
rect 14241 -10 14269 24
rect 14269 -10 14275 24
rect 14315 -10 14337 24
rect 14337 -10 14349 24
rect 14389 -10 14405 24
rect 14405 -10 14423 24
rect 14463 -10 14473 24
rect 14473 -10 14497 24
rect 14537 -10 14541 24
rect 14541 -10 14571 24
rect 14611 -10 14643 24
rect 14643 -10 14645 24
rect 14686 -10 14711 24
rect 14711 -10 14720 24
rect 14761 -10 14779 24
rect 14779 -10 14795 24
rect 14836 -10 14847 24
rect 14847 -10 14870 24
rect 14911 -10 14915 24
rect 14915 -10 14945 24
rect 11346 -71 11380 -57
rect 11346 -91 11348 -71
rect 11348 -91 11380 -71
rect 11420 -91 11454 -57
rect 11494 -71 11528 -57
rect 11567 -71 11601 -57
rect 11640 -71 11674 -57
rect 11494 -91 11527 -71
rect 11527 -91 11528 -71
rect 11567 -91 11598 -71
rect 11598 -91 11601 -71
rect 11640 -91 11669 -71
rect 11669 -91 11674 -71
rect 12322 -782 12350 -768
rect 12350 -782 12356 -768
rect 12399 -782 12418 -768
rect 12418 -782 12433 -768
rect 12475 -782 12486 -768
rect 12486 -782 12509 -768
rect 12551 -782 12554 -768
rect 12554 -782 12585 -768
rect 12627 -782 12656 -768
rect 12656 -782 12661 -768
rect 12703 -782 12724 -768
rect 12724 -782 12737 -768
rect 12322 -802 12356 -782
rect 12399 -802 12433 -782
rect 12475 -802 12509 -782
rect 12551 -802 12585 -782
rect 12627 -802 12661 -782
rect 12703 -802 12737 -782
rect 12322 -853 12350 -840
rect 12350 -853 12356 -840
rect 12399 -853 12418 -840
rect 12418 -853 12433 -840
rect 12475 -853 12486 -840
rect 12486 -853 12509 -840
rect 12551 -853 12554 -840
rect 12554 -853 12585 -840
rect 12627 -853 12656 -840
rect 12656 -853 12661 -840
rect 12703 -853 12724 -840
rect 12724 -853 12737 -840
rect 12322 -874 12356 -853
rect 12399 -874 12433 -853
rect 12475 -874 12509 -853
rect 12551 -874 12585 -853
rect 12627 -874 12661 -853
rect 12703 -874 12737 -853
rect 12322 -924 12350 -912
rect 12350 -924 12356 -912
rect 12399 -924 12418 -912
rect 12418 -924 12433 -912
rect 12475 -924 12486 -912
rect 12486 -924 12509 -912
rect 12551 -924 12554 -912
rect 12554 -924 12585 -912
rect 12627 -924 12656 -912
rect 12656 -924 12661 -912
rect 12703 -924 12724 -912
rect 12724 -924 12737 -912
rect 12322 -946 12356 -924
rect 12399 -946 12433 -924
rect 12475 -946 12509 -924
rect 12551 -946 12585 -924
rect 12627 -946 12661 -924
rect 12703 -946 12737 -924
<< metal1 >>
rect 7820 9819 8157 9825
rect 7820 9813 7995 9819
rect 7820 9779 7826 9813
rect 7860 9779 7942 9813
rect 7976 9779 7995 9813
rect 7820 9767 7995 9779
rect 8047 9767 8105 9819
rect 7820 9739 8157 9767
rect 7820 9705 7826 9739
rect 7860 9705 7942 9739
rect 7976 9728 8157 9739
rect 7976 9705 7995 9728
rect 7820 9676 7995 9705
rect 8047 9676 8105 9728
rect 7820 9665 8157 9676
rect 7820 9631 7826 9665
rect 7860 9631 7942 9665
rect 7976 9637 8157 9665
rect 7976 9631 7995 9637
rect 7820 9591 7995 9631
rect 7820 9557 7826 9591
rect 7860 9557 7942 9591
rect 7976 9585 7995 9591
rect 8047 9585 8105 9637
rect 7976 9557 8157 9585
rect 7820 9546 8157 9557
rect 7820 9517 7995 9546
rect 7820 9483 7826 9517
rect 7860 9483 7942 9517
rect 7976 9494 7995 9517
rect 8047 9494 8105 9546
rect 7976 9483 8157 9494
rect 7820 9455 8157 9483
rect 7820 9443 7995 9455
rect 7820 9409 7826 9443
rect 7860 9409 7942 9443
rect 7976 9409 7995 9443
rect 7820 9403 7995 9409
rect 8047 9403 8105 9455
rect 7820 9397 8157 9403
rect 9212 9819 9513 9825
rect 9212 9767 9213 9819
rect 9265 9767 9305 9819
rect 9357 9813 9397 9819
rect 9391 9779 9397 9813
rect 9357 9767 9397 9779
rect 9449 9813 9513 9819
rect 9449 9779 9473 9813
rect 9507 9779 9513 9813
rect 9449 9767 9513 9779
rect 9212 9739 9513 9767
rect 9212 9728 9357 9739
rect 9212 9676 9213 9728
rect 9265 9676 9305 9728
rect 9391 9728 9473 9739
rect 9391 9705 9397 9728
rect 9357 9676 9397 9705
rect 9449 9705 9473 9728
rect 9507 9705 9513 9739
rect 9449 9676 9513 9705
rect 9212 9665 9513 9676
rect 9212 9637 9357 9665
rect 9212 9585 9213 9637
rect 9265 9585 9305 9637
rect 9391 9637 9473 9665
rect 9391 9631 9397 9637
rect 9357 9591 9397 9631
rect 9212 9557 9357 9585
rect 9391 9585 9397 9591
rect 9449 9631 9473 9637
rect 9507 9631 9513 9665
rect 9449 9591 9513 9631
rect 9449 9585 9473 9591
rect 9391 9557 9473 9585
rect 9507 9557 9513 9591
rect 9212 9546 9513 9557
rect 9212 9494 9213 9546
rect 9265 9494 9305 9546
rect 9357 9517 9397 9546
rect 9212 9483 9357 9494
rect 9391 9494 9397 9517
rect 9449 9517 9513 9546
rect 9449 9494 9473 9517
rect 9391 9483 9473 9494
rect 9507 9483 9513 9517
rect 9212 9455 9513 9483
rect 9212 9403 9213 9455
rect 9265 9403 9305 9455
rect 9357 9443 9397 9455
rect 9391 9409 9397 9443
rect 9357 9403 9397 9409
rect 9449 9443 9513 9455
rect 9449 9409 9473 9443
rect 9507 9409 9513 9443
rect 9449 9403 9513 9409
rect 9212 9397 9513 9403
rect 788 8791 4773 8803
rect 788 8779 911 8791
rect 788 8745 800 8779
rect 834 8757 911 8779
rect 945 8757 983 8791
rect 1017 8757 1055 8791
rect 1089 8757 1127 8791
rect 1161 8757 1199 8791
rect 1233 8757 1271 8791
rect 1305 8757 1343 8791
rect 1377 8757 1415 8791
rect 1449 8757 1487 8791
rect 1521 8757 1559 8791
rect 1593 8757 1631 8791
rect 1665 8757 1703 8791
rect 1737 8757 1775 8791
rect 1809 8757 1847 8791
rect 1881 8757 1919 8791
rect 1953 8757 1991 8791
rect 2025 8757 2063 8791
rect 2097 8757 2135 8791
rect 2169 8757 2207 8791
rect 2241 8757 2279 8791
rect 2313 8757 2351 8791
rect 2385 8757 2423 8791
rect 2457 8757 2495 8791
rect 2529 8757 2567 8791
rect 2601 8757 2639 8791
rect 2673 8757 2711 8791
rect 2745 8757 2783 8791
rect 2817 8757 2855 8791
rect 2889 8757 2927 8791
rect 2961 8757 2999 8791
rect 3033 8757 3071 8791
rect 3105 8757 3143 8791
rect 3177 8757 3215 8791
rect 3249 8757 3287 8791
rect 3321 8757 3359 8791
rect 3393 8757 3431 8791
rect 3465 8757 3503 8791
rect 3537 8757 3575 8791
rect 3609 8757 3647 8791
rect 3681 8757 3719 8791
rect 3753 8757 3791 8791
rect 3825 8757 3863 8791
rect 3897 8757 3935 8791
rect 3969 8757 4007 8791
rect 4041 8757 4079 8791
rect 4113 8757 4151 8791
rect 4185 8757 4223 8791
rect 4257 8757 4295 8791
rect 4329 8757 4367 8791
rect 4401 8757 4439 8791
rect 4473 8757 4511 8791
rect 4545 8757 4583 8791
rect 4617 8757 4655 8791
rect 4689 8757 4727 8791
rect 4761 8757 4773 8791
tri 4773 8766 4810 8803 sw
rect 834 8745 4773 8757
rect 788 8711 992 8745
tri 992 8711 1026 8745 nw
tri 4697 8711 4731 8745 ne
rect 788 8707 945 8711
rect 788 8673 800 8707
rect 834 8673 945 8707
rect 788 8664 945 8673
tri 945 8664 992 8711 nw
rect 8575 8695 8603 8723
rect 788 8635 911 8664
rect 788 8601 800 8635
rect 834 8630 911 8635
tri 911 8630 945 8664 nw
tri 4833 8630 4867 8664 nw
tri 6246 8630 6280 8664 ne
rect 6280 8630 6405 8664
rect 834 8601 876 8630
rect 788 8595 876 8601
tri 876 8595 911 8630 nw
tri 6280 8595 6315 8630 ne
rect 6315 8595 6405 8630
rect 788 8586 867 8595
tri 867 8586 876 8595 nw
rect 1158 8589 1224 8595
rect 788 8563 846 8586
tri 846 8565 867 8586 nw
rect 788 8529 800 8563
rect 834 8529 846 8563
rect 788 8491 846 8529
rect 788 8457 800 8491
rect 834 8457 846 8491
rect 788 8419 846 8457
rect 788 8385 800 8419
rect 834 8385 846 8419
rect 788 8347 846 8385
rect 788 8313 800 8347
rect 834 8313 846 8347
rect 788 8275 846 8313
rect 788 8241 800 8275
rect 834 8241 846 8275
tri 584 8227 589 8232 ne
rect 589 8227 618 8232
tri 589 8220 596 8227 ne
rect 596 8220 618 8227
tri 596 8208 608 8220 ne
rect 608 8208 618 8220
tri 608 8203 613 8208 ne
rect 613 8203 618 8208
tri 613 8198 618 8203 ne
rect 788 8203 846 8241
rect 788 8169 800 8203
rect 834 8169 846 8203
tri 497 8136 515 8154 ne
rect 515 8136 522 8154
tri 515 8131 520 8136 ne
rect 520 8131 522 8136
tri 520 8129 522 8131 ne
rect 788 8131 846 8169
rect 788 8097 800 8131
rect 834 8097 846 8131
tri 408 8073 415 8080 ne
rect 415 8073 433 8080
tri 415 8064 424 8073 ne
rect 424 8064 433 8073
tri 424 8059 429 8064 ne
rect 429 8059 433 8064
tri 429 8055 433 8059 ne
rect 788 8059 846 8097
rect -730 7981 -724 8033
rect -672 7981 -659 8033
rect -607 7981 -594 8033
rect -542 7981 -529 8033
rect -477 7981 -464 8033
rect -412 7981 -399 8033
rect -347 7981 -334 8033
rect -282 7981 -276 8033
rect -730 7961 -276 7981
rect -730 7909 -724 7961
rect -672 7909 -659 7961
rect -607 7909 -594 7961
rect -542 7909 -529 7961
rect -477 7909 -464 7961
rect -412 7909 -399 7961
rect -347 7909 -334 7961
rect -282 7909 -276 7961
rect -730 7889 -276 7909
rect -730 7837 -724 7889
rect -672 7837 -659 7889
rect -607 7837 -594 7889
rect -542 7837 -529 7889
rect -477 7837 -464 7889
rect -412 7837 -399 7889
rect -347 7837 -334 7889
rect -282 7837 -276 7889
rect -730 7817 -276 7837
rect -730 7765 -724 7817
rect -672 7765 -659 7817
rect -607 7765 -594 7817
rect -542 7765 -529 7817
rect -477 7765 -464 7817
rect -412 7765 -399 7817
rect -347 7765 -334 7817
rect -282 7765 -276 7817
rect -730 7745 -276 7765
rect -730 7693 -724 7745
rect -672 7693 -659 7745
rect -607 7693 -594 7745
rect -542 7693 -529 7745
rect -477 7693 -464 7745
rect -412 7693 -399 7745
rect -347 7693 -334 7745
rect -282 7693 -276 7745
rect 788 8025 800 8059
rect 834 8025 846 8059
rect 788 7987 846 8025
rect 788 7953 800 7987
rect 834 7953 846 7987
rect 788 7915 846 7953
rect 788 7881 800 7915
rect 834 7881 846 7915
rect 788 7843 846 7881
rect 788 7809 800 7843
rect 834 7809 846 7843
rect 788 7771 846 7809
rect 788 7737 800 7771
rect 834 7737 846 7771
rect 788 7699 846 7737
rect 788 7665 800 7699
rect 834 7665 846 7699
rect 788 7627 846 7665
rect 788 7593 800 7627
rect 834 7593 846 7627
rect 788 7555 846 7593
rect 788 7521 800 7555
rect 834 7521 846 7555
rect 788 7483 846 7521
tri 159 7449 170 7460 ne
rect 170 7449 193 7460
tri 170 7428 191 7449 ne
rect 191 7428 193 7449
tri 191 7426 193 7428 ne
rect 788 7449 800 7483
rect 834 7449 846 7483
rect 788 7411 846 7449
rect 788 7377 800 7411
rect 834 7377 846 7411
rect 788 7339 846 7377
rect -730 7335 -275 7336
rect -730 7283 -724 7335
rect -672 7283 -658 7335
rect -606 7283 -593 7335
rect -541 7283 -528 7335
rect -476 7283 -463 7335
rect -411 7283 -398 7335
rect -346 7283 -333 7335
rect -281 7283 -275 7335
rect -730 7255 -275 7283
rect -730 7203 -724 7255
rect -672 7203 -658 7255
rect -606 7203 -593 7255
rect -541 7203 -528 7255
rect -476 7203 -463 7255
rect -411 7203 -398 7255
rect -346 7203 -333 7255
rect -281 7203 -275 7255
rect -730 7175 -275 7203
rect -730 7123 -724 7175
rect -672 7123 -658 7175
rect -606 7123 -593 7175
rect -541 7123 -528 7175
rect -476 7123 -463 7175
rect -411 7123 -398 7175
rect -346 7123 -333 7175
rect -281 7123 -275 7175
rect -730 7122 -275 7123
rect 788 7305 800 7339
rect 834 7305 846 7339
rect 788 7267 846 7305
rect 788 7233 800 7267
rect 834 7233 846 7267
rect 788 7195 846 7233
rect 1210 8543 1224 8589
rect 1276 8586 1288 8595
rect 1340 8586 1352 8595
rect 1404 8586 1416 8595
rect 1468 8586 1480 8595
rect 1532 8586 1544 8595
rect 1596 8586 4514 8595
rect 1279 8552 1288 8586
rect 1351 8552 1352 8586
rect 1532 8552 1533 8586
rect 1596 8552 1605 8586
rect 1639 8552 1677 8586
rect 1711 8552 1749 8586
rect 1783 8552 1821 8586
rect 1855 8552 1893 8586
rect 1927 8552 1965 8586
rect 1999 8552 2037 8586
rect 2071 8552 2109 8586
rect 2143 8552 2181 8586
rect 2215 8552 2253 8586
rect 2287 8552 2325 8586
rect 2359 8552 2397 8586
rect 2431 8552 2469 8586
rect 2503 8552 2541 8586
rect 2575 8552 2613 8586
rect 2647 8552 2685 8586
rect 2719 8552 2757 8586
rect 2791 8552 2829 8586
rect 2863 8552 2901 8586
rect 2935 8552 2973 8586
rect 3007 8552 3045 8586
rect 3079 8552 3117 8586
rect 3151 8552 3189 8586
rect 3223 8552 3261 8586
rect 3295 8552 3333 8586
rect 3367 8552 3405 8586
rect 3439 8552 3477 8586
rect 3511 8552 3549 8586
rect 3583 8552 3621 8586
rect 3655 8552 3693 8586
rect 3727 8552 3765 8586
rect 3799 8552 3837 8586
rect 3871 8552 3909 8586
rect 3943 8552 3981 8586
rect 4015 8552 4053 8586
rect 4087 8552 4125 8586
rect 4159 8552 4197 8586
rect 4231 8552 4269 8586
rect 4303 8552 4341 8586
rect 4375 8580 4514 8586
rect 4375 8552 4474 8580
rect 1276 8543 1288 8552
rect 1340 8543 1352 8552
rect 1404 8543 1416 8552
rect 1468 8543 1480 8552
rect 1532 8543 1544 8552
rect 1596 8546 4474 8552
rect 4508 8546 4514 8580
rect 1596 8543 4514 8546
rect 1158 8525 1210 8537
tri 1210 8514 1239 8543 nw
tri 4437 8514 4466 8543 ne
rect 4466 8514 4514 8543
tri 4466 8512 4468 8514 ne
rect 4468 8508 4514 8514
rect 1158 8462 1167 8473
rect 1201 8462 1210 8473
rect 1158 8461 1210 8462
rect 1279 8472 2049 8483
rect 2101 8472 2113 8483
rect 2165 8472 2177 8483
rect 2229 8472 2241 8483
rect 2293 8472 2305 8483
rect 1279 8438 1294 8472
rect 1328 8438 1366 8472
rect 1400 8438 1438 8472
rect 1472 8438 1510 8472
rect 1544 8438 1582 8472
rect 1616 8438 1654 8472
rect 1688 8438 1726 8472
rect 1760 8438 1798 8472
rect 1832 8438 1870 8472
rect 1904 8438 1942 8472
rect 1976 8438 2014 8472
rect 2048 8438 2049 8472
rect 2229 8438 2230 8472
rect 2293 8438 2302 8472
rect 1279 8431 2049 8438
rect 2101 8431 2113 8438
rect 2165 8431 2177 8438
rect 2229 8431 2241 8438
rect 2293 8431 2305 8438
rect 2357 8431 2369 8483
rect 2421 8431 2433 8483
rect 2485 8431 2497 8483
rect 2549 8472 2561 8483
rect 2613 8472 2625 8483
rect 2677 8472 2689 8483
rect 2741 8472 2753 8483
rect 2805 8472 4220 8483
rect 2552 8438 2561 8472
rect 2624 8438 2625 8472
rect 2805 8438 2806 8472
rect 2840 8438 2878 8472
rect 2912 8438 2950 8472
rect 2984 8438 3022 8472
rect 3056 8438 3094 8472
rect 3128 8438 3166 8472
rect 3200 8438 3238 8472
rect 3272 8438 3310 8472
rect 3344 8438 3382 8472
rect 3416 8438 3454 8472
rect 3488 8438 3526 8472
rect 3560 8438 3598 8472
rect 3632 8438 3670 8472
rect 3704 8438 3742 8472
rect 3776 8438 3814 8472
rect 3848 8438 3886 8472
rect 3920 8438 3958 8472
rect 3992 8438 4030 8472
rect 4064 8438 4102 8472
rect 4136 8438 4174 8472
rect 4208 8438 4220 8472
rect 2549 8431 2561 8438
rect 2613 8431 2625 8438
rect 2677 8431 2689 8438
rect 2741 8431 2753 8438
rect 2805 8431 4220 8438
rect 4468 8474 4474 8508
rect 4508 8474 4514 8508
tri 6315 8505 6405 8595 ne
tri 6655 8505 6814 8664 nw
tri 8156 8656 8164 8664 ne
rect 8164 8656 8190 8664
tri 8164 8630 8190 8656 ne
rect 8607 8630 8615 8656
tri 8615 8630 8641 8656 nw
tri 13133 8630 13159 8656 ne
rect 13159 8630 13167 8656
tri 8607 8622 8615 8630 nw
tri 13159 8622 13167 8630 ne
rect 4468 8436 4514 8474
rect 1158 8397 1167 8409
rect 1201 8397 1210 8409
rect 1158 8333 1167 8345
rect 1201 8333 1210 8345
rect 4324 8415 4370 8427
rect 4324 8381 4330 8415
rect 4364 8381 4370 8415
rect 4324 8338 4370 8381
rect 1158 8280 1210 8281
rect 1158 8269 1167 8280
rect 1201 8269 1210 8280
rect 1281 8272 1288 8324
rect 1340 8272 1352 8324
rect 1404 8272 1416 8324
rect 1468 8316 1480 8324
rect 1532 8316 1544 8324
rect 1596 8316 4220 8324
rect 1472 8282 1480 8316
rect 1616 8282 1654 8316
rect 1688 8282 1726 8316
rect 1760 8282 1798 8316
rect 1832 8282 1870 8316
rect 1904 8282 1942 8316
rect 1976 8282 2014 8316
rect 2048 8282 2086 8316
rect 2120 8282 2158 8316
rect 2192 8282 2230 8316
rect 2264 8282 2302 8316
rect 2336 8282 2374 8316
rect 2408 8282 2446 8316
rect 2480 8282 2518 8316
rect 2552 8282 2590 8316
rect 2624 8282 2662 8316
rect 2696 8282 2734 8316
rect 2768 8282 2806 8316
rect 2840 8282 2878 8316
rect 2912 8282 2950 8316
rect 2984 8282 3022 8316
rect 3056 8282 3094 8316
rect 3128 8282 3166 8316
rect 3200 8282 3238 8316
rect 3272 8282 3310 8316
rect 3344 8282 3382 8316
rect 3416 8282 3454 8316
rect 3488 8282 3526 8316
rect 3560 8282 3598 8316
rect 3632 8282 3670 8316
rect 3704 8282 3742 8316
rect 3776 8282 3814 8316
rect 3848 8282 3886 8316
rect 3920 8282 3958 8316
rect 3992 8282 4030 8316
rect 4064 8282 4102 8316
rect 4136 8282 4174 8316
rect 4208 8282 4220 8316
rect 1468 8272 1480 8282
rect 1532 8272 1544 8282
rect 1596 8272 4220 8282
rect 4324 8304 4330 8338
rect 4364 8304 4370 8338
rect 1158 8208 1210 8217
rect 1158 8205 1167 8208
rect 1201 8205 1210 8208
tri 4321 8269 4324 8272 se
rect 4324 8269 4370 8304
rect 4468 8402 4474 8436
rect 4508 8402 4514 8436
rect 4468 8364 4514 8402
rect 4468 8330 4474 8364
rect 4508 8330 4514 8364
rect 4468 8292 4514 8330
tri 4370 8269 4373 8272 sw
rect 4321 8263 4373 8269
rect 4321 8199 4373 8211
rect 1158 8141 1210 8153
rect 1279 8160 2049 8169
rect 2101 8160 2113 8169
rect 2165 8160 2177 8169
rect 2229 8160 2241 8169
rect 2293 8160 2305 8169
rect 1279 8126 1294 8160
rect 1328 8126 1366 8160
rect 1400 8126 1438 8160
rect 1472 8126 1510 8160
rect 1544 8126 1582 8160
rect 1616 8126 1654 8160
rect 1688 8126 1726 8160
rect 1760 8126 1798 8160
rect 1832 8126 1870 8160
rect 1904 8126 1942 8160
rect 1976 8126 2014 8160
rect 2048 8126 2049 8160
rect 2229 8126 2230 8160
rect 2293 8126 2302 8160
rect 1279 8117 2049 8126
rect 2101 8117 2113 8126
rect 2165 8117 2177 8126
rect 2229 8117 2241 8126
rect 2293 8117 2305 8126
rect 2357 8117 2369 8169
rect 2421 8117 2433 8169
rect 2485 8117 2497 8169
rect 2549 8160 2561 8169
rect 2613 8160 2625 8169
rect 2677 8160 2689 8169
rect 2741 8160 2753 8169
rect 2805 8160 4220 8169
rect 2552 8126 2561 8160
rect 2624 8126 2625 8160
rect 2805 8126 2806 8160
rect 2840 8126 2878 8160
rect 2912 8126 2950 8160
rect 2984 8126 3022 8160
rect 3056 8126 3094 8160
rect 3128 8126 3166 8160
rect 3200 8126 3238 8160
rect 3272 8126 3310 8160
rect 3344 8126 3382 8160
rect 3416 8126 3454 8160
rect 3488 8126 3526 8160
rect 3560 8126 3598 8160
rect 3632 8126 3670 8160
rect 3704 8126 3742 8160
rect 3776 8126 3814 8160
rect 3848 8126 3886 8160
rect 3920 8126 3958 8160
rect 3992 8126 4030 8160
rect 4064 8126 4102 8160
rect 4136 8126 4174 8160
rect 4208 8126 4220 8160
rect 4321 8141 4373 8147
tri 4321 8138 4324 8141 ne
rect 2549 8117 2561 8126
rect 2613 8117 2625 8126
rect 2677 8117 2689 8126
rect 2741 8117 2753 8126
rect 2805 8117 4220 8126
rect 1158 8077 1210 8089
rect 1158 8013 1210 8025
rect 4324 8107 4370 8141
tri 4370 8138 4373 8141 nw
rect 4468 8258 4474 8292
rect 4508 8258 4514 8292
rect 4468 8220 4514 8258
rect 4468 8186 4474 8220
rect 4508 8186 4514 8220
rect 14143 8367 14195 8373
rect 14143 8300 14195 8315
rect 14143 8233 14195 8248
rect 4468 8148 4514 8186
rect 4324 8073 4330 8107
rect 4364 8073 4370 8107
rect 4324 8030 4370 8073
rect 1281 7964 1288 8016
rect 1340 7964 1352 8016
rect 1404 7964 1416 8016
rect 1468 8004 1480 8016
rect 1532 8004 1544 8016
rect 1596 8004 4220 8016
rect 1472 7970 1480 8004
rect 1616 7970 1654 8004
rect 1688 7970 1726 8004
rect 1760 7970 1798 8004
rect 1832 7970 1870 8004
rect 1904 7970 1942 8004
rect 1976 7970 2014 8004
rect 2048 7970 2086 8004
rect 2120 7970 2158 8004
rect 2192 7970 2230 8004
rect 2264 7970 2302 8004
rect 2336 7970 2374 8004
rect 2408 7970 2446 8004
rect 2480 7970 2518 8004
rect 2552 7970 2590 8004
rect 2624 7970 2662 8004
rect 2696 7970 2734 8004
rect 2768 7970 2806 8004
rect 2840 7970 2878 8004
rect 2912 7970 2950 8004
rect 2984 7970 3022 8004
rect 3056 7970 3094 8004
rect 3128 7970 3166 8004
rect 3200 7970 3238 8004
rect 3272 7970 3310 8004
rect 3344 7970 3382 8004
rect 3416 7970 3454 8004
rect 3488 7970 3526 8004
rect 3560 7970 3598 8004
rect 3632 7970 3670 8004
rect 3704 7970 3742 8004
rect 3776 7970 3814 8004
rect 3848 7970 3886 8004
rect 3920 7970 3958 8004
rect 3992 7970 4030 8004
rect 4064 7970 4102 8004
rect 4136 7970 4174 8004
rect 4208 7970 4220 8004
rect 1468 7964 1480 7970
rect 1532 7964 1544 7970
rect 1596 7964 4220 7970
rect 4324 7996 4330 8030
rect 4364 7996 4370 8030
rect 1158 7958 1167 7961
rect 1201 7958 1210 7961
rect 1158 7949 1210 7958
rect 1158 7886 1167 7897
rect 1201 7886 1210 7897
rect 1158 7885 1210 7886
rect 4324 7953 4370 7996
rect 4324 7919 4330 7953
rect 4364 7919 4370 7953
rect 4324 7876 4370 7919
rect 1158 7821 1167 7833
rect 1201 7821 1210 7833
rect 1279 7848 2069 7857
rect 1279 7814 1294 7848
rect 1328 7814 1366 7848
rect 1400 7814 1438 7848
rect 1472 7814 1510 7848
rect 1544 7814 1582 7848
rect 1616 7814 1654 7848
rect 1688 7814 1726 7848
rect 1760 7814 1798 7848
rect 1832 7814 1870 7848
rect 1904 7814 1942 7848
rect 1976 7814 2014 7848
rect 2048 7814 2069 7848
rect 1279 7805 2069 7814
rect 2121 7805 2133 7857
rect 2185 7848 2197 7857
rect 2249 7848 2261 7857
rect 2313 7848 2325 7857
rect 2377 7848 2389 7857
rect 2441 7848 2453 7857
rect 2192 7814 2197 7848
rect 2441 7814 2446 7848
rect 2185 7805 2197 7814
rect 2249 7805 2261 7814
rect 2313 7805 2325 7814
rect 2377 7805 2389 7814
rect 2441 7805 2453 7814
rect 2505 7805 2517 7857
rect 2569 7805 2581 7857
rect 2633 7805 2645 7857
rect 2697 7805 2709 7857
rect 2761 7848 2773 7857
rect 2825 7848 2837 7857
rect 2889 7848 4220 7857
rect 2768 7814 2773 7848
rect 2912 7814 2950 7848
rect 2984 7814 3022 7848
rect 3056 7814 3094 7848
rect 3128 7814 3166 7848
rect 3200 7814 3238 7848
rect 3272 7814 3310 7848
rect 3344 7814 3382 7848
rect 3416 7814 3454 7848
rect 3488 7814 3526 7848
rect 3560 7814 3598 7848
rect 3632 7814 3670 7848
rect 3704 7814 3742 7848
rect 3776 7814 3814 7848
rect 3848 7814 3886 7848
rect 3920 7814 3958 7848
rect 3992 7814 4030 7848
rect 4064 7814 4102 7848
rect 4136 7814 4174 7848
rect 4208 7814 4220 7848
rect 2761 7805 2773 7814
rect 2825 7805 2837 7814
rect 2889 7805 4220 7814
rect 4324 7842 4330 7876
rect 4364 7842 4370 7876
rect 1158 7757 1167 7769
rect 1201 7757 1210 7769
rect 1158 7704 1210 7705
rect 1158 7693 1167 7704
rect 1201 7693 1210 7704
rect 4324 7799 4370 7842
rect 4324 7765 4330 7799
rect 4364 7765 4370 7799
rect 4324 7721 4370 7765
rect 1278 7649 1288 7701
rect 1340 7649 1352 7701
rect 1404 7649 1416 7701
rect 1468 7692 1480 7701
rect 1532 7692 1544 7701
rect 1596 7692 4220 7701
rect 1472 7658 1480 7692
rect 1616 7658 1654 7692
rect 1688 7658 1726 7692
rect 1760 7658 1798 7692
rect 1832 7658 1870 7692
rect 1904 7658 1942 7692
rect 1976 7658 2014 7692
rect 2048 7658 2086 7692
rect 2120 7658 2158 7692
rect 2192 7658 2230 7692
rect 2264 7658 2302 7692
rect 2336 7658 2374 7692
rect 2408 7658 2446 7692
rect 2480 7658 2518 7692
rect 2552 7658 2590 7692
rect 2624 7658 2662 7692
rect 2696 7658 2734 7692
rect 2768 7658 2806 7692
rect 2840 7658 2878 7692
rect 2912 7658 2950 7692
rect 2984 7658 3022 7692
rect 3056 7658 3094 7692
rect 3128 7658 3166 7692
rect 3200 7658 3238 7692
rect 3272 7658 3310 7692
rect 3344 7658 3382 7692
rect 3416 7658 3454 7692
rect 3488 7658 3526 7692
rect 3560 7658 3598 7692
rect 3632 7658 3670 7692
rect 3704 7658 3742 7692
rect 3776 7658 3814 7692
rect 3848 7658 3886 7692
rect 3920 7658 3958 7692
rect 3992 7658 4030 7692
rect 4064 7658 4102 7692
rect 4136 7658 4174 7692
rect 4208 7658 4220 7692
rect 1468 7649 1480 7658
rect 1532 7649 1544 7658
rect 1596 7649 4220 7658
rect 4324 7687 4330 7721
rect 4364 7687 4370 7721
rect 1158 7632 1210 7641
rect 1158 7629 1167 7632
rect 1201 7629 1210 7632
rect 1158 7565 1210 7577
rect 4324 7643 4370 7687
rect 4324 7609 4330 7643
rect 4364 7609 4370 7643
rect 4324 7565 4370 7609
rect 1158 7501 1210 7513
rect 1279 7536 2069 7545
rect 1279 7502 1294 7536
rect 1328 7502 1366 7536
rect 1400 7502 1438 7536
rect 1472 7502 1510 7536
rect 1544 7502 1582 7536
rect 1616 7502 1654 7536
rect 1688 7502 1726 7536
rect 1760 7502 1798 7536
rect 1832 7502 1870 7536
rect 1904 7502 1942 7536
rect 1976 7502 2014 7536
rect 2048 7502 2069 7536
rect 1279 7493 2069 7502
rect 2121 7493 2133 7545
rect 2185 7536 2197 7545
rect 2249 7536 2261 7545
rect 2313 7536 2325 7545
rect 2377 7536 2389 7545
rect 2441 7536 2453 7545
rect 2192 7502 2197 7536
rect 2441 7502 2446 7536
rect 2185 7493 2197 7502
rect 2249 7493 2261 7502
rect 2313 7493 2325 7502
rect 2377 7493 2389 7502
rect 2441 7493 2453 7502
rect 2505 7493 2517 7545
rect 2569 7493 2581 7545
rect 2633 7493 2645 7545
rect 2697 7493 2709 7545
rect 2761 7536 2773 7545
rect 2825 7536 2837 7545
rect 2889 7536 4220 7545
rect 2768 7502 2773 7536
rect 2912 7502 2950 7536
rect 2984 7502 3022 7536
rect 3056 7502 3094 7536
rect 3128 7502 3166 7536
rect 3200 7502 3238 7536
rect 3272 7502 3310 7536
rect 3344 7502 3382 7536
rect 3416 7502 3454 7536
rect 3488 7502 3526 7536
rect 3560 7502 3598 7536
rect 3632 7502 3670 7536
rect 3704 7502 3742 7536
rect 3776 7502 3814 7536
rect 3848 7502 3886 7536
rect 3920 7502 3958 7536
rect 3992 7502 4030 7536
rect 4064 7502 4102 7536
rect 4136 7502 4174 7536
rect 4208 7502 4220 7536
rect 2761 7493 2773 7502
rect 2825 7493 2837 7502
rect 2889 7493 4220 7502
rect 4324 7531 4330 7565
rect 4364 7531 4370 7565
rect 4324 7487 4370 7531
tri 1210 7453 1220 7463 sw
rect 4324 7453 4330 7487
rect 4364 7453 4370 7487
rect 1210 7449 1220 7453
rect 1158 7437 1220 7449
rect 1210 7428 1220 7437
tri 1220 7428 1245 7453 sw
rect 4324 7441 4370 7453
rect 4468 8114 4474 8148
rect 4508 8114 4514 8148
rect 4468 8076 4514 8114
rect 4468 8042 4474 8076
rect 4508 8042 4514 8076
rect 4468 8004 4514 8042
rect 4468 7970 4474 8004
rect 4508 7970 4514 8004
rect 4468 7932 4514 7970
rect 4468 7898 4474 7932
rect 4508 7898 4514 7932
rect 4468 7860 4514 7898
rect 4468 7826 4474 7860
rect 4508 7826 4514 7860
rect 4468 7788 4514 7826
rect 4468 7754 4474 7788
rect 4508 7754 4514 7788
rect 4468 7716 4514 7754
rect 4930 8186 5032 8192
rect 4930 8134 4955 8186
rect 5007 8134 5032 8186
rect 4930 8110 5032 8134
rect 4930 8058 4955 8110
rect 5007 8058 5032 8110
rect 4930 8034 5032 8058
rect 4930 7982 4955 8034
rect 5007 7982 5032 8034
rect 4930 7958 5032 7982
rect 4930 7906 4955 7958
rect 5007 7906 5032 7958
rect 4930 7882 5032 7906
rect 4930 7830 4955 7882
rect 5007 7830 5032 7882
rect 4930 7806 5032 7830
rect 4930 7754 4955 7806
rect 5007 7754 5032 7806
rect 14143 8166 14195 8181
rect 14143 8099 14195 8114
rect 14143 8032 14195 8047
rect 14143 7965 14195 7980
rect 14143 7897 14195 7913
rect 14143 7829 14195 7845
rect 14143 7771 14195 7777
rect 4930 7748 5032 7754
rect 4468 7682 4474 7716
rect 4508 7682 4514 7716
rect 4468 7644 4514 7682
rect 4468 7610 4474 7644
rect 4508 7610 4514 7644
rect 4468 7572 4514 7610
rect 4468 7538 4474 7572
rect 4508 7538 4514 7572
rect 4468 7500 4514 7538
rect 4468 7466 4474 7500
rect 4508 7466 4514 7500
rect 4468 7428 4514 7466
rect 1210 7394 1245 7428
tri 1245 7394 1279 7428 sw
rect 4468 7394 4474 7428
rect 4508 7394 4514 7428
rect 1210 7389 1279 7394
tri 1279 7389 1284 7394 sw
rect 1210 7385 1288 7389
rect 1158 7382 1167 7385
rect 1201 7382 1288 7385
rect 1158 7373 1288 7382
rect 1210 7337 1288 7373
rect 1340 7337 1352 7389
rect 1404 7337 1416 7389
rect 1468 7380 1480 7389
rect 1532 7380 1544 7389
rect 1596 7380 4220 7389
rect 1472 7346 1480 7380
rect 1616 7346 1654 7380
rect 1688 7346 1726 7380
rect 1760 7346 1798 7380
rect 1832 7346 1870 7380
rect 1904 7346 1942 7380
rect 1976 7346 2014 7380
rect 2048 7346 2086 7380
rect 2120 7346 2158 7380
rect 2192 7346 2230 7380
rect 2264 7346 2302 7380
rect 2336 7346 2374 7380
rect 2408 7346 2446 7380
rect 2480 7346 2518 7380
rect 2552 7346 2590 7380
rect 2624 7346 2662 7380
rect 2696 7346 2734 7380
rect 2768 7346 2806 7380
rect 2840 7346 2878 7380
rect 2912 7346 2950 7380
rect 2984 7346 3022 7380
rect 3056 7346 3094 7380
rect 3128 7346 3166 7380
rect 3200 7346 3238 7380
rect 3272 7346 3310 7380
rect 3344 7346 3382 7380
rect 3416 7346 3454 7380
rect 3488 7346 3526 7380
rect 3560 7346 3598 7380
rect 3632 7346 3670 7380
rect 3704 7346 3742 7380
rect 3776 7346 3814 7380
rect 3848 7346 3886 7380
rect 3920 7346 3958 7380
rect 3992 7346 4030 7380
rect 4064 7346 4102 7380
rect 4136 7346 4174 7380
rect 4208 7346 4220 7380
rect 1468 7337 1480 7346
rect 1532 7337 1544 7346
rect 1596 7337 4220 7346
tri 4220 7337 4272 7389 sw
rect 1210 7321 4272 7337
tri 4272 7321 4288 7337 sw
rect 1158 7310 1167 7321
rect 1201 7310 1284 7321
rect 1158 7272 1284 7310
rect 1158 7238 1167 7272
rect 1201 7269 1284 7272
rect 1336 7269 1349 7321
rect 1401 7269 1414 7321
rect 1466 7269 1479 7321
rect 1531 7269 1544 7321
rect 1596 7309 4288 7321
tri 4288 7309 4300 7321 sw
rect 1596 7275 4300 7309
tri 4300 7275 4334 7309 sw
tri 4434 7275 4468 7309 se
rect 4468 7275 4514 7394
rect 13764 7374 14044 7465
rect 1596 7269 4514 7275
rect 1201 7266 4514 7269
rect 1201 7238 1300 7266
rect 1158 7232 1300 7238
rect 1334 7232 1372 7266
rect 1406 7232 1444 7266
rect 1478 7232 1516 7266
rect 1550 7232 1588 7266
rect 1622 7232 1660 7266
rect 1694 7232 1732 7266
rect 1766 7232 1804 7266
rect 1838 7232 1876 7266
rect 1910 7232 1948 7266
rect 1982 7232 2020 7266
rect 2054 7232 2092 7266
rect 2126 7232 2164 7266
rect 2198 7232 2236 7266
rect 2270 7232 2308 7266
rect 2342 7232 2380 7266
rect 2414 7232 2452 7266
rect 2486 7232 2524 7266
rect 2558 7232 2596 7266
rect 2630 7232 2668 7266
rect 2702 7232 2740 7266
rect 2774 7232 2812 7266
rect 2846 7232 2884 7266
rect 2918 7232 2956 7266
rect 2990 7232 3028 7266
rect 3062 7232 3100 7266
rect 3134 7232 3172 7266
rect 3206 7232 3244 7266
rect 3278 7232 3316 7266
rect 3350 7232 3388 7266
rect 3422 7232 3460 7266
rect 3494 7232 3532 7266
rect 3566 7232 3604 7266
rect 3638 7232 3676 7266
rect 3710 7232 3748 7266
rect 3782 7232 3820 7266
rect 3854 7232 3892 7266
rect 3926 7232 3964 7266
rect 3998 7232 4036 7266
rect 4070 7232 4108 7266
rect 4142 7232 4180 7266
rect 4214 7232 4252 7266
rect 4286 7232 4324 7266
rect 4358 7232 4396 7266
rect 4430 7232 4468 7266
rect 4502 7232 4514 7266
rect 1158 7223 4514 7232
rect 13392 7322 13398 7374
rect 13450 7322 13472 7374
rect 13524 7322 13545 7374
rect 13597 7322 13618 7374
rect 13670 7322 13691 7374
rect 13743 7322 13764 7374
rect 13816 7322 14044 7374
rect 13392 7302 14044 7322
rect 13392 7250 13398 7302
rect 13450 7250 13472 7302
rect 13524 7250 13545 7302
rect 13597 7250 13618 7302
rect 13670 7250 13691 7302
rect 13743 7250 13764 7302
rect 13816 7250 14044 7302
rect 13392 7230 14044 7250
rect 788 7161 800 7195
rect 834 7161 846 7195
rect 13392 7178 13398 7230
rect 13450 7178 13472 7230
rect 13524 7178 13545 7230
rect 13597 7178 13618 7230
rect 13670 7178 13691 7230
rect 13743 7178 13764 7230
rect 13816 7178 14044 7230
rect 788 7124 846 7161
tri 846 7124 886 7164 sw
rect 13392 7158 14044 7178
rect 788 7090 886 7124
tri 886 7090 920 7124 sw
tri 4697 7090 4731 7124 se
rect 788 7078 4731 7090
rect 788 7044 829 7078
rect 863 7044 901 7078
rect 935 7044 973 7078
rect 1007 7044 1045 7078
rect 1079 7044 1117 7078
rect 1151 7044 1189 7078
rect 1223 7044 1261 7078
rect 1295 7044 1333 7078
rect 1367 7044 1405 7078
rect 1439 7044 1477 7078
rect 1511 7044 1549 7078
rect 1583 7044 1621 7078
rect 1655 7044 1693 7078
rect 1727 7044 1765 7078
rect 1799 7044 1837 7078
rect 1871 7044 1909 7078
rect 1943 7044 1981 7078
rect 2015 7044 2053 7078
rect 2087 7044 2125 7078
rect 2159 7044 2197 7078
rect 2231 7044 2269 7078
rect 2303 7044 2341 7078
rect 2375 7044 2413 7078
rect 2447 7044 2485 7078
rect 2519 7044 2557 7078
rect 2591 7044 2629 7078
rect 2663 7044 2701 7078
rect 2735 7044 2773 7078
rect 2807 7044 2845 7078
rect 2879 7044 2917 7078
rect 2951 7044 2989 7078
rect 3023 7044 3061 7078
rect 3095 7044 3133 7078
rect 3167 7044 3205 7078
rect 3239 7044 3277 7078
rect 3311 7044 3349 7078
rect 3383 7044 3421 7078
rect 3455 7044 3493 7078
rect 3527 7044 3565 7078
rect 3599 7044 3637 7078
rect 3671 7044 3709 7078
rect 3743 7044 3781 7078
rect 3815 7044 3853 7078
rect 3887 7044 3925 7078
rect 3959 7044 3997 7078
rect 4031 7044 4069 7078
rect 4103 7044 4141 7078
rect 4175 7044 4213 7078
rect 4247 7044 4285 7078
rect 4319 7044 4357 7078
rect 4391 7044 4429 7078
rect 4463 7044 4501 7078
rect 4535 7044 4573 7078
rect 4607 7044 4645 7078
rect 4679 7044 4731 7078
rect 13392 7106 13398 7158
rect 13450 7106 13472 7158
rect 13524 7106 13545 7158
rect 13597 7106 13618 7158
rect 13670 7106 13691 7158
rect 13743 7106 13764 7158
rect 13816 7106 14044 7158
rect 13392 7086 14044 7106
tri 756 7006 788 7038 se
rect 788 7032 4737 7044
rect 788 7006 1091 7032
tri 1091 7006 1117 7032 nw
tri 4273 7012 4293 7032 ne
rect 4293 7012 4737 7032
tri 4293 7006 4299 7012 ne
rect 4299 7006 4737 7012
tri 722 6972 756 7006 se
rect 756 6972 1057 7006
tri 1057 6972 1091 7006 nw
tri 4299 6992 4313 7006 ne
rect 4313 6992 4424 7006
tri 687 6937 722 6972 se
rect 722 6937 1022 6972
tri 1022 6937 1057 6972 nw
rect 2059 6940 2065 6992
rect 2117 6940 2129 6992
rect 2181 6972 3802 6992
tri 3802 6972 3822 6992 sw
tri 4313 6972 4333 6992 ne
rect 4333 6972 4424 6992
rect 4458 6972 4507 7006
rect 4541 6972 4590 7006
rect 4624 6972 4672 7006
rect 4706 6972 4737 7006
rect 2181 6940 3822 6972
tri 3822 6940 3854 6972 sw
tri 4333 6940 4365 6972 ne
rect 4365 6940 4737 6972
rect 13392 7034 13398 7086
rect 13450 7034 13472 7086
rect 13524 7034 13545 7086
rect 13597 7034 13618 7086
rect 13670 7034 13691 7086
rect 13743 7034 13764 7086
rect 13816 7034 14044 7086
rect 13392 7014 14044 7034
rect 13392 6962 13398 7014
rect 13450 6962 13472 7014
rect 13524 6962 13545 7014
rect 13597 6962 13618 7014
rect 13670 6962 13691 7014
rect 13743 6962 13764 7014
rect 13816 6962 14044 7014
tri 3780 6937 3783 6940 ne
rect 3783 6937 3854 6940
tri 3854 6937 3857 6940 sw
tri 4365 6937 4368 6940 ne
rect 4368 6937 4737 6940
tri 144 6934 147 6937 se
rect 147 6934 1019 6937
tri 1019 6934 1022 6937 nw
tri 3783 6934 3786 6937 ne
rect 3786 6934 3857 6937
tri 3857 6934 3860 6937 sw
tri 4368 6934 4371 6937 ne
rect 4371 6934 4737 6937
tri 110 6900 144 6934 se
rect 144 6900 985 6934
tri 985 6900 1019 6934 nw
tri 3786 6930 3790 6934 ne
rect 3790 6930 3860 6934
tri 3860 6930 3864 6934 sw
tri 3790 6918 3802 6930 ne
rect 3802 6918 3864 6930
tri 3802 6908 3812 6918 ne
tri 83 6873 110 6900 se
rect 110 6891 976 6900
tri 976 6891 985 6900 nw
rect 110 6873 149 6891
tri 149 6873 167 6891 nw
rect 83 6861 137 6873
tri 137 6861 149 6873 nw
tri 79 6827 83 6831 se
rect 83 6827 129 6861
tri 129 6853 137 6861 nw
tri 49 6797 79 6827 se
rect 79 6797 129 6827
rect -126 6791 129 6797
rect -74 6739 129 6791
rect -126 6727 129 6739
rect -855 6721 -803 6727
rect -74 6713 129 6727
rect 193 6840 245 6846
tri 245 6827 258 6840 sw
rect 245 6821 258 6827
tri 258 6821 264 6827 sw
rect 245 6806 264 6821
tri 264 6806 279 6821 sw
rect 245 6788 3605 6806
rect 193 6776 3605 6788
rect 245 6754 3605 6776
rect 3657 6754 3669 6806
rect 3721 6754 3727 6806
rect 245 6735 260 6754
tri 260 6735 279 6754 nw
rect 245 6729 254 6735
tri 254 6729 260 6735 nw
rect 193 6718 245 6724
tri 245 6720 254 6729 nw
tri 3469 6720 3475 6726 se
rect 3475 6720 3639 6726
tri 3468 6719 3469 6720 se
rect 3469 6719 3639 6720
tri 295 6718 296 6719 se
rect 296 6718 870 6719
tri 294 6717 295 6718 se
rect 295 6717 870 6718
tri 129 6713 133 6717 sw
tri 290 6713 294 6717 se
rect 294 6716 870 6717
tri 870 6716 873 6719 sw
tri 3465 6716 3468 6719 se
rect 3468 6716 3639 6719
rect 294 6713 2180 6716
rect -74 6679 133 6713
tri 133 6679 167 6713 sw
tri 256 6679 290 6713 se
rect 290 6679 308 6713
rect 342 6679 382 6713
rect 416 6679 456 6713
rect 490 6679 530 6713
rect 564 6679 604 6713
rect 638 6679 678 6713
rect 712 6679 751 6713
rect 785 6679 824 6713
rect 858 6700 2180 6713
rect 858 6679 1837 6700
rect -74 6675 167 6679
rect -126 6669 167 6675
tri 167 6669 177 6679 sw
tri 246 6669 256 6679 se
rect 256 6669 1837 6679
rect -855 6657 -803 6669
rect -855 6601 -849 6605
rect -815 6601 -803 6605
rect -855 6599 -803 6601
rect -855 6594 -808 6599
tri -808 6594 -803 6599 nw
tri 83 6594 158 6669 ne
rect 158 6663 177 6669
tri 177 6663 183 6669 sw
tri 240 6663 246 6669 se
rect 246 6663 1837 6669
rect 158 6648 1837 6663
rect 1889 6648 1905 6700
rect 1957 6648 1973 6700
rect 2025 6648 2040 6700
rect 2092 6648 2107 6700
rect 2159 6648 2180 6700
tri 3401 6652 3465 6716 se
rect 3465 6674 3639 6716
rect 3691 6674 3703 6726
rect 3755 6674 3761 6726
rect 3465 6652 3475 6674
tri 3475 6652 3497 6674 nw
rect 158 6630 2180 6648
tri 3379 6630 3401 6652 se
rect 3401 6630 3453 6652
tri 3453 6630 3475 6652 nw
rect 158 6594 937 6630
tri 937 6594 973 6630 nw
tri 3378 6629 3379 6630 se
rect 3379 6629 3452 6630
tri 3452 6629 3453 6630 nw
tri 3365 6616 3378 6629 se
rect 3378 6616 3439 6629
tri 3439 6616 3452 6629 nw
rect -855 6555 -809 6594
tri -809 6593 -808 6594 nw
tri 158 6593 159 6594 ne
rect 159 6593 925 6594
tri 159 6589 163 6593 ne
rect 163 6589 925 6593
tri 163 6575 177 6589 ne
rect 177 6575 308 6589
tri 177 6555 197 6575 ne
rect 197 6555 308 6575
rect 342 6555 382 6589
rect 416 6555 456 6589
rect 490 6555 530 6589
rect 564 6555 604 6589
rect 638 6555 678 6589
rect 712 6555 751 6589
rect 785 6555 824 6589
rect 858 6582 925 6589
tri 925 6582 937 6594 nw
rect 1007 6582 2280 6588
rect 858 6555 891 6582
rect -855 6521 -849 6555
rect -815 6521 -809 6555
tri 197 6548 204 6555 ne
rect 204 6548 891 6555
tri 891 6548 925 6582 nw
rect 1007 6548 1019 6582
rect 1053 6548 1135 6582
rect 1169 6548 2280 6582
tri 204 6547 205 6548 ne
rect 205 6547 890 6548
tri 890 6547 891 6548 nw
rect -855 6475 -809 6521
rect -855 6441 -849 6475
rect -815 6441 -809 6475
rect 1007 6536 2280 6548
rect 2332 6536 2344 6588
rect 2396 6536 2408 6588
rect 2460 6536 2466 6588
rect 1007 6510 2466 6536
rect 1007 6498 2280 6510
rect 1007 6464 1019 6498
rect 1053 6464 1135 6498
rect 1169 6464 2280 6498
rect 1007 6458 2280 6464
rect 2332 6458 2344 6510
rect 2396 6458 2408 6510
rect 2460 6458 2466 6510
rect 2539 6551 3324 6554
rect 2539 6546 2978 6551
rect 3030 6546 3050 6551
rect 3102 6546 3122 6551
rect 3174 6546 3194 6551
rect 3246 6546 3266 6551
rect 2539 6512 2551 6546
rect 2585 6512 2627 6546
rect 2661 6512 2703 6546
rect 2737 6512 2779 6546
rect 2813 6512 2854 6546
rect 2888 6512 2929 6546
rect 2963 6512 2978 6546
rect 3038 6512 3050 6546
rect 3113 6512 3122 6546
rect 3188 6512 3194 6546
rect 3263 6512 3266 6546
rect 2539 6499 2978 6512
rect 3030 6499 3050 6512
rect 3102 6499 3122 6512
rect 3174 6499 3194 6512
rect 3246 6499 3266 6512
rect 3318 6499 3324 6551
rect 2539 6479 3324 6499
rect 2539 6472 2978 6479
rect 3030 6472 3050 6479
rect 3102 6472 3122 6479
rect 3174 6472 3194 6479
rect 3246 6472 3266 6479
rect -855 6395 -809 6441
rect -855 6361 -849 6395
rect -815 6361 -809 6395
rect 2539 6438 2551 6472
rect 2585 6438 2627 6472
rect 2661 6438 2703 6472
rect 2737 6438 2779 6472
rect 2813 6438 2854 6472
rect 2888 6438 2929 6472
rect 2963 6438 2978 6472
rect 3038 6438 3050 6472
rect 3113 6438 3122 6472
rect 3188 6438 3194 6472
rect 3263 6438 3266 6472
rect 2539 6427 2978 6438
rect 3030 6427 3050 6438
rect 3102 6427 3122 6438
rect 3174 6427 3194 6438
rect 3246 6427 3266 6438
rect 3318 6427 3324 6479
rect 2539 6407 3324 6427
rect 2539 6398 2978 6407
rect 3030 6398 3050 6407
rect 3102 6398 3122 6407
rect 3174 6398 3194 6407
rect 3246 6398 3266 6407
rect -855 6315 -809 6361
rect -855 6281 -849 6315
rect -815 6281 -809 6315
rect -855 6234 -809 6281
rect 1007 6379 1336 6385
rect 1007 6345 1019 6379
rect 1053 6345 1135 6379
rect 1169 6364 1336 6379
tri 1336 6364 1357 6385 sw
rect 2539 6364 2551 6398
rect 2585 6364 2627 6398
rect 2661 6364 2703 6398
rect 2737 6364 2779 6398
rect 2813 6364 2854 6398
rect 2888 6364 2929 6398
rect 2963 6364 2978 6398
rect 3038 6364 3050 6398
rect 3113 6364 3122 6398
rect 3188 6364 3194 6398
rect 3263 6364 3266 6398
rect 1169 6360 1357 6364
tri 1357 6360 1361 6364 sw
rect 1169 6345 2298 6360
rect 1007 6308 2298 6345
rect 2350 6308 2362 6360
rect 2414 6308 2426 6360
rect 2478 6308 2484 6360
rect 1007 6295 2484 6308
rect 1007 6261 1019 6295
rect 1053 6261 1135 6295
rect 1169 6282 2484 6295
rect 1169 6261 2298 6282
rect 1007 6255 2298 6261
tri 1282 6250 1287 6255 ne
rect 1287 6250 2298 6255
rect -855 6200 -849 6234
rect -815 6200 -809 6234
tri 1287 6230 1307 6250 ne
rect 1307 6230 2298 6250
rect 2350 6230 2362 6282
rect 2414 6230 2426 6282
rect 2478 6230 2484 6282
rect 2539 6355 2978 6364
rect 3030 6355 3050 6364
rect 3102 6355 3122 6364
rect 3174 6355 3194 6364
rect 3246 6355 3266 6364
rect 3318 6355 3324 6407
rect 2539 6335 3324 6355
rect 2539 6324 2978 6335
rect 3030 6324 3050 6335
rect 3102 6324 3122 6335
rect 3174 6324 3194 6335
rect 3246 6324 3266 6335
rect 2539 6290 2551 6324
rect 2585 6290 2627 6324
rect 2661 6290 2703 6324
rect 2737 6290 2779 6324
rect 2813 6290 2854 6324
rect 2888 6290 2929 6324
rect 2963 6290 2978 6324
rect 3038 6290 3050 6324
rect 3113 6290 3122 6324
rect 3188 6290 3194 6324
rect 3263 6290 3266 6324
rect 2539 6283 2978 6290
rect 3030 6283 3050 6290
rect 3102 6283 3122 6290
rect 3174 6283 3194 6290
rect 3246 6283 3266 6290
rect 3318 6283 3324 6335
rect 2539 6263 3324 6283
rect 2539 6250 2978 6263
rect 3030 6250 3050 6263
rect 3102 6250 3122 6263
rect 3174 6250 3194 6263
rect 3246 6250 3266 6263
rect 2539 6216 2551 6250
rect 2585 6216 2627 6250
rect 2661 6216 2703 6250
rect 2737 6216 2779 6250
rect 2813 6216 2854 6250
rect 2888 6216 2929 6250
rect 2963 6216 2978 6250
rect 3038 6216 3050 6250
rect 3113 6216 3122 6250
rect 3188 6216 3194 6250
rect 3263 6216 3266 6250
rect -855 6153 -809 6200
rect -855 6119 -849 6153
rect -815 6119 -809 6153
tri 756 6193 775 6212 sw
rect 2539 6211 2978 6216
rect 3030 6211 3050 6216
rect 3102 6211 3122 6216
rect 3174 6211 3194 6216
rect 3246 6211 3266 6216
rect 3318 6211 3324 6263
rect 2539 6208 3324 6211
rect 756 6190 775 6193
tri 775 6190 778 6193 sw
rect 756 6178 778 6190
tri 778 6178 790 6190 sw
tri 944 6178 956 6190 se
rect 956 6178 962 6190
rect 756 6150 962 6178
tri 944 6138 956 6150 ne
rect 956 6138 962 6150
rect 1014 6138 1026 6190
rect 1078 6138 1084 6190
rect -855 6107 -809 6119
tri 2771 5841 2805 5875 ne
rect 2805 5871 2857 5877
rect 2805 5807 2857 5819
rect 1994 5704 2000 5756
rect 2052 5704 2064 5756
rect 2116 5749 2160 5756
tri 2160 5749 2167 5756 sw
rect 2805 5749 2857 5755
rect 2116 5704 2167 5749
tri 2167 5704 2212 5749 sw
tri 2138 5669 2173 5704 ne
rect 2173 5669 2212 5704
tri 2212 5669 2247 5704 sw
rect 2473 5669 2479 5721
rect 2531 5669 2543 5721
rect 2595 5669 2601 5721
tri 2173 5635 2207 5669 ne
rect 2207 5635 2247 5669
tri 2247 5635 2281 5669 sw
tri 2515 5635 2549 5669 ne
tri 2207 5633 2209 5635 ne
rect 2209 5633 2281 5635
tri 1585 5601 1617 5633 ne
rect 1617 5601 1619 5633
tri 2209 5630 2212 5633 ne
rect 2212 5630 2281 5633
tri 2281 5630 2286 5635 sw
tri 2212 5601 2241 5630 ne
rect 2241 5601 2286 5630
tri 2286 5601 2315 5630 sw
tri 1617 5599 1619 5601 ne
tri 2241 5599 2243 5601 ne
rect 2243 5599 2315 5601
tri 2315 5599 2317 5601 sw
tri 2243 5583 2259 5599 ne
rect 2259 5583 2317 5599
tri 2317 5583 2333 5599 sw
tri 2259 5571 2271 5583 ne
rect 2271 5571 2333 5583
tri 1492 5549 1514 5571 ne
rect 1514 5549 1526 5571
tri 2271 5556 2286 5571 ne
rect 2286 5556 2333 5571
tri 2333 5556 2360 5583 sw
tri 2286 5549 2293 5556 ne
rect 2293 5549 2360 5556
tri 2360 5549 2367 5556 sw
tri 1514 5542 1521 5549 ne
rect 1521 5542 1526 5549
tri 2293 5542 2300 5549 ne
rect 2300 5542 2367 5549
tri 2367 5542 2374 5549 sw
tri 1521 5539 1524 5542 ne
rect 1524 5539 1526 5542
tri 2300 5539 2303 5542 ne
rect 2303 5539 2374 5542
tri 2374 5539 2377 5542 sw
tri 1524 5537 1526 5539 ne
tri 2303 5537 2305 5539 ne
rect 2305 5537 2377 5539
tri 2305 5534 2308 5537 ne
rect 2308 5534 2377 5537
tri 2377 5534 2382 5539 sw
tri 2308 5516 2326 5534 ne
rect 2326 5516 2382 5534
rect -768 5488 -740 5516
tri 2326 5515 2327 5516 ne
rect 2327 5515 2382 5516
rect 1365 5487 1393 5515
tri 2327 5503 2339 5515 ne
rect 2339 5503 2382 5515
tri 2382 5503 2413 5534 sw
tri 2339 5487 2355 5503 ne
rect 2355 5487 2413 5503
tri 2355 5482 2360 5487 ne
rect 2360 5482 2413 5487
tri 2413 5482 2434 5503 sw
tri 2360 5476 2366 5482 ne
rect 2366 5476 2434 5482
tri 2434 5476 2440 5482 sw
tri 2366 5472 2370 5476 ne
rect 2370 5472 2440 5476
tri 2440 5472 2444 5476 sw
tri 2370 5465 2377 5472 ne
rect 2377 5465 2444 5472
rect -228 5437 -200 5465
tri 2377 5438 2404 5465 ne
rect 2404 5438 2444 5465
tri 2444 5438 2478 5472 sw
tri 2404 5437 2405 5438 ne
rect 2405 5437 2478 5438
tri 2405 5415 2427 5437 ne
rect 2427 5415 2478 5437
tri 2478 5415 2501 5438 sw
tri 2427 5413 2429 5415 ne
rect 2429 5414 2501 5415
tri 2501 5414 2502 5415 sw
rect 2429 5413 2502 5414
tri 2429 5408 2434 5413 ne
rect 2434 5408 2502 5413
tri 2434 5403 2439 5408 ne
rect 2439 5403 2502 5408
tri -429 5377 -415 5391 se
rect 71 5385 79 5403
tri 79 5385 97 5403 nw
tri 2439 5392 2450 5403 ne
rect 71 5383 77 5385
tri 77 5383 79 5385 nw
rect 71 5381 75 5383
tri 75 5381 77 5383 nw
tri 71 5377 75 5381 nw
tri -449 5357 -429 5377 se
rect -429 5357 -415 5377
tri -369 5357 -351 5375 sw
tri -457 5301 -447 5311 ne
rect -447 5301 -423 5311
tri -447 5279 -425 5301 ne
rect -425 5279 -423 5301
rect -383 5305 -357 5311
tri -357 5305 -351 5311 nw
rect -383 5301 -361 5305
tri -361 5301 -357 5305 nw
rect -383 5298 -364 5301
tri -364 5298 -361 5301 nw
tri -383 5279 -364 5298 nw
tri -425 5277 -423 5279 ne
rect -590 5199 -586 5251
rect 434 5213 462 5241
tri 2432 5213 2450 5231 se
rect 2450 5213 2502 5403
tri 2430 5211 2432 5213 se
rect 2432 5211 2502 5213
tri 2427 5208 2430 5211 se
rect 2430 5209 2502 5211
rect 2430 5208 2493 5209
tri 844 5203 849 5208 nw
tri 2422 5203 2427 5208 se
rect 2427 5203 2493 5208
tri 2419 5200 2422 5203 se
rect 2422 5200 2493 5203
tri 2493 5200 2502 5209 nw
tri 2418 5199 2419 5200 se
rect 2419 5199 2489 5200
tri 2390 5171 2418 5199 se
rect 2418 5196 2489 5199
tri 2489 5196 2493 5200 nw
rect 2418 5171 2464 5196
tri 2464 5171 2489 5196 nw
tri 2527 5174 2549 5196 se
rect 2549 5174 2601 5669
rect 3085 5599 3137 5601
rect 3365 5549 3417 6616
tri 3417 6594 3439 6616 nw
rect 3712 6371 3764 6377
tri 3678 6332 3712 6366 se
rect 3448 6319 3712 6332
rect 3448 6307 3764 6319
rect 3448 6280 3712 6307
rect 3448 6249 3519 6280
tri 3519 6249 3550 6280 nw
tri 3681 6249 3712 6280 ne
rect 3712 6249 3764 6255
rect 3448 5737 3500 6249
tri 3500 6230 3519 6249 nw
rect 3448 5673 3500 5685
rect 3448 5615 3500 5621
rect 3721 6187 3773 6193
rect 3721 6123 3773 6135
tri 3417 5549 3451 5583 sw
tri 2935 5539 2938 5542 se
tri 2930 5534 2935 5539 se
rect 2935 5534 2938 5539
tri 2971 5534 2976 5539 sw
rect 3365 5497 3541 5549
rect 3593 5497 3605 5549
rect 3657 5497 3663 5549
tri 3289 5472 3293 5476 sw
tri 3717 5472 3721 5476 se
rect 3721 5472 3773 6071
rect 3812 5708 3864 6918
tri 4371 6900 4405 6934 ne
rect 4405 6900 4424 6934
rect 4458 6900 4507 6934
rect 4541 6900 4590 6934
rect 4624 6900 4672 6934
rect 4706 6900 4737 6934
tri 4405 6894 4411 6900 ne
rect 4411 6894 4737 6900
tri 4411 6891 4414 6894 ne
rect 4414 6891 4737 6894
rect 13764 6893 14044 6962
tri 4414 6873 4432 6891 ne
rect 4432 6873 4737 6891
tri 4432 6867 4438 6873 ne
rect 4438 6867 4737 6873
tri 4438 6861 4444 6867 ne
rect 4444 6861 4737 6867
tri 4444 6853 4452 6861 ne
rect 4452 6853 4502 6861
tri 4452 6827 4478 6853 ne
rect 4478 6827 4502 6853
rect 4536 6827 4576 6861
rect 4610 6827 4649 6861
rect 4683 6827 4737 6861
tri 11383 6831 11404 6852 se
tri 4478 6821 4484 6827 ne
rect 4484 6821 4737 6827
tri 4484 6775 4530 6821 ne
rect 4530 6775 4737 6821
tri 7913 6803 7941 6831 se
tri 11355 6803 11383 6831 se
rect 11383 6803 11404 6831
tri 7907 6797 7913 6803 se
rect 7913 6797 7941 6803
tri 8800 6797 8806 6803 sw
tri 11349 6797 11355 6803 se
rect 11355 6797 11404 6803
tri 4530 6769 4536 6775 ne
rect 4536 6769 4737 6775
rect 8800 6769 8806 6797
tri 8806 6769 8834 6797 sw
tri 11321 6769 11349 6797 se
rect 11349 6769 11404 6797
tri 4536 6735 4570 6769 ne
rect 4570 6735 4596 6769
rect 4630 6735 4668 6769
rect 4702 6735 4737 6769
tri 4570 6729 4576 6735 ne
rect 4576 6729 4737 6735
tri 4576 6719 4586 6729 ne
rect 4586 6719 4737 6729
tri 4586 6716 4589 6719 ne
rect 4589 6716 4737 6719
tri 4589 6630 4675 6716 ne
rect 4675 6630 4737 6716
tri 4675 6629 4676 6630 ne
rect 4676 6629 4737 6630
rect 4046 6602 4549 6629
tri 4549 6602 4576 6629 sw
tri 4676 6602 4703 6629 ne
rect 4703 6602 4737 6629
rect 4046 6594 4576 6602
rect 4046 6560 4058 6594
rect 4092 6560 4174 6594
rect 4208 6568 4576 6594
tri 4576 6568 4610 6602 sw
tri 4703 6568 4737 6602 ne
tri 4833 6568 4841 6576 sw
tri 8182 6568 8190 6576 se
rect 4208 6560 4610 6568
rect 4046 6547 4610 6560
tri 4610 6547 4631 6568 sw
rect 4833 6547 4841 6568
tri 4841 6547 4862 6568 sw
tri 8161 6547 8182 6568 se
rect 8182 6547 8190 6568
rect 4046 6542 4631 6547
tri 4631 6542 4636 6547 sw
rect 4833 6542 4862 6547
tri 4862 6542 4867 6547 sw
tri 8156 6542 8161 6547 se
rect 8161 6542 8190 6547
tri 8607 6568 8615 6576 sw
tri 11589 6568 11597 6576 se
rect 8607 6547 8615 6568
tri 8615 6547 8636 6568 sw
tri 11568 6547 11589 6568 se
rect 11589 6547 11597 6568
rect 8607 6542 8636 6547
tri 8636 6542 8641 6547 sw
tri 11563 6542 11568 6547 se
rect 11568 6542 11597 6547
tri 11699 6542 11733 6576 sw
rect 4046 6510 4636 6542
rect 4046 6476 4058 6510
rect 4092 6476 4174 6510
rect 4208 6476 4636 6510
rect 4046 6475 4636 6476
tri 4636 6475 4703 6542 sw
rect 4046 6455 4703 6475
tri 4493 6440 4508 6455 ne
rect 4508 6440 4703 6455
tri 4508 6406 4542 6440 ne
rect 4542 6406 4703 6440
tri 4833 6406 4867 6440 nw
tri 8156 6406 8190 6440 ne
tri 8607 6406 8641 6440 nw
tri 11563 6406 11597 6440 ne
tri 11699 6406 11733 6440 nw
tri 4542 6385 4563 6406 ne
rect 4563 6385 4703 6406
tri 4563 6377 4571 6385 ne
rect 3895 6197 3901 6249
rect 3953 6197 3965 6249
rect 4017 6197 4023 6249
rect 3895 6193 3977 6197
tri 3977 6193 3981 6197 nw
rect 3895 6179 3963 6193
tri 3963 6179 3977 6193 nw
rect 3895 6005 3947 6179
tri 3947 6163 3963 6179 nw
rect 4046 6167 4351 6179
tri 4351 6167 4363 6179 sw
rect 4046 6161 4363 6167
rect 4046 6127 4058 6161
rect 4092 6127 4174 6161
rect 4208 6127 4363 6161
rect 4046 6117 4363 6127
tri 4363 6117 4413 6167 sw
rect 4046 6077 4413 6117
rect 4046 6043 4058 6077
rect 4092 6043 4174 6077
rect 4208 6074 4413 6077
tri 4413 6074 4456 6117 sw
rect 4208 6043 4456 6074
rect 4046 6037 4456 6043
tri 4456 6037 4493 6074 sw
tri 3947 6005 3948 6006 sw
rect 4046 6005 4493 6037
rect 3895 5989 3948 6005
tri 3948 5989 3964 6005 sw
tri 4295 5989 4311 6005 ne
rect 4311 5989 4493 6005
tri 4493 5989 4541 6037 sw
rect 3895 5984 3964 5989
tri 3964 5984 3969 5989 sw
tri 4311 5984 4316 5989 ne
rect 4316 5984 4541 5989
tri 3895 5961 3918 5984 ne
rect 3918 5961 3969 5984
tri 3969 5961 3992 5984 sw
tri 4316 5961 4339 5984 ne
rect 4339 5961 4541 5984
tri 3918 5955 3924 5961 ne
rect 3924 5955 4088 5961
tri 4339 5955 4345 5961 ne
rect 4345 5955 4541 5961
tri 3924 5949 3930 5955 ne
rect 3930 5949 4036 5955
tri 3930 5910 3969 5949 ne
rect 3969 5910 4036 5949
tri 3969 5891 3988 5910 ne
rect 3988 5903 4036 5910
tri 4345 5949 4351 5955 ne
rect 4351 5949 4541 5955
rect 3988 5891 4088 5903
tri 4351 5891 4409 5949 ne
tri 3988 5843 4036 5891 ne
rect 4036 5833 4088 5839
tri 3812 5705 3815 5708 ne
rect 3815 5705 3864 5708
tri 3864 5705 3889 5730 sw
tri 3815 5656 3864 5705 ne
rect 3864 5656 3889 5705
tri 3864 5631 3889 5656 ne
tri 3889 5631 3963 5705 sw
rect 4409 5633 4541 5949
rect 4571 6013 4703 6385
tri 11370 6185 11398 6213 ne
rect 11398 6185 11404 6213
tri 7907 6179 7913 6185 ne
rect 7913 6179 7941 6185
tri 11398 6179 11404 6185 ne
tri 7913 6151 7941 6179 ne
rect 13764 6021 14044 6089
rect 4571 5961 4577 6013
rect 4629 5961 4645 6013
rect 4697 5961 4703 6013
rect 4571 5935 4703 5961
rect 4571 5883 4577 5935
rect 4629 5883 4645 5935
rect 4697 5883 4703 5935
rect 13392 5969 13398 6021
rect 13450 5969 13472 6021
rect 13524 5969 13545 6021
rect 13597 5969 13618 6021
rect 13670 5969 13691 6021
rect 13743 5969 13764 6021
rect 13816 5969 14044 6021
rect 13392 5949 14044 5969
rect 13392 5897 13398 5949
rect 13450 5897 13472 5949
rect 13524 5897 13545 5949
rect 13597 5897 13618 5949
rect 13670 5897 13691 5949
rect 13743 5897 13764 5949
rect 13816 5897 14044 5949
tri 3889 5583 3937 5631 ne
rect 3937 5583 3963 5631
tri 3963 5583 4011 5631 sw
tri 3937 5557 3963 5583 ne
rect 3963 5557 4011 5583
tri 4011 5557 4037 5583 sw
rect 4409 5581 4415 5633
rect 4467 5581 4483 5633
rect 4535 5581 4541 5633
rect 13392 5877 14044 5897
rect 13392 5825 13398 5877
rect 13450 5825 13472 5877
rect 13524 5825 13545 5877
rect 13597 5825 13618 5877
rect 13670 5825 13691 5877
rect 13743 5825 13764 5877
rect 13816 5825 14044 5877
rect 13392 5805 14044 5825
rect 13392 5753 13398 5805
rect 13450 5753 13472 5805
rect 13524 5753 13545 5805
rect 13597 5753 13618 5805
rect 13670 5753 13691 5805
rect 13743 5753 13764 5805
rect 13816 5753 14044 5805
rect 13392 5733 14044 5753
rect 13392 5681 13398 5733
rect 13450 5681 13472 5733
rect 13524 5681 13545 5733
rect 13597 5681 13618 5733
rect 13670 5681 13691 5733
rect 13743 5681 13764 5733
rect 13816 5681 14044 5733
rect 13392 5661 14044 5681
rect 13392 5609 13398 5661
rect 13450 5609 13472 5661
rect 13524 5609 13545 5661
rect 13597 5609 13618 5661
rect 13670 5609 13691 5661
rect 13743 5609 13764 5661
rect 13816 5609 14044 5661
tri 3963 5549 3971 5557 ne
rect 3971 5549 4037 5557
tri 4037 5549 4045 5557 sw
rect 4409 5555 4541 5581
tri 3971 5497 4023 5549 ne
rect 4023 5503 4045 5549
tri 4045 5503 4091 5549 sw
rect 4409 5503 4415 5555
rect 4467 5503 4483 5555
rect 4535 5503 4541 5555
tri 4720 5517 4742 5539 se
rect 13764 5517 14044 5609
tri 4706 5503 4720 5517 se
rect 4720 5503 4742 5517
rect 4023 5497 4091 5503
tri 4091 5497 4097 5503 sw
tri 4700 5497 4706 5503 se
rect 4706 5497 4742 5503
tri 4023 5483 4037 5497 ne
rect 4037 5483 4097 5497
tri 4097 5483 4111 5497 sw
tri 4686 5483 4700 5497 se
rect 4700 5483 4742 5497
tri 4037 5482 4038 5483 ne
rect 4038 5482 4111 5483
tri 4111 5482 4112 5483 sw
tri 4685 5482 4686 5483 se
rect 4686 5482 4742 5483
tri 4038 5476 4044 5482 ne
rect 4044 5476 4112 5482
tri 4112 5476 4118 5482 sw
tri 4679 5476 4685 5482 se
rect 4685 5476 4742 5482
tri 2976 5442 3006 5472 sw
rect 3289 5442 3293 5472
tri 3293 5442 3323 5472 sw
tri 3687 5442 3717 5472 se
rect 3717 5442 3773 5472
tri 4044 5442 4078 5476 ne
rect 4078 5442 4118 5476
tri 4118 5442 4152 5476 sw
tri 4645 5442 4679 5476 se
rect 4679 5442 4742 5476
rect 2976 5438 3006 5442
tri 3006 5438 3010 5442 sw
tri 4078 5438 4082 5442 ne
rect 4082 5438 4152 5442
tri 4152 5438 4156 5442 sw
tri 4641 5438 4645 5442 se
rect 4645 5438 4742 5442
tri 4082 5415 4105 5438 ne
rect 4105 5415 4156 5438
tri 4156 5415 4179 5438 sw
tri 4618 5415 4641 5438 se
rect 4641 5415 4742 5438
tri 3289 5413 3291 5415 nw
tri 4105 5413 4107 5415 ne
rect 4107 5413 4179 5415
tri 4179 5413 4181 5415 sw
tri 4616 5413 4618 5415 se
rect 4618 5413 4742 5415
tri 4107 5409 4111 5413 ne
rect 4111 5409 4181 5413
tri 4181 5409 4185 5413 sw
tri 4612 5409 4616 5413 se
rect 4616 5409 4742 5413
tri 4111 5385 4135 5409 ne
rect 4135 5385 4185 5409
tri 4185 5385 4209 5409 sw
tri 4588 5385 4612 5409 se
rect 4612 5385 4742 5409
tri 3197 5383 3199 5385 sw
tri 4135 5383 4137 5385 ne
rect 4137 5383 4209 5385
tri 2758 5381 2760 5383 ne
rect 2812 5351 2814 5383
tri 2814 5351 2846 5383 nw
rect 3197 5351 3199 5383
tri 3199 5351 3231 5383 sw
tri 4137 5351 4169 5383 ne
rect 4169 5351 4209 5383
tri 4209 5351 4243 5385 sw
tri 4554 5351 4588 5385 se
rect 4588 5351 4742 5385
tri 2812 5349 2814 5351 nw
rect 2929 5305 2950 5351
rect 3057 5298 3080 5350
rect 3189 5301 3219 5305
tri 3219 5301 3223 5305 nw
rect 3189 5294 3212 5301
tri 3212 5294 3219 5301 nw
rect 3485 5299 3491 5351
rect 3543 5299 3555 5351
rect 3607 5346 3696 5351
tri 3696 5346 3701 5351 sw
tri 4169 5346 4174 5351 ne
rect 4174 5346 4243 5351
tri 4243 5346 4248 5351 sw
tri 4549 5346 4554 5351 se
rect 4554 5346 4742 5351
rect 3607 5335 3701 5346
tri 3701 5335 3712 5346 sw
rect 3607 5309 3712 5335
tri 3712 5309 3738 5335 sw
rect 3607 5299 3738 5309
tri 3647 5294 3652 5299 ne
rect 3652 5294 3738 5299
rect 3778 5294 3784 5346
rect 3836 5294 3848 5346
rect 3900 5294 3906 5346
tri 4174 5335 4185 5346 ne
rect 4185 5341 4248 5346
tri 4248 5341 4253 5346 sw
tri 4544 5341 4549 5346 se
rect 4549 5341 4742 5346
rect 4185 5335 4253 5341
tri 4253 5335 4259 5341 sw
tri 4538 5335 4544 5341 se
rect 4544 5335 4742 5341
tri 4185 5301 4219 5335 ne
rect 4219 5301 4259 5335
tri 4259 5301 4293 5335 sw
tri 4504 5301 4538 5335 se
rect 4538 5301 4579 5335
rect 4613 5301 4651 5335
rect 4685 5301 4742 5335
tri 3189 5271 3212 5294 nw
tri 3652 5271 3675 5294 ne
rect 3675 5271 3738 5294
tri 3675 5260 3686 5271 ne
rect 3266 5200 3268 5252
tri 2524 5171 2527 5174 se
rect 2527 5171 2598 5174
tri 2598 5171 2601 5174 nw
tri 2376 5157 2390 5171 se
rect 2390 5157 2450 5171
tri 2450 5157 2464 5171 nw
tri 2510 5157 2524 5171 se
rect 2524 5157 2584 5171
tri 2584 5157 2598 5171 nw
tri 2356 5137 2376 5157 se
rect 2376 5137 2430 5157
tri 2430 5137 2450 5157 nw
tri 2490 5137 2510 5157 se
rect 2510 5137 2564 5157
tri 2564 5137 2584 5157 nw
tri 2350 5131 2356 5137 se
rect 2356 5131 2424 5137
tri 2424 5131 2430 5137 nw
tri 2484 5131 2490 5137 se
rect 2490 5131 2558 5137
tri 2558 5131 2564 5137 nw
tri 2346 5127 2350 5131 se
rect 2350 5127 2420 5131
tri 2420 5127 2424 5131 nw
tri 2480 5127 2484 5131 se
rect 2484 5127 2554 5131
tri 2554 5127 2558 5131 nw
tri 2913 5127 2917 5131 ne
tri 2333 5114 2346 5127 se
rect 2346 5123 2416 5127
tri 2416 5123 2420 5127 nw
tri 2476 5123 2480 5127 se
rect 2480 5123 2541 5127
rect 2346 5114 2407 5123
tri 2407 5114 2416 5123 nw
tri 2467 5114 2476 5123 se
rect 2476 5114 2541 5123
tri 2541 5114 2554 5127 nw
tri 14 5063 25 5074 se
tri -9 5040 14 5063 se
rect 14 5040 25 5063
tri 71 5063 82 5074 sw
rect 71 5062 82 5063
tri 82 5062 83 5063 sw
rect 2154 5062 2160 5114
rect 2212 5062 2224 5114
rect 2276 5097 2390 5114
tri 2390 5097 2407 5114 nw
tri 2450 5097 2467 5114 se
rect 2467 5097 2524 5114
tri 2524 5097 2541 5114 nw
rect 2276 5063 2356 5097
tri 2356 5063 2390 5097 nw
tri 2416 5063 2450 5097 se
rect 2450 5063 2490 5097
tri 2490 5063 2524 5097 nw
rect 2276 5062 2355 5063
tri 2355 5062 2356 5063 nw
tri 2415 5062 2416 5063 se
rect 2416 5062 2489 5063
tri 2489 5062 2490 5063 nw
rect 71 5054 83 5062
tri 83 5054 91 5062 sw
tri 2407 5054 2415 5062 se
rect 2415 5054 2481 5062
tri 2481 5054 2489 5062 nw
rect 71 5040 91 5054
tri 91 5040 105 5054 sw
tri 2393 5040 2407 5054 se
rect 2407 5040 2467 5054
tri 2467 5040 2481 5054 nw
tri 2643 5040 2657 5054 se
tri 2376 5023 2393 5040 se
rect 2393 5023 2450 5040
tri 2450 5023 2467 5040 nw
tri 2626 5023 2643 5040 se
rect 2643 5023 2657 5040
tri 2342 4989 2376 5023 se
rect 2376 5020 2447 5023
tri 2447 5020 2450 5023 nw
tri 2623 5020 2626 5023 se
rect 2626 5020 2657 5023
tri 2703 5023 2734 5054 sw
tri 3189 5023 3220 5054 sw
rect 2703 5020 2734 5023
tri 2734 5020 2737 5023 sw
rect 3189 5020 3220 5023
tri 3220 5020 3223 5023 sw
rect 2376 4989 2416 5020
tri 2416 4989 2447 5020 nw
tri 2302 4949 2342 4989 se
rect 2342 4949 2376 4989
tri 2376 4949 2416 4989 nw
tri 2268 4915 2302 4949 se
rect 2302 4915 2342 4949
tri 2342 4915 2376 4949 nw
tri 2246 4893 2268 4915 se
rect 2268 4893 2320 4915
tri 2320 4893 2342 4915 nw
rect 1953 4841 1959 4893
rect 2011 4841 2023 4893
rect 2075 4875 2302 4893
tri 2302 4875 2320 4893 nw
rect 2075 4841 2268 4875
tri 2268 4841 2302 4875 nw
tri 3426 4813 3451 4838 se
tri 3427 4727 3429 4729 ne
rect 3429 4727 3451 4729
tri 3429 4705 3451 4727 ne
rect 2691 4673 2711 4701
rect 2908 4639 3054 4645
rect 470 4570 498 4598
rect 2960 4587 3002 4639
rect 1789 4559 1817 4587
rect 2908 4573 3054 4587
rect 2960 4521 3002 4573
rect 2908 4506 3054 4521
rect 2960 4454 3002 4506
rect 2908 4448 3054 4454
tri 3652 4376 3686 4410 se
rect 3686 4376 3738 5271
rect 3824 5245 3857 5294
tri 3857 5245 3906 5294 nw
tri 4219 5261 4259 5301 ne
rect 4259 5295 4293 5301
tri 4293 5295 4299 5301 sw
tri 4498 5295 4504 5301 se
rect 4504 5295 4742 5301
rect 4259 5261 4299 5295
tri 4299 5261 4333 5295 sw
tri 4259 5257 4263 5261 ne
rect 4263 5257 4333 5261
tri 4460 5257 4498 5295 se
rect 4498 5257 4742 5295
tri 4263 5256 4264 5257 ne
rect 4264 5256 4333 5257
tri 4264 5245 4275 5256 ne
rect 4275 5245 4333 5256
tri 3824 5212 3857 5245 nw
tri 4275 5239 4281 5245 ne
tri 3932 5123 3936 5127 ne
rect 3971 5122 3975 5127
tri 3971 5118 3975 5122 ne
tri 3975 5118 3984 5127 nw
tri 3852 5024 3856 5028 ne
rect 3895 5023 3899 5028
tri 3899 5023 3904 5028 nw
rect 3895 5020 3896 5023
tri 3896 5020 3899 5023 nw
tri 3895 5019 3896 5020 nw
tri 4127 4702 4152 4727 nw
tri 4011 4626 4014 4629 ne
rect 4014 4626 4024 4629
tri 4014 4616 4024 4626 ne
rect 4050 4626 4060 4629
tri 4060 4626 4063 4629 nw
tri 4050 4616 4060 4626 nw
rect 4281 4611 4333 5245
tri 4456 5253 4459 5256 se
rect 4459 5253 4742 5257
rect 4456 5245 4742 5253
rect 4456 5211 4466 5245
rect 4500 5211 4556 5245
rect 4590 5211 4646 5245
rect 4680 5211 4742 5245
rect 4456 5171 4742 5211
rect 4456 5137 4466 5171
rect 4500 5137 4556 5171
rect 4590 5137 4646 5171
rect 4680 5137 4742 5171
rect 4456 5097 4742 5137
rect 4456 5063 4466 5097
rect 4500 5063 4556 5097
rect 4590 5063 4646 5097
rect 4680 5063 4742 5097
rect 4456 5023 4742 5063
rect 13983 5273 14035 5279
rect 13983 5206 14035 5221
rect 13983 5139 14035 5154
rect 13983 5072 14035 5087
rect 4456 4989 4466 5023
rect 4500 4989 4556 5023
rect 4590 4989 4646 5023
rect 4680 4989 4742 5023
rect 4456 4949 4742 4989
rect 4456 4915 4466 4949
rect 4500 4915 4556 4949
rect 4590 4915 4646 4949
rect 4680 4915 4742 4949
rect 4456 4875 4742 4915
rect 4456 4841 4466 4875
rect 4500 4841 4556 4875
rect 4590 4841 4646 4875
rect 4680 4841 4742 4875
rect 4456 4801 4742 4841
rect 4456 4767 4466 4801
rect 4500 4767 4556 4801
rect 4590 4767 4646 4801
rect 4680 4767 4742 4801
rect 4456 4727 4742 4767
rect 4456 4693 4466 4727
rect 4500 4693 4556 4727
rect 4590 4693 4646 4727
rect 4680 4693 4742 4727
rect 4456 4685 4742 4693
tri 4456 4682 4459 4685 ne
rect 4459 4681 4742 4685
tri 4460 4632 4509 4681 ne
rect 4509 4632 4742 4681
tri 4509 4626 4515 4632 ne
rect 4515 4626 4742 4632
tri 4515 4592 4549 4626 ne
rect 4549 4592 4579 4626
rect 4613 4592 4651 4626
rect 4685 4592 4742 4626
tri 4549 4586 4555 4592 ne
rect 4555 4586 4742 4592
rect 4281 4547 4333 4559
rect 4281 4489 4333 4495
tri 4555 4489 4652 4586 ne
rect 4652 4489 4742 4586
tri 4652 4416 4725 4489 ne
rect 4725 4416 4742 4489
rect 4930 5047 5032 5053
rect 4930 4995 4955 5047
rect 5007 4995 5032 5047
rect 4930 4975 5032 4995
rect 4930 4923 4955 4975
rect 5007 4923 5032 4975
rect 4930 4902 5032 4923
rect 4930 4850 4955 4902
rect 5007 4850 5032 4902
rect 4930 4829 5032 4850
rect 4930 4777 4955 4829
rect 5007 4777 5032 4829
rect 4930 4756 5032 4777
rect 4930 4704 4955 4756
rect 5007 4704 5032 4756
rect 4930 4683 5032 4704
rect 4930 4631 4955 4683
rect 5007 4631 5032 4683
rect 13983 5005 14035 5020
rect 13983 4938 14035 4953
rect 13983 4871 14035 4886
rect 13983 4803 14035 4819
rect 13983 4735 14035 4751
rect 13983 4667 14035 4683
tri 5115 4647 5118 4650 ne
tri 8751 4647 8754 4650 ne
tri 8800 4647 8803 4650 nw
rect 4930 4610 5032 4631
rect 4930 4558 4955 4610
rect 5007 4587 5032 4610
tri 5032 4587 5060 4615 sw
tri 7913 4587 7941 4615 se
rect 13983 4609 14035 4615
rect 5007 4581 5060 4587
tri 5060 4581 5066 4587 sw
tri 7907 4581 7913 4587 se
rect 7913 4581 7941 4587
tri 8800 4581 8806 4587 sw
rect 5007 4558 5032 4581
rect 4930 4537 5032 4558
rect 8800 4553 8806 4581
tri 8806 4553 8834 4581 sw
rect 4930 4485 4955 4537
rect 5007 4485 5032 4537
rect 4930 4479 5032 4485
rect 3441 4324 3738 4376
rect 4369 4410 4589 4416
tri 4725 4410 4731 4416 ne
rect 4731 4410 4742 4416
rect 4421 4358 4537 4410
rect 5075 4358 5081 4410
rect 5133 4358 5145 4410
rect 5197 4358 5658 4410
rect 5710 4358 5722 4410
rect 5774 4358 5780 4410
tri 8607 4358 8609 4360 sw
tri 14903 4358 14905 4360 se
rect 4369 4346 4589 4358
rect 8607 4352 8609 4358
tri 8609 4352 8615 4358 sw
tri 14897 4352 14903 4358 se
rect 14903 4352 14905 4358
rect 3441 4314 3517 4324
tri 3517 4314 3527 4324 nw
rect -651 3961 -626 3970
tri -626 3961 -617 3970 nw
tri 2768 3961 2777 3970 ne
rect 2777 3961 2802 3970
rect -651 3954 -633 3961
tri -633 3954 -626 3961 nw
tri 2777 3954 2784 3961 ne
rect 2784 3954 2802 3961
tri -651 3936 -633 3954 nw
tri 2784 3936 2802 3954 ne
rect -493 3863 -476 3915
rect 2755 3863 2759 3915
tri -215 3842 -212 3845 ne
rect -212 3842 -181 3845
tri -212 3828 -198 3842 ne
rect -198 3828 -181 3842
rect 2332 3842 2363 3845
tri 2363 3842 2366 3845 nw
tri 266 3828 270 3832 ne
rect 270 3828 272 3832
tri -198 3825 -195 3828 ne
rect -195 3825 -181 3828
tri 270 3826 272 3828 ne
tri 695 3826 697 3828 sw
rect -618 3773 -616 3825
tri -195 3817 -187 3825 ne
rect -187 3817 -181 3825
rect 695 3825 697 3826
tri 697 3825 698 3826 sw
tri -187 3815 -185 3817 ne
rect -185 3815 -181 3817
tri 641 3815 643 3817 se
tri -185 3811 -181 3815 ne
tri 637 3811 641 3815 se
rect 641 3811 643 3815
tri 636 3810 637 3811 se
rect 637 3810 643 3811
tri 634 3808 636 3810 se
rect 636 3808 643 3810
rect -257 3756 -255 3808
tri 620 3794 634 3808 se
rect 634 3794 643 3808
rect 695 3815 698 3825
tri 698 3815 708 3825 sw
rect 2332 3815 2336 3842
tri 2336 3815 2363 3842 nw
rect 695 3811 708 3815
tri 708 3811 712 3815 sw
rect 2332 3812 2333 3815
tri 2333 3812 2336 3815 nw
tri 2332 3811 2333 3812 nw
rect 695 3810 712 3811
tri 712 3810 713 3811 sw
rect 695 3804 713 3810
tri 713 3804 719 3810 sw
rect 695 3794 719 3804
tri 719 3794 729 3804 sw
rect 2406 3752 2408 3804
tri -730 3632 -722 3640 se
tri -735 3627 -730 3632 se
rect -730 3627 -722 3632
tri -739 3623 -735 3627 se
rect -735 3623 -722 3627
tri -741 3621 -739 3623 se
rect -739 3621 -722 3623
tri -765 3597 -741 3621 se
rect -741 3597 -722 3621
tri -766 3596 -765 3597 se
rect -765 3596 -722 3597
tri -767 3595 -766 3596 se
rect -766 3595 -722 3596
rect -662 3623 -659 3627
tri -659 3623 -655 3627 sw
rect -662 3621 -655 3623
tri -655 3621 -653 3623 sw
rect -662 3597 -653 3621
tri -653 3597 -629 3621 sw
rect -662 3596 -629 3597
tri -629 3596 -628 3597 sw
rect -662 3594 -628 3596
tri -628 3594 -626 3596 sw
rect -662 3582 -626 3594
tri -626 3582 -614 3594 sw
rect -662 3562 -614 3582
tri -614 3562 -594 3582 sw
tri -508 3562 -488 3582 se
tri -442 3562 -422 3582 sw
rect -662 3561 -594 3562
tri -594 3561 -593 3562 sw
rect 1260 3378 1407 3381
tri 1407 3378 1410 3381 nw
tri 1749 3378 1752 3381 ne
rect 1752 3378 1783 3381
rect 1260 3344 1373 3378
tri 1373 3344 1407 3378 nw
tri 1752 3347 1783 3378 ne
rect 1829 3378 1860 3381
tri 1860 3378 1863 3381 nw
tri 2455 3378 2458 3381 ne
rect 2458 3378 2489 3381
tri 1829 3347 1860 3378 nw
tri 2458 3347 2489 3378 ne
rect 2535 3378 2566 3381
tri 2566 3378 2569 3381 nw
tri 2740 3378 2743 3381 ne
rect 2743 3378 2768 3381
tri 2535 3347 2566 3378 nw
tri 2743 3353 2768 3378 ne
rect 2814 3378 2845 3381
tri 2845 3378 2848 3381 nw
rect 2814 3353 2820 3378
tri 2820 3353 2845 3378 nw
tri 2814 3347 2820 3353 nw
rect 1260 3342 1371 3344
tri 1371 3342 1373 3344 nw
rect 1260 3340 1369 3342
tri 1369 3340 1371 3342 nw
rect 1260 3338 1367 3340
tri 1367 3338 1369 3340 nw
tri 1485 3338 1487 3340 se
rect 1487 3338 1493 3340
rect 1260 3337 1366 3338
tri 1366 3337 1367 3338 nw
rect 1260 3330 1359 3337
tri 1359 3330 1366 3337 nw
tri 1863 3330 1870 3337 se
rect 1870 3330 2243 3337
rect 1260 3324 1353 3330
tri 1353 3324 1359 3330 nw
tri 1857 3324 1863 3330 se
rect 1863 3324 2243 3330
rect 1260 3306 1335 3324
tri 1335 3306 1353 3324 nw
rect 1260 3299 1328 3306
tri 1328 3299 1335 3306 nw
rect 1857 3305 2243 3324
rect 1260 3286 1315 3299
tri 1315 3286 1328 3299 nw
rect 1857 3295 1925 3305
rect 1518 3286 1544 3294
tri 1544 3286 1552 3294 nw
rect 1260 3274 1303 3286
tri 1303 3274 1315 3286 nw
rect 1518 3274 1532 3286
tri 1532 3274 1544 3286 nw
rect 1260 3265 1294 3274
tri 1294 3265 1303 3274 nw
rect 1518 3265 1523 3274
tri 1523 3265 1532 3274 nw
rect 1260 3264 1293 3265
tri 1293 3264 1294 3265 nw
rect 1518 3264 1522 3265
tri 1522 3264 1523 3265 nw
rect -615 3252 -598 3264
tri -598 3252 -586 3264 nw
rect 1260 3259 1288 3264
tri 1288 3259 1293 3264 nw
tri 1518 3260 1522 3264 nw
tri -511 3252 -504 3259 ne
rect -504 3252 -483 3259
rect 1260 3258 1287 3259
tri 1287 3258 1288 3259 nw
rect -615 3250 -600 3252
tri -600 3250 -598 3252 nw
tri -504 3250 -502 3252 ne
rect -502 3250 -483 3252
rect -615 3240 -610 3250
tri -610 3240 -600 3250 nw
tri -502 3240 -492 3250 ne
rect -492 3240 -483 3250
rect -658 3234 -616 3240
tri -616 3234 -610 3240 nw
tri -492 3236 -488 3240 ne
rect -488 3236 -483 3240
rect -443 3252 -426 3258
tri -426 3252 -420 3258 nw
rect 1260 3252 1281 3258
tri 1281 3252 1287 3258 nw
rect -443 3250 -428 3252
tri -428 3250 -426 3252 nw
rect 1260 3250 1279 3252
tri 1279 3250 1281 3252 nw
rect -443 3236 -442 3250
tri -442 3236 -428 3250 nw
rect 1260 3236 1265 3250
tri 1265 3236 1279 3250 nw
rect 1909 3292 1925 3295
tri 1925 3292 1938 3305 nw
tri 2151 3292 2164 3305 ne
rect 2164 3295 2243 3305
rect 2164 3292 2191 3295
rect 1909 3286 1919 3292
tri 1919 3286 1925 3292 nw
tri 2164 3286 2170 3292 ne
rect 2170 3286 2191 3292
tri 1909 3276 1919 3286 nw
tri 2170 3276 2180 3286 ne
rect 2180 3276 2191 3286
tri 2180 3274 2182 3276 ne
rect 2182 3274 2191 3276
tri 2182 3265 2191 3274 ne
rect 1260 3234 1263 3236
tri 1263 3234 1265 3236 nw
rect -658 3223 -627 3234
tri -627 3223 -616 3234 nw
tri 1260 3231 1263 3234 nw
rect 1857 3231 1909 3243
tri -767 3200 -744 3223 ne
rect -744 3200 -711 3223
tri -744 3195 -739 3200 ne
rect -739 3195 -711 3200
tri -739 3194 -738 3195 ne
rect -738 3194 -711 3195
tri -738 3192 -736 3194 ne
rect -736 3192 -711 3194
rect -658 3200 -650 3223
tri -650 3200 -627 3223 nw
tri 1023 3200 1046 3223 ne
rect 1046 3200 1104 3223
rect -658 3195 -655 3200
tri -655 3195 -650 3200 nw
tri 1046 3195 1051 3200 ne
rect 1051 3195 1104 3200
rect -658 3194 -656 3195
tri -656 3194 -655 3195 nw
tri 1051 3194 1052 3195 ne
rect 1052 3194 1104 3195
tri 1672 3200 1673 3201 sw
rect 1672 3195 1673 3200
tri 1673 3195 1678 3200 sw
rect 1672 3194 1678 3195
tri 1678 3194 1679 3195 sw
tri -658 3192 -656 3194 nw
tri 1052 3192 1054 3194 ne
rect 1054 3192 1104 3194
tri -736 3177 -721 3192 ne
rect -721 3187 -711 3192
tri -721 3177 -711 3187 nw
tri 1054 3177 1069 3192 ne
rect 1069 3177 1104 3192
tri 1069 3173 1073 3177 ne
rect 1073 3173 1104 3177
rect 1857 3173 1909 3179
rect 2599 3291 2610 3343
rect 2191 3231 2243 3243
rect 2191 3173 2243 3179
tri 1073 3170 1076 3173 ne
rect 1076 3170 1104 3173
tri 1076 3142 1104 3170 ne
rect 2318 3166 2370 3236
rect 2639 3166 2691 3236
tri 3411 3200 3441 3230 se
rect 3441 3200 3493 4314
tri 3493 4290 3517 4314 nw
rect 4421 4294 4537 4346
tri 4833 4326 4859 4352 sw
tri 8164 4326 8190 4352 se
rect 8607 4326 8615 4352
tri 8615 4326 8641 4352 sw
tri 14888 4343 14897 4352 se
rect 14897 4343 14905 4352
tri 13739 4341 13741 4343 ne
tri 14886 4341 14888 4343 se
rect 14888 4341 14905 4343
tri 14871 4326 14886 4341 se
rect 14886 4326 14905 4341
tri 15012 4326 15023 4337 sw
rect 4833 4318 4859 4326
tri 4859 4318 4867 4326 sw
tri 8156 4318 8164 4326 se
rect 8164 4318 8190 4326
tri 13165 4318 13173 4326 ne
rect 13173 4318 13267 4326
rect 4369 4288 4589 4294
rect 5915 4293 6186 4318
tri 13173 4314 13177 4318 ne
rect 13177 4314 13267 4318
tri 13267 4314 13279 4326 nw
tri 14943 4314 14955 4326 ne
rect 14955 4314 15023 4326
tri 3770 4269 3778 4277 se
tri 3746 4245 3770 4269 se
rect 3770 4245 3778 4269
tri 3744 4243 3746 4245 se
rect 3746 4243 3778 4245
rect 5915 4241 5921 4293
rect 5973 4241 6025 4293
rect 6077 4241 6128 4293
rect 6180 4241 6186 4293
tri 13177 4292 13199 4314 ne
rect 13199 4280 13205 4314
rect 13239 4280 13245 4314
tri 13245 4292 13267 4314 nw
tri 14955 4292 14977 4314 ne
tri 11953 4245 11977 4269 se
rect 11977 4245 12928 4269
tri 6665 4242 6668 4245 ne
tri 6714 4242 6717 4245 nw
tri 6991 4242 6994 4245 ne
tri 7040 4242 7043 4245 nw
tri 7317 4242 7320 4245 ne
tri 7366 4242 7369 4245 nw
tri 11024 4242 11027 4245 ne
tri 11073 4242 11076 4245 nw
tri 11950 4242 11953 4245 se
rect 11953 4242 12928 4245
tri 4209 4217 4214 4222 sw
rect 4209 4208 4214 4217
tri 4214 4208 4223 4217 sw
rect 5915 4216 6186 4241
tri 11925 4217 11950 4242 se
rect 11950 4217 12928 4242
rect 12980 4217 12992 4269
rect 13044 4217 13050 4269
rect 13199 4242 13245 4280
rect 14977 4280 14983 4314
rect 15017 4280 15023 4314
tri 11924 4216 11925 4217 se
rect 11925 4216 11990 4217
tri 11916 4208 11924 4216 se
rect 11924 4208 11990 4216
tri 11990 4208 11999 4217 nw
rect 13199 4208 13205 4242
rect 13239 4208 13245 4242
rect 13546 4217 13552 4269
rect 13604 4217 13616 4269
rect 13668 4241 14669 4269
tri 14669 4241 14697 4269 sw
rect 14977 4241 15023 4280
rect 13668 4223 14697 4241
tri 14697 4223 14715 4241 sw
rect 13668 4217 13674 4223
tri 13674 4217 13680 4223 nw
tri 14649 4217 14655 4223 ne
rect 14655 4217 14715 4223
tri 14715 4217 14721 4223 sw
rect 4209 4207 4223 4208
tri 4223 4207 4224 4208 sw
tri 11915 4207 11916 4208 se
rect 11916 4207 11989 4208
tri 11989 4207 11990 4208 nw
rect 3583 4188 3608 4197
tri 3608 4188 3617 4197 nw
rect 4209 4192 4224 4207
tri 4224 4192 4239 4207 sw
tri 11904 4196 11915 4207 se
rect 11915 4196 11978 4207
tri 11978 4196 11989 4207 nw
rect 4209 4189 4239 4192
tri 4239 4189 4242 4192 sw
rect 4209 4188 4242 4189
tri 4242 4188 4243 4189 sw
rect 3583 4180 3600 4188
tri 3600 4180 3608 4188 nw
rect 3583 4170 3590 4180
tri 3590 4170 3600 4180 nw
tri 3583 4163 3590 4170 nw
rect 10312 4144 10318 4196
rect 10370 4144 10382 4196
rect 10434 4192 11974 4196
tri 11974 4192 11978 4196 nw
rect 10434 4189 11971 4192
tri 11971 4189 11974 4192 nw
rect 10434 4188 11970 4189
tri 11970 4188 11971 4189 nw
rect 10434 4180 11962 4188
tri 11962 4180 11970 4188 nw
rect 10434 4170 11952 4180
tri 11952 4170 11962 4180 nw
rect 13199 4170 13245 4208
tri 14655 4207 14665 4217 ne
rect 14665 4207 14721 4217
tri 14721 4207 14731 4217 sw
rect 14977 4207 14983 4241
rect 15017 4207 15023 4241
tri 14665 4205 14667 4207 ne
rect 14667 4205 14731 4207
tri 14731 4205 14733 4207 sw
tri 14667 4203 14669 4205 ne
rect 14669 4203 14733 4205
tri 14669 4192 14680 4203 ne
rect 14680 4192 14733 4203
tri 14680 4189 14683 4192 ne
rect 14683 4189 14733 4192
tri 14683 4188 14684 4189 ne
rect 14684 4188 14733 4189
tri 14684 4186 14686 4188 ne
rect 14686 4186 14733 4188
rect 10434 4144 11926 4170
tri 11926 4144 11952 4170 nw
rect 13199 4136 13205 4170
rect 13239 4136 13245 4170
rect 13199 4098 13245 4136
tri 4209 4064 4230 4085 sw
rect 13199 4064 13205 4098
rect 13239 4064 13245 4098
rect 4209 4057 4230 4064
tri 4230 4057 4237 4064 sw
rect 4209 4051 4237 4057
tri 4237 4051 4243 4057 sw
tri 10797 4026 10800 4029 sw
rect 13199 4026 13245 4064
rect 10797 4024 10800 4026
tri 10800 4024 10802 4026 sw
rect 4209 4018 4233 4023
tri 4233 4018 4238 4023 nw
rect 10797 4018 10802 4024
tri 10802 4018 10808 4024 sw
rect 11452 4018 11880 4024
rect 4209 4004 4219 4018
tri 4219 4004 4233 4018 nw
rect 4209 4001 4216 4004
tri 4216 4001 4219 4004 nw
tri 10125 4001 10128 4004 ne
rect 10128 4001 10159 4004
rect 10797 4001 10808 4018
tri 10808 4001 10825 4018 sw
tri 4209 3994 4216 4001 nw
tri 10128 3994 10135 4001 ne
rect 10135 3994 10159 4001
tri 10135 3984 10145 3994 ne
rect 10145 3984 10159 3994
tri 10709 3984 10726 4001 ne
rect 10726 3984 10743 4001
rect 10797 3999 10825 4001
tri 10825 3999 10827 4001 sw
tri 10145 3970 10159 3984 ne
tri 10726 3970 10740 3984 ne
rect 10740 3970 10743 3984
tri 10740 3967 10743 3970 ne
rect 11452 3984 11464 4018
rect 11498 3984 11538 4018
rect 11572 3984 11612 4018
rect 11646 3984 11686 4018
rect 11720 3984 11760 4018
rect 11794 3984 11834 4018
rect 11868 3984 11880 4018
rect 4302 3896 4308 3948
rect 4360 3896 4372 3948
rect 4424 3926 4430 3948
tri 4430 3926 4452 3948 sw
rect 4424 3897 5619 3926
tri 10743 3902 10746 3905 ne
rect 10746 3902 10777 3905
tri 10746 3897 10751 3902 ne
rect 10751 3897 10777 3902
rect 4424 3896 5623 3897
tri 5615 3892 5619 3896 ne
rect 5619 3892 5623 3896
tri 10751 3892 10756 3897 ne
rect 10756 3892 10777 3897
tri 10756 3871 10777 3892 ne
rect 11452 3902 11880 3984
rect 11452 3868 11464 3902
rect 11498 3868 11538 3902
rect 11572 3868 11612 3902
rect 11646 3868 11686 3902
rect 11720 3868 11760 3902
rect 11794 3868 11834 3902
rect 11868 3868 11880 3902
tri 7543 3842 7547 3846 ne
rect 7547 3842 7577 3846
tri 7547 3815 7574 3842 ne
rect 7574 3815 7577 3842
tri 7574 3812 7577 3815 ne
tri 8450 3776 8456 3782 se
rect 8456 3776 9400 3782
tri 8444 3770 8450 3776 se
rect 8450 3770 9400 3776
tri 8441 3767 8444 3770 se
rect 8444 3767 9400 3770
tri 8432 3758 8441 3767 se
rect 8441 3758 9400 3767
tri 8430 3756 8432 3758 se
rect 8432 3756 8474 3758
rect 4228 3735 4241 3756
tri 4241 3735 4262 3756 nw
tri 8409 3735 8430 3756 se
rect 8430 3735 8474 3756
rect 4228 3724 4230 3735
tri 4230 3724 4241 3735 nw
tri 8006 3724 8017 3735 se
tri 8398 3724 8409 3735 se
rect 8409 3724 8474 3735
rect 8508 3724 8547 3758
rect 8581 3724 8620 3758
rect 8654 3724 8693 3758
rect 8727 3724 8766 3758
rect 8800 3724 8839 3758
rect 8873 3724 8912 3758
rect 8946 3724 8984 3758
rect 9018 3724 9056 3758
rect 9090 3724 9128 3758
rect 9162 3724 9200 3758
rect 9234 3724 9272 3758
rect 9306 3724 9344 3758
rect 9378 3724 9400 3758
tri 4228 3722 4230 3724 nw
tri 8004 3722 8006 3724 se
rect 8006 3722 8017 3724
tri 7993 3711 8004 3722 se
rect 8004 3711 8017 3722
tri 8385 3711 8398 3724 se
rect 8398 3711 9400 3724
tri 8378 3704 8385 3711 se
rect 8385 3704 9400 3711
tri 8375 3701 8378 3704 se
rect 8378 3701 9400 3704
tri 8357 3683 8375 3701 se
rect 8375 3683 9400 3701
rect 4447 3678 4476 3683
tri 4476 3678 4481 3683 nw
tri 8352 3678 8357 3683 se
rect 8357 3678 9400 3683
rect 11452 3678 11880 3868
rect 11952 4018 12380 4024
rect 11952 3984 11964 4018
rect 11998 3984 12038 4018
rect 12072 3984 12112 4018
rect 12146 3984 12186 4018
rect 12220 3984 12260 4018
rect 12294 3984 12334 4018
rect 12368 3984 12380 4018
rect 11952 3902 12380 3984
rect 11952 3868 11964 3902
rect 11998 3868 12038 3902
rect 12072 3868 12112 3902
rect 12146 3868 12186 3902
rect 12220 3868 12260 3902
rect 12294 3868 12334 3902
rect 12368 3868 12380 3902
rect 11952 3810 12380 3868
rect 12453 4018 13061 4024
rect 12453 3984 12465 4018
rect 12499 3984 12539 4018
rect 12573 3984 12613 4018
rect 12647 3984 12687 4018
rect 12721 3984 12761 4018
rect 12795 3984 12835 4018
rect 12869 3984 13061 4018
rect 12453 3951 13061 3984
rect 12453 3902 12939 3951
rect 12453 3868 12465 3902
rect 12499 3868 12539 3902
rect 12573 3868 12613 3902
rect 12647 3868 12687 3902
rect 12721 3868 12761 3902
rect 12795 3868 12835 3902
rect 12869 3899 12939 3902
rect 12991 3899 13003 3951
rect 13055 3899 13061 3951
rect 12869 3868 13061 3899
rect 12453 3862 13061 3868
rect 13199 3992 13205 4026
rect 13239 3992 13245 4026
rect 13428 4180 14615 4186
tri 14686 4185 14687 4186 ne
rect 13428 4146 13509 4180
rect 13543 4146 13583 4180
rect 13617 4146 13657 4180
rect 13691 4146 13731 4180
rect 13765 4146 13805 4180
rect 13839 4146 13879 4180
rect 13913 4146 13953 4180
rect 13987 4146 14027 4180
rect 14061 4146 14101 4180
rect 14135 4146 14175 4180
rect 14209 4146 14249 4180
rect 14283 4146 14323 4180
rect 14357 4146 14397 4180
rect 14431 4146 14470 4180
rect 14504 4146 14543 4180
rect 14577 4146 14615 4180
rect 13428 4140 14615 4146
rect 13428 4134 13508 4140
tri 13508 4134 13514 4140 nw
rect 13428 4129 13503 4134
tri 13503 4129 13508 4134 nw
rect 13480 4109 13483 4129
tri 13483 4109 13503 4129 nw
tri 14667 4109 14687 4129 se
rect 14687 4109 14733 4186
tri 13480 4106 13483 4109 nw
tri 14664 4106 14667 4109 se
rect 14667 4106 14721 4109
tri 14655 4097 14664 4106 se
rect 14664 4097 14721 4106
tri 14721 4097 14733 4109 nw
rect 14977 4168 15023 4207
rect 14977 4134 14983 4168
rect 15017 4134 15023 4168
rect 13428 4073 13437 4077
rect 13471 4073 13480 4077
rect 13428 4065 13480 4073
rect 13599 4091 13978 4097
rect 13599 4057 13686 4091
rect 13802 4057 13850 4091
rect 13884 4057 13932 4091
rect 13966 4057 13978 4091
rect 13599 4051 13720 4057
tri 13686 4022 13715 4051 ne
rect 13715 4039 13720 4051
rect 13772 4051 13978 4057
rect 14156 4095 14719 4097
tri 14719 4095 14721 4097 nw
rect 14977 4095 15023 4134
rect 14156 4091 14685 4095
rect 14156 4057 14168 4091
rect 14202 4057 14249 4091
rect 14283 4057 14330 4091
rect 14364 4057 14411 4091
rect 14445 4057 14492 4091
rect 14526 4061 14685 4091
tri 14685 4061 14719 4095 nw
rect 14977 4061 14983 4095
rect 15017 4061 15023 4095
rect 14526 4057 14675 4061
rect 14156 4051 14675 4057
tri 14675 4051 14685 4061 nw
rect 13772 4039 13778 4051
rect 13715 4027 13778 4039
rect 13715 4022 13720 4027
tri 13715 4017 13720 4022 ne
rect 13428 4007 13437 4013
tri 13428 4004 13431 4007 ne
rect 13199 3954 13245 3992
rect 13199 3920 13205 3954
rect 13239 3920 13245 3954
rect 13199 3882 13245 3920
rect 13199 3848 13205 3882
rect 13239 3848 13245 3882
tri 12380 3810 12384 3814 sw
rect 13199 3810 13245 3848
rect 11952 3776 12384 3810
tri 12384 3776 12418 3810 sw
rect 13199 3776 13205 3810
rect 13239 3776 13245 3810
rect 11952 3770 12418 3776
tri 12418 3770 12424 3776 sw
rect 11952 3767 12424 3770
tri 12424 3767 12427 3770 sw
rect 11952 3755 12427 3767
tri 11952 3742 11965 3755 ne
rect 11965 3742 12427 3755
tri 12427 3742 12452 3767 sw
tri 11965 3738 11969 3742 ne
rect 11969 3738 12452 3742
tri 12452 3738 12456 3742 sw
rect 13199 3738 13245 3776
tri 11969 3709 11998 3738 ne
rect 11998 3709 12456 3738
tri 12456 3709 12485 3738 sw
tri 11998 3707 12000 3709 ne
rect 12000 3707 12939 3709
tri 12000 3704 12003 3707 ne
rect 12003 3704 12939 3707
tri 12003 3701 12006 3704 ne
rect 12006 3701 12939 3704
tri 12006 3700 12007 3701 ne
rect 12007 3700 12939 3701
tri 11880 3678 11902 3700 sw
tri 12007 3678 12029 3700 ne
rect 12029 3678 12939 3700
rect 4447 3672 4470 3678
tri 4470 3672 4476 3678 nw
tri 8346 3672 8352 3678 se
rect 8352 3673 9400 3678
rect 8352 3672 9119 3673
rect 4447 3669 4467 3672
tri 4467 3669 4470 3672 nw
tri 8343 3669 8346 3672 se
rect 8346 3669 9119 3672
rect 4447 3666 4464 3669
tri 4464 3666 4467 3669 nw
tri 8340 3666 8343 3669 se
rect 8343 3666 9119 3669
tri 4447 3649 4464 3666 nw
tri 8327 3653 8340 3666 se
rect 8340 3655 9119 3666
rect 8340 3653 8464 3655
rect 9113 3621 9119 3655
rect 9171 3621 9194 3673
rect 9246 3621 9268 3673
rect 9320 3621 9342 3673
rect 9394 3621 9400 3673
rect 9113 3609 9400 3621
rect 9113 3557 9119 3609
rect 9171 3557 9194 3609
rect 9246 3557 9268 3609
rect 9320 3557 9342 3609
rect 9394 3557 9400 3609
rect 10241 3626 10247 3678
rect 10299 3626 10315 3678
rect 10367 3626 10383 3678
rect 10435 3626 10451 3678
rect 10503 3626 10519 3678
rect 10571 3626 10587 3678
rect 10639 3626 10654 3678
rect 10706 3626 10712 3678
rect 10241 3606 10712 3626
rect 10241 3554 10247 3606
rect 10299 3554 10315 3606
rect 10367 3554 10383 3606
rect 10435 3554 10451 3606
rect 10503 3554 10519 3606
rect 10571 3554 10587 3606
rect 10639 3554 10654 3606
rect 10706 3554 10712 3606
rect 11452 3672 11902 3678
tri 11902 3672 11908 3678 sw
tri 12029 3672 12035 3678 ne
rect 12035 3672 12939 3678
rect 11452 3669 11908 3672
tri 11908 3669 11911 3672 sw
tri 12035 3669 12038 3672 ne
rect 12038 3669 12939 3672
rect 11452 3666 11911 3669
tri 11911 3666 11914 3669 sw
tri 12038 3666 12041 3669 ne
rect 12041 3666 12939 3669
rect 11452 3657 11914 3666
tri 11914 3657 11923 3666 sw
tri 12041 3657 12050 3666 ne
rect 12050 3657 12939 3666
rect 12991 3657 13003 3709
rect 13055 3657 13061 3709
rect 13199 3704 13205 3738
rect 13239 3704 13245 3738
rect 13199 3666 13245 3704
rect 11452 3644 11923 3657
tri 11923 3644 11936 3657 sw
rect 11452 3632 11936 3644
tri 11936 3632 11948 3644 sw
rect 13199 3632 13205 3666
rect 13239 3632 13245 3666
rect 11452 3623 11948 3632
tri 11948 3623 11957 3632 sw
rect 11452 3621 11957 3623
tri 11957 3621 11959 3623 sw
rect 11452 3604 11959 3621
tri 11959 3604 11976 3621 sw
rect 11452 3552 12930 3604
rect 12982 3552 12994 3604
rect 13046 3552 13052 3604
rect 13199 3594 13245 3632
rect 13199 3560 13205 3594
rect 13239 3560 13245 3594
rect 13199 3522 13245 3560
rect 13113 3514 13165 3520
rect 5450 3487 5502 3493
tri 5449 3450 5450 3451 se
tri 5445 3446 5449 3450 se
rect 5449 3446 5450 3450
rect 4176 3440 4228 3446
tri 4228 3417 4257 3446 sw
tri 5416 3417 5445 3446 se
rect 5445 3435 5450 3446
rect 5445 3423 5502 3435
tri 5710 3452 5725 3467 sw
rect 5710 3450 5725 3452
tri 5725 3450 5727 3452 sw
rect 13113 3450 13165 3462
rect 5710 3433 5727 3450
tri 5727 3433 5744 3450 sw
rect 5445 3417 5450 3423
rect 4228 3388 5450 3417
rect 4176 3376 5450 3388
rect 4228 3371 5450 3376
rect 5708 3404 5715 3408
tri 5715 3404 5719 3408 nw
rect 5708 3399 5710 3404
tri 5710 3399 5715 3404 nw
tri 6563 3371 6569 3377 sw
rect 4228 3365 5502 3371
tri 6505 3365 6511 3371 se
rect 4228 3354 4251 3365
tri 4251 3354 4262 3365 nw
tri 6494 3354 6505 3365 se
rect 6505 3354 6511 3365
rect 6563 3365 6569 3371
tri 6569 3365 6575 3371 sw
rect 6563 3364 6575 3365
tri 6575 3364 6576 3365 sw
rect 6563 3354 6576 3364
tri 6576 3354 6586 3364 sw
rect 4228 3344 4241 3354
tri 4241 3344 4251 3354 nw
rect 4228 3342 4239 3344
tri 4239 3342 4241 3344 nw
tri 4228 3331 4239 3342 nw
rect 4176 3318 4228 3324
tri 6776 3308 6779 3311 se
tri 6494 3306 6496 3308 ne
rect 6496 3306 6512 3308
tri 6496 3290 6512 3306 ne
rect 6563 3306 6595 3308
tri 6595 3306 6597 3308 nw
tri 6774 3306 6776 3308 se
rect 6776 3306 6779 3308
rect 5210 3259 5238 3287
rect 6563 3286 6575 3306
tri 6575 3286 6595 3306 nw
tri 6754 3286 6774 3306 se
rect 6774 3286 6779 3306
rect 6563 3277 6566 3286
tri 6566 3277 6575 3286 nw
tri 6745 3277 6754 3286 se
rect 6754 3277 6779 3286
tri 6825 3306 6830 3311 sw
rect 6825 3292 6830 3306
tri 6830 3292 6844 3306 sw
rect 6825 3286 6844 3292
tri 6844 3286 6850 3292 sw
rect 11452 3291 12913 3292
rect 6825 3277 6850 3286
tri 6850 3277 6859 3286 sw
tri 6563 3274 6566 3277 nw
rect 8762 3259 8790 3287
rect 11452 3286 12100 3291
tri 3407 3196 3411 3200 se
rect 3411 3196 3493 3200
rect 3441 3170 3493 3196
rect 11452 3252 11464 3286
rect 11498 3252 11537 3286
rect 11571 3252 11610 3286
rect 11644 3252 11683 3286
rect 11717 3252 11756 3286
rect 11790 3252 11828 3286
rect 11862 3252 11900 3286
rect 11934 3252 11972 3286
rect 12006 3252 12044 3286
rect 12078 3252 12100 3286
rect 11452 3239 12100 3252
rect 12152 3239 12169 3291
rect 12221 3286 12238 3291
rect 12290 3286 12307 3291
rect 12359 3286 12376 3291
rect 12428 3286 12445 3291
rect 12497 3286 12514 3291
rect 12566 3286 12583 3291
rect 12635 3286 12651 3291
rect 12703 3286 12719 3291
rect 12222 3252 12238 3286
rect 12294 3252 12307 3286
rect 12366 3252 12376 3286
rect 12438 3252 12445 3286
rect 12703 3252 12712 3286
rect 12221 3239 12238 3252
rect 12290 3239 12307 3252
rect 12359 3239 12376 3252
rect 12428 3239 12445 3252
rect 12497 3239 12514 3252
rect 12566 3239 12583 3252
rect 12635 3239 12651 3252
rect 12703 3239 12719 3252
rect 12771 3239 12787 3291
rect 12839 3239 12855 3291
rect 12907 3239 12913 3291
rect 11452 3203 12913 3239
rect 11452 3170 12100 3203
rect 1789 3124 1817 3152
tri 3407 3142 3409 3144 ne
rect 3409 3142 3441 3144
tri 3409 3136 3415 3142 ne
rect 3415 3136 3441 3142
tri 3415 3131 3420 3136 ne
rect 3420 3131 3441 3136
rect 11452 3136 11464 3170
rect 11498 3136 11537 3170
rect 11571 3136 11610 3170
rect 11644 3136 11683 3170
rect 11717 3136 11756 3170
rect 11790 3136 11828 3170
rect 11862 3136 11900 3170
rect 11934 3136 11972 3170
rect 12006 3136 12044 3170
rect 12078 3151 12100 3170
rect 12152 3151 12169 3203
rect 12221 3170 12238 3203
rect 12290 3170 12307 3203
rect 12359 3170 12376 3203
rect 12428 3170 12445 3203
rect 12497 3194 12514 3203
rect 12566 3194 12583 3203
rect 12635 3194 12651 3203
rect 12703 3194 12719 3203
rect 12222 3151 12238 3170
rect 12294 3151 12307 3170
rect 12366 3151 12376 3170
rect 12438 3151 12445 3170
rect 12703 3160 12712 3194
rect 12497 3151 12514 3160
rect 12566 3151 12583 3160
rect 12635 3151 12651 3160
rect 12703 3151 12719 3160
rect 12771 3151 12787 3203
rect 12839 3151 12855 3203
rect 12907 3151 12913 3203
rect 12078 3136 12116 3151
rect 12150 3136 12188 3151
rect 12222 3136 12260 3151
rect 12294 3136 12332 3151
rect 12366 3136 12404 3151
rect 12438 3136 12913 3151
tri 3420 3128 3423 3131 ne
rect 3423 3128 3441 3131
tri 3423 3124 3427 3128 ne
rect 3427 3124 3441 3128
tri 3427 3112 3439 3124 ne
rect 3439 3112 3441 3124
tri 3439 3110 3441 3112 ne
rect 6592 3130 6615 3131
tri 6615 3130 6616 3131 nw
rect 11452 3130 12913 3136
rect 6592 3128 6613 3130
tri 6613 3128 6615 3130 nw
tri 12026 3128 12028 3130 ne
rect 12028 3128 12913 3130
rect 6592 3112 6597 3128
tri 6597 3112 6613 3128 nw
tri 12028 3112 12044 3128 ne
rect 12044 3115 12913 3128
rect 12044 3112 12100 3115
rect 6592 3110 6595 3112
tri 6595 3110 6597 3112 nw
tri 12044 3110 12046 3112 ne
rect 12046 3110 12100 3112
tri 6592 3107 6595 3110 nw
tri 12046 3107 12049 3110 ne
rect 12049 3107 12100 3110
tri 12049 3106 12050 3107 ne
rect 12050 3106 12100 3107
tri 12050 3102 12054 3106 ne
rect 12054 3102 12100 3106
tri 2691 3075 2718 3102 sw
tri 12054 3075 12081 3102 ne
rect 12081 3075 12100 3102
tri 1260 3068 1267 3075 sw
rect 2691 3068 2718 3075
tri 2718 3068 2725 3075 sw
tri 12081 3068 12088 3075 ne
rect 12088 3068 12100 3075
rect 1260 3063 1267 3068
tri 1267 3063 1272 3068 sw
tri 12088 3066 12090 3068 ne
rect 12090 3066 12100 3068
rect 1627 3064 1679 3066
tri 12090 3064 12092 3066 ne
rect 12092 3064 12100 3066
tri 12092 3063 12093 3064 ne
rect 12093 3063 12100 3064
rect 12152 3063 12169 3115
rect 12221 3063 12238 3115
rect 12290 3063 12307 3115
rect 12359 3063 12376 3115
rect 12428 3063 12445 3115
rect 12497 3102 12514 3115
rect 12566 3102 12583 3115
rect 12635 3102 12651 3115
rect 12703 3102 12719 3115
rect 12703 3068 12712 3102
rect 12497 3063 12514 3068
rect 12566 3063 12583 3068
rect 12635 3063 12651 3068
rect 12703 3063 12719 3068
rect 12771 3063 12787 3115
rect 12839 3063 12855 3115
rect 12907 3063 12913 3115
rect -618 2994 -616 3046
rect -257 3011 -255 3063
rect 1260 3062 1272 3063
tri 1272 3062 1273 3063 sw
tri 12093 3062 12094 3063 ne
rect 12094 3062 12913 3063
rect 1260 3055 1273 3062
tri 1273 3055 1280 3062 sw
rect 1260 3039 1280 3055
tri 1280 3039 1296 3055 sw
rect 2691 3039 2696 3040
tri 2696 3039 2697 3040 nw
rect 1260 3025 1296 3039
tri 1296 3025 1310 3039 sw
rect 2691 3038 2695 3039
tri 2695 3038 2696 3039 nw
rect 2318 3034 2370 3038
tri 2691 3034 2695 3038 nw
rect 1260 3024 1310 3025
tri 1310 3024 1311 3025 sw
tri 620 3016 628 3024 ne
rect 628 3016 644 3024
tri 628 3011 633 3016 ne
rect 633 3011 644 3016
tri 633 3007 637 3011 ne
rect 637 3007 644 3011
tri -194 2994 -181 3007 se
tri 637 3000 644 3007 ne
rect 695 3016 721 3024
tri 721 3016 729 3024 nw
rect 1260 3016 1311 3024
tri 1311 3016 1319 3024 sw
rect 695 3011 716 3016
tri 716 3011 721 3016 nw
rect 1260 3011 1319 3016
tri 1319 3011 1324 3016 sw
rect 695 3007 712 3011
tri 712 3007 716 3011 nw
rect 1260 3007 1324 3011
tri 1324 3007 1328 3011 sw
rect 695 3000 705 3007
tri 705 3000 712 3007 nw
tri -206 2982 -194 2994 se
rect -194 2982 -181 2994
tri 695 2990 705 3000 nw
rect 1260 2990 1328 3007
tri 1328 2990 1345 3007 sw
rect 1260 2989 1345 2990
tri 1345 2989 1346 2990 sw
tri 270 2986 273 2989 se
rect 1260 2986 1346 2989
tri 1346 2986 1349 2989 sw
rect 9018 2986 9400 2988
tri -215 2973 -206 2982 se
rect -206 2973 -181 2982
rect 1260 2982 1349 2986
tri 1349 2982 1353 2986 sw
rect 1260 2973 1353 2982
tri 1353 2973 1362 2982 sw
rect 1260 2966 1362 2973
tri 1362 2966 1369 2973 sw
rect 1260 2961 1369 2966
tri 1369 2961 1374 2966 sw
rect -493 2903 -476 2955
rect 4717 2941 4769 2947
tri 270 2937 273 2940 ne
rect 6886 2928 6914 2956
rect 9018 2934 9024 2986
rect 9076 2934 9104 2986
rect 9156 2934 9184 2986
rect 9236 2934 9263 2986
rect 9315 2934 9342 2986
rect 9394 2934 9400 2986
rect 9018 2910 9400 2934
rect 9018 2891 9024 2910
tri -651 2880 -649 2882 sw
rect -651 2848 -649 2880
tri -649 2848 -617 2880 sw
rect 4717 2877 4769 2889
tri 8956 2880 8967 2891 ne
rect 8967 2880 9024 2891
tri 8967 2846 9001 2880 ne
rect 9001 2858 9024 2880
rect 9076 2858 9104 2910
rect 9156 2858 9184 2910
rect 9236 2858 9263 2910
rect 9315 2858 9342 2910
rect 9394 2858 9400 2910
rect 9001 2846 9400 2858
tri 9001 2836 9011 2846 ne
rect 9011 2836 9400 2846
tri 9011 2829 9018 2836 ne
rect 9018 2834 9400 2836
rect 4717 2819 4769 2825
rect 1627 2799 1679 2801
rect 2318 2799 2370 2801
rect 9018 2782 9024 2834
rect 9076 2782 9104 2834
rect 9156 2782 9184 2834
rect 9236 2782 9263 2834
rect 9315 2782 9342 2834
rect 9394 2782 9400 2834
rect 3186 2747 3238 2766
rect 9018 2758 9400 2782
tri 3238 2747 3246 2755 sw
tri 3371 2747 3379 2755 se
rect 3186 2728 3246 2747
tri 3246 2728 3265 2747 sw
tri 3352 2728 3371 2747 se
rect 3371 2728 3379 2747
rect 3186 2721 3265 2728
tri 3265 2721 3272 2728 sw
tri 3345 2721 3352 2728 se
rect 3352 2721 3379 2728
rect 3186 2675 3238 2721
rect 9018 2706 9024 2758
rect 9076 2706 9104 2758
rect 9156 2706 9184 2758
rect 9236 2706 9263 2758
rect 9315 2706 9342 2758
rect 9394 2706 9400 2758
rect 9018 2704 9400 2706
rect 11552 2956 12364 2962
rect 11552 2904 11553 2956
rect 11605 2904 11623 2956
rect 11675 2904 11693 2956
rect 11750 2922 11792 2956
rect 11826 2922 11868 2956
rect 11902 2922 11943 2956
rect 11977 2922 12018 2956
rect 12052 2922 12093 2956
rect 12127 2922 12168 2956
rect 12202 2922 12243 2956
rect 12277 2922 12318 2956
rect 12352 2922 12364 2956
rect 11745 2904 12364 2922
rect 11552 2891 12364 2904
rect 11552 2839 11553 2891
rect 11605 2839 11623 2891
rect 11675 2839 11693 2891
rect 11745 2880 12364 2891
rect 11750 2846 11792 2880
rect 11826 2846 11868 2880
rect 11902 2846 11943 2880
rect 11977 2846 12018 2880
rect 12052 2846 12093 2880
rect 12127 2846 12168 2880
rect 12202 2846 12243 2880
rect 12277 2846 12318 2880
rect 12352 2846 12364 2880
rect 11745 2839 12364 2846
rect 11552 2826 12364 2839
rect 11552 2774 11553 2826
rect 11605 2774 11623 2826
rect 11675 2774 11693 2826
rect 11745 2804 12364 2826
rect 11552 2770 11564 2774
rect 11598 2770 11640 2774
rect 11674 2770 11716 2774
rect 11750 2770 11792 2804
rect 11826 2770 11868 2804
rect 11902 2770 11943 2804
rect 11977 2770 12018 2804
rect 12052 2770 12093 2804
rect 12127 2770 12168 2804
rect 12202 2770 12243 2804
rect 12277 2770 12318 2804
rect 12352 2770 12364 2804
rect 11552 2761 12364 2770
rect 11552 2709 11553 2761
rect 11605 2709 11623 2761
rect 11675 2709 11693 2761
rect 11745 2728 12364 2761
rect 11552 2696 11564 2709
rect 11598 2696 11640 2709
rect 11674 2696 11716 2709
rect 4229 2675 4249 2689
tri 4249 2675 4263 2689 nw
tri 2771 2673 2773 2675 se
rect 1973 2671 2025 2673
rect 2639 2671 2691 2673
tri 2769 2671 2771 2673 se
rect 2771 2671 2773 2673
tri 2756 2658 2769 2671 se
rect 2769 2658 2773 2671
tri 2750 2652 2756 2658 se
rect 2756 2652 2773 2658
rect 4229 2658 4232 2675
tri 4232 2658 4249 2675 nw
tri 4229 2655 4232 2658 nw
tri 2741 2643 2750 2652 se
rect 2750 2643 2773 2652
rect 11552 2644 11553 2696
rect 11605 2644 11623 2696
rect 11675 2644 11693 2696
rect 11750 2694 11792 2728
rect 11826 2694 11868 2728
rect 11902 2694 11943 2728
rect 11977 2694 12018 2728
rect 12052 2694 12093 2728
rect 12127 2694 12168 2728
rect 12202 2694 12243 2728
rect 12277 2694 12318 2728
rect 12352 2694 12364 2728
rect 11745 2652 12364 2694
rect 11552 2631 11564 2644
rect 11598 2631 11640 2644
rect 11674 2631 11716 2644
rect 6754 2593 6782 2621
rect 8762 2572 8790 2600
rect 11552 2579 11553 2631
rect 11605 2579 11623 2631
rect 11675 2579 11693 2631
rect 11750 2618 11792 2652
rect 11826 2618 11868 2652
rect 11902 2618 11943 2652
rect 11977 2618 12018 2652
rect 12052 2618 12093 2652
rect 12127 2618 12168 2652
rect 12202 2618 12243 2652
rect 12277 2618 12318 2652
rect 12352 2618 12364 2652
rect 11745 2579 12364 2618
rect 11552 2576 12364 2579
rect 11552 2566 11564 2576
rect 11598 2566 11640 2576
rect 11674 2566 11716 2576
rect 11552 2514 11553 2566
rect 11605 2514 11623 2566
rect 11675 2514 11693 2566
rect 11750 2542 11792 2576
rect 11826 2542 11868 2576
rect 11902 2542 11943 2576
rect 11977 2542 12018 2576
rect 12052 2542 12093 2576
rect 12127 2542 12168 2576
rect 12202 2542 12243 2576
rect 12277 2542 12318 2576
rect 12352 2542 12364 2576
tri 13105 2544 13113 2552 se
rect 13113 2544 13165 3398
rect 11745 2514 12364 2542
tri 13100 2539 13105 2544 se
rect 13105 2539 13165 2544
tri 13077 2516 13100 2539 se
rect 13100 2516 13165 2539
rect 328 2480 356 2508
rect 11552 2500 12364 2514
tri 13066 2505 13077 2516 se
rect 13077 2505 13165 2516
rect 11552 2448 11553 2500
rect 11605 2448 11623 2500
rect 11675 2448 11693 2500
rect 11750 2466 11792 2500
rect 11826 2466 11868 2500
rect 11902 2466 11943 2500
rect 11977 2466 12018 2500
rect 12052 2466 12093 2500
rect 12127 2466 12168 2500
rect 12202 2466 12243 2500
rect 12277 2466 12318 2500
rect 12352 2466 12364 2500
tri 13053 2492 13066 2505 se
rect 13066 2492 13165 2505
rect 11745 2448 12364 2466
rect 11552 2434 12364 2448
rect 11552 2382 11553 2434
rect 11605 2382 11623 2434
rect 11675 2382 11693 2434
rect 11745 2424 12364 2434
rect 11750 2390 11792 2424
rect 11826 2390 11868 2424
rect 11902 2390 11943 2424
rect 11977 2390 12018 2424
rect 12052 2390 12093 2424
rect 12127 2390 12168 2424
rect 12202 2390 12243 2424
rect 12277 2390 12318 2424
rect 12352 2390 12364 2424
rect 11745 2382 12364 2390
tri 2748 2358 2754 2364 se
rect 2754 2358 2755 2364
rect 11552 2348 12364 2382
rect 4171 2261 4177 2313
rect 4229 2261 4241 2313
rect 4293 2261 5144 2313
rect 5196 2261 5208 2313
rect 5260 2261 5266 2313
rect 7595 2300 7862 2323
rect 7595 2248 7601 2300
rect 7653 2248 7703 2300
rect 7755 2248 7804 2300
rect 7856 2248 7862 2300
rect 9490 2313 9522 2318
rect 11552 2314 11564 2348
rect 11598 2314 11640 2348
rect 11674 2314 11716 2348
rect 11750 2314 11792 2348
rect 11826 2314 11868 2348
rect 11902 2314 11943 2348
rect 11977 2314 12018 2348
rect 12052 2314 12093 2348
rect 12127 2314 12168 2348
rect 12202 2314 12243 2348
rect 12277 2314 12318 2348
rect 12352 2314 12364 2348
rect 12453 2486 13165 2492
rect 12453 2452 12465 2486
rect 12499 2452 12539 2486
rect 12573 2452 12613 2486
rect 12647 2452 12687 2486
rect 12721 2452 12761 2486
rect 12795 2452 12835 2486
rect 12869 2452 13165 2486
rect 12453 2378 13165 2452
rect 12453 2370 13146 2378
rect 12453 2336 12465 2370
rect 12499 2336 12539 2370
rect 12573 2336 12613 2370
rect 12647 2336 12687 2370
rect 12721 2336 12761 2370
rect 12795 2336 12835 2370
rect 12869 2359 13146 2370
tri 13146 2359 13165 2378 nw
rect 13199 3488 13205 3522
rect 13239 3488 13245 3522
rect 13199 3450 13245 3488
rect 13199 3416 13205 3450
rect 13239 3416 13245 3450
rect 13199 3378 13245 3416
rect 13199 3344 13205 3378
rect 13239 3344 13245 3378
rect 13199 3306 13245 3344
rect 13199 3272 13205 3306
rect 13239 3272 13245 3306
rect 13199 3234 13245 3272
rect 13199 3200 13205 3234
rect 13239 3200 13245 3234
rect 13431 4000 13437 4007
rect 13471 4007 13480 4013
rect 13471 4000 13477 4007
tri 13477 4004 13480 4007 nw
rect 13431 3961 13477 4000
rect 13772 4023 13778 4027
tri 13778 4023 13806 4051 nw
rect 13772 4022 13777 4023
tri 13777 4022 13778 4023 nw
tri 13923 4022 13924 4023 se
rect 13924 4022 14606 4023
tri 14606 4022 14607 4023 sw
rect 14977 4022 15023 4061
tri 13772 4017 13777 4022 nw
tri 13918 4017 13923 4022 se
rect 13923 4017 14607 4022
tri 13912 4011 13918 4017 se
rect 13918 4011 14607 4017
tri 14607 4011 14618 4022 sw
tri 13889 3988 13912 4011 se
rect 13912 3988 14618 4011
tri 14618 3988 14641 4011 sw
rect 14977 3988 14983 4022
rect 15017 3988 15023 4022
tri 13881 3980 13889 3988 se
rect 13889 3980 14641 3988
tri 14641 3980 14649 3988 sw
rect 13720 3969 13772 3975
tri 13870 3969 13881 3980 se
rect 13881 3969 13944 3980
tri 13944 3969 13955 3980 nw
tri 14589 3969 14600 3980 ne
rect 14600 3969 14649 3980
rect 13431 3927 13437 3961
rect 13471 3927 13477 3961
tri 13850 3949 13870 3969 se
rect 13870 3949 13924 3969
tri 13924 3949 13944 3969 nw
tri 14600 3952 14617 3969 ne
rect 14617 3967 14649 3969
tri 14649 3967 14662 3980 sw
rect 14617 3952 14662 3967
tri 13846 3945 13850 3949 se
rect 13850 3945 13920 3949
tri 13920 3945 13924 3949 nw
tri 13841 3940 13846 3945 se
rect 13846 3940 13920 3945
tri 13839 3938 13841 3940 se
rect 13841 3938 13920 3940
tri 13829 3928 13839 3938 se
rect 13839 3928 13920 3938
rect 13431 3888 13477 3927
rect 13431 3854 13437 3888
rect 13471 3854 13477 3888
rect 13431 3815 13477 3854
rect 13431 3781 13437 3815
rect 13471 3781 13477 3815
rect 13549 3922 13601 3928
rect 13549 3858 13601 3870
rect 13549 3800 13601 3806
tri 13549 3797 13552 3800 ne
rect 13431 3742 13477 3781
rect 13431 3708 13437 3742
rect 13471 3708 13477 3742
rect 13552 3767 13598 3800
tri 13598 3797 13601 3800 nw
rect 13708 3922 13920 3928
rect 13708 3916 13868 3922
rect 13708 3882 13714 3916
rect 13748 3882 13868 3916
rect 13708 3870 13868 3882
rect 13708 3851 13920 3870
rect 13708 3842 13868 3851
rect 13708 3808 13714 3842
rect 13748 3808 13868 3842
rect 13708 3799 13868 3808
rect 13552 3733 13558 3767
rect 13592 3733 13598 3767
rect 13708 3780 13920 3799
rect 13708 3767 13868 3780
tri 13677 3733 13708 3764 se
rect 13708 3733 13714 3767
rect 13748 3733 13868 3767
rect 13552 3721 13598 3733
tri 13669 3725 13677 3733 se
rect 13677 3728 13868 3733
rect 13677 3725 13920 3728
tri 13665 3721 13669 3725 se
rect 13669 3721 13920 3725
rect 13980 3944 14035 3950
rect 13980 3892 13983 3944
rect 13980 3880 14035 3892
rect 13980 3828 13983 3880
rect 13980 3816 14035 3828
rect 13980 3764 13983 3816
rect 13980 3758 14035 3764
rect 13980 3753 14030 3758
tri 14030 3753 14035 3758 nw
rect 14063 3944 14115 3950
rect 14063 3855 14115 3892
rect 14143 3946 14574 3952
tri 14617 3951 14618 3952 ne
rect 14195 3940 14574 3946
rect 14195 3906 14534 3940
rect 14568 3906 14574 3940
rect 14195 3894 14574 3906
rect 14143 3868 14574 3894
rect 14195 3861 14574 3868
rect 14195 3827 14534 3861
rect 14568 3827 14574 3861
rect 14195 3816 14574 3827
rect 14143 3810 14574 3816
tri 14452 3803 14459 3810 ne
rect 14459 3803 14574 3810
rect 14063 3765 14115 3803
tri 14459 3781 14481 3803 ne
rect 14481 3781 14574 3803
tri 14481 3779 14483 3781 ne
rect 14483 3779 14534 3781
tri 13663 3719 13665 3721 se
rect 13665 3719 13729 3721
tri 13729 3719 13731 3721 nw
tri 13653 3709 13663 3719 se
rect 13663 3709 13719 3719
tri 13719 3709 13729 3719 nw
rect 13431 3669 13477 3708
tri 13645 3701 13653 3709 se
rect 13653 3707 13717 3709
tri 13717 3707 13719 3709 nw
rect 13653 3701 13711 3707
tri 13711 3701 13717 3707 nw
tri 13622 3678 13645 3701 se
rect 13645 3678 13688 3701
tri 13688 3678 13711 3701 nw
tri 13977 3684 13980 3687 se
rect 13980 3684 14026 3753
tri 14026 3749 14030 3753 nw
tri 13616 3672 13622 3678 se
rect 13622 3672 13682 3678
tri 13682 3672 13688 3678 nw
rect 13431 3635 13437 3669
rect 13471 3635 13477 3669
tri 13603 3659 13616 3672 se
rect 13616 3659 13669 3672
tri 13669 3659 13682 3672 nw
tri 13601 3657 13603 3659 se
rect 13603 3657 13667 3659
tri 13667 3657 13669 3659 nw
tri 13588 3644 13601 3657 se
rect 13601 3644 13654 3657
tri 13654 3644 13667 3657 nw
tri 13582 3638 13588 3644 se
rect 13588 3638 13648 3644
tri 13648 3638 13654 3644 nw
rect 13431 3596 13477 3635
tri 13567 3623 13582 3638 se
rect 13582 3623 13633 3638
tri 13633 3623 13648 3638 nw
rect 13742 3632 13748 3684
rect 13800 3632 13812 3684
rect 13864 3632 13870 3684
tri 13971 3678 13977 3684 se
rect 13977 3678 14026 3684
tri 13960 3667 13971 3678 se
rect 13971 3667 14026 3678
tri 13742 3623 13751 3632 ne
rect 13751 3623 13870 3632
tri 13565 3621 13567 3623 se
rect 13567 3621 13631 3623
tri 13631 3621 13633 3623 nw
tri 13751 3621 13753 3623 ne
rect 13753 3621 13870 3623
rect 13431 3562 13437 3596
rect 13471 3562 13477 3596
rect 13431 3523 13477 3562
rect 13431 3489 13437 3523
rect 13471 3489 13477 3523
rect 13431 3450 13477 3489
rect 13431 3416 13437 3450
rect 13471 3416 13477 3450
rect 13431 3376 13477 3416
rect 13431 3342 13437 3376
rect 13471 3342 13477 3376
rect 13431 3302 13477 3342
rect 13431 3268 13437 3302
rect 13471 3268 13477 3302
rect 13431 3230 13477 3268
tri 13557 3613 13565 3621 se
rect 13565 3613 13614 3621
rect 13557 3604 13614 3613
tri 13614 3604 13631 3621 nw
tri 13753 3604 13770 3621 ne
rect 13770 3604 13870 3621
rect 13557 3597 13607 3604
tri 13607 3597 13614 3604 nw
tri 13770 3597 13777 3604 ne
rect 13777 3597 13870 3604
rect 13557 3364 13603 3597
tri 13603 3593 13607 3597 nw
tri 13777 3593 13781 3597 ne
rect 13781 3593 13830 3597
tri 13781 3563 13811 3593 ne
rect 13811 3563 13830 3593
rect 13864 3563 13870 3597
tri 13811 3550 13824 3563 ne
rect 13824 3521 13870 3563
rect 13824 3487 13830 3521
rect 13864 3487 13870 3521
rect 13824 3445 13870 3487
rect 13824 3411 13830 3445
rect 13864 3411 13870 3445
rect 13824 3399 13870 3411
tri 13954 3661 13960 3667 se
rect 13960 3661 14018 3667
rect 13954 3659 14018 3661
tri 14018 3659 14026 3667 nw
rect 13954 3657 14016 3659
tri 14016 3657 14018 3659 nw
rect 13954 3644 14003 3657
tri 14003 3644 14016 3657 nw
tri 13951 3404 13954 3407 se
rect 13954 3404 14000 3644
tri 14000 3641 14003 3644 nw
tri 14060 3641 14063 3644 se
rect 14063 3641 14115 3713
rect 14143 3773 14418 3779
rect 14195 3733 14418 3773
tri 14483 3747 14515 3779 ne
rect 14515 3747 14534 3779
rect 14568 3747 14574 3781
tri 14515 3734 14528 3747 ne
rect 14195 3730 14226 3733
tri 14226 3730 14229 3733 nw
tri 14338 3730 14341 3733 ne
rect 14341 3730 14418 3733
rect 14195 3721 14217 3730
tri 14217 3721 14226 3730 nw
tri 14341 3721 14350 3730 ne
rect 14350 3721 14418 3730
rect 14143 3709 14205 3721
tri 14205 3709 14217 3721 nw
tri 14350 3709 14362 3721 ne
rect 14362 3709 14418 3721
rect 14195 3707 14203 3709
tri 14203 3707 14205 3709 nw
tri 14362 3707 14364 3709 ne
rect 14364 3707 14418 3709
rect 14195 3701 14197 3707
tri 14197 3701 14203 3707 nw
tri 14364 3701 14370 3707 ne
rect 14370 3701 14418 3707
tri 14195 3699 14197 3701 nw
tri 14370 3699 14372 3701 ne
rect 14143 3651 14195 3657
rect 14256 3678 14302 3690
tri 14250 3644 14256 3650 se
rect 14256 3644 14262 3678
rect 14296 3644 14302 3678
tri 14047 3628 14060 3641 se
rect 14060 3628 14115 3641
rect 14047 3622 14115 3628
tri 14229 3623 14250 3644 se
rect 14250 3623 14302 3644
rect 14047 3621 14114 3622
tri 14114 3621 14115 3622 nw
tri 14227 3621 14229 3623 se
rect 14229 3621 14302 3623
tri 14000 3404 14008 3412 sw
rect 14047 3408 14099 3621
tri 14099 3606 14114 3621 nw
tri 14212 3606 14227 3621 se
rect 14227 3606 14302 3621
tri 14193 3587 14212 3606 se
rect 14212 3587 14302 3606
tri 14190 3584 14193 3587 se
rect 14193 3584 14302 3587
tri 14188 3582 14190 3584 se
rect 14190 3582 14302 3584
tri 14175 3569 14188 3582 se
rect 14188 3569 14262 3582
rect 14135 3563 14262 3569
rect 14187 3548 14262 3563
rect 14296 3548 14302 3582
rect 14187 3511 14302 3548
rect 14135 3499 14302 3511
rect 14187 3486 14302 3499
rect 14187 3452 14262 3486
rect 14296 3452 14302 3486
rect 14187 3447 14302 3452
rect 14135 3440 14302 3447
rect 14372 3678 14418 3701
rect 14372 3644 14378 3678
rect 14412 3644 14418 3678
rect 14372 3582 14418 3644
rect 14372 3548 14378 3582
rect 14412 3548 14418 3582
rect 14372 3486 14418 3548
rect 14372 3452 14378 3486
rect 14412 3452 14418 3486
rect 14528 3701 14574 3747
rect 14528 3667 14534 3701
rect 14568 3667 14574 3701
rect 14528 3621 14574 3667
rect 14528 3587 14534 3621
rect 14568 3587 14574 3621
rect 14528 3541 14574 3587
rect 14528 3507 14534 3541
rect 14568 3507 14574 3541
tri 14524 3477 14528 3481 se
rect 14528 3477 14574 3507
rect 14372 3440 14418 3452
tri 14487 3440 14524 3477 se
rect 14524 3461 14574 3477
rect 14524 3440 14551 3461
tri 14485 3438 14487 3440 se
rect 14487 3438 14551 3440
tri 14551 3438 14574 3461 nw
tri 14483 3436 14485 3438 se
rect 14485 3436 14534 3438
tri 14099 3408 14127 3436 sw
tri 14468 3421 14483 3436 se
rect 14483 3421 14534 3436
tri 14534 3421 14551 3438 nw
rect 14468 3413 14526 3421
tri 14526 3413 14534 3421 nw
rect 14468 3408 14521 3413
tri 14521 3408 14526 3413 nw
tri 14613 3408 14618 3413 se
rect 14618 3408 14662 3952
tri 14047 3404 14051 3408 ne
rect 14051 3404 14127 3408
tri 14127 3404 14131 3408 sw
rect 14468 3404 14517 3408
tri 14517 3404 14521 3408 nw
tri 14609 3404 14613 3408 se
rect 14613 3404 14662 3408
tri 13946 3399 13951 3404 se
rect 13951 3399 14008 3404
tri 13923 3376 13946 3399 se
rect 13946 3388 14008 3399
tri 14008 3388 14024 3404 sw
tri 14051 3388 14067 3404 ne
rect 14067 3388 14131 3404
tri 14131 3388 14147 3404 sw
rect 13946 3376 14024 3388
tri 14024 3376 14036 3388 sw
rect 13557 3330 13563 3364
rect 13597 3330 13603 3364
rect 13909 3370 14039 3376
rect 13909 3336 13921 3370
rect 13955 3336 13993 3370
rect 14027 3336 14039 3370
rect 14067 3336 14073 3388
rect 14125 3336 14137 3388
rect 14189 3336 14195 3388
rect 13909 3330 14039 3336
rect 13557 3292 13603 3330
rect 13557 3258 13563 3292
rect 13597 3258 13603 3292
rect 13557 3246 13603 3258
rect 13707 3296 14425 3302
rect 13707 3284 13875 3296
rect 13707 3250 13719 3284
rect 13753 3250 13835 3284
rect 13869 3250 13875 3284
rect 13707 3244 13875 3250
rect 13927 3284 14425 3296
rect 13927 3250 14263 3284
rect 14297 3250 14379 3284
rect 14413 3250 14425 3284
rect 13927 3244 14425 3250
rect 13707 3232 14425 3244
tri 13813 3230 13815 3232 ne
rect 13815 3230 13973 3232
tri 13815 3218 13827 3230 ne
rect 13827 3218 13973 3230
tri 13973 3218 13987 3232 nw
tri 13827 3201 13844 3218 ne
rect 13844 3206 13961 3218
tri 13961 3206 13973 3218 nw
rect 13844 3204 13956 3206
rect 13844 3201 13875 3204
rect 13199 3162 13245 3200
rect 13199 3128 13205 3162
rect 13239 3128 13245 3162
rect 13437 3149 13443 3201
rect 13495 3149 13507 3201
rect 13559 3195 13797 3201
tri 13844 3198 13847 3201 ne
rect 13559 3161 13617 3195
rect 13651 3161 13751 3195
rect 13785 3161 13797 3195
rect 13559 3155 13797 3161
tri 13844 3155 13847 3158 se
rect 13847 3155 13875 3201
rect 13559 3149 13565 3155
tri 13565 3149 13571 3155 nw
tri 13838 3149 13844 3155 se
rect 13844 3152 13875 3155
rect 13927 3201 13956 3204
tri 13956 3201 13961 3206 nw
rect 13927 3155 13953 3201
tri 13953 3198 13956 3201 nw
tri 13953 3155 13956 3158 sw
rect 13927 3152 13956 3155
rect 13844 3149 13956 3152
tri 13956 3149 13962 3155 sw
rect 14011 3152 14017 3204
rect 14069 3152 14081 3204
rect 14133 3195 14424 3204
rect 14148 3161 14202 3195
rect 14236 3161 14290 3195
rect 14324 3161 14378 3195
rect 14412 3161 14424 3195
rect 14133 3152 14424 3161
tri 13835 3146 13838 3149 se
rect 13838 3146 13962 3149
tri 13962 3146 13965 3149 sw
rect 13199 3089 13245 3128
tri 13813 3124 13835 3146 se
rect 13835 3124 13965 3146
tri 13965 3124 13987 3146 sw
rect 13707 3112 14425 3124
rect 13199 3055 13205 3089
rect 13239 3055 13245 3089
rect 13199 3016 13245 3055
rect 13199 2982 13205 3016
rect 13239 2982 13245 3016
rect 13199 2943 13245 2982
rect 13557 3097 13603 3109
rect 13557 3063 13563 3097
rect 13597 3063 13603 3097
rect 13557 3025 13603 3063
rect 13707 3106 13875 3112
rect 13707 3072 13719 3106
rect 13753 3072 13835 3106
rect 13869 3072 13875 3106
rect 13707 3060 13875 3072
rect 13927 3106 14425 3112
rect 13927 3072 14263 3106
rect 14297 3072 14379 3106
rect 14413 3072 14425 3106
rect 13927 3060 14425 3072
rect 13707 3054 14425 3060
rect 14468 3094 14514 3404
tri 14514 3401 14517 3404 nw
tri 14606 3401 14609 3404 se
rect 14609 3401 14662 3404
tri 14593 3388 14606 3401 se
rect 14606 3388 14662 3401
tri 14570 3365 14593 3388 se
rect 14593 3383 14662 3388
rect 14593 3365 14644 3383
tri 14644 3365 14662 3383 nw
rect 14977 3949 15023 3988
rect 14977 3915 14983 3949
rect 15017 3915 15023 3949
rect 14977 3876 15023 3915
rect 14977 3842 14983 3876
rect 15017 3842 15023 3876
rect 14977 3803 15023 3842
rect 14977 3769 14983 3803
rect 15017 3769 15023 3803
rect 14977 3730 15023 3769
rect 14977 3696 14983 3730
rect 15017 3696 15023 3730
rect 14977 3657 15023 3696
rect 14977 3623 14983 3657
rect 15017 3623 15023 3657
rect 14977 3584 15023 3623
rect 14977 3550 14983 3584
rect 15017 3550 15023 3584
rect 14977 3511 15023 3550
rect 14977 3477 14983 3511
rect 15017 3477 15023 3511
rect 14977 3438 15023 3477
rect 14977 3404 14983 3438
rect 15017 3404 15023 3438
rect 14977 3365 15023 3404
tri 14550 3345 14570 3365 se
rect 14570 3345 14624 3365
tri 14624 3345 14644 3365 nw
rect 14550 3336 14615 3345
tri 14615 3336 14624 3345 nw
rect 14550 3331 14610 3336
tri 14610 3331 14615 3336 nw
rect 14977 3331 14983 3365
rect 15017 3331 15023 3365
rect 14550 3324 14596 3331
rect 14550 3290 14556 3324
rect 14590 3290 14596 3324
tri 14596 3317 14610 3331 nw
rect 14550 3252 14596 3290
rect 14550 3218 14556 3252
rect 14590 3218 14596 3252
rect 14550 3206 14596 3218
rect 14977 3292 15023 3331
rect 14977 3258 14983 3292
rect 15017 3258 15023 3292
rect 14977 3219 15023 3258
rect 14468 3060 14474 3094
rect 14508 3060 14514 3094
rect 13557 2991 13563 3025
rect 13597 2991 13603 3025
rect 13557 2973 13603 2991
rect 13979 3016 14073 3025
rect 14125 3016 14137 3025
rect 13979 2982 13991 3016
rect 14025 2982 14073 3016
tri 13603 2973 13607 2977 sw
rect 13979 2973 14073 2982
rect 14125 2973 14137 2982
rect 14189 2973 14195 3025
rect 14468 3022 14514 3060
rect 14468 2988 14474 3022
rect 14508 2988 14514 3022
rect 13557 2966 13607 2973
tri 13607 2966 13614 2973 sw
tri 14461 2966 14468 2973 se
rect 14468 2966 14514 2988
rect 13557 2961 13614 2966
tri 13614 2961 13619 2966 sw
tri 14456 2961 14461 2966 se
rect 14461 2961 14514 2966
rect 13557 2957 13619 2961
tri 13619 2957 13623 2961 sw
tri 14452 2957 14456 2961 se
rect 14456 2957 14514 2961
tri 13557 2955 13559 2957 ne
rect 13559 2955 13623 2957
tri 13559 2947 13567 2955 ne
rect 13567 2953 13623 2955
tri 13623 2953 13627 2957 sw
tri 14448 2953 14452 2957 se
rect 14452 2953 14514 2957
rect 13567 2947 13627 2953
rect 13199 2909 13205 2943
rect 13239 2909 13245 2943
tri 13567 2927 13587 2947 ne
rect 13587 2945 13627 2947
tri 13627 2945 13635 2953 sw
tri 14440 2945 14448 2953 se
rect 14448 2945 14488 2953
rect 13587 2927 14488 2945
tri 14488 2927 14514 2953 nw
rect 14977 3185 14983 3219
rect 15017 3185 15023 3219
rect 14977 3146 15023 3185
rect 14977 3112 14983 3146
rect 15017 3112 15023 3146
rect 14977 3073 15023 3112
rect 14977 3039 14983 3073
rect 15017 3039 15023 3073
rect 14977 3000 15023 3039
rect 14977 2966 14983 3000
rect 15017 2966 15023 3000
rect 14977 2927 15023 2966
tri 13587 2917 13597 2927 ne
rect 13597 2917 14478 2927
tri 14478 2917 14488 2927 nw
rect 13199 2893 13245 2909
tri 13245 2893 13269 2917 sw
tri 13597 2911 13603 2917 ne
rect 13603 2911 14472 2917
tri 14472 2911 14478 2917 nw
tri 14971 2911 14977 2917 se
rect 14977 2911 14983 2927
tri 14953 2893 14971 2911 se
rect 14971 2893 14983 2911
rect 15017 2893 15023 2927
rect 13199 2883 13269 2893
tri 13269 2883 13279 2893 sw
tri 14943 2883 14953 2893 se
rect 14953 2883 15023 2893
rect 13199 2877 15023 2883
rect 13199 2870 13277 2877
rect 13199 2836 13205 2870
rect 13239 2843 13277 2870
rect 13311 2843 13352 2877
rect 13386 2843 13427 2877
rect 13461 2843 13502 2877
rect 13536 2843 13577 2877
rect 13611 2843 13652 2877
rect 13686 2843 13727 2877
rect 13761 2843 13801 2877
rect 13835 2843 13875 2877
rect 13909 2843 13949 2877
rect 13983 2843 14023 2877
rect 14057 2843 14097 2877
rect 14131 2843 14171 2877
rect 14205 2843 14245 2877
rect 14279 2843 14319 2877
rect 14353 2843 14393 2877
rect 14427 2843 14467 2877
rect 14501 2843 14541 2877
rect 14575 2843 14615 2877
rect 14649 2843 14689 2877
rect 14723 2843 14763 2877
rect 14797 2843 14837 2877
rect 14871 2843 14911 2877
rect 14945 2854 15023 2877
rect 14945 2843 14983 2854
rect 13239 2837 14983 2843
rect 13239 2836 13262 2837
rect 13199 2820 13262 2836
tri 13262 2820 13279 2837 nw
tri 14943 2820 14960 2837 ne
rect 14960 2820 14983 2837
rect 15017 2820 15023 2854
rect 13199 2819 13261 2820
tri 13261 2819 13262 2820 nw
tri 14960 2819 14961 2820 ne
rect 14961 2819 15023 2820
rect 13199 2797 13245 2819
tri 13245 2803 13261 2819 nw
tri 14961 2803 14977 2819 ne
tri 13348 2799 13349 2800 se
rect 13349 2799 13908 2800
rect 13199 2763 13205 2797
rect 13239 2763 13245 2797
tri 13330 2781 13348 2799 se
rect 13348 2781 13908 2799
tri 13315 2766 13330 2781 se
rect 13330 2766 13908 2781
rect 13199 2724 13245 2763
tri 13304 2755 13315 2766 se
rect 13315 2755 13908 2766
tri 13296 2747 13304 2755 se
rect 13304 2748 13908 2755
rect 13960 2748 13972 2800
rect 14024 2748 14030 2800
rect 14977 2781 15023 2819
rect 13304 2747 13370 2748
tri 13370 2747 13371 2748 nw
rect 14977 2747 14983 2781
rect 15017 2747 15023 2781
rect 13199 2690 13205 2724
rect 13239 2690 13245 2724
rect 13199 2651 13245 2690
rect 13199 2617 13205 2651
rect 13239 2617 13245 2651
rect 13199 2578 13245 2617
rect 13199 2544 13205 2578
rect 13239 2544 13245 2578
rect 13199 2505 13245 2544
rect 13199 2471 13205 2505
rect 13239 2471 13245 2505
rect 13199 2432 13245 2471
rect 13199 2398 13205 2432
rect 13239 2398 13245 2432
rect 13199 2359 13245 2398
rect 12869 2336 13117 2359
rect 12453 2330 13117 2336
tri 13117 2330 13146 2359 nw
rect 7595 2225 7862 2248
rect 9090 2278 9280 2293
rect 9090 2226 9091 2278
rect 9143 2226 9159 2278
rect 9211 2226 9227 2278
rect 9279 2226 9280 2278
tri 8875 2213 8880 2218 se
tri 8854 2192 8875 2213 se
rect 8875 2192 8880 2213
tri 9075 2192 9090 2207 se
rect 9090 2193 9280 2226
rect 9090 2192 9091 2193
tri 9073 2190 9075 2192 se
rect 9075 2190 9091 2192
tri 9062 2179 9073 2190 se
rect 9073 2179 9091 2190
tri 9059 2176 9062 2179 se
rect 9062 2176 9091 2179
tri 9049 2166 9059 2176 se
rect 9059 2166 9091 2176
tri 9023 2140 9049 2166 se
rect 9049 2141 9091 2166
rect 9143 2141 9159 2193
rect 9211 2141 9227 2193
rect 9279 2141 9280 2193
rect 9490 2261 9496 2313
rect 9548 2261 9582 2313
rect 9634 2261 9640 2313
rect 9490 2249 9640 2261
rect 9490 2197 9496 2249
rect 9548 2197 9582 2249
rect 9634 2197 9640 2249
rect 11552 2272 12364 2314
rect 11552 2238 11564 2272
rect 11598 2238 11640 2272
rect 11674 2238 11716 2272
rect 11750 2238 11792 2272
rect 11826 2238 11868 2272
rect 11902 2238 11943 2272
rect 11977 2238 12018 2272
rect 12052 2238 12093 2272
rect 12127 2238 12168 2272
rect 12202 2238 12243 2272
rect 12277 2238 12318 2272
rect 12352 2238 12364 2272
rect 11552 2232 12364 2238
rect 13199 2325 13205 2359
rect 13239 2325 13245 2359
rect 13199 2286 13245 2325
rect 13199 2252 13205 2286
rect 13239 2252 13245 2286
rect 13199 2213 13245 2252
rect 9490 2190 9522 2197
rect 9049 2140 9280 2141
tri 9008 2125 9023 2140 se
rect 9023 2125 9280 2140
rect 13199 2179 13205 2213
rect 13239 2179 13245 2213
rect 13199 2140 13245 2179
tri 9004 2121 9008 2125 se
rect 9008 2121 9280 2125
tri 4366 2106 4381 2121 se
rect 4381 2106 5267 2121
tri 4365 2105 4366 2106 se
rect 4366 2105 5267 2106
tri 4354 2094 4365 2105 se
rect 4365 2094 5267 2105
tri 4335 2075 4354 2094 se
rect 4354 2075 5267 2094
rect 8924 2119 9280 2121
tri 9817 2119 9823 2125 sw
rect 8924 2075 9068 2119
rect 9090 2107 9280 2119
tri 4327 2067 4335 2075 se
rect 4335 2067 5267 2075
tri 4293 2033 4327 2067 se
rect 4327 2033 5267 2067
rect 9090 2055 9091 2107
rect 9143 2055 9159 2107
rect 9211 2055 9227 2107
rect 9279 2055 9280 2107
rect 9090 2049 9280 2055
tri 4288 2028 4293 2033 se
rect 4293 2028 5267 2033
tri 4281 2021 4288 2028 se
rect 4288 2021 4397 2028
tri 4397 2021 4404 2028 nw
tri 5155 2021 5162 2028 ne
rect 5162 2021 5267 2028
tri 4278 2018 4281 2021 se
rect 4281 2018 4394 2021
tri 4394 2018 4397 2021 nw
tri 5162 2018 5165 2021 ne
rect 5165 2018 5267 2021
rect 3715 2012 3767 2018
tri 1495 1935 1502 1942 ne
rect 1502 1935 1507 1942
rect 2542 1936 3270 1988
rect 3322 1936 3388 1988
rect 3440 1936 3446 1988
rect 2542 1910 3446 1936
rect 2542 1858 3270 1910
rect 3322 1858 3388 1910
rect 3440 1858 3446 1910
rect 3715 1948 3767 1960
rect 1940 1748 1968 1776
rect -225 1614 -197 1642
tri 2095 1410 2098 1413 se
tri 2087 1402 2095 1410 se
rect 2095 1402 2098 1410
tri 2090 1367 2098 1375 ne
rect 2098 1367 2108 1375
rect 2154 1374 2182 1402
rect 2516 1361 2525 1413
rect 2862 1364 2864 1416
tri -977 1230 -949 1258 sw
rect -977 1228 -949 1230
tri -949 1228 -947 1230 sw
rect -977 1224 -947 1228
tri -947 1224 -943 1228 sw
rect -317 1125 217 1224
rect -311 1118 -259 1125
tri -259 1118 -252 1125 nw
rect -311 1084 -293 1118
tri -293 1084 -259 1118 nw
rect -311 1082 -295 1084
tri -295 1082 -293 1084 nw
rect -311 1080 -297 1082
tri -297 1080 -295 1082 nw
rect -311 1073 -304 1080
tri -304 1073 -297 1080 nw
rect -311 1072 -305 1073
tri -305 1072 -304 1073 nw
tri -311 1066 -305 1072 nw
tri 3691 869 3715 893 se
rect 3715 871 3767 1896
rect 4163 2012 4370 2018
rect 4215 1994 4370 2012
tri 4370 1994 4394 2018 nw
tri 5165 1994 5189 2018 ne
rect 5189 1994 5267 2018
rect 4215 1960 4336 1994
tri 4336 1960 4370 1994 nw
tri 5189 1960 5223 1994 ne
rect 5223 1960 5267 1994
rect 4163 1957 4333 1960
tri 4333 1957 4336 1960 nw
tri 5223 1957 5226 1960 ne
rect 5226 1957 5267 1960
rect 4163 1954 4330 1957
tri 4330 1954 4333 1957 nw
rect 4163 1949 4325 1954
tri 4325 1949 4330 1954 nw
rect 4482 1951 4534 1957
tri 5226 1954 5229 1957 ne
rect 5229 1954 5267 1957
rect 4163 1948 4324 1949
tri 4324 1948 4325 1949 nw
rect 4215 1921 4297 1948
tri 4297 1921 4324 1948 nw
rect 4215 1896 4266 1921
rect 4163 1890 4266 1896
tri 4266 1890 4297 1921 nw
tri 5229 1949 5234 1954 ne
rect 5234 1949 5267 1954
tri 5234 1948 5235 1949 ne
rect 5235 1948 5267 1949
tri 5235 1921 5262 1948 ne
rect 5262 1921 5267 1948
tri 5262 1916 5267 1921 ne
rect 9110 1916 9280 2049
rect 13199 2106 13205 2140
rect 13239 2106 13245 2140
rect 13199 2067 13245 2106
rect 13199 2033 13205 2067
rect 13239 2033 13245 2067
rect 13199 1994 13245 2033
rect 13199 1960 13205 1994
rect 13239 1960 13245 1994
rect 13199 1921 13245 1960
rect 4482 1888 4534 1899
rect 4482 1887 5726 1888
rect 4534 1836 5726 1887
rect 13199 1887 13205 1921
rect 13239 1887 13245 1921
tri 8556 1880 8558 1882 se
rect 8558 1880 8562 1882
tri 8552 1876 8556 1880 se
rect 8556 1876 8562 1880
tri 8686 1880 8688 1882 sw
rect 8686 1876 8688 1880
tri 8688 1876 8692 1880 sw
rect 8686 1875 8692 1876
tri 8692 1875 8693 1876 sw
rect 5854 1858 5876 1860
tri 5876 1858 5878 1860 nw
rect 5854 1848 5866 1858
tri 5866 1848 5876 1858 nw
rect 13199 1848 13245 1887
tri 5854 1836 5866 1848 nw
rect 4482 1829 4534 1835
tri 7607 1829 7614 1836 sw
rect 7607 1814 7614 1829
tri 7614 1814 7629 1829 sw
rect 13199 1814 13205 1848
rect 13239 1814 13245 1848
rect 7607 1806 7629 1814
tri 7629 1806 7637 1814 sw
rect 7607 1804 7637 1806
tri 7637 1804 7639 1806 sw
tri 6982 1802 6984 1804 ne
rect 6984 1802 7016 1804
rect 7607 1802 7639 1804
tri 7639 1802 7641 1804 sw
tri 6984 1775 7011 1802 ne
rect 7011 1775 7016 1802
tri 7011 1770 7016 1775 ne
rect 13199 1775 13245 1814
rect 5628 1741 5633 1770
tri 5633 1741 5662 1770 nw
tri 5729 1741 5758 1770 ne
rect 5758 1741 5763 1770
tri 5628 1736 5633 1741 nw
tri 5758 1736 5763 1741 ne
rect 5809 1741 5814 1770
tri 5814 1741 5843 1770 nw
tri 6600 1742 6618 1760 se
rect 7607 1750 7635 1756
tri 7635 1750 7641 1756 nw
tri 7387 1742 7395 1750 se
tri 7386 1741 7387 1742 se
rect 7387 1741 7395 1742
tri 5809 1736 5814 1741 nw
tri 7382 1737 7386 1741 se
rect 7386 1737 7395 1741
rect 7607 1741 7626 1750
tri 7626 1741 7635 1750 nw
rect 13199 1741 13205 1775
rect 13239 1741 13245 1775
rect 7607 1737 7622 1741
tri 7622 1737 7626 1741 nw
rect 7607 1736 7621 1737
tri 7621 1736 7622 1737 nw
rect 7607 1732 7617 1736
tri 7617 1732 7621 1736 nw
rect 7607 1729 7614 1732
tri 7614 1729 7617 1732 nw
tri 7607 1722 7614 1729 nw
rect 5976 1702 5998 1714
tri 5998 1702 6010 1714 nw
tri 7041 1702 7052 1713 sw
rect 13199 1702 13245 1741
rect 5976 1682 5978 1702
tri 5978 1682 5998 1702 nw
rect 7041 1692 7052 1702
tri 7052 1692 7062 1702 sw
tri 7361 1682 7364 1685 ne
rect 7364 1682 7395 1685
tri 5976 1680 5978 1682 nw
tri 7364 1680 7366 1682 ne
rect 7366 1680 7395 1682
tri 7366 1678 7368 1680 ne
rect 7368 1678 7395 1680
tri 6612 1670 6620 1678 se
tri 7368 1670 7376 1678 ne
rect 7376 1670 7395 1678
tri 7376 1668 7378 1670 ne
rect 7378 1668 7395 1670
tri 7378 1658 7388 1668 ne
rect 7388 1658 7395 1668
tri 7388 1657 7389 1658 ne
rect 7389 1657 7395 1658
rect 6026 1631 6072 1657
tri 7389 1656 7390 1657 ne
rect 7390 1656 7395 1657
tri 7390 1651 7395 1656 ne
rect 8086 1668 8106 1682
tri 8106 1668 8120 1682 nw
rect 13199 1668 13205 1702
rect 13239 1668 13245 1702
rect 8086 1658 8096 1668
tri 8096 1658 8106 1668 nw
rect 8086 1656 8094 1658
tri 8094 1656 8096 1658 nw
rect 8086 1651 8089 1656
tri 8089 1651 8094 1656 nw
tri 8086 1648 8089 1651 nw
rect 6746 1646 6798 1648
rect 6929 1646 6981 1648
rect 6026 1629 6104 1631
tri 6104 1629 6106 1631 nw
tri 6250 1629 6252 1631 ne
rect 6252 1629 6284 1631
rect 6026 1626 6101 1629
tri 6101 1626 6104 1629 nw
tri 6252 1626 6255 1629 ne
rect 6255 1626 6284 1629
rect 13199 1629 13245 1668
tri 6004 1595 6026 1617 se
rect 6026 1599 6074 1626
tri 6074 1599 6101 1626 nw
tri 6255 1624 6257 1626 ne
rect 6257 1624 6284 1626
tri 8672 1624 8674 1626 ne
rect 8674 1624 8706 1626
tri 6257 1599 6282 1624 ne
rect 6282 1599 6284 1624
rect 6026 1598 6073 1599
tri 6073 1598 6074 1599 nw
tri 6282 1598 6283 1599 ne
rect 6283 1598 6284 1599
rect 6026 1595 6072 1598
tri 6072 1597 6073 1598 nw
tri 6283 1597 6284 1598 ne
rect 6418 1599 6427 1624
tri 6427 1599 6452 1624 nw
tri 6566 1599 6591 1624 ne
rect 6591 1599 6620 1624
tri 8674 1599 8699 1624 ne
rect 8699 1599 8706 1624
rect 6418 1598 6426 1599
tri 6426 1598 6427 1599 nw
tri 6591 1598 6592 1599 ne
rect 6592 1598 6620 1599
rect 8034 1598 8086 1599
tri 8699 1598 8700 1599 ne
rect 8700 1598 8706 1599
rect 6418 1597 6425 1598
tri 6425 1597 6426 1598 nw
tri 6592 1597 6593 1598 ne
rect 6593 1597 6620 1598
tri 5998 1589 6004 1595 se
rect 6004 1589 6072 1595
rect 6418 1595 6423 1597
tri 6423 1595 6425 1597 nw
tri 6593 1595 6595 1597 ne
rect 6595 1595 6620 1597
tri 8700 1595 8703 1598 ne
rect 8703 1595 8706 1598
rect 6418 1592 6420 1595
tri 6420 1592 6423 1595 nw
tri 6595 1592 6598 1595 ne
rect 6598 1592 6620 1595
tri 8703 1592 8706 1595 ne
rect 13199 1595 13205 1629
rect 13239 1595 13245 1629
tri 6418 1590 6420 1592 nw
tri 6598 1590 6600 1592 ne
rect 6600 1590 6620 1592
rect 5462 1537 5468 1589
rect 5520 1537 5532 1589
rect 5584 1584 5590 1589
tri 5996 1587 5998 1589 se
rect 5998 1587 6072 1589
tri 5590 1584 5593 1587 sw
tri 5993 1584 5996 1587 se
rect 5996 1584 6072 1587
tri 6600 1584 6606 1590 ne
rect 6606 1584 6620 1590
rect 5584 1583 5593 1584
tri 5593 1583 5594 1584 sw
tri 5992 1583 5993 1584 se
rect 5993 1583 6072 1584
tri 6606 1583 6607 1584 ne
rect 6607 1583 6620 1584
rect 5584 1537 6072 1583
tri 6607 1570 6620 1583 ne
tri 8444 1556 8458 1570 ne
rect 8458 1556 8478 1570
tri 8458 1540 8474 1556 ne
rect 8474 1540 8478 1556
rect 7149 1537 7180 1540
tri 7180 1537 7183 1540 nw
tri 8474 1537 8477 1540 ne
rect 8477 1537 8478 1540
rect 7149 1536 7179 1537
tri 7179 1536 7180 1537 nw
tri 8477 1536 8478 1537 ne
rect 13199 1556 13245 1595
rect 7149 1522 7165 1536
tri 7165 1522 7179 1536 nw
rect 13199 1522 13205 1556
rect 13239 1522 13245 1556
rect 7149 1511 7154 1522
tri 7154 1511 7165 1522 nw
rect 7149 1510 7153 1511
tri 7153 1510 7154 1511 nw
tri 7149 1506 7153 1510 nw
rect 5394 1496 5446 1502
tri 8323 1483 8324 1484 se
tri 8290 1450 8323 1483 se
rect 8323 1450 8324 1483
rect 13199 1483 13245 1522
tri 9013 1459 9022 1468 sw
tri 8359 1451 8367 1459 se
rect 8359 1450 8367 1451
tri 8367 1450 8376 1459 sw
rect 9013 1450 9022 1459
tri 9022 1450 9031 1459 sw
rect 5394 1430 5446 1444
rect 9013 1449 9031 1450
tri 9031 1449 9032 1450 sw
rect 13199 1449 13205 1483
rect 13239 1449 13245 1483
rect 9013 1447 9032 1449
tri 9032 1447 9034 1449 sw
rect 9013 1438 9034 1447
tri 9034 1438 9043 1447 sw
rect 9013 1437 9043 1438
tri 9043 1437 9044 1438 sw
rect 9013 1435 9044 1437
tri 9044 1435 9046 1437 sw
tri 8966 1434 8967 1435 se
rect 9013 1434 9046 1435
tri 9046 1434 9047 1435 sw
rect 5310 1372 5362 1388
rect 13199 1410 13245 1449
tri 7524 1386 7542 1404 sw
tri 8493 1386 8511 1404 se
rect 5394 1372 5446 1378
tri 6618 1376 6628 1386 sw
rect 7524 1376 7542 1386
tri 7542 1376 7552 1386 sw
tri 8483 1376 8493 1386 se
rect 8493 1376 8511 1386
rect 6618 1372 6628 1376
tri 6628 1372 6632 1376 sw
rect 6618 1365 6632 1372
tri 6632 1365 6639 1372 sw
rect 7524 1370 7552 1376
tri 7552 1370 7558 1376 sw
tri 8477 1370 8483 1376 se
rect 8483 1370 8511 1376
rect 13199 1376 13205 1410
rect 13239 1376 13245 1410
rect 8797 1365 8849 1371
rect 6618 1364 6639 1365
tri 6639 1364 6640 1365 sw
rect 6618 1361 6640 1364
tri 6640 1361 6643 1364 sw
rect 6618 1352 6643 1361
tri 6643 1352 6652 1361 sw
tri 9687 1337 9689 1339 se
rect 9689 1337 9716 1339
tri 9653 1303 9687 1337 se
rect 9687 1303 9716 1337
tri 9652 1302 9653 1303 se
rect 9653 1302 9716 1303
tri 9646 1296 9652 1302 se
rect 9652 1296 9716 1302
rect 7595 1244 7601 1296
rect 7653 1244 7669 1296
rect 7721 1244 7737 1296
rect 7789 1244 7804 1296
rect 7856 1244 7862 1296
rect 9771 1287 9777 1339
rect 9829 1287 9842 1339
rect 9771 1275 9842 1287
rect 5825 1210 5853 1238
rect 9771 1223 9777 1275
rect 9829 1223 9842 1275
rect 9771 1211 9842 1223
rect 9771 1159 9777 1211
rect 9829 1159 9842 1211
rect 10086 1159 10092 1339
tri 12467 1291 12469 1293 ne
rect 12469 1291 12501 1293
tri 12469 1264 12496 1291 ne
rect 12496 1264 12501 1291
tri 12496 1259 12501 1264 ne
rect 12503 1286 12509 1338
rect 12561 1286 12584 1338
rect 12636 1286 12659 1338
rect 12711 1286 12717 1338
rect 12503 1270 12717 1286
rect 12503 1218 12509 1270
rect 12561 1218 12584 1270
rect 12636 1218 12659 1270
rect 12711 1218 12717 1270
rect 13199 1337 13245 1376
rect 13199 1303 13205 1337
rect 13239 1303 13245 1337
rect 13199 1264 13245 1303
rect 12503 1202 12717 1218
rect 12503 1150 12509 1202
rect 12561 1150 12584 1202
rect 12636 1150 12659 1202
rect 12711 1150 12717 1202
rect 12503 1134 12717 1150
rect 12503 1082 12509 1134
rect 12561 1082 12584 1134
rect 12636 1082 12659 1134
rect 12711 1082 12717 1134
rect 13021 1239 13073 1246
rect 13021 1175 13073 1187
tri 12999 1015 13021 1037 se
rect 13021 1015 13073 1123
rect 6393 1014 6417 1015
tri 6417 1014 6418 1015 nw
tri 12998 1014 12999 1015 se
rect 12999 1014 13069 1015
rect 6393 1011 6414 1014
tri 6414 1011 6417 1014 nw
tri 11175 1011 11178 1014 ne
rect 11178 1011 11209 1014
tri 12995 1011 12998 1014 se
rect 12998 1011 13069 1014
tri 13069 1011 13073 1015 nw
rect 13199 1230 13205 1264
rect 13239 1230 13245 1264
rect 13199 1191 13245 1230
rect 13199 1157 13205 1191
rect 13239 1157 13245 1191
rect 13199 1118 13245 1157
rect 13199 1084 13205 1118
rect 13239 1084 13245 1118
tri 13281 2732 13296 2747 se
rect 13296 2732 13355 2747
tri 13355 2732 13370 2747 nw
rect 13281 2721 13344 2732
tri 13344 2721 13355 2732 nw
rect 13281 1239 13333 2721
tri 13333 2710 13344 2721 nw
rect 14977 2708 15023 2747
rect 13281 1175 13333 1187
rect 13281 1117 13333 1123
rect 13433 2692 14745 2698
rect 13433 2658 13511 2692
rect 13545 2658 13586 2692
rect 13620 2658 13661 2692
rect 13695 2658 13736 2692
rect 13770 2658 13811 2692
rect 13845 2658 13886 2692
rect 13920 2658 13961 2692
rect 13995 2658 14036 2692
rect 14070 2658 14111 2692
rect 14145 2658 14186 2692
rect 14220 2658 14261 2692
rect 14295 2658 14335 2692
rect 14369 2658 14409 2692
rect 14443 2658 14483 2692
rect 14517 2658 14557 2692
rect 14591 2658 14631 2692
rect 14665 2658 14745 2692
rect 13433 2652 14745 2658
rect 13433 2635 13496 2652
tri 13496 2635 13513 2652 nw
tri 14121 2635 14138 2652 ne
rect 14138 2635 14745 2652
rect 13433 2622 13483 2635
tri 13483 2622 13496 2635 nw
tri 14138 2622 14151 2635 ne
rect 14151 2622 14745 2635
rect 13433 2620 13481 2622
tri 13481 2620 13483 2622 nw
rect 13433 2592 13479 2620
tri 13479 2618 13481 2620 nw
rect 13433 2558 13439 2592
rect 13473 2558 13479 2592
rect 13433 2492 13479 2558
rect 13672 2570 13722 2622
rect 13774 2570 13786 2622
rect 13838 2570 13850 2622
rect 13902 2570 13915 2622
rect 13967 2620 13990 2622
tri 13990 2620 13992 2622 sw
tri 14151 2620 14153 2622 ne
rect 14153 2620 14745 2622
rect 13967 2618 13992 2620
tri 13992 2618 13994 2620 sw
tri 14153 2618 14155 2620 ne
rect 13967 2586 13994 2618
tri 13994 2586 14026 2618 sw
rect 14155 2586 14705 2620
rect 14739 2586 14745 2620
rect 13967 2573 14026 2586
tri 14026 2573 14039 2586 sw
rect 14155 2573 14745 2586
rect 13967 2570 14039 2573
rect 13672 2539 14039 2570
tri 14039 2539 14073 2573 sw
rect 14155 2539 14167 2573
rect 14201 2539 14240 2573
rect 14274 2539 14312 2573
rect 14346 2539 14384 2573
rect 14418 2539 14456 2573
rect 14490 2539 14528 2573
rect 14562 2539 14600 2573
rect 14634 2546 14745 2573
rect 14634 2539 14705 2546
rect 13433 2458 13439 2492
rect 13473 2458 13479 2492
rect 13433 2382 13479 2458
rect 13433 2348 13439 2382
rect 13473 2348 13479 2382
rect 13433 2310 13479 2348
rect 13433 2276 13439 2310
rect 13473 2276 13479 2310
rect 13433 2238 13479 2276
rect 13433 2204 13439 2238
rect 13473 2204 13479 2238
rect 13433 2166 13479 2204
rect 13433 2132 13439 2166
rect 13473 2132 13479 2166
rect 13433 2094 13479 2132
rect 13433 2060 13439 2094
rect 13473 2060 13479 2094
rect 13433 2021 13479 2060
rect 13433 1987 13439 2021
rect 13473 1987 13479 2021
rect 13433 1948 13479 1987
rect 13433 1914 13439 1948
rect 13473 1914 13479 1948
rect 13433 1875 13479 1914
rect 13433 1841 13439 1875
rect 13473 1841 13479 1875
rect 13433 1802 13479 1841
rect 13433 1768 13439 1802
rect 13473 1768 13479 1802
rect 13433 1729 13479 1768
rect 13433 1695 13439 1729
rect 13473 1695 13479 1729
rect 13433 1656 13479 1695
rect 13433 1622 13439 1656
rect 13473 1622 13479 1656
rect 13433 1583 13479 1622
rect 13433 1549 13439 1583
rect 13473 1549 13479 1583
rect 13433 1510 13479 1549
rect 13433 1476 13439 1510
rect 13473 1476 13479 1510
rect 13433 1437 13479 1476
rect 13433 1403 13439 1437
rect 13473 1403 13479 1437
rect 13433 1364 13479 1403
rect 13433 1330 13439 1364
rect 13473 1330 13479 1364
rect 13433 1291 13479 1330
rect 13433 1257 13439 1291
rect 13473 1257 13479 1291
rect 13433 1218 13479 1257
rect 13433 1184 13439 1218
rect 13473 1184 13479 1218
rect 13433 1145 13479 1184
rect 13199 1045 13245 1084
rect 13199 1011 13205 1045
rect 13239 1011 13245 1045
rect 6393 1006 6409 1011
tri 6409 1006 6414 1011 nw
tri 11178 1006 11183 1011 ne
rect 11183 1006 11209 1011
tri 12990 1006 12995 1011 se
rect 12995 1006 13064 1011
tri 13064 1006 13069 1011 nw
rect 6393 999 6402 1006
tri 6402 999 6409 1006 nw
tri 11183 999 11190 1006 ne
rect 11190 999 11209 1006
tri 12983 999 12990 1006 se
rect 12990 999 13057 1006
tri 13057 999 13064 1006 nw
tri 6393 990 6402 999 nw
tri 11190 990 11199 999 ne
rect 11199 990 11209 999
tri 12976 992 12983 999 se
rect 12983 992 13050 999
tri 13050 992 13057 999 nw
tri 11199 980 11209 990 ne
rect 11304 980 13038 992
tri 13038 980 13050 992 nw
rect 11304 972 13030 980
tri 13030 972 13038 980 nw
rect 13199 972 13245 1011
tri 6625 960 6636 971 se
tri 6241 958 6243 960 sw
tri 6623 958 6625 960 se
rect 6625 958 6636 960
rect 11304 958 13016 972
tri 13016 958 13030 972 nw
rect 6241 938 6243 958
tri 6243 938 6263 958 sw
tri 6603 938 6623 958 se
rect 6623 938 6636 958
rect 6241 937 6263 938
tri 6263 937 6264 938 sw
tri 6602 937 6603 938 se
rect 6603 937 6636 938
rect 6664 938 6678 958
tri 6678 938 6698 958 nw
tri 11101 938 11121 958 ne
rect 11121 938 11135 958
rect 6664 937 6677 938
tri 6677 937 6678 938 nw
tri 11121 937 11122 938 ne
rect 11122 937 11135 938
rect 6241 935 6264 937
tri 6264 935 6266 937 sw
rect 6664 935 6675 937
tri 6675 935 6677 937 nw
tri 11122 935 11124 937 ne
rect 11124 935 11135 937
rect 6664 932 6672 935
tri 6672 932 6675 935 nw
tri 11124 932 11127 935 ne
rect 11127 932 11135 935
rect 6664 927 6667 932
tri 6667 927 6672 932 nw
tri 11127 927 11132 932 ne
rect 11132 927 11135 932
rect 6664 926 6666 927
tri 6666 926 6667 927 nw
tri 11132 926 11133 927 ne
rect 11133 926 11135 927
tri 6664 924 6666 926 nw
tri 11133 924 11135 926 ne
rect 11304 940 12998 958
tri 12998 940 13016 958 nw
rect 11304 938 11388 940
tri 11388 938 11390 940 nw
rect 13199 938 13205 972
rect 13239 938 13245 972
rect 11304 932 11382 938
tri 11382 932 11388 938 nw
rect 11304 927 11377 932
tri 11377 927 11382 932 nw
rect 11304 926 11376 927
tri 11376 926 11377 927 nw
rect 11304 924 11374 926
tri 11374 924 11376 926 nw
rect 6233 908 6241 912
tri 6241 908 6245 912 nw
rect 3715 869 3765 871
tri 3765 869 3767 871 nw
tri 6666 869 6693 896 se
tri 3687 865 3691 869 se
rect 3691 865 3761 869
tri 3761 865 3765 869 nw
tri 6662 865 6666 869 se
rect 6666 865 6693 869
tri 3684 862 3687 865 se
rect 3687 862 3758 865
tri 3758 862 3761 865 nw
tri 6659 862 6662 865 se
rect 6662 862 6693 865
rect 6719 868 6745 869
tri 6745 868 6746 869 nw
rect 6719 865 6742 868
tri 6742 865 6745 868 nw
tri 6924 865 6927 868 ne
rect 6927 865 6949 868
tri 3682 860 3684 862 se
rect 3684 860 3756 862
tri 3756 860 3758 862 nw
rect 3682 858 3754 860
tri 3754 858 3756 860 nw
rect 6719 858 6735 865
tri 6735 858 6742 865 nw
tri 6927 858 6934 865 ne
rect 6934 858 6949 865
rect 3682 857 3753 858
tri 3753 857 3754 858 nw
rect 6719 857 6734 858
tri 6734 857 6735 858 nw
tri 6934 857 6935 858 ne
rect 6935 857 6949 858
rect 3682 853 3749 857
tri 3749 853 3753 857 nw
rect 6719 853 6730 857
tri 6730 853 6734 857 nw
tri 6935 853 6939 857 ne
rect 6939 853 6949 857
rect 3682 844 3740 853
tri 3740 844 3749 853 nw
rect 6719 844 6721 853
tri 6721 844 6730 853 nw
tri 6939 844 6948 853 ne
rect 6948 844 6949 853
rect 3682 839 3735 844
tri 3735 839 3740 844 nw
tri 3670 765 3682 777 se
rect 3682 765 3734 839
tri 3734 838 3735 839 nw
tri 6772 838 6773 839 se
rect 6773 838 6785 839
rect 9628 838 9656 866
tri 6771 837 6772 838 se
rect 6772 837 6785 838
tri 6757 823 6771 837 se
rect 6771 823 6785 837
tri 3784 803 3804 823 se
tri 6744 810 6757 823 se
rect 6757 810 6785 823
tri 3776 795 3784 803 se
rect 3784 795 3804 803
tri 3636 731 3670 765 se
rect 3670 731 3734 765
tri 3628 723 3636 731 se
rect 3636 723 3734 731
rect 846 671 852 723
rect 904 671 916 723
rect 968 721 3734 723
rect 968 720 3733 721
tri 3733 720 3734 721 nw
rect 968 719 3732 720
tri 3732 719 3733 720 nw
tri 3896 719 3897 720 sw
rect 968 710 3723 719
tri 3723 710 3732 719 nw
rect 3896 710 3897 719
tri 3897 710 3906 719 sw
rect 968 708 3721 710
tri 3721 708 3723 710 nw
rect 3896 708 3906 710
tri 3906 708 3908 710 sw
rect 968 707 3720 708
tri 3720 707 3721 708 nw
rect 3896 707 3908 708
tri 3908 707 3909 708 sw
rect 968 693 3706 707
tri 3706 693 3720 707 nw
rect 3896 693 3909 707
tri 3909 693 3923 707 sw
rect 968 686 3699 693
tri 3699 686 3706 693 nw
rect 3896 686 3923 693
tri 3923 686 3930 693 sw
tri 7688 686 7694 692 sw
rect 968 671 3684 686
tri 3684 671 3699 686 nw
rect 8595 646 8599 648
tri 8599 646 8601 648 nw
tri 8595 642 8599 646 nw
tri 7003 621 7007 625 se
tri 6994 612 7003 621 se
rect 7003 612 7007 621
rect 11304 621 11356 924
tri 11356 906 11374 924 nw
rect 13199 899 13245 938
rect 13199 865 13205 899
rect 13239 865 13245 899
tri 6996 573 7007 584 ne
tri 7161 562 7162 563 se
tri 7160 561 7161 562 se
rect 7161 561 7162 562
tri 7148 549 7160 561 se
rect 7160 549 7162 561
tri 7142 543 7148 549 se
rect 7148 543 7162 549
rect 11304 557 11356 569
tri 7155 515 7158 518 ne
rect 7158 515 7162 518
tri 7158 511 7162 515 ne
rect 11304 499 11356 505
rect 11490 837 12803 850
rect 11490 803 11502 837
rect 11536 803 11576 837
rect 11610 803 11650 837
rect 11684 803 11724 837
rect 11758 803 11798 837
rect 11832 803 11872 837
rect 11906 803 11946 837
rect 11980 803 12020 837
rect 12054 803 12094 837
rect 12128 803 12168 837
rect 12202 803 12242 837
rect 12276 803 12316 837
rect 12350 803 12390 837
rect 12424 803 12464 837
rect 12498 803 12538 837
rect 12572 803 12611 837
rect 12645 803 12684 837
rect 12718 803 12757 837
rect 12791 803 12803 837
rect 11490 765 12803 803
rect 11490 731 11502 765
rect 11536 731 11576 765
rect 11610 731 11650 765
rect 11684 731 11724 765
rect 11758 731 11798 765
rect 11832 731 11872 765
rect 11906 731 11946 765
rect 11980 731 12020 765
rect 12054 731 12094 765
rect 12128 731 12168 765
rect 12202 731 12242 765
rect 12276 731 12316 765
rect 12350 731 12390 765
rect 12424 731 12464 765
rect 12498 731 12538 765
rect 12572 731 12611 765
rect 12645 731 12684 765
rect 12718 731 12757 765
rect 12791 731 12803 765
rect 11490 693 12803 731
rect 11490 659 11502 693
rect 11536 659 11576 693
rect 11610 659 11650 693
rect 11684 659 11724 693
rect 11758 659 11798 693
rect 11832 659 11872 693
rect 11906 659 11946 693
rect 11980 659 12020 693
rect 12054 659 12094 693
rect 12128 659 12168 693
rect 12202 659 12242 693
rect 12276 659 12316 693
rect 12350 659 12390 693
rect 12424 659 12464 693
rect 12498 659 12538 693
rect 12572 659 12611 693
rect 12645 659 12684 693
rect 12718 659 12757 693
rect 12791 659 12803 693
rect 11490 621 12803 659
rect 11490 587 11502 621
rect 11536 587 11576 621
rect 11610 587 11650 621
rect 11684 587 11724 621
rect 11758 587 11798 621
rect 11832 587 11872 621
rect 11906 587 11946 621
rect 11980 587 12020 621
rect 12054 587 12094 621
rect 12128 587 12168 621
rect 12202 587 12242 621
rect 12276 587 12316 621
rect 12350 587 12390 621
rect 12424 587 12464 621
rect 12498 587 12538 621
rect 12572 587 12611 621
rect 12645 587 12684 621
rect 12718 587 12757 621
rect 12791 587 12803 621
rect 11490 549 12803 587
rect 11490 515 11502 549
rect 11536 515 11576 549
rect 11610 515 11650 549
rect 11684 515 11724 549
rect 11758 515 11798 549
rect 11832 515 11872 549
rect 11906 515 11946 549
rect 11980 515 12020 549
rect 12054 515 12094 549
rect 12128 515 12168 549
rect 12202 515 12242 549
rect 12276 515 12316 549
rect 12350 515 12390 549
rect 12424 515 12464 549
rect 12498 515 12538 549
rect 12572 515 12611 549
rect 12645 515 12684 549
rect 12718 515 12757 549
rect 12791 515 12803 549
rect 7627 477 7656 482
tri 7656 477 7661 482 nw
tri 10959 477 10964 482 ne
rect 10964 477 10993 482
rect 7627 457 7636 477
tri 7636 457 7656 477 nw
tri 10964 462 10979 477 ne
rect 10979 462 10993 477
tri 5267 448 5276 457 ne
rect 5276 448 5301 457
tri 7627 448 7636 457 nw
rect 9667 456 9670 462
tri 9670 456 9676 462 nw
tri 10979 456 10985 462 ne
rect 10985 456 10993 462
tri 10985 450 10991 456 ne
rect 10991 450 10993 456
tri 7672 448 7674 450 se
tri 10991 448 10993 450 ne
rect 11490 477 12803 515
tri 5276 443 5281 448 ne
rect 5281 443 5301 448
tri 5281 427 5297 443 ne
rect 5297 427 5301 443
tri 5297 423 5301 427 ne
tri 7670 446 7672 448 se
rect 7672 446 7674 448
tri 4137 405 4145 413 se
tri 4121 389 4137 405 se
rect 4137 389 4145 405
rect 7670 402 7674 446
rect 11490 443 11502 477
rect 11536 443 11576 477
rect 11610 443 11650 477
rect 11684 443 11724 477
rect 11758 443 11798 477
rect 11832 443 11872 477
rect 11906 443 11946 477
rect 11980 443 12020 477
rect 12054 443 12094 477
rect 12128 443 12168 477
rect 12202 443 12242 477
rect 12276 443 12316 477
rect 12350 443 12390 477
rect 12424 443 12464 477
rect 12498 443 12538 477
rect 12572 443 12611 477
rect 12645 443 12684 477
rect 12718 443 12757 477
rect 12791 443 12803 477
rect 11490 405 12803 443
rect 4562 386 4614 392
tri 8063 354 8066 357 ne
rect 8066 354 8097 357
tri 8066 350 8070 354 ne
rect 8070 350 8097 354
tri 8070 344 8076 350 ne
rect 8076 344 8097 350
tri 8076 343 8077 344 ne
rect 8077 343 8097 344
tri 8521 343 8522 344 ne
rect 8522 343 8527 344
tri 8077 342 8078 343 ne
rect 8078 342 8097 343
tri 8522 342 8523 343 ne
rect 8523 342 8527 343
tri 8078 338 8082 342 ne
rect 8082 338 8097 342
tri 8523 338 8527 342 ne
rect 9965 338 9974 390
rect 11490 371 11502 405
rect 11536 371 11576 405
rect 11610 371 11650 405
rect 11684 371 11724 405
rect 11758 371 11798 405
rect 11832 371 11872 405
rect 11906 371 11946 405
rect 11980 371 12020 405
rect 12054 371 12094 405
rect 12128 371 12168 405
rect 12202 371 12242 405
rect 12276 371 12316 405
rect 12350 371 12390 405
rect 12424 371 12464 405
rect 12498 371 12538 405
rect 12572 371 12611 405
rect 12645 371 12684 405
rect 12718 371 12757 405
rect 12791 371 12803 405
rect 10523 354 10554 357
tri 10554 354 10557 357 nw
rect 10523 350 10550 354
tri 10550 350 10554 354 nw
rect 10102 343 10107 344
tri 10107 343 10108 344 nw
rect 10523 343 10543 350
tri 10543 343 10550 350 nw
rect 10102 342 10106 343
tri 10106 342 10107 343 nw
rect 10523 342 10542 343
tri 10542 342 10543 343 nw
tri 10102 338 10106 342 nw
tri 8082 334 8086 338 ne
rect 8086 334 8097 338
rect 4562 333 4614 334
tri 4614 333 4615 334 sw
tri 8086 333 8087 334 ne
rect 8087 333 8097 334
rect 4562 322 4615 333
tri 4283 300 4288 305 ne
rect 4288 300 4307 305
tri 4288 299 4289 300 ne
rect 4289 299 4307 300
tri 4289 281 4307 299 ne
tri 3722 270 3729 277 se
rect 3729 270 3739 277
tri 3715 263 3722 270 se
rect 3722 263 3739 270
rect 4614 300 4615 322
tri 4615 300 4648 333 sw
tri 8087 323 8097 333 ne
rect 10523 334 10534 342
tri 10534 334 10542 342 nw
rect 10523 333 10533 334
tri 10533 333 10534 334 nw
tri 10523 323 10533 333 nw
rect 4614 270 5951 300
rect 4562 264 5951 270
rect 7893 266 7913 318
tri 9595 306 9598 309 se
tri 5917 263 5918 264 ne
rect 5918 263 5951 264
tri 5918 261 5920 263 ne
rect 5920 261 5951 263
tri 5920 254 5927 261 ne
rect 5927 254 5951 261
tri 9595 257 9598 260 ne
rect 9598 257 9604 309
rect 9656 257 9668 309
rect 9720 257 9726 309
rect 10722 264 10727 316
rect 10958 282 10960 334
rect 11490 333 12803 371
tri 11237 300 11254 317 sw
rect 11237 299 11254 300
tri 11254 299 11255 300 sw
rect 11490 299 11502 333
rect 11536 299 11576 333
rect 11610 299 11650 333
rect 11684 299 11724 333
rect 11758 299 11798 333
rect 11832 299 11872 333
rect 11906 299 11946 333
rect 11980 299 12020 333
rect 12054 299 12094 333
rect 12128 299 12168 333
rect 12202 299 12242 333
rect 12276 299 12316 333
rect 12350 299 12390 333
rect 12424 299 12464 333
rect 12498 299 12538 333
rect 12572 299 12611 333
rect 12645 299 12684 333
rect 12718 299 12757 333
rect 12791 299 12803 333
rect 11237 293 11255 299
tri 11255 293 11261 299 sw
tri 11486 282 11490 286 se
rect 11490 282 12803 299
tri 11485 281 11486 282 se
rect 11486 281 12803 282
tri 11482 278 11485 281 se
rect 11485 278 12803 281
tri 11474 270 11482 278 se
rect 11482 270 12803 278
tri 11468 264 11474 270 se
rect 11474 264 12803 270
tri 11465 261 11468 264 se
rect 11468 261 12803 264
tri 11461 257 11465 261 se
rect 11465 257 11502 261
tri 11458 254 11461 257 se
rect 11461 254 11502 257
tri 5927 240 5941 254 ne
rect 5941 240 5951 254
tri 3714 227 3727 240 ne
rect 3727 227 3748 240
tri 5941 230 5951 240 ne
rect 5997 240 6017 254
tri 6017 240 6031 254 nw
tri 11444 240 11458 254 se
rect 11458 240 11502 254
tri 3727 225 3729 227 ne
rect 3729 225 3748 227
rect 5997 227 6004 240
tri 6004 227 6017 240 nw
tri 11431 227 11444 240 se
rect 11444 227 11502 240
rect 11536 227 11576 261
rect 11610 227 11650 261
rect 11684 227 11724 261
rect 11758 227 11798 261
rect 11832 227 11872 261
rect 11906 227 11946 261
rect 11980 227 12020 261
rect 12054 227 12094 261
rect 12128 227 12168 261
rect 12202 227 12242 261
rect 12276 227 12316 261
rect 12350 227 12390 261
rect 12424 227 12464 261
rect 12498 227 12538 261
rect 12572 227 12611 261
rect 12645 227 12684 261
rect 12718 227 12757 261
rect 12791 227 12803 261
rect 5997 225 6002 227
tri 6002 225 6004 227 nw
tri 11429 225 11431 227 se
rect 11431 225 12803 227
tri 5997 220 6002 225 nw
tri 11424 220 11429 225 se
rect 11429 220 12803 225
tri 11417 213 11424 220 se
rect 11424 213 12803 220
tri 5493 210 5496 213 se
rect 5496 210 5548 213
tri 11414 210 11417 213 se
rect 11417 210 12803 213
tri 5491 208 5493 210 se
rect 5493 208 5496 210
tri 11412 208 11414 210 se
rect 11414 208 12803 210
tri 5490 207 5491 208 se
rect 5491 207 5496 208
tri 11411 207 11412 208 se
rect 11412 207 12803 208
rect 3680 206 3687 207
tri 3687 206 3688 207 sw
tri 3947 206 3948 207 se
rect 3948 206 3955 207
tri 11410 206 11411 207 se
rect 11411 206 12803 207
rect 3680 189 3688 206
tri 3688 189 3705 206 sw
tri 3930 189 3947 206 se
rect 3947 189 3955 206
tri 11393 189 11410 206 se
rect 11410 189 12803 206
rect 3680 186 3705 189
tri 3705 186 3708 189 sw
tri 3927 186 3930 189 se
rect 3930 186 3955 189
tri 11390 186 11393 189 se
rect 11393 186 11502 189
tri 11383 179 11390 186 se
rect 11390 179 11502 186
tri 3635 159 3655 179 ne
rect 3655 159 3657 179
rect 3976 159 3978 179
tri 3978 159 3998 179 nw
tri 11381 177 11383 179 se
rect 11383 177 11502 179
tri 5462 159 5480 177 ne
rect 5480 159 5496 177
tri 5480 155 5484 159 ne
rect 5484 155 5496 159
tri 11359 155 11381 177 se
rect 11381 155 11502 177
rect 11536 155 11576 189
rect 11610 155 11650 189
rect 11684 155 11724 189
rect 11758 155 11798 189
rect 11832 155 11872 189
rect 11906 155 11946 189
rect 11980 155 12020 189
rect 12054 155 12094 189
rect 12128 155 12168 189
rect 12202 155 12242 189
rect 12276 155 12316 189
rect 12350 155 12390 189
rect 12424 155 12464 189
rect 12498 155 12538 189
rect 12572 155 12611 189
rect 12645 155 12684 189
rect 12718 155 12757 189
rect 12791 155 12803 189
tri 5484 143 5496 155 ne
tri 11347 143 11359 155 se
rect 11359 143 12803 155
tri 11339 135 11347 143 se
rect 11347 135 12803 143
tri 11338 134 11339 135 se
rect 11339 134 12803 135
tri 11321 117 11338 134 se
rect 11338 117 12803 134
tri 11311 107 11321 117 se
rect 11321 107 11502 117
rect 11109 83 11502 107
rect 11536 83 11576 117
rect 11610 83 11650 117
rect 11684 83 11724 117
rect 11758 83 11798 117
rect 11832 83 11872 117
rect 11906 83 11946 117
rect 11980 83 12020 117
rect 12054 83 12094 117
rect 12128 83 12168 117
rect 12202 83 12242 117
rect 12276 83 12316 117
rect 12350 83 12390 117
rect 12424 83 12464 117
rect 12498 83 12538 117
rect 12572 83 12611 117
rect 12645 83 12684 117
rect 12718 83 12757 117
rect 12791 83 12803 117
rect 11109 70 12803 83
rect 13199 826 13245 865
rect 13199 792 13205 826
rect 13239 792 13245 826
rect 13199 753 13245 792
rect 13199 719 13205 753
rect 13239 719 13245 753
rect 13199 680 13245 719
rect 13199 646 13205 680
rect 13239 646 13245 680
rect 13199 607 13245 646
rect 13199 573 13205 607
rect 13239 573 13245 607
rect 13199 534 13245 573
rect 13199 500 13205 534
rect 13239 500 13245 534
rect 13199 461 13245 500
rect 13199 427 13205 461
rect 13239 427 13245 461
rect 13199 388 13245 427
rect 13199 354 13205 388
rect 13239 354 13245 388
rect 13199 315 13245 354
rect 13199 281 13205 315
rect 13239 281 13245 315
rect 13199 242 13245 281
rect 13199 208 13205 242
rect 13239 208 13245 242
rect 13199 169 13245 208
rect 13199 135 13205 169
rect 13239 135 13245 169
rect 13199 96 13245 135
rect 13433 1111 13439 1145
rect 13473 1111 13479 1145
rect 13433 1072 13479 1111
rect 13433 1038 13439 1072
rect 13473 1038 13479 1072
rect 13433 999 13479 1038
rect 13433 965 13439 999
rect 13473 965 13479 999
rect 13433 926 13479 965
rect 13433 892 13439 926
rect 13473 892 13479 926
rect 13433 853 13479 892
rect 13433 819 13439 853
rect 13473 819 13479 853
rect 13433 780 13479 819
rect 13433 746 13439 780
rect 13473 746 13479 780
rect 13433 707 13479 746
rect 13433 673 13439 707
rect 13473 673 13479 707
rect 13433 634 13479 673
rect 13433 600 13439 634
rect 13473 600 13479 634
rect 13433 561 13479 600
rect 13433 527 13439 561
rect 13473 527 13479 561
rect 13433 488 13479 527
rect 13433 454 13439 488
rect 13473 454 13479 488
rect 13545 2516 13597 2528
rect 13545 2482 13554 2516
rect 13588 2482 13597 2516
rect 13545 2443 13597 2482
rect 13545 2409 13554 2443
rect 13588 2409 13597 2443
rect 13545 2370 13597 2409
rect 13545 2336 13554 2370
rect 13588 2336 13597 2370
rect 13545 2297 13597 2336
rect 13545 2263 13554 2297
rect 13588 2263 13597 2297
rect 13545 2224 13597 2263
rect 13545 2190 13554 2224
rect 13588 2190 13597 2224
rect 13545 2150 13597 2190
rect 13545 2116 13554 2150
rect 13588 2116 13597 2150
rect 13545 2101 13597 2116
rect 13545 2042 13554 2049
rect 13588 2042 13597 2049
rect 13545 2037 13597 2042
rect 13545 1968 13554 1985
rect 13588 1968 13597 1985
rect 13545 1928 13597 1968
rect 13545 1894 13554 1928
rect 13588 1894 13597 1928
rect 13545 1854 13597 1894
rect 13545 1820 13554 1854
rect 13588 1820 13597 1854
rect 13545 1780 13597 1820
rect 13545 1746 13554 1780
rect 13588 1746 13597 1780
rect 13545 1706 13597 1746
rect 13545 1672 13554 1706
rect 13588 1672 13597 1706
rect 13545 1632 13597 1672
rect 13545 1598 13554 1632
rect 13588 1598 13597 1632
rect 13545 1558 13597 1598
rect 13545 1524 13554 1558
rect 13588 1524 13597 1558
rect 13545 1484 13597 1524
rect 13545 1450 13554 1484
rect 13588 1450 13597 1484
rect 13545 1410 13597 1450
rect 13672 2519 14073 2539
tri 14073 2519 14093 2539 sw
rect 13672 2417 14093 2519
rect 13672 2383 13684 2417
rect 13718 2383 13757 2417
rect 13791 2383 13830 2417
rect 13864 2383 13903 2417
rect 13937 2383 13975 2417
rect 14009 2383 14047 2417
rect 14081 2383 14093 2417
rect 13672 2105 14093 2383
rect 13672 2071 13684 2105
rect 13718 2071 13757 2105
rect 13791 2071 13830 2105
rect 13864 2071 13903 2105
rect 13937 2071 13975 2105
rect 14009 2071 14047 2105
rect 14081 2071 14093 2105
rect 13672 1793 14093 2071
rect 13672 1759 13684 1793
rect 13718 1759 13757 1793
rect 13791 1759 13830 1793
rect 13864 1759 13903 1793
rect 13937 1759 13975 1793
rect 14009 1759 14047 1793
rect 14081 1759 14093 1793
rect 13672 1481 14093 1759
rect 13672 1447 13684 1481
rect 13718 1447 13757 1481
rect 13791 1447 13830 1481
rect 13864 1447 13903 1481
rect 13937 1447 13975 1481
rect 14009 1447 14047 1481
rect 14081 1447 14093 1481
rect 13672 1441 14093 1447
rect 14155 2512 14705 2539
rect 14739 2512 14745 2546
rect 14155 2472 14745 2512
rect 14155 2438 14705 2472
rect 14739 2438 14745 2472
rect 14155 2398 14745 2438
rect 14155 2364 14705 2398
rect 14739 2364 14745 2398
rect 14155 2324 14745 2364
rect 14155 2290 14705 2324
rect 14739 2290 14745 2324
rect 14155 2261 14745 2290
rect 14155 2227 14167 2261
rect 14201 2227 14240 2261
rect 14274 2227 14312 2261
rect 14346 2227 14384 2261
rect 14418 2227 14456 2261
rect 14490 2227 14528 2261
rect 14562 2227 14600 2261
rect 14634 2250 14745 2261
rect 14634 2227 14705 2250
rect 14155 2216 14705 2227
rect 14739 2216 14745 2250
rect 14155 2176 14745 2216
rect 14155 2142 14705 2176
rect 14739 2142 14745 2176
rect 14155 2102 14745 2142
rect 14155 2068 14705 2102
rect 14739 2068 14745 2102
rect 14155 2028 14745 2068
rect 14155 1994 14705 2028
rect 14739 1994 14745 2028
rect 14155 1954 14745 1994
rect 14155 1949 14705 1954
rect 14155 1915 14167 1949
rect 14201 1915 14240 1949
rect 14274 1915 14312 1949
rect 14346 1915 14384 1949
rect 14418 1915 14456 1949
rect 14490 1915 14528 1949
rect 14562 1915 14600 1949
rect 14634 1920 14705 1949
rect 14739 1920 14745 1954
rect 14634 1915 14745 1920
rect 14155 1880 14745 1915
rect 14155 1846 14705 1880
rect 14739 1846 14745 1880
rect 14155 1806 14745 1846
rect 14155 1772 14705 1806
rect 14739 1772 14745 1806
rect 14155 1732 14745 1772
rect 14155 1698 14705 1732
rect 14739 1698 14745 1732
rect 14155 1658 14745 1698
rect 14155 1637 14705 1658
rect 14155 1603 14167 1637
rect 14201 1603 14240 1637
rect 14274 1603 14312 1637
rect 14346 1603 14384 1637
rect 14418 1603 14456 1637
rect 14490 1603 14528 1637
rect 14562 1603 14600 1637
rect 14634 1624 14705 1637
rect 14739 1624 14745 1658
rect 14634 1603 14745 1624
rect 14155 1584 14745 1603
rect 14155 1550 14705 1584
rect 14739 1550 14745 1584
rect 14155 1511 14745 1550
rect 14155 1477 14705 1511
rect 14739 1477 14745 1511
rect 13545 1376 13554 1410
rect 13588 1376 13597 1410
rect 13545 1336 13597 1376
rect 13545 1302 13554 1336
rect 13588 1302 13597 1336
rect 13545 1262 13597 1302
rect 13545 1228 13554 1262
rect 13588 1228 13597 1262
rect 13545 1188 13597 1228
rect 13545 1154 13554 1188
rect 13588 1154 13597 1188
rect 14155 1438 14745 1477
rect 14155 1404 14705 1438
rect 14739 1404 14745 1438
rect 14155 1365 14745 1404
rect 14155 1331 14705 1365
rect 14739 1331 14745 1365
rect 14155 1325 14745 1331
rect 14155 1291 14167 1325
rect 14201 1291 14240 1325
rect 14274 1291 14312 1325
rect 14346 1291 14384 1325
rect 14418 1291 14456 1325
rect 14490 1291 14528 1325
rect 14562 1291 14600 1325
rect 14634 1292 14745 1325
rect 14634 1291 14705 1292
rect 14155 1258 14705 1291
rect 14739 1258 14745 1292
rect 14155 1219 14745 1258
rect 14155 1185 14705 1219
rect 14739 1185 14745 1219
rect 13545 1114 13597 1154
rect 13545 1080 13554 1114
rect 13588 1080 13597 1114
rect 13545 1040 13597 1080
rect 13545 1006 13554 1040
rect 13588 1006 13597 1040
rect 13545 966 13597 1006
rect 13545 932 13554 966
rect 13588 932 13597 966
rect 13545 892 13597 932
rect 13545 858 13554 892
rect 13588 858 13597 892
rect 13545 818 13597 858
rect 13545 784 13554 818
rect 13588 784 13597 818
rect 13545 744 13597 784
rect 13545 710 13554 744
rect 13588 710 13597 744
rect 13545 670 13597 710
rect 13545 636 13554 670
rect 13588 636 13597 670
rect 13545 596 13597 636
rect 13545 562 13554 596
rect 13588 562 13597 596
rect 13545 522 13597 562
rect 13545 488 13554 522
rect 13588 488 13597 522
rect 13672 1173 14093 1179
rect 13672 1169 13725 1173
rect 13777 1169 14093 1173
rect 13672 1135 13684 1169
rect 13718 1135 13725 1169
rect 13791 1135 13830 1169
rect 13864 1135 13903 1169
rect 13937 1135 13975 1169
rect 14009 1135 14047 1169
rect 14081 1135 14093 1169
rect 13672 1121 13725 1135
rect 13777 1121 14093 1135
rect 13672 1061 14093 1121
rect 13672 1009 13725 1061
rect 13777 1009 14093 1061
rect 13672 948 14093 1009
rect 13672 896 13725 948
rect 13777 896 14093 948
rect 13672 857 14093 896
rect 13672 823 13684 857
rect 13718 835 13757 857
rect 13718 823 13725 835
rect 13791 823 13830 857
rect 13864 823 13903 857
rect 13937 823 13975 857
rect 14009 823 14047 857
rect 14081 823 14093 857
rect 13672 783 13725 823
rect 13777 783 14093 823
rect 13672 722 14093 783
rect 13672 670 13725 722
rect 13777 670 14093 722
rect 13672 609 14093 670
rect 13672 557 13725 609
rect 13777 557 14093 609
rect 13672 545 14093 557
rect 13672 511 13684 545
rect 13718 511 13757 545
rect 13791 511 13830 545
rect 13864 511 13903 545
rect 13937 511 13975 545
rect 14009 511 14047 545
rect 14081 511 14093 545
rect 13672 505 14093 511
rect 14155 1146 14745 1185
rect 14155 1112 14705 1146
rect 14739 1112 14745 1146
rect 14155 1073 14745 1112
rect 14155 1039 14705 1073
rect 14739 1039 14745 1073
rect 14155 1013 14745 1039
rect 14155 979 14167 1013
rect 14201 979 14240 1013
rect 14274 979 14312 1013
rect 14346 979 14384 1013
rect 14418 979 14456 1013
rect 14490 979 14528 1013
rect 14562 979 14600 1013
rect 14634 1000 14745 1013
rect 14634 979 14705 1000
rect 14155 966 14705 979
rect 14739 966 14745 1000
rect 14155 927 14745 966
rect 14155 893 14705 927
rect 14739 893 14745 927
rect 14155 854 14745 893
rect 14155 820 14705 854
rect 14739 820 14745 854
rect 14155 781 14745 820
rect 14155 747 14705 781
rect 14739 747 14745 781
rect 14155 708 14745 747
rect 14155 701 14705 708
rect 14155 667 14167 701
rect 14201 667 14240 701
rect 14274 667 14312 701
rect 14346 667 14384 701
rect 14418 667 14456 701
rect 14490 667 14528 701
rect 14562 667 14600 701
rect 14634 674 14705 701
rect 14739 674 14745 708
rect 14634 667 14745 674
rect 14155 635 14745 667
rect 14155 601 14705 635
rect 14739 601 14745 635
rect 14155 562 14745 601
rect 14155 528 14705 562
rect 14739 528 14745 562
rect 13545 476 13597 488
rect 14155 489 14745 528
rect 13433 415 13479 454
rect 13433 381 13439 415
rect 13473 381 13479 415
rect 13433 343 13479 381
rect 14155 455 14705 489
rect 14739 455 14745 489
rect 14155 416 14745 455
rect 14155 389 14705 416
rect 14155 355 14167 389
rect 14201 355 14240 389
rect 14274 355 14312 389
rect 14346 355 14384 389
rect 14418 355 14456 389
rect 14490 355 14528 389
rect 14562 355 14600 389
rect 14634 382 14705 389
rect 14739 382 14745 416
rect 14634 355 14745 382
tri 13479 343 13484 348 sw
tri 14150 343 14155 348 se
rect 14155 343 14745 355
rect 13433 342 13484 343
rect 13433 262 13439 342
rect 13473 314 13484 342
tri 13484 314 13513 343 sw
tri 14121 314 14150 343 se
rect 14150 314 14705 343
rect 13491 262 13508 314
rect 13560 262 13577 314
rect 13629 262 13646 314
rect 13698 262 13714 314
rect 13766 270 13782 314
rect 13834 270 13850 314
rect 13902 270 13918 314
rect 13970 309 14705 314
rect 14739 309 14745 343
rect 13970 270 14745 309
rect 13769 262 13782 270
rect 13843 262 13850 270
rect 13917 262 13918 270
rect 13433 242 13513 262
rect 13547 242 13587 262
rect 13621 242 13661 262
rect 13695 242 13735 262
rect 13769 242 13809 262
rect 13843 242 13883 262
rect 13917 242 13958 262
rect 13433 190 13439 242
rect 13491 190 13508 242
rect 13560 190 13577 242
rect 13629 190 13646 242
rect 13698 190 13714 242
rect 13769 236 13782 242
rect 13843 236 13850 242
rect 13917 236 13918 242
rect 13992 236 14033 270
rect 14067 236 14108 270
rect 14142 236 14183 270
rect 14217 236 14258 270
rect 14292 236 14333 270
rect 14367 236 14408 270
rect 14442 236 14483 270
rect 14517 236 14558 270
rect 14592 236 14633 270
rect 14667 236 14745 270
rect 13766 190 13782 236
rect 13834 190 13850 236
rect 13902 190 13918 236
rect 13970 190 14745 236
rect 13433 170 14745 190
rect 13433 118 13439 170
rect 13491 118 13508 170
rect 13560 118 13577 170
rect 13629 118 13646 170
rect 13698 118 13714 170
rect 13766 118 13782 170
rect 13834 118 13850 170
rect 13902 118 13918 170
rect 13970 118 14745 170
rect 14977 2674 14983 2708
rect 15017 2674 15023 2708
rect 14977 2635 15023 2674
rect 14977 2601 14983 2635
rect 15017 2601 15023 2635
rect 14977 2562 15023 2601
rect 14977 2528 14983 2562
rect 15017 2528 15023 2562
rect 14977 2489 15023 2528
rect 14977 2455 14983 2489
rect 15017 2455 15023 2489
rect 14977 2416 15023 2455
rect 14977 2382 14983 2416
rect 15017 2382 15023 2416
rect 14977 2343 15023 2382
rect 14977 2309 14983 2343
rect 15017 2309 15023 2343
rect 14977 2270 15023 2309
rect 14977 2236 14983 2270
rect 15017 2236 15023 2270
rect 14977 2197 15023 2236
rect 14977 2163 14983 2197
rect 15017 2163 15023 2197
rect 14977 2124 15023 2163
rect 14977 2090 14983 2124
rect 15017 2090 15023 2124
rect 14977 2051 15023 2090
rect 14977 2017 14983 2051
rect 15017 2017 15023 2051
rect 14977 1978 15023 2017
rect 14977 1944 14983 1978
rect 15017 1944 15023 1978
rect 14977 1905 15023 1944
rect 14977 1871 14983 1905
rect 15017 1871 15023 1905
rect 14977 1832 15023 1871
rect 14977 1798 14983 1832
rect 15017 1798 15023 1832
rect 14977 1759 15023 1798
rect 14977 1725 14983 1759
rect 15017 1725 15023 1759
rect 14977 1686 15023 1725
rect 14977 1652 14983 1686
rect 15017 1652 15023 1686
rect 14977 1613 15023 1652
rect 14977 1579 14983 1613
rect 15017 1579 15023 1613
rect 14977 1540 15023 1579
rect 14977 1506 14983 1540
rect 15017 1506 15023 1540
rect 14977 1467 15023 1506
rect 14977 1433 14983 1467
rect 15017 1433 15023 1467
rect 14977 1394 15023 1433
rect 14977 1360 14983 1394
rect 15017 1360 15023 1394
rect 14977 1321 15023 1360
rect 14977 1287 14983 1321
rect 15017 1287 15023 1321
rect 14977 1248 15023 1287
rect 14977 1214 14983 1248
rect 15017 1214 15023 1248
rect 14977 1176 15023 1214
rect 14977 1142 14983 1176
rect 15017 1142 15023 1176
rect 14977 1104 15023 1142
rect 14977 1070 14983 1104
rect 15017 1070 15023 1104
rect 14977 1032 15023 1070
rect 14977 998 14983 1032
rect 15017 998 15023 1032
rect 14977 960 15023 998
rect 14977 926 14983 960
rect 15017 926 15023 960
rect 14977 888 15023 926
rect 14977 854 14983 888
rect 15017 854 15023 888
rect 14977 816 15023 854
rect 14977 782 14983 816
rect 15017 782 15023 816
rect 14977 744 15023 782
rect 14977 710 14983 744
rect 15017 710 15023 744
rect 14977 672 15023 710
rect 14977 638 14983 672
rect 15017 638 15023 672
rect 14977 600 15023 638
rect 14977 566 14983 600
rect 15017 566 15023 600
rect 14977 528 15023 566
rect 14977 494 14983 528
rect 15017 494 15023 528
rect 14977 456 15023 494
rect 14977 422 14983 456
rect 15017 422 15023 456
rect 14977 384 15023 422
rect 14977 350 14983 384
rect 15017 350 15023 384
rect 14977 312 15023 350
rect 14977 278 14983 312
rect 15017 278 15023 312
rect 14977 240 15023 278
rect 14977 206 14983 240
rect 15017 206 15023 240
rect 14977 168 15023 206
rect 14977 134 14983 168
rect 15017 134 15023 168
rect 11109 62 11852 70
tri 11852 62 11860 70 nw
rect 13199 62 13205 96
rect 13239 62 13245 96
rect 14977 96 15023 134
tri 13245 62 13247 64 sw
tri 14975 62 14977 64 se
rect 14977 62 14983 96
rect 15017 62 15023 96
rect 11109 24 11814 62
tri 11814 24 11852 62 nw
rect 13199 30 13247 62
tri 13247 30 13279 62 sw
tri 14943 30 14975 62 se
rect 14975 30 15023 62
rect 13199 24 15023 30
rect 11109 21 11811 24
tri 11811 21 11814 24 nw
rect 11109 15 11780 21
rect 7596 -43 7602 9
rect 7654 -43 7703 9
rect 7755 -43 7803 9
rect 7855 -43 7861 9
rect 7596 -55 7861 -43
rect 7596 -107 7602 -55
rect 7654 -107 7703 -55
rect 7755 -107 7803 -55
rect 7855 -107 7861 -55
rect 11109 -19 11346 15
rect 11380 -19 11420 15
rect 11454 -19 11494 15
rect 11528 -19 11567 15
rect 11601 -19 11640 15
rect 11674 -10 11780 15
tri 11780 -10 11811 21 nw
rect 13199 -10 13279 24
rect 13313 -10 13353 24
rect 13387 -10 13427 24
rect 13461 -10 13501 24
rect 13535 -10 13575 24
rect 13609 -10 13649 24
rect 13683 -10 13723 24
rect 13757 -10 13797 24
rect 13831 -10 13871 24
rect 13905 -10 13945 24
rect 13979 -10 14019 24
rect 14053 -10 14093 24
rect 14127 -10 14167 24
rect 14201 -10 14241 24
rect 14275 -10 14315 24
rect 14349 -10 14389 24
rect 14423 -10 14463 24
rect 14497 -10 14537 24
rect 14571 -10 14611 24
rect 14645 -10 14686 24
rect 14720 -10 14761 24
rect 14795 -10 14836 24
rect 14870 -10 14911 24
rect 14945 -10 15023 24
rect 11674 -16 11774 -10
tri 11774 -16 11780 -10 nw
rect 13199 -16 15023 -10
rect 11674 -19 11693 -16
rect 11109 -57 11693 -19
rect 11109 -91 11346 -57
rect 11380 -91 11420 -57
rect 11454 -91 11494 -57
rect 11528 -91 11567 -57
rect 11601 -91 11640 -57
rect 11674 -91 11693 -57
rect 11109 -97 11693 -91
tri 11693 -97 11774 -16 nw
rect 11109 -107 11683 -97
tri 11683 -107 11693 -97 nw
tri -797 -472 -763 -438 nw
rect 12310 -768 12749 -762
rect 12310 -802 12322 -768
rect 12356 -802 12399 -768
rect 12433 -802 12475 -768
rect 12509 -802 12551 -768
rect 12585 -802 12627 -768
rect 12661 -802 12703 -768
rect 12737 -802 12749 -768
rect 12310 -840 12749 -802
rect 12310 -874 12322 -840
rect 12356 -874 12399 -840
rect 12433 -874 12475 -840
rect 12509 -874 12551 -840
rect 12585 -874 12627 -840
rect 12661 -874 12703 -840
rect 12737 -874 12749 -840
rect 12310 -912 12749 -874
rect -76 -954 -48 -926
rect 12310 -946 12322 -912
rect 12356 -946 12399 -912
rect 12433 -946 12475 -912
rect 12509 -946 12551 -912
rect 12585 -946 12627 -912
rect 12661 -946 12703 -912
rect 12737 -946 12749 -912
rect 12310 -952 12749 -946
rect 8711 -2433 8717 -2381
rect 8769 -2433 8781 -2381
rect 8833 -2433 8839 -2381
rect 13260 -7040 13288 -7012
rect 14429 -7926 14457 -7898
rect 13634 -7974 13662 -7946
rect 14072 -8266 14100 -8238
rect 13265 -8570 13293 -8542
rect 13244 -8912 13272 -8884
rect 13347 -9239 13375 -9211
rect 14822 -10026 14874 -10020
rect 14822 -10090 14874 -10078
rect 14822 -10148 14874 -10142
<< via1 >>
rect 7995 9767 8047 9819
rect 8105 9767 8157 9819
rect 7995 9676 8047 9728
rect 8105 9676 8157 9728
rect 7995 9585 8047 9637
rect 8105 9585 8157 9637
rect 7995 9494 8047 9546
rect 8105 9494 8157 9546
rect 7995 9403 8047 9455
rect 8105 9403 8157 9455
rect 9213 9767 9265 9819
rect 9305 9767 9357 9819
rect 9397 9767 9449 9819
rect 9213 9676 9265 9728
rect 9305 9676 9357 9728
rect 9397 9676 9449 9728
rect 9213 9585 9265 9637
rect 9305 9585 9357 9637
rect 9397 9585 9449 9637
rect 9213 9494 9265 9546
rect 9305 9494 9357 9546
rect 9397 9494 9449 9546
rect 9213 9403 9265 9455
rect 9305 9403 9357 9455
rect 9397 9403 9449 9455
rect 1158 8586 1210 8589
rect -724 7981 -672 8033
rect -659 7981 -607 8033
rect -594 7981 -542 8033
rect -529 7981 -477 8033
rect -464 7981 -412 8033
rect -399 7981 -347 8033
rect -334 7981 -282 8033
rect -724 7909 -672 7961
rect -659 7909 -607 7961
rect -594 7909 -542 7961
rect -529 7909 -477 7961
rect -464 7909 -412 7961
rect -399 7909 -347 7961
rect -334 7909 -282 7961
rect -724 7837 -672 7889
rect -659 7837 -607 7889
rect -594 7837 -542 7889
rect -529 7837 -477 7889
rect -464 7837 -412 7889
rect -399 7837 -347 7889
rect -334 7837 -282 7889
rect -724 7765 -672 7817
rect -659 7765 -607 7817
rect -594 7765 -542 7817
rect -529 7765 -477 7817
rect -464 7765 -412 7817
rect -399 7765 -347 7817
rect -334 7765 -282 7817
rect -724 7693 -672 7745
rect -659 7693 -607 7745
rect -594 7693 -542 7745
rect -529 7693 -477 7745
rect -464 7693 -412 7745
rect -399 7693 -347 7745
rect -334 7693 -282 7745
rect -724 7283 -672 7335
rect -658 7283 -606 7335
rect -593 7283 -541 7335
rect -528 7283 -476 7335
rect -463 7283 -411 7335
rect -398 7283 -346 7335
rect -333 7283 -281 7335
rect -724 7203 -672 7255
rect -658 7203 -606 7255
rect -593 7203 -541 7255
rect -528 7203 -476 7255
rect -463 7203 -411 7255
rect -398 7203 -346 7255
rect -333 7203 -281 7255
rect -724 7123 -672 7175
rect -658 7123 -606 7175
rect -593 7123 -541 7175
rect -528 7123 -476 7175
rect -463 7123 -411 7175
rect -398 7123 -346 7175
rect -333 7123 -281 7175
rect 1158 8552 1173 8586
rect 1173 8552 1207 8586
rect 1207 8552 1210 8586
rect 1158 8537 1210 8552
rect 1224 8586 1276 8595
rect 1288 8586 1340 8595
rect 1352 8586 1404 8595
rect 1416 8586 1468 8595
rect 1480 8586 1532 8595
rect 1544 8586 1596 8595
rect 1224 8552 1245 8586
rect 1245 8552 1276 8586
rect 1288 8552 1317 8586
rect 1317 8552 1340 8586
rect 1352 8552 1389 8586
rect 1389 8552 1404 8586
rect 1416 8552 1423 8586
rect 1423 8552 1461 8586
rect 1461 8552 1468 8586
rect 1480 8552 1495 8586
rect 1495 8552 1532 8586
rect 1544 8552 1567 8586
rect 1567 8552 1596 8586
rect 1224 8543 1276 8552
rect 1288 8543 1340 8552
rect 1352 8543 1404 8552
rect 1416 8543 1468 8552
rect 1480 8543 1532 8552
rect 1544 8543 1596 8552
rect 1158 8496 1210 8525
rect 1158 8473 1167 8496
rect 1167 8473 1201 8496
rect 1201 8473 1210 8496
rect 1158 8424 1210 8461
rect 2049 8472 2101 8483
rect 2113 8472 2165 8483
rect 2177 8472 2229 8483
rect 2241 8472 2293 8483
rect 2305 8472 2357 8483
rect 2049 8438 2086 8472
rect 2086 8438 2101 8472
rect 2113 8438 2120 8472
rect 2120 8438 2158 8472
rect 2158 8438 2165 8472
rect 2177 8438 2192 8472
rect 2192 8438 2229 8472
rect 2241 8438 2264 8472
rect 2264 8438 2293 8472
rect 2305 8438 2336 8472
rect 2336 8438 2357 8472
rect 2049 8431 2101 8438
rect 2113 8431 2165 8438
rect 2177 8431 2229 8438
rect 2241 8431 2293 8438
rect 2305 8431 2357 8438
rect 2369 8472 2421 8483
rect 2369 8438 2374 8472
rect 2374 8438 2408 8472
rect 2408 8438 2421 8472
rect 2369 8431 2421 8438
rect 2433 8472 2485 8483
rect 2433 8438 2446 8472
rect 2446 8438 2480 8472
rect 2480 8438 2485 8472
rect 2433 8431 2485 8438
rect 2497 8472 2549 8483
rect 2561 8472 2613 8483
rect 2625 8472 2677 8483
rect 2689 8472 2741 8483
rect 2753 8472 2805 8483
rect 2497 8438 2518 8472
rect 2518 8438 2549 8472
rect 2561 8438 2590 8472
rect 2590 8438 2613 8472
rect 2625 8438 2662 8472
rect 2662 8438 2677 8472
rect 2689 8438 2696 8472
rect 2696 8438 2734 8472
rect 2734 8438 2741 8472
rect 2753 8438 2768 8472
rect 2768 8438 2805 8472
rect 2497 8431 2549 8438
rect 2561 8431 2613 8438
rect 2625 8431 2677 8438
rect 2689 8431 2741 8438
rect 2753 8431 2805 8438
rect 1158 8409 1167 8424
rect 1167 8409 1201 8424
rect 1201 8409 1210 8424
rect 1158 8390 1167 8397
rect 1167 8390 1201 8397
rect 1201 8390 1210 8397
rect 1158 8352 1210 8390
rect 1158 8345 1167 8352
rect 1167 8345 1201 8352
rect 1201 8345 1210 8352
rect 1158 8318 1167 8333
rect 1167 8318 1201 8333
rect 1201 8318 1210 8333
rect 1158 8281 1210 8318
rect 1288 8272 1340 8324
rect 1352 8316 1404 8324
rect 1352 8282 1366 8316
rect 1366 8282 1400 8316
rect 1400 8282 1404 8316
rect 1352 8272 1404 8282
rect 1416 8316 1468 8324
rect 1480 8316 1532 8324
rect 1544 8316 1596 8324
rect 1416 8282 1438 8316
rect 1438 8282 1468 8316
rect 1480 8282 1510 8316
rect 1510 8282 1532 8316
rect 1544 8282 1582 8316
rect 1582 8282 1596 8316
rect 1416 8272 1468 8282
rect 1480 8272 1532 8282
rect 1544 8272 1596 8282
rect 1158 8246 1167 8269
rect 1167 8246 1201 8269
rect 1201 8246 1210 8269
rect 1158 8217 1210 8246
rect 1158 8174 1167 8205
rect 1167 8174 1201 8205
rect 1201 8174 1210 8205
rect 1158 8153 1210 8174
rect 4321 8261 4373 8263
rect 4321 8227 4330 8261
rect 4330 8227 4364 8261
rect 4364 8227 4373 8261
rect 4321 8211 4373 8227
rect 4321 8184 4373 8199
rect 1158 8136 1210 8141
rect 1158 8102 1167 8136
rect 1167 8102 1201 8136
rect 1201 8102 1210 8136
rect 2049 8160 2101 8169
rect 2113 8160 2165 8169
rect 2177 8160 2229 8169
rect 2241 8160 2293 8169
rect 2305 8160 2357 8169
rect 2049 8126 2086 8160
rect 2086 8126 2101 8160
rect 2113 8126 2120 8160
rect 2120 8126 2158 8160
rect 2158 8126 2165 8160
rect 2177 8126 2192 8160
rect 2192 8126 2229 8160
rect 2241 8126 2264 8160
rect 2264 8126 2293 8160
rect 2305 8126 2336 8160
rect 2336 8126 2357 8160
rect 2049 8117 2101 8126
rect 2113 8117 2165 8126
rect 2177 8117 2229 8126
rect 2241 8117 2293 8126
rect 2305 8117 2357 8126
rect 2369 8160 2421 8169
rect 2369 8126 2374 8160
rect 2374 8126 2408 8160
rect 2408 8126 2421 8160
rect 2369 8117 2421 8126
rect 2433 8160 2485 8169
rect 2433 8126 2446 8160
rect 2446 8126 2480 8160
rect 2480 8126 2485 8160
rect 2433 8117 2485 8126
rect 2497 8160 2549 8169
rect 2561 8160 2613 8169
rect 2625 8160 2677 8169
rect 2689 8160 2741 8169
rect 2753 8160 2805 8169
rect 2497 8126 2518 8160
rect 2518 8126 2549 8160
rect 2561 8126 2590 8160
rect 2590 8126 2613 8160
rect 2625 8126 2662 8160
rect 2662 8126 2677 8160
rect 2689 8126 2696 8160
rect 2696 8126 2734 8160
rect 2734 8126 2741 8160
rect 2753 8126 2768 8160
rect 2768 8126 2805 8160
rect 4321 8150 4330 8184
rect 4330 8150 4364 8184
rect 4364 8150 4373 8184
rect 4321 8147 4373 8150
rect 2497 8117 2549 8126
rect 2561 8117 2613 8126
rect 2625 8117 2677 8126
rect 2689 8117 2741 8126
rect 2753 8117 2805 8126
rect 1158 8089 1210 8102
rect 1158 8064 1210 8077
rect 1158 8030 1167 8064
rect 1167 8030 1201 8064
rect 1201 8030 1210 8064
rect 1158 8025 1210 8030
rect 14143 8315 14195 8367
rect 14143 8248 14195 8300
rect 1158 7992 1210 8013
rect 1158 7961 1167 7992
rect 1167 7961 1201 7992
rect 1201 7961 1210 7992
rect 1288 7964 1340 8016
rect 1352 8004 1404 8016
rect 1352 7970 1366 8004
rect 1366 7970 1400 8004
rect 1400 7970 1404 8004
rect 1352 7964 1404 7970
rect 1416 8004 1468 8016
rect 1480 8004 1532 8016
rect 1544 8004 1596 8016
rect 1416 7970 1438 8004
rect 1438 7970 1468 8004
rect 1480 7970 1510 8004
rect 1510 7970 1532 8004
rect 1544 7970 1582 8004
rect 1582 7970 1596 8004
rect 1416 7964 1468 7970
rect 1480 7964 1532 7970
rect 1544 7964 1596 7970
rect 1158 7920 1210 7949
rect 1158 7897 1167 7920
rect 1167 7897 1201 7920
rect 1201 7897 1210 7920
rect 1158 7848 1210 7885
rect 1158 7833 1167 7848
rect 1167 7833 1201 7848
rect 1201 7833 1210 7848
rect 1158 7814 1167 7821
rect 1167 7814 1201 7821
rect 1201 7814 1210 7821
rect 1158 7776 1210 7814
rect 2069 7848 2121 7857
rect 2069 7814 2086 7848
rect 2086 7814 2120 7848
rect 2120 7814 2121 7848
rect 2069 7805 2121 7814
rect 2133 7848 2185 7857
rect 2197 7848 2249 7857
rect 2261 7848 2313 7857
rect 2325 7848 2377 7857
rect 2389 7848 2441 7857
rect 2453 7848 2505 7857
rect 2133 7814 2158 7848
rect 2158 7814 2185 7848
rect 2197 7814 2230 7848
rect 2230 7814 2249 7848
rect 2261 7814 2264 7848
rect 2264 7814 2302 7848
rect 2302 7814 2313 7848
rect 2325 7814 2336 7848
rect 2336 7814 2374 7848
rect 2374 7814 2377 7848
rect 2389 7814 2408 7848
rect 2408 7814 2441 7848
rect 2453 7814 2480 7848
rect 2480 7814 2505 7848
rect 2133 7805 2185 7814
rect 2197 7805 2249 7814
rect 2261 7805 2313 7814
rect 2325 7805 2377 7814
rect 2389 7805 2441 7814
rect 2453 7805 2505 7814
rect 2517 7848 2569 7857
rect 2517 7814 2518 7848
rect 2518 7814 2552 7848
rect 2552 7814 2569 7848
rect 2517 7805 2569 7814
rect 2581 7848 2633 7857
rect 2581 7814 2590 7848
rect 2590 7814 2624 7848
rect 2624 7814 2633 7848
rect 2581 7805 2633 7814
rect 2645 7848 2697 7857
rect 2645 7814 2662 7848
rect 2662 7814 2696 7848
rect 2696 7814 2697 7848
rect 2645 7805 2697 7814
rect 2709 7848 2761 7857
rect 2773 7848 2825 7857
rect 2837 7848 2889 7857
rect 2709 7814 2734 7848
rect 2734 7814 2761 7848
rect 2773 7814 2806 7848
rect 2806 7814 2825 7848
rect 2837 7814 2840 7848
rect 2840 7814 2878 7848
rect 2878 7814 2889 7848
rect 2709 7805 2761 7814
rect 2773 7805 2825 7814
rect 2837 7805 2889 7814
rect 1158 7769 1167 7776
rect 1167 7769 1201 7776
rect 1201 7769 1210 7776
rect 1158 7742 1167 7757
rect 1167 7742 1201 7757
rect 1201 7742 1210 7757
rect 1158 7705 1210 7742
rect 1158 7670 1167 7693
rect 1167 7670 1201 7693
rect 1201 7670 1210 7693
rect 1158 7641 1210 7670
rect 1288 7649 1340 7701
rect 1352 7692 1404 7701
rect 1352 7658 1366 7692
rect 1366 7658 1400 7692
rect 1400 7658 1404 7692
rect 1352 7649 1404 7658
rect 1416 7692 1468 7701
rect 1480 7692 1532 7701
rect 1544 7692 1596 7701
rect 1416 7658 1438 7692
rect 1438 7658 1468 7692
rect 1480 7658 1510 7692
rect 1510 7658 1532 7692
rect 1544 7658 1582 7692
rect 1582 7658 1596 7692
rect 1416 7649 1468 7658
rect 1480 7649 1532 7658
rect 1544 7649 1596 7658
rect 1158 7598 1167 7629
rect 1167 7598 1201 7629
rect 1201 7598 1210 7629
rect 1158 7577 1210 7598
rect 1158 7560 1210 7565
rect 1158 7526 1167 7560
rect 1167 7526 1201 7560
rect 1201 7526 1210 7560
rect 1158 7513 1210 7526
rect 1158 7488 1210 7501
rect 2069 7536 2121 7545
rect 2069 7502 2086 7536
rect 2086 7502 2120 7536
rect 2120 7502 2121 7536
rect 2069 7493 2121 7502
rect 2133 7536 2185 7545
rect 2197 7536 2249 7545
rect 2261 7536 2313 7545
rect 2325 7536 2377 7545
rect 2389 7536 2441 7545
rect 2453 7536 2505 7545
rect 2133 7502 2158 7536
rect 2158 7502 2185 7536
rect 2197 7502 2230 7536
rect 2230 7502 2249 7536
rect 2261 7502 2264 7536
rect 2264 7502 2302 7536
rect 2302 7502 2313 7536
rect 2325 7502 2336 7536
rect 2336 7502 2374 7536
rect 2374 7502 2377 7536
rect 2389 7502 2408 7536
rect 2408 7502 2441 7536
rect 2453 7502 2480 7536
rect 2480 7502 2505 7536
rect 2133 7493 2185 7502
rect 2197 7493 2249 7502
rect 2261 7493 2313 7502
rect 2325 7493 2377 7502
rect 2389 7493 2441 7502
rect 2453 7493 2505 7502
rect 2517 7536 2569 7545
rect 2517 7502 2518 7536
rect 2518 7502 2552 7536
rect 2552 7502 2569 7536
rect 2517 7493 2569 7502
rect 2581 7536 2633 7545
rect 2581 7502 2590 7536
rect 2590 7502 2624 7536
rect 2624 7502 2633 7536
rect 2581 7493 2633 7502
rect 2645 7536 2697 7545
rect 2645 7502 2662 7536
rect 2662 7502 2696 7536
rect 2696 7502 2697 7536
rect 2645 7493 2697 7502
rect 2709 7536 2761 7545
rect 2773 7536 2825 7545
rect 2837 7536 2889 7545
rect 2709 7502 2734 7536
rect 2734 7502 2761 7536
rect 2773 7502 2806 7536
rect 2806 7502 2825 7536
rect 2837 7502 2840 7536
rect 2840 7502 2878 7536
rect 2878 7502 2889 7536
rect 2709 7493 2761 7502
rect 2773 7493 2825 7502
rect 2837 7493 2889 7502
rect 1158 7454 1167 7488
rect 1167 7454 1201 7488
rect 1201 7454 1210 7488
rect 1158 7449 1210 7454
rect 1158 7416 1210 7437
rect 4955 8134 5007 8186
rect 4955 8058 5007 8110
rect 4955 7982 5007 8034
rect 4955 7906 5007 7958
rect 4955 7830 5007 7882
rect 4955 7754 5007 7806
rect 14143 8181 14195 8233
rect 14143 8114 14195 8166
rect 14143 8047 14195 8099
rect 14143 7980 14195 8032
rect 14143 7913 14195 7965
rect 14143 7845 14195 7897
rect 14143 7777 14195 7829
rect 1158 7385 1167 7416
rect 1167 7385 1201 7416
rect 1201 7385 1210 7416
rect 1288 7380 1340 7389
rect 1158 7344 1210 7373
rect 1158 7321 1167 7344
rect 1167 7321 1201 7344
rect 1201 7321 1210 7344
rect 1288 7346 1294 7380
rect 1294 7346 1328 7380
rect 1328 7346 1340 7380
rect 1288 7337 1340 7346
rect 1352 7380 1404 7389
rect 1352 7346 1366 7380
rect 1366 7346 1400 7380
rect 1400 7346 1404 7380
rect 1352 7337 1404 7346
rect 1416 7380 1468 7389
rect 1480 7380 1532 7389
rect 1544 7380 1596 7389
rect 1416 7346 1438 7380
rect 1438 7346 1468 7380
rect 1480 7346 1510 7380
rect 1510 7346 1532 7380
rect 1544 7346 1582 7380
rect 1582 7346 1596 7380
rect 1416 7337 1468 7346
rect 1480 7337 1532 7346
rect 1544 7337 1596 7346
rect 1284 7269 1336 7321
rect 1349 7269 1401 7321
rect 1414 7269 1466 7321
rect 1479 7269 1531 7321
rect 1544 7269 1596 7321
rect 13398 7322 13450 7374
rect 13472 7322 13524 7374
rect 13545 7322 13597 7374
rect 13618 7322 13670 7374
rect 13691 7322 13743 7374
rect 13764 7322 13816 7374
rect 13398 7250 13450 7302
rect 13472 7250 13524 7302
rect 13545 7250 13597 7302
rect 13618 7250 13670 7302
rect 13691 7250 13743 7302
rect 13764 7250 13816 7302
rect 13398 7178 13450 7230
rect 13472 7178 13524 7230
rect 13545 7178 13597 7230
rect 13618 7178 13670 7230
rect 13691 7178 13743 7230
rect 13764 7178 13816 7230
rect 13398 7106 13450 7158
rect 13472 7106 13524 7158
rect 13545 7106 13597 7158
rect 13618 7106 13670 7158
rect 13691 7106 13743 7158
rect 13764 7106 13816 7158
rect 2065 6940 2117 6992
rect 2129 6940 2181 6992
rect 13398 7034 13450 7086
rect 13472 7034 13524 7086
rect 13545 7034 13597 7086
rect 13618 7034 13670 7086
rect 13691 7034 13743 7086
rect 13764 7034 13816 7086
rect 13398 6962 13450 7014
rect 13472 6962 13524 7014
rect 13545 6962 13597 7014
rect 13618 6962 13670 7014
rect 13691 6962 13743 7014
rect 13764 6962 13816 7014
rect -126 6739 -74 6791
rect -855 6715 -803 6721
rect -855 6681 -849 6715
rect -849 6681 -815 6715
rect -815 6681 -803 6715
rect -855 6669 -803 6681
rect -126 6675 -74 6727
rect 193 6788 245 6840
rect 193 6724 245 6776
rect 3605 6754 3657 6806
rect 3669 6754 3721 6806
rect -855 6635 -803 6657
rect -855 6605 -849 6635
rect -849 6605 -815 6635
rect -815 6605 -803 6635
rect 1837 6648 1889 6700
rect 1905 6648 1957 6700
rect 1973 6648 2025 6700
rect 2040 6648 2092 6700
rect 2107 6648 2159 6700
rect 3639 6674 3691 6726
rect 3703 6674 3755 6726
rect 2280 6536 2332 6588
rect 2344 6536 2396 6588
rect 2408 6536 2460 6588
rect 2280 6458 2332 6510
rect 2344 6458 2396 6510
rect 2408 6458 2460 6510
rect 2978 6546 3030 6551
rect 3050 6546 3102 6551
rect 3122 6546 3174 6551
rect 3194 6546 3246 6551
rect 2978 6512 3004 6546
rect 3004 6512 3030 6546
rect 3050 6512 3079 6546
rect 3079 6512 3102 6546
rect 3122 6512 3154 6546
rect 3154 6512 3174 6546
rect 3194 6512 3229 6546
rect 3229 6512 3246 6546
rect 2978 6499 3030 6512
rect 3050 6499 3102 6512
rect 3122 6499 3174 6512
rect 3194 6499 3246 6512
rect 3266 6499 3318 6551
rect 2978 6472 3030 6479
rect 3050 6472 3102 6479
rect 3122 6472 3174 6479
rect 3194 6472 3246 6479
rect 2978 6438 3004 6472
rect 3004 6438 3030 6472
rect 3050 6438 3079 6472
rect 3079 6438 3102 6472
rect 3122 6438 3154 6472
rect 3154 6438 3174 6472
rect 3194 6438 3229 6472
rect 3229 6438 3246 6472
rect 2978 6427 3030 6438
rect 3050 6427 3102 6438
rect 3122 6427 3174 6438
rect 3194 6427 3246 6438
rect 3266 6427 3318 6479
rect 2978 6398 3030 6407
rect 3050 6398 3102 6407
rect 3122 6398 3174 6407
rect 3194 6398 3246 6407
rect 2978 6364 3004 6398
rect 3004 6364 3030 6398
rect 3050 6364 3079 6398
rect 3079 6364 3102 6398
rect 3122 6364 3154 6398
rect 3154 6364 3174 6398
rect 3194 6364 3229 6398
rect 3229 6364 3246 6398
rect 2298 6308 2350 6360
rect 2362 6308 2414 6360
rect 2426 6308 2478 6360
rect 2298 6230 2350 6282
rect 2362 6230 2414 6282
rect 2426 6230 2478 6282
rect 2978 6355 3030 6364
rect 3050 6355 3102 6364
rect 3122 6355 3174 6364
rect 3194 6355 3246 6364
rect 3266 6355 3318 6407
rect 2978 6324 3030 6335
rect 3050 6324 3102 6335
rect 3122 6324 3174 6335
rect 3194 6324 3246 6335
rect 2978 6290 3004 6324
rect 3004 6290 3030 6324
rect 3050 6290 3079 6324
rect 3079 6290 3102 6324
rect 3122 6290 3154 6324
rect 3154 6290 3174 6324
rect 3194 6290 3229 6324
rect 3229 6290 3246 6324
rect 2978 6283 3030 6290
rect 3050 6283 3102 6290
rect 3122 6283 3174 6290
rect 3194 6283 3246 6290
rect 3266 6283 3318 6335
rect 2978 6250 3030 6263
rect 3050 6250 3102 6263
rect 3122 6250 3174 6263
rect 3194 6250 3246 6263
rect 2978 6216 3004 6250
rect 3004 6216 3030 6250
rect 3050 6216 3079 6250
rect 3079 6216 3102 6250
rect 3122 6216 3154 6250
rect 3154 6216 3174 6250
rect 3194 6216 3229 6250
rect 3229 6216 3246 6250
rect 2978 6211 3030 6216
rect 3050 6211 3102 6216
rect 3122 6211 3174 6216
rect 3194 6211 3246 6216
rect 3266 6211 3318 6263
rect 962 6138 1014 6190
rect 1026 6138 1078 6190
rect 2805 5819 2857 5871
rect 2000 5704 2052 5756
rect 2064 5704 2116 5756
rect 2805 5755 2857 5807
rect 2479 5669 2531 5721
rect 2543 5669 2595 5721
rect 3712 6319 3764 6371
rect 3712 6255 3764 6307
rect 3448 5685 3500 5737
rect 3448 5621 3500 5673
rect 3721 6135 3773 6187
rect 3721 6071 3773 6123
rect 3541 5497 3593 5549
rect 3605 5497 3657 5549
rect 3901 6197 3953 6249
rect 3965 6197 4017 6249
rect 4036 5903 4088 5955
rect 4036 5839 4088 5891
rect 4577 5961 4629 6013
rect 4645 5961 4697 6013
rect 4577 5883 4629 5935
rect 4645 5883 4697 5935
rect 13398 5969 13450 6021
rect 13472 5969 13524 6021
rect 13545 5969 13597 6021
rect 13618 5969 13670 6021
rect 13691 5969 13743 6021
rect 13764 5969 13816 6021
rect 13398 5897 13450 5949
rect 13472 5897 13524 5949
rect 13545 5897 13597 5949
rect 13618 5897 13670 5949
rect 13691 5897 13743 5949
rect 13764 5897 13816 5949
rect 4415 5581 4467 5633
rect 4483 5581 4535 5633
rect 13398 5825 13450 5877
rect 13472 5825 13524 5877
rect 13545 5825 13597 5877
rect 13618 5825 13670 5877
rect 13691 5825 13743 5877
rect 13764 5825 13816 5877
rect 13398 5753 13450 5805
rect 13472 5753 13524 5805
rect 13545 5753 13597 5805
rect 13618 5753 13670 5805
rect 13691 5753 13743 5805
rect 13764 5753 13816 5805
rect 13398 5681 13450 5733
rect 13472 5681 13524 5733
rect 13545 5681 13597 5733
rect 13618 5681 13670 5733
rect 13691 5681 13743 5733
rect 13764 5681 13816 5733
rect 13398 5609 13450 5661
rect 13472 5609 13524 5661
rect 13545 5609 13597 5661
rect 13618 5609 13670 5661
rect 13691 5609 13743 5661
rect 13764 5609 13816 5661
rect 4415 5503 4467 5555
rect 4483 5503 4535 5555
rect 3491 5299 3543 5351
rect 3555 5299 3607 5351
rect 3784 5294 3836 5346
rect 3848 5294 3900 5346
rect 2160 5062 2212 5114
rect 2224 5062 2276 5114
rect 1959 4841 2011 4893
rect 2023 4841 2075 4893
rect 2908 4587 2960 4639
rect 3002 4587 3054 4639
rect 2908 4521 2960 4573
rect 3002 4521 3054 4573
rect 2908 4454 2960 4506
rect 3002 4454 3054 4506
rect 13983 5221 14035 5273
rect 13983 5154 14035 5206
rect 13983 5087 14035 5139
rect 4281 4559 4333 4611
rect 4281 4495 4333 4547
rect 4955 4995 5007 5047
rect 4955 4923 5007 4975
rect 4955 4850 5007 4902
rect 4955 4777 5007 4829
rect 4955 4704 5007 4756
rect 4955 4631 5007 4683
rect 13983 5020 14035 5072
rect 13983 4953 14035 5005
rect 13983 4886 14035 4938
rect 13983 4819 14035 4871
rect 13983 4751 14035 4803
rect 13983 4683 14035 4735
rect 13983 4615 14035 4667
rect 4955 4558 5007 4610
rect 4955 4485 5007 4537
rect 4369 4358 4421 4410
rect 4537 4358 4589 4410
rect 5081 4358 5133 4410
rect 5145 4358 5197 4410
rect 5658 4358 5710 4410
rect 5722 4358 5774 4410
rect 1857 3243 1909 3295
rect 1857 3179 1909 3231
rect 2191 3243 2243 3295
rect 2191 3179 2243 3231
rect 4369 4294 4421 4346
rect 4537 4294 4589 4346
rect 5921 4241 5973 4293
rect 6025 4241 6077 4293
rect 6128 4241 6180 4293
rect 12928 4217 12980 4269
rect 12992 4217 13044 4269
rect 13552 4217 13604 4269
rect 13616 4217 13668 4269
rect 10318 4144 10370 4196
rect 10382 4144 10434 4196
rect 4308 3896 4360 3948
rect 4372 3896 4424 3948
rect 12939 3899 12991 3951
rect 13003 3899 13055 3951
rect 13428 4107 13480 4129
rect 13428 4077 13437 4107
rect 13437 4077 13471 4107
rect 13471 4077 13480 4107
rect 13428 4034 13480 4065
rect 13720 4057 13768 4091
rect 13768 4057 13772 4091
rect 13428 4013 13437 4034
rect 13437 4013 13471 4034
rect 13471 4013 13480 4034
rect 13720 4039 13772 4057
rect 9119 3621 9171 3673
rect 9194 3621 9246 3673
rect 9268 3621 9320 3673
rect 9342 3621 9394 3673
rect 9119 3557 9171 3609
rect 9194 3557 9246 3609
rect 9268 3557 9320 3609
rect 9342 3557 9394 3609
rect 10247 3626 10299 3678
rect 10315 3626 10367 3678
rect 10383 3626 10435 3678
rect 10451 3626 10503 3678
rect 10519 3626 10571 3678
rect 10587 3626 10639 3678
rect 10654 3626 10706 3678
rect 10247 3554 10299 3606
rect 10315 3554 10367 3606
rect 10383 3554 10435 3606
rect 10451 3554 10503 3606
rect 10519 3554 10571 3606
rect 10587 3554 10639 3606
rect 10654 3554 10706 3606
rect 12939 3657 12991 3709
rect 13003 3657 13055 3709
rect 12930 3552 12982 3604
rect 12994 3552 13046 3604
rect 4176 3388 4228 3440
rect 5450 3435 5502 3487
rect 13113 3462 13165 3514
rect 4176 3324 4228 3376
rect 5450 3371 5502 3423
rect 13113 3398 13165 3450
rect 12100 3286 12152 3291
rect 12100 3252 12116 3286
rect 12116 3252 12150 3286
rect 12150 3252 12152 3286
rect 12100 3239 12152 3252
rect 12169 3286 12221 3291
rect 12238 3286 12290 3291
rect 12307 3286 12359 3291
rect 12376 3286 12428 3291
rect 12445 3286 12497 3291
rect 12514 3286 12566 3291
rect 12583 3286 12635 3291
rect 12651 3286 12703 3291
rect 12719 3286 12771 3291
rect 12169 3252 12188 3286
rect 12188 3252 12221 3286
rect 12238 3252 12260 3286
rect 12260 3252 12290 3286
rect 12307 3252 12332 3286
rect 12332 3252 12359 3286
rect 12376 3252 12404 3286
rect 12404 3252 12428 3286
rect 12445 3252 12480 3286
rect 12480 3252 12497 3286
rect 12514 3252 12558 3286
rect 12558 3252 12566 3286
rect 12583 3252 12592 3286
rect 12592 3252 12635 3286
rect 12651 3252 12669 3286
rect 12669 3252 12703 3286
rect 12719 3252 12746 3286
rect 12746 3252 12771 3286
rect 12169 3239 12221 3252
rect 12238 3239 12290 3252
rect 12307 3239 12359 3252
rect 12376 3239 12428 3252
rect 12445 3239 12497 3252
rect 12514 3239 12566 3252
rect 12583 3239 12635 3252
rect 12651 3239 12703 3252
rect 12719 3239 12771 3252
rect 12787 3286 12839 3291
rect 12787 3252 12789 3286
rect 12789 3252 12823 3286
rect 12823 3252 12839 3286
rect 12787 3239 12839 3252
rect 12855 3286 12907 3291
rect 12855 3252 12866 3286
rect 12866 3252 12900 3286
rect 12900 3252 12907 3286
rect 12855 3239 12907 3252
rect 12100 3170 12152 3203
rect 12100 3151 12116 3170
rect 12116 3151 12150 3170
rect 12150 3151 12152 3170
rect 12169 3170 12221 3203
rect 12238 3170 12290 3203
rect 12307 3170 12359 3203
rect 12376 3170 12428 3203
rect 12445 3194 12497 3203
rect 12514 3194 12566 3203
rect 12583 3194 12635 3203
rect 12651 3194 12703 3203
rect 12719 3194 12771 3203
rect 12169 3151 12188 3170
rect 12188 3151 12221 3170
rect 12238 3151 12260 3170
rect 12260 3151 12290 3170
rect 12307 3151 12332 3170
rect 12332 3151 12359 3170
rect 12376 3151 12404 3170
rect 12404 3151 12428 3170
rect 12445 3160 12480 3194
rect 12480 3160 12497 3194
rect 12514 3160 12558 3194
rect 12558 3160 12566 3194
rect 12583 3160 12592 3194
rect 12592 3160 12635 3194
rect 12651 3160 12669 3194
rect 12669 3160 12703 3194
rect 12719 3160 12746 3194
rect 12746 3160 12771 3194
rect 12445 3151 12497 3160
rect 12514 3151 12566 3160
rect 12583 3151 12635 3160
rect 12651 3151 12703 3160
rect 12719 3151 12771 3160
rect 12787 3194 12839 3203
rect 12787 3160 12789 3194
rect 12789 3160 12823 3194
rect 12823 3160 12839 3194
rect 12787 3151 12839 3160
rect 12855 3194 12907 3203
rect 12855 3160 12866 3194
rect 12866 3160 12900 3194
rect 12900 3160 12907 3194
rect 12855 3151 12907 3160
rect 12100 3063 12152 3115
rect 12169 3063 12221 3115
rect 12238 3063 12290 3115
rect 12307 3063 12359 3115
rect 12376 3063 12428 3115
rect 12445 3102 12497 3115
rect 12514 3102 12566 3115
rect 12583 3102 12635 3115
rect 12651 3102 12703 3115
rect 12719 3102 12771 3115
rect 12445 3068 12480 3102
rect 12480 3068 12497 3102
rect 12514 3068 12558 3102
rect 12558 3068 12566 3102
rect 12583 3068 12592 3102
rect 12592 3068 12635 3102
rect 12651 3068 12669 3102
rect 12669 3068 12703 3102
rect 12719 3068 12746 3102
rect 12746 3068 12771 3102
rect 12445 3063 12497 3068
rect 12514 3063 12566 3068
rect 12583 3063 12635 3068
rect 12651 3063 12703 3068
rect 12719 3063 12771 3068
rect 12787 3102 12839 3115
rect 12787 3068 12789 3102
rect 12789 3068 12823 3102
rect 12823 3068 12839 3102
rect 12787 3063 12839 3068
rect 12855 3102 12907 3115
rect 12855 3068 12866 3102
rect 12866 3068 12900 3102
rect 12900 3068 12907 3102
rect 12855 3063 12907 3068
rect 4717 2889 4769 2941
rect 9024 2934 9076 2986
rect 9104 2934 9156 2986
rect 9184 2934 9236 2986
rect 9263 2934 9315 2986
rect 9342 2934 9394 2986
rect 4717 2825 4769 2877
rect 9024 2858 9076 2910
rect 9104 2858 9156 2910
rect 9184 2858 9236 2910
rect 9263 2858 9315 2910
rect 9342 2858 9394 2910
rect 9024 2782 9076 2834
rect 9104 2782 9156 2834
rect 9184 2782 9236 2834
rect 9263 2782 9315 2834
rect 9342 2782 9394 2834
rect 9024 2706 9076 2758
rect 9104 2706 9156 2758
rect 9184 2706 9236 2758
rect 9263 2706 9315 2758
rect 9342 2706 9394 2758
rect 11553 2922 11564 2956
rect 11564 2922 11598 2956
rect 11598 2922 11605 2956
rect 11553 2904 11605 2922
rect 11623 2922 11640 2956
rect 11640 2922 11674 2956
rect 11674 2922 11675 2956
rect 11623 2904 11675 2922
rect 11693 2922 11716 2956
rect 11716 2922 11745 2956
rect 11693 2904 11745 2922
rect 11553 2880 11605 2891
rect 11553 2846 11564 2880
rect 11564 2846 11598 2880
rect 11598 2846 11605 2880
rect 11553 2839 11605 2846
rect 11623 2880 11675 2891
rect 11623 2846 11640 2880
rect 11640 2846 11674 2880
rect 11674 2846 11675 2880
rect 11623 2839 11675 2846
rect 11693 2880 11745 2891
rect 11693 2846 11716 2880
rect 11716 2846 11745 2880
rect 11693 2839 11745 2846
rect 11553 2804 11605 2826
rect 11553 2774 11564 2804
rect 11564 2774 11598 2804
rect 11598 2774 11605 2804
rect 11623 2804 11675 2826
rect 11623 2774 11640 2804
rect 11640 2774 11674 2804
rect 11674 2774 11675 2804
rect 11693 2804 11745 2826
rect 11693 2774 11716 2804
rect 11716 2774 11745 2804
rect 11553 2728 11605 2761
rect 11553 2709 11564 2728
rect 11564 2709 11598 2728
rect 11598 2709 11605 2728
rect 11623 2728 11675 2761
rect 11623 2709 11640 2728
rect 11640 2709 11674 2728
rect 11674 2709 11675 2728
rect 11693 2728 11745 2761
rect 11693 2709 11716 2728
rect 11716 2709 11745 2728
rect 11553 2694 11564 2696
rect 11564 2694 11598 2696
rect 11598 2694 11605 2696
rect 11553 2652 11605 2694
rect 11553 2644 11564 2652
rect 11564 2644 11598 2652
rect 11598 2644 11605 2652
rect 11623 2694 11640 2696
rect 11640 2694 11674 2696
rect 11674 2694 11675 2696
rect 11623 2652 11675 2694
rect 11623 2644 11640 2652
rect 11640 2644 11674 2652
rect 11674 2644 11675 2652
rect 11693 2694 11716 2696
rect 11716 2694 11745 2696
rect 11693 2652 11745 2694
rect 11693 2644 11716 2652
rect 11716 2644 11745 2652
rect 11553 2618 11564 2631
rect 11564 2618 11598 2631
rect 11598 2618 11605 2631
rect 11553 2579 11605 2618
rect 11623 2618 11640 2631
rect 11640 2618 11674 2631
rect 11674 2618 11675 2631
rect 11623 2579 11675 2618
rect 11693 2618 11716 2631
rect 11716 2618 11745 2631
rect 11693 2579 11745 2618
rect 11553 2542 11564 2566
rect 11564 2542 11598 2566
rect 11598 2542 11605 2566
rect 11553 2514 11605 2542
rect 11623 2542 11640 2566
rect 11640 2542 11674 2566
rect 11674 2542 11675 2566
rect 11623 2514 11675 2542
rect 11693 2542 11716 2566
rect 11716 2542 11745 2566
rect 11693 2514 11745 2542
rect 11553 2466 11564 2500
rect 11564 2466 11598 2500
rect 11598 2466 11605 2500
rect 11553 2448 11605 2466
rect 11623 2466 11640 2500
rect 11640 2466 11674 2500
rect 11674 2466 11675 2500
rect 11623 2448 11675 2466
rect 11693 2466 11716 2500
rect 11716 2466 11745 2500
rect 11693 2448 11745 2466
rect 11553 2424 11605 2434
rect 11553 2390 11564 2424
rect 11564 2390 11598 2424
rect 11598 2390 11605 2424
rect 11553 2382 11605 2390
rect 11623 2424 11675 2434
rect 11623 2390 11640 2424
rect 11640 2390 11674 2424
rect 11674 2390 11675 2424
rect 11623 2382 11675 2390
rect 11693 2424 11745 2434
rect 11693 2390 11716 2424
rect 11716 2390 11745 2424
rect 11693 2382 11745 2390
rect 4177 2261 4229 2313
rect 4241 2261 4293 2313
rect 5144 2261 5196 2313
rect 5208 2261 5260 2313
rect 7601 2248 7653 2300
rect 7703 2248 7755 2300
rect 7804 2248 7856 2300
rect 13720 3975 13772 4027
rect 13549 3916 13601 3922
rect 13549 3882 13558 3916
rect 13558 3882 13592 3916
rect 13592 3882 13601 3916
rect 13549 3870 13601 3882
rect 13549 3842 13601 3858
rect 13549 3808 13558 3842
rect 13558 3808 13592 3842
rect 13592 3808 13601 3842
rect 13549 3806 13601 3808
rect 13868 3870 13920 3922
rect 13868 3799 13920 3851
rect 13868 3728 13920 3780
rect 13983 3938 14035 3944
rect 13983 3904 13986 3938
rect 13986 3904 14020 3938
rect 14020 3904 14035 3938
rect 13983 3892 14035 3904
rect 13983 3828 14035 3880
rect 13983 3804 14035 3816
rect 13983 3770 13986 3804
rect 13986 3770 14020 3804
rect 14020 3770 14035 3804
rect 13983 3764 14035 3770
rect 14063 3938 14115 3944
rect 14063 3904 14075 3938
rect 14075 3904 14109 3938
rect 14109 3904 14115 3938
rect 14063 3892 14115 3904
rect 14063 3846 14115 3855
rect 14063 3812 14075 3846
rect 14075 3812 14109 3846
rect 14109 3812 14115 3846
rect 14063 3803 14115 3812
rect 14143 3894 14195 3946
rect 14143 3816 14195 3868
rect 14063 3753 14115 3765
rect 13748 3632 13800 3684
rect 13812 3672 13864 3684
rect 13812 3638 13830 3672
rect 13830 3638 13864 3672
rect 13812 3632 13864 3638
rect 14063 3719 14075 3753
rect 14075 3719 14109 3753
rect 14109 3719 14115 3753
rect 14063 3713 14115 3719
rect 14143 3721 14195 3773
rect 14143 3657 14195 3709
rect 14135 3511 14187 3563
rect 14135 3447 14187 3499
rect 14073 3336 14125 3388
rect 14137 3336 14189 3388
rect 13875 3244 13927 3296
rect 13443 3149 13495 3201
rect 13507 3149 13559 3201
rect 13875 3152 13927 3204
rect 14017 3195 14069 3204
rect 14017 3161 14025 3195
rect 14025 3161 14059 3195
rect 14059 3161 14069 3195
rect 14017 3152 14069 3161
rect 14081 3195 14133 3204
rect 14081 3161 14114 3195
rect 14114 3161 14133 3195
rect 14081 3152 14133 3161
rect 13875 3060 13927 3112
rect 14073 3016 14125 3025
rect 14137 3016 14189 3025
rect 14073 2982 14107 3016
rect 14107 2982 14125 3016
rect 14137 2982 14141 3016
rect 14141 2982 14189 3016
rect 14073 2973 14125 2982
rect 14137 2973 14189 2982
rect 13908 2748 13960 2800
rect 13972 2748 14024 2800
rect 9091 2226 9143 2278
rect 9159 2226 9211 2278
rect 9227 2226 9279 2278
rect 9091 2141 9143 2193
rect 9159 2141 9211 2193
rect 9227 2141 9279 2193
rect 9496 2261 9548 2313
rect 9582 2261 9634 2313
rect 9496 2197 9548 2249
rect 9582 2197 9634 2249
rect 9091 2055 9143 2107
rect 9159 2055 9211 2107
rect 9227 2055 9279 2107
rect 3270 1936 3322 1988
rect 3388 1936 3440 1988
rect 3270 1858 3322 1910
rect 3388 1858 3440 1910
rect 3715 1960 3767 2012
rect 3715 1896 3767 1948
rect 4163 1960 4215 2012
rect 4163 1896 4215 1948
rect 4482 1899 4534 1951
rect 4482 1835 4534 1887
rect 5468 1537 5520 1589
rect 5532 1537 5584 1589
rect 5394 1444 5446 1496
rect 5394 1378 5446 1430
rect 7601 1244 7653 1296
rect 7669 1244 7721 1296
rect 7737 1244 7789 1296
rect 7804 1244 7856 1296
rect 9777 1287 9829 1339
rect 9777 1223 9829 1275
rect 9777 1159 9829 1211
rect 9842 1159 10086 1339
rect 12509 1286 12561 1338
rect 12584 1286 12636 1338
rect 12659 1286 12711 1338
rect 12509 1218 12561 1270
rect 12584 1218 12636 1270
rect 12659 1218 12711 1270
rect 12509 1150 12561 1202
rect 12584 1150 12636 1202
rect 12659 1150 12711 1202
rect 12509 1082 12561 1134
rect 12584 1082 12636 1134
rect 12659 1082 12711 1134
rect 13021 1187 13073 1239
rect 13021 1123 13073 1175
rect 13281 1187 13333 1239
rect 13281 1123 13333 1175
rect 13722 2570 13774 2622
rect 13786 2570 13838 2622
rect 13850 2570 13902 2622
rect 13915 2570 13967 2622
rect 852 671 904 723
rect 916 671 968 723
rect 11304 569 11356 621
rect 11304 505 11356 557
rect 4562 334 4614 386
rect 4562 270 4614 322
rect 9604 257 9656 309
rect 9668 257 9720 309
rect 13545 2076 13597 2101
rect 13545 2049 13554 2076
rect 13554 2049 13588 2076
rect 13588 2049 13597 2076
rect 13545 2002 13597 2037
rect 13545 1985 13554 2002
rect 13554 1985 13588 2002
rect 13588 1985 13597 2002
rect 13725 1169 13777 1173
rect 13725 1135 13757 1169
rect 13757 1135 13777 1169
rect 13725 1121 13777 1135
rect 13725 1009 13777 1061
rect 13725 896 13777 948
rect 13725 823 13757 835
rect 13757 823 13777 835
rect 13725 783 13777 823
rect 13725 670 13777 722
rect 13725 557 13777 609
rect 13439 308 13473 314
rect 13473 308 13491 314
rect 13439 262 13491 308
rect 13508 270 13560 314
rect 13508 262 13513 270
rect 13513 262 13547 270
rect 13547 262 13560 270
rect 13577 270 13629 314
rect 13577 262 13587 270
rect 13587 262 13621 270
rect 13621 262 13629 270
rect 13646 270 13698 314
rect 13646 262 13661 270
rect 13661 262 13695 270
rect 13695 262 13698 270
rect 13714 270 13766 314
rect 13782 270 13834 314
rect 13850 270 13902 314
rect 13918 270 13970 314
rect 13714 262 13735 270
rect 13735 262 13766 270
rect 13782 262 13809 270
rect 13809 262 13834 270
rect 13850 262 13883 270
rect 13883 262 13902 270
rect 13918 262 13958 270
rect 13958 262 13970 270
rect 13439 190 13491 242
rect 13508 236 13513 242
rect 13513 236 13547 242
rect 13547 236 13560 242
rect 13508 190 13560 236
rect 13577 236 13587 242
rect 13587 236 13621 242
rect 13621 236 13629 242
rect 13577 190 13629 236
rect 13646 236 13661 242
rect 13661 236 13695 242
rect 13695 236 13698 242
rect 13646 190 13698 236
rect 13714 236 13735 242
rect 13735 236 13766 242
rect 13782 236 13809 242
rect 13809 236 13834 242
rect 13850 236 13883 242
rect 13883 236 13902 242
rect 13918 236 13958 242
rect 13958 236 13970 242
rect 13714 190 13766 236
rect 13782 190 13834 236
rect 13850 190 13902 236
rect 13918 190 13970 236
rect 13439 118 13491 170
rect 13508 118 13560 170
rect 13577 118 13629 170
rect 13646 118 13698 170
rect 13714 118 13766 170
rect 13782 118 13834 170
rect 13850 118 13902 170
rect 13918 118 13970 170
rect 7602 -43 7654 9
rect 7703 -43 7755 9
rect 7803 -43 7855 9
rect 7602 -107 7654 -55
rect 7703 -107 7755 -55
rect 7803 -107 7855 -55
rect 8717 -2433 8769 -2381
rect 8781 -2433 8833 -2381
rect 14822 -10078 14874 -10026
rect 14822 -10142 14874 -10090
<< metal2 >>
rect 7993 9819 8231 9829
rect 7993 9767 7995 9819
rect 8047 9767 8105 9819
rect 8157 9767 8231 9819
rect 7993 9728 8231 9767
rect 7993 9676 7995 9728
rect 8047 9676 8105 9728
rect 8157 9676 8231 9728
rect 7993 9637 8231 9676
rect 7993 9585 7995 9637
rect 8047 9585 8105 9637
rect 8157 9585 8231 9637
rect 7993 9546 8231 9585
rect 7993 9494 7995 9546
rect 8047 9494 8105 9546
rect 8157 9494 8231 9546
rect 7993 9455 8231 9494
rect 7993 9403 7995 9455
rect 8047 9403 8105 9455
rect 8157 9403 8231 9455
tri 7818 8907 7993 9082 se
rect 7993 8982 8231 9403
rect 7993 8907 8156 8982
tri 8156 8907 8231 8982 nw
rect 9212 9819 9450 9825
rect 9212 9767 9213 9819
rect 9265 9767 9305 9819
rect 9357 9767 9397 9819
rect 9449 9767 9450 9819
rect 9212 9728 9450 9767
rect 9212 9676 9213 9728
rect 9265 9676 9305 9728
rect 9357 9676 9397 9728
rect 9449 9676 9450 9728
rect 9212 9637 9450 9676
rect 9212 9585 9213 9637
rect 9265 9585 9305 9637
rect 9357 9585 9397 9637
rect 9449 9585 9450 9637
rect 9212 9546 9450 9585
rect 9212 9494 9213 9546
rect 9265 9494 9305 9546
rect 9357 9494 9397 9546
rect 9449 9494 9450 9546
rect 9212 9455 9450 9494
rect 9212 9403 9213 9455
rect 9265 9403 9305 9455
rect 9357 9403 9397 9455
rect 9449 9403 9450 9455
tri 4107 8878 4136 8907 se
rect 4136 8878 8052 8907
rect 1129 8869 1794 8878
rect 1185 8813 1794 8869
rect 1129 8803 1794 8813
tri 1794 8803 1869 8878 sw
tri 4032 8803 4107 8878 se
rect 4107 8803 8052 8878
tri 8052 8803 8156 8907 nw
rect 1129 8789 1869 8803
rect 1185 8733 1869 8789
rect 1129 8724 1869 8733
tri 1869 8724 1948 8803 sw
tri 3953 8724 4032 8803 se
rect 4032 8724 7918 8803
tri 1730 8628 1826 8724 ne
rect 1826 8628 1948 8724
tri 1948 8628 2044 8724 sw
tri 3857 8628 3953 8724 se
rect 3953 8669 7918 8724
tri 7918 8669 8052 8803 nw
tri 9078 8669 9212 8803 se
rect 9212 8703 9450 9403
rect 9212 8669 9375 8703
rect 3953 8628 4195 8669
tri 4195 8628 4236 8669 nw
tri 9037 8628 9078 8669 se
rect 9078 8628 9375 8669
tri 9375 8628 9450 8703 nw
tri 1826 8615 1839 8628 ne
rect 1839 8615 2044 8628
rect 984 8595 1602 8615
rect 984 8589 1224 8595
rect 984 8537 1158 8589
rect 1210 8543 1224 8589
rect 1276 8543 1288 8595
rect 1340 8593 1352 8595
rect 1404 8593 1416 8595
rect 1468 8593 1480 8595
rect 1532 8593 1544 8595
rect 1596 8593 1602 8595
rect 1351 8543 1352 8593
rect 1532 8543 1541 8593
rect 1210 8537 1295 8543
rect 1351 8537 1377 8543
rect 1433 8537 1459 8543
rect 1515 8537 1541 8543
rect 1597 8537 1602 8593
tri 1839 8569 1885 8615 ne
rect 1885 8569 2044 8615
tri 2044 8569 2103 8628 sw
tri 3798 8569 3857 8628 se
rect 3857 8578 4145 8628
tri 4145 8578 4195 8628 nw
tri 4236 8578 4286 8628 se
rect 4286 8578 9137 8628
rect 3857 8569 4136 8578
tri 4136 8569 4145 8578 nw
tri 4227 8569 4236 8578 se
rect 4236 8569 9137 8578
rect 984 8525 1602 8537
rect 984 8473 1158 8525
rect 1210 8509 1602 8525
rect 1210 8473 1295 8509
rect 984 8461 1295 8473
rect 984 8409 1158 8461
rect 1210 8453 1295 8461
rect 1351 8453 1377 8509
rect 1433 8453 1459 8509
rect 1515 8453 1541 8509
rect 1597 8453 1602 8509
tri 1885 8507 1947 8569 ne
rect 1947 8513 2103 8569
tri 2103 8513 2159 8569 sw
tri 3742 8513 3798 8569 se
rect 3798 8513 4074 8569
rect 1947 8507 2159 8513
tri 2159 8507 2165 8513 sw
tri 3736 8507 3742 8513 se
rect 3742 8507 4074 8513
tri 4074 8507 4136 8569 nw
tri 4165 8507 4227 8569 se
rect 4227 8507 9137 8569
tri 1947 8506 1948 8507 ne
rect 1948 8506 4045 8507
tri 1948 8483 1971 8506 ne
rect 1971 8483 4045 8506
rect 1210 8425 1602 8453
tri 1971 8431 2023 8483 ne
rect 2023 8431 2049 8483
rect 2101 8431 2113 8483
rect 2165 8431 2177 8483
rect 2229 8431 2241 8483
rect 2293 8431 2305 8483
rect 2357 8431 2369 8483
rect 2421 8431 2433 8483
rect 2485 8431 2497 8483
rect 2549 8431 2561 8483
rect 2613 8431 2625 8483
rect 2677 8431 2689 8483
rect 2741 8431 2753 8483
rect 2805 8478 4045 8483
tri 4045 8478 4074 8507 nw
tri 4136 8478 4165 8507 se
rect 4165 8478 9137 8507
rect 2805 8431 3954 8478
rect 1210 8409 1295 8425
rect 984 8397 1295 8409
rect 984 8345 1158 8397
rect 1210 8369 1295 8397
rect 1351 8369 1377 8425
rect 1433 8369 1459 8425
rect 1515 8369 1541 8425
rect 1597 8369 1602 8425
tri 2023 8412 2042 8431 ne
rect 1210 8345 1602 8369
rect 984 8341 1602 8345
rect 984 8333 1295 8341
rect 984 8281 1158 8333
rect 1210 8324 1295 8333
rect 1351 8324 1377 8341
rect 1433 8324 1459 8341
rect 1515 8324 1541 8341
rect 1210 8281 1288 8324
rect 1351 8285 1352 8324
rect 1532 8285 1541 8324
rect 1597 8285 1602 8341
rect 984 8272 1288 8281
rect 1340 8272 1352 8285
rect 1404 8272 1416 8285
rect 1468 8272 1480 8285
rect 1532 8272 1544 8285
rect 1596 8272 1602 8285
rect 984 8269 1602 8272
rect 984 8217 1158 8269
rect 1210 8257 1602 8269
rect 1210 8217 1295 8257
rect 984 8205 1295 8217
rect 984 8153 1158 8205
rect 1210 8201 1295 8205
rect 1351 8201 1377 8257
rect 1433 8201 1459 8257
rect 1515 8201 1541 8257
rect 1597 8201 1602 8257
rect 1210 8173 1602 8201
rect 1210 8153 1295 8173
rect 984 8141 1295 8153
rect 984 8089 1158 8141
rect 1210 8117 1295 8141
rect 1351 8117 1377 8173
rect 1433 8117 1459 8173
rect 1515 8117 1541 8173
rect 1597 8117 1602 8173
rect 2042 8387 3954 8431
tri 3954 8387 4045 8478 nw
tri 4045 8387 4136 8478 se
rect 4136 8390 9137 8478
tri 9137 8390 9375 8628 nw
tri 11756 8513 11807 8564 se
rect 11807 8513 14064 8564
tri 14064 8513 14115 8564 sw
tri 11733 8490 11756 8513 se
rect 11756 8512 14115 8513
rect 11756 8490 11807 8512
tri 11807 8490 11829 8512 nw
tri 14006 8490 14028 8512 ne
rect 14028 8490 14115 8512
tri 11659 8416 11733 8490 se
tri 11733 8416 11807 8490 nw
tri 14028 8455 14063 8490 ne
tri 11633 8390 11659 8416 se
rect 11659 8390 11690 8416
rect 4136 8387 4363 8390
rect 2042 8381 3948 8387
tri 3948 8381 3954 8387 nw
tri 4039 8381 4045 8387 se
rect 4045 8381 4363 8387
rect 2042 8367 3934 8381
tri 3934 8367 3948 8381 nw
tri 4025 8367 4039 8381 se
rect 4039 8367 4363 8381
tri 4363 8367 4386 8390 nw
tri 11616 8373 11633 8390 se
rect 11633 8373 11690 8390
tri 11690 8373 11733 8416 nw
tri 11610 8367 11616 8373 se
rect 11616 8367 11684 8373
tri 11684 8367 11690 8373 nw
rect 2042 8315 3882 8367
tri 3882 8315 3934 8367 nw
tri 3973 8315 4025 8367 se
rect 4025 8315 4311 8367
tri 4311 8315 4363 8367 nw
tri 11585 8342 11610 8367 se
rect 11610 8342 11659 8367
tri 11659 8342 11684 8367 nw
tri 11575 8332 11585 8342 se
rect 11585 8332 11649 8342
tri 11649 8332 11659 8342 nw
rect 11453 8315 11632 8332
tri 11632 8315 11649 8332 nw
rect 2042 8300 3867 8315
tri 3867 8300 3882 8315 nw
tri 3958 8300 3973 8315 se
rect 3973 8300 4296 8315
tri 4296 8300 4311 8315 nw
rect 11453 8300 11617 8315
tri 11617 8300 11632 8315 nw
rect 2042 8290 3857 8300
tri 3857 8290 3867 8300 nw
tri 3948 8290 3958 8300 se
rect 3958 8290 4286 8300
tri 4286 8290 4296 8300 nw
rect 11453 8290 11607 8300
tri 11607 8290 11617 8300 nw
rect 2042 8269 3836 8290
tri 3836 8269 3857 8290 nw
tri 3927 8269 3948 8290 se
rect 3948 8269 4265 8290
tri 4265 8269 4286 8290 nw
rect 11453 8269 11586 8290
tri 11586 8269 11607 8290 nw
rect 2042 8263 2949 8269
tri 2949 8263 2955 8269 nw
tri 3921 8263 3927 8269 se
rect 3927 8263 4259 8269
tri 4259 8263 4265 8269 nw
tri 4301 8263 4307 8269 se
rect 4307 8263 4373 8269
rect 2042 8211 2897 8263
tri 2897 8211 2949 8263 nw
tri 3869 8211 3921 8263 se
rect 3921 8227 4223 8263
tri 4223 8227 4259 8263 nw
tri 4265 8227 4301 8263 se
rect 4301 8227 4321 8263
rect 3921 8225 4221 8227
tri 4221 8225 4223 8227 nw
tri 4263 8225 4265 8227 se
rect 4265 8225 4321 8227
rect 3921 8211 4207 8225
tri 4207 8211 4221 8225 nw
tri 4249 8211 4263 8225 se
rect 4263 8211 4321 8225
rect 2042 8199 2885 8211
tri 2885 8199 2897 8211 nw
tri 3857 8199 3869 8211 se
rect 3869 8199 4195 8211
tri 4195 8199 4207 8211 nw
tri 4237 8199 4249 8211 se
rect 4249 8199 4373 8211
rect 2042 8169 2855 8199
tri 2855 8169 2885 8199 nw
tri 3827 8169 3857 8199 se
rect 3857 8183 4179 8199
tri 4179 8183 4195 8199 nw
tri 4221 8183 4237 8199 se
rect 4237 8183 4321 8199
rect 3857 8169 4143 8183
rect 2042 8117 2049 8169
rect 2101 8117 2113 8169
rect 2165 8117 2177 8169
rect 2229 8117 2241 8169
rect 2293 8117 2305 8169
rect 2357 8117 2369 8169
rect 2421 8117 2433 8169
rect 2485 8117 2497 8169
rect 2549 8117 2561 8169
rect 2613 8117 2625 8169
rect 2677 8117 2689 8169
rect 2741 8117 2753 8169
rect 2805 8147 2833 8169
tri 2833 8147 2855 8169 nw
tri 3805 8147 3827 8169 se
rect 3827 8147 4143 8169
tri 4143 8147 4179 8183 nw
tri 4185 8147 4221 8183 se
rect 4221 8147 4321 8183
rect 11453 8248 11565 8269
tri 11565 8248 11586 8269 nw
rect 11453 8233 11550 8248
tri 11550 8233 11565 8248 nw
rect 11453 8192 11509 8233
tri 11509 8192 11550 8233 nw
rect 2805 8134 2820 8147
tri 2820 8134 2833 8147 nw
tri 3792 8134 3805 8147 se
rect 3805 8141 4137 8147
tri 4137 8141 4143 8147 nw
tri 4179 8141 4185 8147 se
rect 4185 8141 4373 8147
rect 4814 8186 5032 8192
rect 4814 8183 4955 8186
rect 5007 8183 5032 8186
rect 3805 8134 4130 8141
tri 4130 8134 4137 8141 nw
tri 4172 8134 4179 8141 se
rect 4179 8134 4246 8141
tri 4246 8134 4253 8141 nw
rect 2805 8117 2811 8134
tri 2811 8125 2820 8134 nw
tri 3783 8125 3792 8134 se
rect 3792 8125 4110 8134
tri 3775 8117 3783 8125 se
rect 3783 8117 4110 8125
rect 1210 8089 1602 8117
tri 3772 8114 3775 8117 se
rect 3775 8114 4110 8117
tri 4110 8114 4130 8134 nw
tri 4152 8114 4172 8134 se
rect 4172 8114 4226 8134
tri 4226 8114 4246 8134 nw
rect 4870 8127 4894 8183
rect 4950 8134 4955 8183
rect 4950 8127 4974 8134
rect 5030 8127 5032 8183
rect 11453 8181 11498 8192
tri 11498 8181 11509 8192 nw
rect 11453 8166 11483 8181
tri 11483 8166 11498 8181 nw
tri 11453 8136 11483 8166 nw
tri 3768 8110 3772 8114 se
rect 3772 8110 4106 8114
tri 4106 8110 4110 8114 nw
tri 4148 8110 4152 8114 se
rect 4152 8110 4222 8114
tri 4222 8110 4226 8114 nw
rect 4814 8110 5032 8127
rect 984 8077 1295 8089
rect -731 8033 -275 8036
rect -731 7981 -724 8033
rect -672 7981 -659 8033
rect -607 7981 -594 8033
rect -542 7981 -529 8033
rect -477 7981 -464 8033
rect -412 7981 -399 8033
rect -347 7981 -334 8033
rect -282 7981 -275 8033
rect -731 7961 -275 7981
rect -731 7909 -724 7961
rect -672 7909 -659 7961
rect -607 7909 -594 7961
rect -542 7909 -529 7961
rect -477 7909 -464 7961
rect -412 7909 -399 7961
rect -347 7909 -334 7961
rect -282 7909 -275 7961
rect -731 7889 -275 7909
rect -731 7837 -724 7889
rect -672 7837 -659 7889
rect -607 7837 -594 7889
rect -542 7837 -529 7889
rect -477 7837 -464 7889
rect -412 7837 -399 7889
rect -347 7837 -334 7889
rect -282 7837 -275 7889
rect -731 7817 -275 7837
rect -731 7765 -724 7817
rect -672 7765 -659 7817
rect -607 7765 -594 7817
rect -542 7765 -529 7817
rect -477 7765 -464 7817
rect -412 7765 -399 7817
rect -347 7765 -334 7817
rect -282 7765 -275 7817
rect -731 7745 -275 7765
rect -731 7693 -724 7745
rect -672 7693 -659 7745
rect -607 7693 -594 7745
rect -542 7693 -529 7745
rect -477 7693 -464 7745
rect -412 7693 -399 7745
rect -347 7693 -334 7745
rect -282 7693 -275 7745
rect -731 7335 -275 7693
rect -731 7283 -724 7335
rect -672 7283 -658 7335
rect -606 7283 -593 7335
rect -541 7283 -528 7335
rect -476 7283 -463 7335
rect -411 7283 -398 7335
rect -346 7283 -333 7335
rect -281 7283 -275 7335
rect -731 7255 -275 7283
rect 984 8025 1158 8077
rect 1210 8033 1295 8077
rect 1351 8033 1377 8089
rect 1433 8033 1459 8089
rect 1515 8033 1541 8089
rect 1597 8033 1602 8089
tri 3716 8058 3768 8110 se
rect 3768 8109 4105 8110
tri 4105 8109 4106 8110 nw
tri 4147 8109 4148 8110 se
rect 4148 8109 4179 8110
rect 3768 8067 4063 8109
tri 4063 8067 4105 8109 nw
tri 4105 8067 4147 8109 se
rect 4147 8067 4179 8109
tri 4179 8067 4222 8110 nw
rect 3768 8058 4054 8067
tri 4054 8058 4063 8067 nw
tri 4096 8058 4105 8067 se
rect 4105 8058 4170 8067
tri 4170 8058 4179 8067 nw
rect 4814 8060 4955 8110
rect 5007 8060 5032 8110
tri 3705 8047 3716 8058 se
rect 3716 8047 4043 8058
tri 4043 8047 4054 8058 nw
tri 4085 8047 4096 8058 se
rect 4096 8047 4159 8058
tri 4159 8047 4170 8058 nw
tri 3692 8034 3705 8047 se
rect 3705 8035 4031 8047
tri 4031 8035 4043 8047 nw
tri 4073 8035 4085 8047 se
rect 4085 8035 4146 8047
rect 3705 8034 4030 8035
tri 4030 8034 4031 8035 nw
tri 4072 8034 4073 8035 se
rect 4073 8034 4146 8035
tri 4146 8034 4159 8047 nw
tri 3691 8033 3692 8034 se
rect 3692 8033 3989 8034
rect 1210 8025 1602 8033
rect 984 8016 1602 8025
rect 984 8013 1288 8016
rect 984 7961 1158 8013
rect 1210 7964 1288 8013
rect 1340 8005 1352 8016
rect 1404 8005 1416 8016
rect 1468 8005 1480 8016
rect 1532 8005 1544 8016
rect 1596 8005 1602 8016
rect 1351 7964 1352 8005
rect 1532 7964 1541 8005
rect 1210 7961 1295 7964
rect 984 7949 1295 7961
rect 1351 7949 1377 7964
rect 1433 7949 1459 7964
rect 1515 7949 1541 7964
rect 1597 7949 1602 8005
tri 3640 7982 3691 8033 se
rect 3691 7993 3989 8033
tri 3989 7993 4030 8034 nw
tri 4031 7993 4072 8034 se
rect 4072 7993 4105 8034
tri 4105 7993 4146 8034 nw
rect 4870 8004 4894 8060
rect 4950 8058 4955 8060
rect 4950 8034 4974 8058
rect 4950 8004 4955 8034
rect 5030 8004 5032 8060
rect 3691 7982 3978 7993
tri 3978 7982 3989 7993 nw
tri 4020 7982 4031 7993 se
rect 4031 7982 4094 7993
tri 4094 7982 4105 7993 nw
rect 4814 7982 4955 8004
rect 5007 7982 5032 8004
tri 3638 7980 3640 7982 se
rect 3640 7980 3976 7982
tri 3976 7980 3978 7982 nw
tri 4018 7980 4020 7982 se
rect 4020 7980 4092 7982
tri 4092 7980 4094 7982 nw
tri 3623 7965 3638 7980 se
rect 3638 7965 3961 7980
tri 3961 7965 3976 7980 nw
tri 4003 7965 4018 7980 se
rect 4018 7965 4077 7980
tri 4077 7965 4092 7980 nw
tri 3616 7958 3623 7965 se
rect 3623 7961 3957 7965
tri 3957 7961 3961 7965 nw
tri 3999 7961 4003 7965 se
rect 4003 7961 4070 7965
rect 3623 7958 3954 7961
tri 3954 7958 3957 7961 nw
tri 3996 7958 3999 7961 se
rect 3999 7958 4070 7961
tri 4070 7958 4077 7965 nw
rect 4814 7958 5032 7982
tri 3610 7952 3616 7958 se
rect 3616 7952 3948 7958
tri 3948 7952 3954 7958 nw
tri 3990 7952 3996 7958 se
rect 3996 7952 4031 7958
rect 984 7897 1158 7949
rect 1210 7921 1602 7949
rect 1210 7897 1295 7921
rect 984 7885 1295 7897
rect 984 7833 1158 7885
rect 1210 7865 1295 7885
rect 1351 7865 1377 7921
rect 1433 7865 1459 7921
rect 1515 7865 1541 7921
rect 1597 7865 1602 7921
tri 3564 7906 3610 7952 se
rect 3610 7919 3915 7952
tri 3915 7919 3948 7952 nw
tri 3957 7919 3990 7952 se
rect 3990 7919 4031 7952
tri 4031 7919 4070 7958 nw
rect 4814 7937 4955 7958
rect 5007 7937 5032 7958
rect 3610 7906 3902 7919
tri 3902 7906 3915 7919 nw
tri 3944 7906 3957 7919 se
rect 3957 7906 4018 7919
tri 4018 7906 4031 7919 nw
tri 3555 7897 3564 7906 se
rect 3564 7897 3893 7906
tri 3893 7897 3902 7906 nw
tri 3935 7897 3944 7906 se
rect 3944 7897 4009 7906
tri 4009 7897 4018 7906 nw
tri 3540 7882 3555 7897 se
rect 3555 7887 3883 7897
tri 3883 7887 3893 7897 nw
tri 3925 7887 3935 7897 se
rect 3935 7887 3994 7897
rect 3555 7882 3878 7887
tri 3878 7882 3883 7887 nw
tri 3920 7882 3925 7887 se
rect 3925 7882 3994 7887
tri 3994 7882 4009 7897 nw
tri 3525 7867 3540 7882 se
rect 3540 7867 3863 7882
tri 3863 7867 3878 7882 nw
tri 3905 7867 3920 7882 se
rect 3920 7867 3957 7882
rect 1210 7837 1602 7865
rect 1210 7833 1295 7837
rect 984 7821 1295 7833
rect 984 7769 1158 7821
rect 1210 7781 1295 7821
rect 1351 7781 1377 7837
rect 1433 7781 1459 7837
rect 1515 7781 1541 7837
rect 1597 7781 1602 7837
rect 1210 7769 1602 7781
rect 984 7757 1602 7769
rect 984 7705 1158 7757
rect 1210 7753 1602 7757
rect 1210 7705 1295 7753
rect 984 7701 1295 7705
rect 1351 7701 1377 7753
rect 1433 7701 1459 7753
rect 1515 7701 1541 7753
rect 984 7693 1288 7701
rect 1351 7697 1352 7701
rect 1532 7697 1541 7701
rect 1597 7697 1602 7753
rect 984 7641 1158 7693
rect 1210 7649 1288 7693
rect 1340 7669 1352 7697
rect 1404 7669 1416 7697
rect 1468 7669 1480 7697
rect 1532 7669 1544 7697
rect 1596 7669 1602 7697
rect 2042 7857 3841 7867
rect 2042 7805 2069 7857
rect 2121 7805 2133 7857
rect 2185 7805 2197 7857
rect 2249 7805 2261 7857
rect 2313 7805 2325 7857
rect 2377 7805 2389 7857
rect 2441 7805 2453 7857
rect 2505 7805 2517 7857
rect 2569 7805 2581 7857
rect 2633 7805 2645 7857
rect 2697 7805 2709 7857
rect 2761 7805 2773 7857
rect 2825 7805 2837 7857
rect 2889 7845 3841 7857
tri 3841 7845 3863 7867 nw
tri 3883 7845 3905 7867 se
rect 3905 7845 3957 7867
tri 3957 7845 3994 7882 nw
rect 4870 7881 4894 7937
rect 4950 7906 4955 7937
rect 4950 7882 4974 7906
rect 4950 7881 4955 7882
rect 5030 7881 5032 7937
tri 6972 7897 6985 7910 se
rect 2889 7837 3833 7845
tri 3833 7837 3841 7845 nw
tri 3875 7837 3883 7845 se
rect 3883 7837 3942 7845
rect 2889 7830 3826 7837
tri 3826 7830 3833 7837 nw
tri 3868 7830 3875 7837 se
rect 3875 7830 3942 7837
tri 3942 7830 3957 7845 nw
rect 4814 7830 4955 7881
rect 5007 7830 5032 7881
tri 6920 7845 6972 7897 se
rect 6972 7845 6985 7897
tri 6913 7838 6920 7845 se
rect 6920 7838 6985 7845
rect 2889 7829 3825 7830
tri 3825 7829 3826 7830 nw
tri 3867 7829 3868 7830 se
rect 3868 7829 3941 7830
tri 3941 7829 3942 7830 nw
rect 2889 7813 3809 7829
tri 3809 7813 3825 7829 nw
tri 3851 7813 3867 7829 se
rect 3867 7813 3918 7829
rect 2889 7806 3802 7813
tri 3802 7806 3809 7813 nw
tri 3844 7806 3851 7813 se
rect 3851 7806 3918 7813
tri 3918 7806 3941 7829 nw
rect 4814 7813 5032 7830
rect 2889 7805 3767 7806
rect 2042 7771 3767 7805
tri 3767 7771 3802 7806 nw
tri 3809 7771 3844 7806 se
rect 3844 7771 3883 7806
tri 3883 7771 3918 7806 nw
rect 2042 7754 3750 7771
tri 3750 7754 3767 7771 nw
tri 3792 7754 3809 7771 se
rect 3809 7754 3866 7771
tri 3866 7754 3883 7771 nw
rect 4870 7757 4894 7813
rect 4950 7806 4974 7813
rect 4950 7757 4955 7806
rect 5030 7757 5032 7813
rect 4814 7754 4955 7757
rect 5007 7754 5032 7757
rect 2042 7739 3735 7754
tri 3735 7739 3750 7754 nw
tri 3786 7748 3792 7754 se
rect 3792 7748 3860 7754
tri 3860 7748 3866 7754 nw
rect 4814 7748 5032 7754
rect 6470 7837 9707 7838
rect 6470 7781 6479 7837
rect 6535 7781 6561 7837
rect 6617 7781 6643 7837
rect 6699 7781 6725 7837
rect 6781 7781 6807 7837
rect 6863 7781 6888 7837
rect 6944 7781 6969 7837
rect 7025 7781 7050 7837
rect 7106 7781 7131 7837
rect 7187 7781 7212 7837
rect 7268 7781 7293 7837
rect 7349 7781 7374 7837
rect 7430 7781 7455 7837
rect 7511 7781 7536 7837
rect 7592 7781 7617 7837
rect 7673 7781 7698 7837
rect 7754 7781 7779 7837
rect 7835 7781 7860 7837
rect 7916 7781 7941 7837
rect 7997 7781 8022 7837
rect 8078 7781 8103 7837
rect 8159 7781 8184 7837
rect 8240 7781 8265 7837
rect 8321 7781 8346 7837
rect 8402 7781 8427 7837
rect 8483 7781 8508 7837
rect 8564 7781 8589 7837
rect 8645 7781 8670 7837
rect 8726 7781 8751 7837
rect 8807 7781 8832 7837
rect 8888 7781 8913 7837
rect 8969 7781 8994 7837
rect 9050 7781 9075 7837
rect 9131 7781 9156 7837
rect 9212 7781 9237 7837
rect 9293 7781 9318 7837
rect 9374 7781 9399 7837
rect 9455 7781 9480 7837
rect 9536 7781 9561 7837
rect 9617 7781 9642 7837
rect 9698 7781 9707 7837
tri 3777 7739 3786 7748 se
rect 3786 7739 3809 7748
rect 2042 7697 3693 7739
tri 3693 7697 3735 7739 nw
tri 3735 7697 3777 7739 se
rect 3777 7697 3809 7739
tri 3809 7697 3860 7748 nw
rect 6470 7743 9707 7781
rect 2042 7693 3689 7697
tri 3689 7693 3693 7697 nw
tri 3731 7693 3735 7697 se
rect 3735 7693 3774 7697
rect 1351 7649 1352 7669
rect 1532 7649 1541 7669
rect 1210 7641 1295 7649
rect 984 7629 1295 7641
rect 984 7577 1158 7629
rect 1210 7613 1295 7629
rect 1351 7613 1377 7649
rect 1433 7613 1459 7649
rect 1515 7613 1541 7649
rect 1597 7613 1602 7669
rect 1210 7585 1602 7613
rect 1210 7577 1295 7585
rect 984 7565 1295 7577
rect 984 7513 1158 7565
rect 1210 7529 1295 7565
rect 1351 7529 1377 7585
rect 1433 7529 1459 7585
rect 1515 7529 1541 7585
rect 1597 7529 1602 7585
tri 1894 7545 2042 7693 se
rect 2042 7665 3661 7693
tri 3661 7665 3689 7693 nw
tri 3703 7665 3731 7693 se
rect 3731 7665 3774 7693
rect 2042 7623 3619 7665
tri 3619 7623 3661 7665 nw
tri 3700 7662 3703 7665 se
rect 3703 7662 3774 7665
tri 3774 7662 3809 7697 nw
rect 6470 7687 6479 7743
rect 6535 7687 6561 7743
rect 6617 7687 6643 7743
rect 6699 7687 6725 7743
rect 6781 7687 6807 7743
rect 6863 7687 6888 7743
rect 6944 7687 6969 7743
rect 7025 7687 7050 7743
rect 7106 7687 7131 7743
rect 7187 7687 7212 7743
rect 7268 7687 7293 7743
rect 7349 7687 7374 7743
rect 7430 7687 7455 7743
rect 7511 7687 7536 7743
rect 7592 7687 7617 7743
rect 7673 7687 7698 7743
rect 7754 7687 7779 7743
rect 7835 7687 7860 7743
rect 7916 7687 7941 7743
rect 7997 7687 8022 7743
rect 8078 7687 8103 7743
rect 8159 7687 8184 7743
rect 8240 7687 8265 7743
rect 8321 7687 8346 7743
rect 8402 7687 8427 7743
rect 8483 7687 8508 7743
rect 8564 7687 8589 7743
rect 8645 7687 8670 7743
rect 8726 7687 8751 7743
rect 8807 7687 8832 7743
rect 8888 7687 8913 7743
rect 8969 7687 8994 7743
rect 9050 7687 9075 7743
rect 9131 7687 9156 7743
rect 9212 7687 9237 7743
rect 9293 7687 9318 7743
rect 9374 7687 9399 7743
rect 9455 7687 9480 7743
rect 9536 7687 9561 7743
rect 9617 7687 9642 7743
rect 9698 7687 9707 7743
tri 3669 7631 3700 7662 se
rect 3700 7631 3743 7662
tri 3743 7631 3774 7662 nw
tri 4760 7631 4791 7662 se
rect 4791 7631 6136 7662
tri 6136 7631 6167 7662 sw
rect 6470 7649 9707 7687
tri 3661 7623 3669 7631 se
rect 3669 7623 3735 7631
tri 3735 7623 3743 7631 nw
tri 4752 7623 4760 7631 se
rect 4760 7623 6167 7631
rect 2042 7591 3587 7623
tri 3587 7591 3619 7623 nw
tri 3629 7591 3661 7623 se
rect 3661 7591 3682 7623
rect 2042 7570 3566 7591
tri 3566 7570 3587 7591 nw
tri 3608 7570 3629 7591 se
rect 3629 7570 3682 7591
tri 3682 7570 3735 7623 nw
tri 4699 7570 4752 7623 se
rect 4752 7570 6167 7623
tri 6167 7570 6228 7631 sw
rect 6470 7593 6479 7649
rect 6535 7593 6561 7649
rect 6617 7593 6643 7649
rect 6699 7593 6725 7649
rect 6781 7593 6807 7649
rect 6863 7593 6888 7649
rect 6944 7593 6969 7649
rect 7025 7593 7050 7649
rect 7106 7593 7131 7649
rect 7187 7593 7212 7649
rect 7268 7593 7293 7649
rect 7349 7593 7374 7649
rect 7430 7593 7455 7649
rect 7511 7593 7536 7649
rect 7592 7593 7617 7649
rect 7673 7593 7698 7649
rect 7754 7593 7779 7649
rect 7835 7593 7860 7649
rect 7916 7593 7941 7649
rect 7997 7593 8022 7649
rect 8078 7593 8103 7649
rect 8159 7593 8184 7649
rect 8240 7593 8265 7649
rect 8321 7593 8346 7649
rect 8402 7593 8427 7649
rect 8483 7593 8508 7649
rect 8564 7593 8589 7649
rect 8645 7593 8670 7649
rect 8726 7593 8751 7649
rect 8807 7593 8832 7649
rect 8888 7593 8913 7649
rect 8969 7593 8994 7649
rect 9050 7593 9075 7649
rect 9131 7593 9156 7649
rect 9212 7593 9237 7649
rect 9293 7593 9318 7649
rect 9374 7593 9399 7649
rect 9455 7593 9480 7649
rect 9536 7593 9561 7649
rect 9617 7593 9642 7649
rect 9698 7593 9707 7649
rect 2042 7549 3545 7570
tri 3545 7549 3566 7570 nw
tri 3587 7549 3608 7570 se
rect 3608 7549 3661 7570
tri 3661 7549 3682 7570 nw
tri 4678 7549 4699 7570 se
rect 4699 7549 6228 7570
rect 2042 7545 3513 7549
rect 1210 7513 1602 7529
rect 984 7501 1602 7513
rect 984 7449 1158 7501
rect 1210 7449 1295 7501
rect 984 7445 1295 7449
rect 1351 7445 1377 7501
rect 1433 7445 1459 7501
rect 1515 7445 1541 7501
rect 1597 7445 1602 7501
tri 1842 7493 1894 7545 se
rect 1894 7493 2069 7545
rect 2121 7493 2133 7545
rect 2185 7493 2197 7545
rect 2249 7493 2261 7545
rect 2313 7493 2325 7545
rect 2377 7493 2389 7545
rect 2441 7493 2453 7545
rect 2505 7493 2517 7545
rect 2569 7493 2581 7545
rect 2633 7493 2645 7545
rect 2697 7493 2709 7545
rect 2761 7493 2773 7545
rect 2825 7493 2837 7545
rect 2889 7517 3513 7545
tri 3513 7517 3545 7549 nw
tri 3555 7517 3587 7549 se
rect 3587 7517 3605 7549
rect 2889 7493 3489 7517
tri 3489 7493 3513 7517 nw
tri 3531 7493 3555 7517 se
rect 3555 7493 3605 7517
tri 3605 7493 3661 7549 nw
tri 4622 7493 4678 7549 se
rect 4678 7493 6228 7549
tri 6228 7493 6305 7570 sw
rect 6470 7555 9707 7593
rect 6470 7499 6479 7555
rect 6535 7499 6561 7555
rect 6617 7499 6643 7555
rect 6699 7499 6725 7555
rect 6781 7499 6807 7555
rect 6863 7499 6888 7555
rect 6944 7499 6969 7555
rect 7025 7499 7050 7555
rect 7106 7499 7131 7555
rect 7187 7499 7212 7555
rect 7268 7499 7293 7555
rect 7349 7499 7374 7555
rect 7430 7499 7455 7555
rect 7511 7499 7536 7555
rect 7592 7499 7617 7555
rect 7673 7499 7698 7555
rect 7754 7499 7779 7555
rect 7835 7499 7860 7555
rect 7916 7499 7941 7555
rect 7997 7499 8022 7555
rect 8078 7499 8103 7555
rect 8159 7499 8184 7555
rect 8240 7499 8265 7555
rect 8321 7499 8346 7555
rect 8402 7499 8427 7555
rect 8483 7499 8508 7555
rect 8564 7499 8589 7555
rect 8645 7499 8670 7555
rect 8726 7499 8751 7555
rect 8807 7499 8832 7555
rect 8888 7499 8913 7555
rect 8969 7499 8994 7555
rect 9050 7499 9075 7555
rect 9131 7499 9156 7555
rect 9212 7499 9237 7555
rect 9293 7499 9318 7555
rect 9374 7499 9399 7555
rect 9455 7499 9480 7555
rect 9536 7499 9561 7555
rect 9617 7499 9642 7555
rect 9698 7499 9707 7555
rect 6470 7498 9707 7499
tri 9707 7498 9779 7570 nw
rect 984 7437 1602 7445
rect 984 7385 1158 7437
rect 1210 7417 1602 7437
rect 1210 7389 1295 7417
rect 1351 7389 1377 7417
rect 1433 7389 1459 7417
rect 1515 7389 1541 7417
rect 1210 7385 1288 7389
rect 984 7373 1288 7385
rect 984 7321 1158 7373
rect 1210 7337 1288 7373
rect 1351 7361 1352 7389
rect 1532 7361 1541 7389
rect 1597 7361 1602 7417
rect 1340 7337 1352 7361
rect 1404 7337 1416 7361
rect 1468 7337 1480 7361
rect 1532 7337 1544 7361
rect 1596 7337 1602 7361
rect 1210 7333 1602 7337
rect 1210 7321 1295 7333
rect 1351 7321 1377 7333
rect 1433 7321 1459 7333
rect 1515 7321 1541 7333
rect 984 7269 1284 7321
rect 1531 7277 1541 7321
rect 1597 7277 1602 7333
rect 1336 7269 1349 7277
rect 1401 7269 1414 7277
rect 1466 7269 1479 7277
rect 1531 7269 1544 7277
rect 1596 7269 1602 7277
rect 984 7268 1602 7269
tri 1754 7405 1842 7493 se
rect 1842 7475 2042 7493
tri 2042 7475 2060 7493 nw
tri 3513 7475 3531 7493 se
rect 3531 7475 3587 7493
tri 3587 7475 3605 7493 nw
tri 4604 7475 4622 7493 se
rect 4622 7475 6305 7493
rect 1842 7441 2008 7475
tri 2008 7441 2042 7475 nw
tri 3479 7441 3513 7475 se
rect 3513 7441 3553 7475
tri 3553 7441 3587 7475 nw
tri 4570 7441 4604 7475 se
rect 4604 7470 6305 7475
rect 4604 7441 4829 7470
rect 1842 7430 1997 7441
tri 1997 7430 2008 7441 nw
tri 2250 7430 2261 7441 se
rect 2261 7430 3542 7441
tri 3542 7430 3553 7441 nw
tri 4559 7430 4570 7441 se
rect 4570 7430 4829 7441
tri 4829 7430 4869 7470 nw
tri 6058 7430 6098 7470 ne
rect 6098 7459 6305 7470
tri 6305 7459 6339 7493 sw
rect 6098 7430 6339 7459
tri 6339 7430 6368 7459 sw
rect 1842 7405 1959 7430
rect 1754 7392 1959 7405
tri 1959 7392 1997 7430 nw
tri 2212 7392 2250 7430 se
rect 2250 7392 3504 7430
tri 3504 7392 3542 7430 nw
tri 4521 7392 4559 7430 se
rect 4559 7392 4791 7430
tri 4791 7392 4829 7430 nw
tri 5126 7392 5164 7430 se
rect 5164 7421 5408 7430
rect 1754 7374 1941 7392
tri 1941 7374 1959 7392 nw
tri 2194 7374 2212 7392 se
rect 2212 7389 3501 7392
tri 3501 7389 3504 7392 nw
tri 4518 7389 4521 7392 se
rect 4521 7389 4773 7392
rect 2212 7374 2268 7389
tri 2268 7374 2283 7389 nw
tri 4503 7374 4518 7389 se
rect 4518 7374 4773 7389
tri 4773 7374 4791 7392 nw
tri 5108 7374 5126 7392 se
rect 5126 7374 5164 7392
rect 1754 7367 1934 7374
tri 1934 7367 1941 7374 nw
tri 2187 7367 2194 7374 se
rect 2194 7367 2261 7374
tri 2261 7367 2268 7374 nw
tri 4496 7367 4503 7374 se
rect 4503 7367 4735 7374
rect -731 7203 -724 7255
rect -672 7203 -658 7255
rect -606 7203 -593 7255
rect -541 7203 -528 7255
rect -476 7203 -463 7255
rect -411 7203 -398 7255
rect -346 7203 -333 7255
rect -281 7203 -275 7255
rect -731 7175 -275 7203
rect -731 7123 -724 7175
rect -672 7123 -658 7175
rect -606 7123 -593 7175
rect -541 7123 -528 7175
rect -476 7123 -463 7175
rect -411 7123 -398 7175
rect -346 7123 -333 7175
rect -281 7123 -275 7175
rect -731 7122 -275 7123
tri 1733 7122 1754 7143 se
rect 1754 7122 1908 7367
tri 1908 7341 1934 7367 nw
tri 2161 7341 2187 7367 se
rect 2187 7341 2230 7367
tri 2156 7336 2161 7341 se
rect 2161 7336 2230 7341
tri 2230 7336 2261 7367 nw
tri 4465 7336 4496 7367 se
rect 4496 7336 4735 7367
tri 4735 7336 4773 7374 nw
tri 5070 7336 5108 7374 se
rect 5108 7365 5164 7374
rect 5220 7365 5258 7421
rect 5314 7365 5352 7421
tri 6098 7374 6154 7430 ne
rect 6154 7374 6368 7430
tri 6368 7374 6424 7430 sw
rect 9394 7413 10141 7459
rect 5108 7336 5408 7365
tri 6154 7361 6167 7374 ne
rect 6167 7361 6424 7374
tri 6424 7361 6437 7374 sw
tri 2142 7322 2156 7336 se
rect 2156 7322 2216 7336
tri 2216 7322 2230 7336 nw
tri 4451 7322 4465 7336 se
rect 4465 7322 4721 7336
tri 4721 7322 4735 7336 nw
tri 5056 7322 5070 7336 se
rect 5070 7322 5408 7336
tri 6167 7322 6206 7361 ne
rect 6206 7322 8856 7361
tri 2141 7321 2142 7322 se
rect 2142 7321 2215 7322
tri 2215 7321 2216 7322 nw
tri 4450 7321 4451 7322 se
rect 4451 7321 4720 7322
tri 4720 7321 4721 7322 nw
tri 5055 7321 5056 7322 se
rect 5056 7321 5408 7322
tri 2138 7318 2141 7321 se
rect 2141 7318 2212 7321
tri 2212 7318 2215 7321 nw
tri 4447 7318 4450 7321 se
rect 4450 7318 4717 7321
tri 4717 7318 4720 7321 nw
tri 5052 7318 5055 7321 se
rect 5055 7319 5408 7321
rect 5055 7318 5164 7319
tri 2122 7302 2138 7318 se
rect 2138 7302 2196 7318
tri 2196 7302 2212 7318 nw
tri 2688 7302 2704 7318 se
rect 2704 7302 4701 7318
tri 4701 7302 4717 7318 nw
tri 5036 7302 5052 7318 se
rect 5052 7302 5164 7318
tri 2113 7293 2122 7302 se
rect 2122 7293 2187 7302
tri 2187 7293 2196 7302 nw
tri 2679 7293 2688 7302 se
rect 2688 7293 4668 7302
tri 1717 7106 1733 7122 se
rect 1733 7106 1908 7122
tri 1697 7086 1717 7106 se
rect 1717 7086 1908 7106
tri 1690 7079 1697 7086 se
rect 1697 7079 1908 7086
tri 1665 7054 1690 7079 se
rect 1690 7054 1883 7079
tri 1883 7054 1908 7079 nw
tri 2092 7272 2113 7293 se
rect 2113 7272 2166 7293
tri 2166 7272 2187 7293 nw
tri 2658 7272 2679 7293 se
rect 2679 7272 4668 7293
rect 2092 7269 2163 7272
tri 2163 7269 2166 7272 nw
tri 2655 7269 2658 7272 se
rect 2658 7269 4668 7272
tri 4668 7269 4701 7302 nw
tri 5003 7269 5036 7302 se
rect 5036 7269 5164 7302
rect 2092 7268 2162 7269
tri 2162 7268 2163 7269 nw
tri 2654 7268 2655 7269 se
rect 2655 7268 4649 7269
rect 1003 7045 1863 7054
rect 1059 7034 1863 7045
tri 1863 7034 1883 7054 nw
rect 1059 7025 1854 7034
tri 1854 7025 1863 7034 nw
rect 1059 7014 1843 7025
tri 1843 7014 1854 7025 nw
tri 2081 7014 2092 7025 se
rect 2092 7014 2144 7268
tri 2144 7250 2162 7268 nw
tri 2636 7250 2654 7268 se
rect 2654 7250 4649 7268
tri 4649 7250 4668 7269 nw
tri 4984 7250 5003 7269 se
rect 5003 7263 5164 7269
rect 5220 7263 5258 7319
rect 5314 7263 5352 7319
tri 5740 7302 5760 7322 se
tri 6206 7302 6226 7322 ne
rect 6226 7305 8856 7322
rect 8912 7305 8947 7361
rect 9003 7305 9038 7361
rect 9094 7305 9129 7361
rect 9185 7305 9219 7361
rect 9275 7305 9284 7361
rect 6226 7302 9284 7305
tri 5721 7283 5740 7302 se
rect 5740 7283 5760 7302
tri 6226 7283 6245 7302 ne
rect 6245 7283 9284 7302
rect 5003 7250 5408 7263
tri 2616 7230 2636 7250 se
rect 2636 7230 4629 7250
tri 4629 7230 4649 7250 nw
tri 4964 7230 4984 7250 se
rect 4984 7230 5408 7250
tri 2564 7178 2616 7230 se
rect 2616 7178 4577 7230
tri 4577 7178 4629 7230 nw
tri 4912 7178 4964 7230 se
rect 4964 7217 5408 7230
rect 4964 7178 5164 7217
tri 2544 7158 2564 7178 se
rect 2564 7158 4557 7178
tri 4557 7158 4577 7178 nw
tri 4892 7158 4912 7178 se
rect 4912 7161 5164 7178
rect 5220 7161 5258 7217
rect 5314 7161 5352 7217
rect 4912 7158 5408 7161
tri 2508 7122 2544 7158 se
rect 2544 7126 4525 7158
tri 4525 7126 4557 7158 nw
tri 4860 7126 4892 7158 se
rect 4892 7126 5408 7158
rect 2544 7122 2778 7126
tri 2778 7122 2782 7126 nw
tri 4856 7122 4860 7126 se
rect 4860 7122 5408 7126
tri 2492 7106 2508 7122 se
rect 2508 7106 2762 7122
tri 2762 7106 2778 7122 nw
tri 4840 7106 4856 7122 se
rect 4856 7115 5408 7122
rect 4856 7106 5164 7115
tri 2476 7090 2492 7106 se
rect 2492 7090 2746 7106
tri 2746 7090 2762 7106 nw
tri 4824 7090 4840 7106 se
rect 4840 7090 5164 7106
tri 2472 7086 2476 7090 se
rect 2476 7086 2742 7090
tri 2742 7086 2746 7090 nw
tri 3103 7086 3107 7090 se
rect 3107 7086 5164 7090
tri 2436 7050 2472 7086 se
rect 2472 7050 2706 7086
tri 2706 7050 2742 7086 nw
tri 3067 7050 3103 7086 se
rect 3103 7059 5164 7086
rect 5220 7059 5258 7115
rect 5314 7059 5352 7115
rect 3103 7050 5408 7059
tri 2434 7048 2436 7050 se
rect 2436 7048 2704 7050
tri 2704 7048 2706 7050 nw
tri 3065 7048 3067 7050 se
rect 3067 7048 5408 7050
tri 2420 7034 2434 7048 se
rect 2434 7034 2690 7048
tri 2690 7034 2704 7048 nw
tri 3051 7034 3065 7048 se
rect 3065 7034 5408 7048
tri 2412 7026 2420 7034 se
rect 2420 7026 2670 7034
tri 2144 7014 2156 7026 sw
tri 2400 7014 2412 7026 se
rect 2412 7014 2670 7026
tri 2670 7014 2690 7034 nw
tri 3031 7014 3051 7034 se
rect 3051 7014 5408 7034
rect 1059 6992 1821 7014
tri 1821 6992 1843 7014 nw
tri 2059 6992 2081 7014 se
rect 2081 6992 2156 7014
tri 2156 6992 2178 7014 sw
tri 2378 6992 2400 7014 se
rect 2400 6992 2618 7014
rect 1059 6989 1769 6992
rect 1003 6965 1769 6989
rect 1059 6940 1769 6965
tri 1769 6940 1821 6992 nw
rect 2059 6940 2065 6992
rect 2117 6940 2129 6992
rect 2181 6940 2187 6992
tri 2348 6962 2378 6992 se
rect 2378 6962 2618 6992
tri 2618 6962 2670 7014 nw
tri 2979 6962 3031 7014 se
rect 3031 6962 5408 7014
tri 2329 6943 2348 6962 se
rect 2348 6943 2599 6962
tri 2599 6943 2618 6962 nw
tri 2960 6943 2979 6962 se
rect 2979 6943 5408 6962
rect 5592 7274 5970 7283
rect 5592 7218 5593 7274
rect 5649 7218 5673 7274
rect 5729 7218 5753 7274
rect 5809 7218 5833 7274
rect 5889 7218 5913 7274
rect 5969 7218 5970 7274
tri 6245 7250 6278 7283 ne
rect 6278 7250 9284 7283
tri 6278 7230 6298 7250 ne
rect 6298 7230 9284 7250
rect 5592 7186 5970 7218
rect 5592 7130 5593 7186
rect 5649 7130 5673 7186
rect 5729 7130 5753 7186
rect 5809 7130 5833 7186
rect 5889 7130 5913 7186
rect 5969 7130 5970 7186
tri 6298 7178 6350 7230 ne
rect 6350 7225 9284 7230
rect 6350 7178 8856 7225
tri 6350 7169 6359 7178 ne
rect 6359 7169 8856 7178
rect 8912 7169 8947 7225
rect 9003 7169 9038 7225
rect 9094 7169 9129 7225
rect 9185 7169 9219 7225
rect 9275 7169 9284 7225
rect 9394 7357 9403 7413
rect 9459 7357 9490 7413
rect 9546 7357 9577 7413
rect 9633 7357 9664 7413
rect 9720 7357 9750 7413
rect 9806 7357 10141 7413
rect 9394 7321 10141 7357
rect 9394 7265 9403 7321
rect 9459 7265 9490 7321
rect 9546 7265 9577 7321
rect 9633 7265 9664 7321
rect 9720 7265 9750 7321
rect 9806 7265 10141 7321
rect 9394 7229 10141 7265
rect 9394 7173 9403 7229
rect 9459 7173 9490 7229
rect 9546 7173 9577 7229
rect 9633 7173 9664 7229
rect 9720 7173 9750 7229
rect 9806 7173 10141 7229
rect 5592 7097 5970 7130
rect 5592 7041 5593 7097
rect 5649 7041 5673 7097
rect 5729 7041 5753 7097
rect 5809 7041 5833 7097
rect 5889 7041 5913 7097
rect 5969 7041 5970 7097
rect 9394 7137 10141 7173
rect 9394 7081 9403 7137
rect 9459 7081 9490 7137
rect 9546 7081 9577 7137
rect 9633 7081 9664 7137
rect 9720 7081 9750 7137
rect 9806 7081 10141 7137
rect 9394 7079 10141 7081
rect 10519 7079 10793 7459
rect 13389 7322 13398 7374
rect 13450 7322 13472 7374
rect 13524 7322 13545 7374
rect 13597 7322 13618 7374
rect 13670 7322 13691 7374
rect 13743 7322 13764 7374
rect 13816 7322 13822 7374
rect 13389 7302 13822 7322
rect 13389 7250 13398 7302
rect 13450 7250 13472 7302
rect 13524 7250 13545 7302
rect 13597 7250 13618 7302
rect 13670 7250 13691 7302
rect 13743 7250 13764 7302
rect 13816 7250 13822 7302
rect 13389 7230 13822 7250
rect 13389 7178 13398 7230
rect 13450 7178 13472 7230
rect 13524 7178 13545 7230
rect 13597 7178 13618 7230
rect 13670 7178 13691 7230
rect 13743 7178 13764 7230
rect 13816 7178 13822 7230
rect 13389 7158 13822 7178
rect 13389 7106 13398 7158
rect 13450 7106 13472 7158
rect 13524 7106 13545 7158
rect 13597 7106 13618 7158
rect 13670 7106 13691 7158
rect 13743 7106 13764 7158
rect 13816 7106 13822 7158
rect 13389 7086 13822 7106
rect 5592 7008 5970 7041
rect 5592 6952 5593 7008
rect 5649 6952 5673 7008
rect 5729 6952 5753 7008
rect 5809 6952 5833 7008
rect 5889 6952 5913 7008
rect 5969 6952 5970 7008
rect 5592 6943 5970 6952
rect 13389 7034 13398 7086
rect 13450 7034 13472 7086
rect 13524 7034 13545 7086
rect 13597 7034 13618 7086
rect 13670 7034 13691 7086
rect 13743 7034 13764 7086
rect 13816 7034 13822 7086
rect 13389 7014 13822 7034
rect 13389 6962 13398 7014
rect 13450 6962 13472 7014
rect 13524 6962 13545 7014
rect 13597 6962 13618 7014
rect 13670 6962 13691 7014
rect 13743 6962 13764 7014
rect 13816 6962 13822 7014
tri 13383 6943 13389 6949 se
rect 13389 6943 13822 6962
tri 2326 6940 2329 6943 se
rect 2329 6940 2548 6943
rect 1059 6909 1729 6940
rect 1003 6900 1729 6909
tri 1729 6900 1769 6940 nw
tri 2286 6900 2326 6940 se
rect 2326 6900 2548 6940
tri 2278 6892 2286 6900 se
rect 2286 6892 2548 6900
tri 2548 6892 2599 6943 nw
tri 2909 6892 2960 6943 se
rect 2960 6923 5408 6943
tri 5811 6942 5812 6943 ne
tri 13382 6942 13383 6943 se
rect 13383 6942 13822 6943
tri 13363 6923 13382 6942 se
rect 13382 6923 13822 6942
rect 2960 6892 3143 6923
tri 3143 6892 3174 6923 nw
tri 13332 6892 13363 6923 se
rect 13363 6892 13822 6923
tri 2274 6888 2278 6892 se
rect 2278 6888 2544 6892
tri 2544 6888 2548 6892 nw
tri 2905 6888 2909 6892 se
rect 2909 6888 3107 6892
rect 2274 6856 2512 6888
tri 2512 6856 2544 6888 nw
tri 2873 6856 2905 6888 se
rect 2905 6856 3107 6888
tri 3107 6856 3143 6892 nw
rect 193 6840 245 6846
tri -694 6791 -688 6797 se
rect -688 6791 -74 6797
tri -746 6739 -694 6791 se
rect -694 6739 -126 6791
tri -758 6727 -746 6739 se
rect -746 6727 -74 6739
rect -855 6721 -126 6727
rect -803 6675 -126 6721
rect 193 6776 245 6788
rect 193 6718 245 6724
rect -803 6669 -74 6675
rect -855 6657 -655 6669
rect -803 6648 -655 6657
tri -655 6648 -634 6669 nw
rect -803 6605 -704 6648
rect -855 6599 -704 6605
tri -704 6599 -655 6648 nw
rect 1792 6646 1801 6702
rect 1857 6700 1905 6702
rect 1961 6700 2008 6702
rect 2064 6700 2111 6702
rect 1889 6648 1905 6700
rect 1961 6648 1973 6700
rect 2092 6648 2107 6700
rect 1857 6646 1905 6648
rect 1961 6646 2008 6648
rect 2064 6646 2111 6648
rect 2167 6646 2176 6702
rect 2274 6588 2466 6856
tri 2466 6810 2512 6856 nw
tri 2827 6810 2873 6856 se
rect 2873 6810 3057 6856
tri 2823 6806 2827 6810 se
rect 2827 6806 3057 6810
tri 3057 6806 3107 6856 nw
rect 3465 6834 4731 6892
tri 13274 6834 13332 6892 se
rect 13332 6834 13822 6892
rect 3465 6806 3529 6834
tri 3529 6806 3557 6834 nw
tri 13246 6806 13274 6834 se
rect 13274 6806 13822 6834
tri 2814 6797 2823 6806 se
rect 2823 6797 3005 6806
tri 2771 6754 2814 6797 se
rect 2814 6754 3005 6797
tri 3005 6754 3057 6806 nw
tri 2743 6726 2771 6754 se
rect 2771 6726 2977 6754
tri 2977 6726 3005 6754 nw
rect 2274 6536 2280 6588
rect 2332 6536 2344 6588
rect 2396 6536 2408 6588
rect 2460 6536 2466 6588
rect 2274 6510 2466 6536
rect 2274 6458 2280 6510
rect 2332 6458 2344 6510
rect 2396 6458 2408 6510
rect 2460 6458 2466 6510
tri 2728 6711 2743 6726 se
rect 2743 6711 2962 6726
tri 2962 6711 2977 6726 nw
rect 2728 6702 2953 6711
tri 2953 6702 2962 6711 nw
rect 2728 6674 2925 6702
tri 2925 6674 2953 6702 nw
rect 2728 6646 2897 6674
tri 2897 6646 2925 6674 nw
tri 2723 6458 2728 6463 se
rect 2728 6458 2894 6646
tri 2894 6643 2897 6646 nw
tri 2692 6427 2723 6458 se
rect 2723 6427 2894 6458
tri 2672 6407 2692 6427 se
rect 2692 6407 2894 6427
tri 2625 6360 2672 6407 se
rect 2672 6360 2894 6407
rect 2292 6308 2298 6360
rect 2350 6308 2362 6360
rect 2414 6308 2426 6360
rect 2478 6308 2894 6360
rect 2292 6301 2894 6308
rect 2292 6283 2876 6301
tri 2876 6283 2894 6301 nw
rect 2972 6551 3324 6554
rect 2972 6499 2978 6551
rect 3030 6546 3050 6551
rect 3102 6546 3122 6551
rect 3174 6546 3194 6551
rect 3246 6546 3266 6551
rect 3043 6499 3050 6546
rect 3246 6499 3247 6546
rect 3318 6499 3324 6551
rect 2972 6490 2987 6499
rect 3043 6490 3074 6499
rect 3130 6490 3161 6499
rect 3217 6490 3247 6499
rect 3303 6490 3324 6499
rect 2972 6479 3324 6490
rect 2972 6427 2978 6479
rect 3030 6456 3050 6479
rect 3102 6456 3122 6479
rect 3174 6456 3194 6479
rect 3246 6456 3266 6479
rect 3043 6427 3050 6456
rect 3246 6427 3247 6456
rect 3318 6427 3324 6479
rect 2972 6407 2987 6427
rect 3043 6407 3074 6427
rect 3130 6407 3161 6427
rect 3217 6407 3247 6427
rect 3303 6407 3324 6427
rect 2972 6355 2978 6407
rect 3043 6400 3050 6407
rect 3246 6400 3247 6407
rect 3030 6366 3050 6400
rect 3102 6366 3122 6400
rect 3174 6366 3194 6400
rect 3246 6366 3266 6400
rect 3043 6355 3050 6366
rect 3246 6355 3247 6366
rect 3318 6355 3324 6407
rect 2972 6335 2987 6355
rect 3043 6335 3074 6355
rect 3130 6335 3161 6355
rect 3217 6335 3247 6355
rect 3303 6335 3324 6355
rect 2972 6283 2978 6335
rect 3043 6310 3050 6335
rect 3246 6310 3247 6335
rect 3030 6283 3050 6310
rect 3102 6283 3122 6310
rect 3174 6283 3194 6310
rect 3246 6283 3266 6310
rect 3318 6283 3324 6335
rect 2292 6282 2856 6283
rect 2292 6230 2298 6282
rect 2350 6230 2362 6282
rect 2414 6230 2426 6282
rect 2478 6263 2856 6282
tri 2856 6263 2876 6283 nw
rect 2972 6276 3324 6283
rect 2972 6263 2987 6276
rect 3043 6263 3074 6276
rect 3130 6263 3161 6276
rect 3217 6263 3247 6276
rect 3303 6263 3324 6276
rect 2478 6230 2823 6263
tri 2823 6230 2856 6263 nw
rect 2972 6211 2978 6263
rect 3043 6220 3050 6263
rect 3246 6220 3247 6263
rect 3030 6211 3050 6220
rect 3102 6211 3122 6220
rect 3174 6211 3194 6220
rect 3246 6211 3266 6220
rect 3318 6211 3324 6263
rect 2972 6208 3324 6211
rect 956 6138 962 6190
rect 1014 6138 1026 6190
rect 1078 6138 1084 6190
tri 956 6135 959 6138 ne
rect 959 6135 1084 6138
tri 959 6123 971 6135 ne
rect 971 6123 1084 6135
tri 971 6086 1008 6123 ne
rect 1008 6043 1084 6123
tri 1008 6041 1010 6043 ne
rect 1010 6041 1084 6043
tri 1010 6021 1030 6041 ne
rect 1030 6021 1084 6041
tri 1084 6021 1104 6041 sw
tri 1030 6013 1038 6021 ne
rect 1038 6013 1104 6021
tri 1104 6013 1112 6021 sw
tri 1038 5978 1073 6013 ne
rect 1073 5978 1112 6013
tri 1112 5978 1147 6013 sw
tri 1073 5967 1084 5978 ne
rect 1084 5967 1147 5978
tri 1084 5961 1090 5967 ne
rect 1090 5961 1147 5967
tri 1147 5961 1164 5978 sw
rect 3465 5976 3523 6806
tri 3523 6800 3529 6806 nw
rect 3599 6754 3605 6806
rect 3657 6754 3669 6806
rect 3721 6754 4731 6806
tri 13194 6754 13246 6806 se
rect 13246 6754 13822 6806
tri 13166 6726 13194 6754 se
rect 13194 6726 13822 6754
rect 3633 6674 3639 6726
rect 3691 6674 3703 6726
rect 3755 6674 4731 6726
tri 13115 6675 13166 6726 se
rect 13166 6675 13822 6726
tri 3619 6601 3659 6641 se
rect 3659 6601 4731 6641
rect 3619 6589 4731 6601
rect 8847 6619 8856 6675
rect 8912 6619 8947 6675
rect 9003 6619 9038 6675
rect 9094 6619 9129 6675
rect 9185 6619 9219 6675
rect 9275 6619 13822 6675
rect 8847 6595 13822 6619
tri 3523 5976 3547 6000 sw
tri 3465 5961 3480 5976 ne
rect 3480 5961 3547 5976
tri 3547 5961 3562 5976 sw
rect 3619 5961 3671 6589
tri 3671 6535 3725 6589 nw
rect 8847 6539 8856 6595
rect 8912 6539 8947 6595
rect 9003 6539 9038 6595
rect 9094 6539 9129 6595
rect 9185 6539 9219 6595
rect 9275 6539 13822 6595
rect 8847 6515 13822 6539
rect 8847 6459 8856 6515
rect 8912 6459 8947 6515
rect 9003 6459 9038 6515
rect 9094 6459 9129 6515
rect 9185 6459 9219 6515
rect 9275 6459 13822 6515
rect 8847 6435 13822 6459
tri 4287 6377 4303 6393 se
rect 4303 6377 4731 6393
rect 3712 6371 3764 6377
tri 4276 6366 4287 6377 se
rect 4287 6366 4731 6377
rect 8847 6379 8856 6435
rect 8912 6379 8947 6435
rect 9003 6379 9038 6435
rect 9094 6379 9129 6435
rect 9185 6379 9219 6435
rect 9275 6379 13822 6435
rect 8847 6376 13822 6379
tri 3764 6332 3798 6366 sw
tri 4242 6332 4276 6366 se
rect 4276 6341 4731 6366
tri 13089 6341 13124 6376 ne
rect 13124 6341 13822 6376
rect 4276 6332 4316 6341
tri 4316 6332 4325 6341 nw
tri 13124 6332 13133 6341 ne
rect 13133 6332 13822 6341
rect 3764 6319 4264 6332
rect 3712 6307 4264 6319
rect 3764 6280 4264 6307
tri 4264 6280 4316 6332 nw
tri 13133 6308 13157 6332 ne
rect 13157 6308 13822 6332
tri 4375 6280 4403 6308 se
rect 4403 6280 4731 6308
rect 3712 6249 3764 6255
tri 3764 6249 3795 6280 nw
tri 4344 6249 4375 6280 se
rect 4375 6256 4731 6280
tri 13157 6256 13209 6308 ne
rect 13209 6256 13822 6308
rect 4375 6249 4418 6256
tri 4418 6249 4425 6256 nw
tri 13209 6249 13216 6256 ne
rect 13216 6249 13822 6256
rect 3895 6197 3901 6249
rect 3953 6197 3965 6249
rect 4017 6197 4366 6249
tri 4366 6197 4418 6249 nw
tri 13216 6228 13237 6249 ne
rect 13237 6228 13822 6249
tri 4454 6197 4485 6228 se
rect 4485 6197 4731 6228
tri 4450 6193 4454 6197 se
rect 4454 6193 4731 6197
rect 3721 6187 3773 6193
tri 3773 6169 3797 6193 sw
tri 4426 6169 4450 6193 se
rect 4450 6176 4731 6193
tri 13237 6176 13289 6228 ne
rect 13289 6176 13822 6228
rect 4450 6169 4500 6176
tri 4500 6169 4507 6176 nw
tri 13289 6169 13296 6176 ne
rect 13296 6169 13822 6176
rect 3773 6148 4479 6169
tri 4479 6148 4500 6169 nw
tri 13296 6148 13317 6169 ne
rect 13317 6148 13822 6169
rect 3773 6135 4458 6148
rect 3721 6127 4458 6135
tri 4458 6127 4479 6148 nw
tri 4519 6127 4540 6148 se
rect 4540 6127 4731 6148
rect 3721 6123 4448 6127
rect 3773 6117 4448 6123
tri 4448 6117 4458 6127 nw
tri 4509 6117 4519 6127 se
rect 4519 6117 4731 6127
tri 13317 6117 13348 6148 ne
rect 13348 6117 13822 6148
rect 3773 6076 3774 6117
tri 3774 6076 3815 6117 nw
tri 4468 6076 4509 6117 se
rect 4509 6090 4731 6117
tri 13348 6090 13375 6117 ne
rect 13375 6090 13822 6117
rect 4509 6076 4550 6090
tri 4550 6076 4564 6090 nw
tri 13375 6076 13389 6090 ne
tri 3773 6075 3774 6076 nw
tri 4467 6075 4468 6076 se
rect 4468 6075 4540 6076
rect 3721 6065 3773 6071
tri 4458 6066 4467 6075 se
rect 4467 6066 4540 6075
tri 4540 6066 4550 6076 nw
tri 4457 6065 4458 6066 se
rect 4458 6065 4533 6066
tri 4451 6059 4457 6065 se
rect 4457 6059 4533 6065
tri 4533 6059 4540 6066 nw
rect 3894 6040 4514 6059
tri 4514 6040 4533 6059 nw
rect 3894 6021 4495 6040
tri 4495 6021 4514 6040 nw
rect 5592 6031 5970 6040
rect 3894 6013 4487 6021
tri 4487 6013 4495 6021 nw
rect 3894 6001 4475 6013
tri 4475 6001 4487 6013 nw
rect 3894 5968 3947 6001
tri 3947 5968 3980 6001 nw
tri 3671 5961 3678 5968 sw
tri 1090 5955 1096 5961 ne
rect 1096 5955 1164 5961
tri 1164 5955 1170 5961 sw
tri 3480 5955 3486 5961 ne
rect 3486 5955 3562 5961
tri 3562 5955 3568 5961 sw
rect 3619 5955 3678 5961
tri 3678 5955 3684 5961 sw
tri 1096 5904 1147 5955 ne
rect 1147 5904 1170 5955
tri 1170 5904 1221 5955 sw
tri 3486 5904 3537 5955 ne
rect 3537 5946 3568 5955
tri 3568 5946 3577 5955 sw
rect 3619 5946 3684 5955
tri 3684 5946 3693 5955 sw
rect 3537 5904 3577 5946
tri 3577 5904 3619 5946 sw
tri 3619 5904 3661 5946 ne
rect 3661 5904 3693 5946
tri 1147 5903 1148 5904 ne
rect 1148 5903 1221 5904
tri 1221 5903 1222 5904 sw
tri 3537 5903 3538 5904 ne
rect 3538 5903 3619 5904
tri 3619 5903 3620 5904 sw
tri 3661 5903 3662 5904 ne
rect 3662 5903 3693 5904
tri 3693 5903 3736 5946 sw
tri 1148 5891 1160 5903 ne
rect 1160 5894 1222 5903
tri 1222 5894 1231 5903 sw
tri 3538 5894 3547 5903 ne
rect 3547 5894 3620 5903
tri 3620 5894 3629 5903 sw
tri 3662 5894 3671 5903 ne
rect 3671 5894 3736 5903
rect 1160 5891 1231 5894
tri 1231 5891 1234 5894 sw
tri 3547 5891 3550 5894 ne
rect 3550 5891 3629 5894
tri 3629 5891 3632 5894 sw
tri 3671 5891 3674 5894 ne
rect 3674 5891 3736 5894
tri 3736 5891 3748 5903 sw
tri 1160 5871 1180 5891 ne
rect 1180 5883 1234 5891
tri 1234 5883 1242 5891 sw
tri 3550 5883 3558 5891 ne
rect 3558 5883 3632 5891
tri 3632 5883 3640 5891 sw
tri 3674 5883 3682 5891 ne
rect 3682 5883 3748 5891
rect 1180 5877 1242 5883
tri 1242 5877 1248 5883 sw
tri 3558 5877 3564 5883 ne
rect 3564 5877 3640 5883
rect 1180 5871 1248 5877
tri 1248 5871 1254 5877 sw
rect 2805 5871 2857 5877
tri 1180 5830 1221 5871 ne
rect 1221 5830 1254 5871
tri 1254 5830 1295 5871 sw
tri 1221 5819 1232 5830 ne
rect 1232 5819 1295 5830
tri 1295 5819 1306 5830 sw
tri 2857 5853 2881 5877 sw
tri 3564 5853 3588 5877 ne
rect 3588 5872 3640 5877
tri 3640 5872 3651 5883 sw
tri 3682 5872 3693 5883 ne
rect 3693 5872 3748 5883
tri 3748 5872 3767 5891 sw
rect 3588 5853 3651 5872
rect 2857 5839 3532 5853
tri 3532 5839 3546 5853 sw
tri 3588 5839 3602 5853 ne
rect 3602 5839 3651 5853
tri 3651 5839 3684 5872 sw
tri 3693 5839 3726 5872 ne
rect 3726 5839 3767 5872
tri 3767 5839 3800 5872 sw
rect 2857 5838 3546 5839
tri 3546 5838 3547 5839 sw
tri 3602 5838 3603 5839 ne
rect 3603 5838 3684 5839
rect 2857 5829 3547 5838
tri 3547 5829 3556 5838 sw
tri 3603 5829 3612 5838 ne
rect 3612 5830 3684 5838
tri 3684 5830 3693 5839 sw
tri 3726 5830 3735 5839 ne
rect 3735 5830 3800 5839
rect 3612 5829 3693 5830
tri 3693 5829 3694 5830 sw
tri 3735 5829 3736 5830 ne
rect 3736 5829 3800 5830
tri 3800 5829 3810 5839 sw
rect 2857 5825 3556 5829
tri 3556 5825 3560 5829 sw
tri 3612 5825 3616 5829 ne
rect 3616 5825 3694 5829
tri 3694 5825 3698 5829 sw
tri 3736 5825 3740 5829 ne
rect 3740 5825 3810 5829
tri 3810 5825 3814 5829 sw
rect 2857 5819 3560 5825
tri 1232 5807 1244 5819 ne
rect 1244 5807 1306 5819
tri 1306 5807 1318 5819 sw
rect 2805 5812 3560 5819
tri 3560 5812 3573 5825 sw
tri 3616 5812 3629 5825 ne
rect 3629 5812 3698 5825
tri 3698 5812 3711 5825 sw
tri 3740 5812 3753 5825 ne
rect 3753 5812 3814 5825
rect 2805 5807 3573 5812
tri 1244 5756 1295 5807 ne
rect 1295 5756 1318 5807
tri 1318 5756 1369 5807 sw
tri 1295 5749 1302 5756 ne
rect 1302 5749 2000 5756
tri 1302 5730 1321 5749 ne
rect 1321 5730 2000 5749
tri 1321 5719 1332 5730 ne
rect 1332 5719 2000 5730
tri 405 5704 420 5719 sw
tri 1332 5704 1347 5719 ne
rect 1347 5704 2000 5719
rect 2052 5704 2064 5756
rect 2116 5704 2122 5756
rect 2857 5805 3573 5807
tri 3573 5805 3580 5812 sw
tri 3629 5805 3636 5812 ne
rect 3636 5805 3711 5812
tri 3711 5805 3718 5812 sw
tri 3753 5805 3760 5812 ne
rect 3760 5805 3814 5812
tri 3814 5805 3834 5825 sw
rect 3894 5805 3946 5968
tri 3946 5967 3947 5968 nw
rect 4571 5961 4577 6013
rect 4629 5961 4645 6013
rect 4697 5961 4703 6013
rect 4036 5955 4088 5961
rect 4036 5891 4088 5903
tri 3946 5805 3950 5809 sw
rect 2857 5801 3580 5805
tri 2857 5767 2891 5801 nw
tri 3510 5767 3544 5801 ne
rect 3544 5767 3580 5801
tri 3544 5755 3556 5767 ne
rect 3556 5756 3580 5767
tri 3580 5756 3629 5805 sw
tri 3636 5774 3667 5805 ne
rect 3667 5798 3718 5805
tri 3718 5798 3725 5805 sw
tri 3760 5798 3767 5805 ne
rect 3767 5798 3834 5805
tri 3834 5798 3841 5805 sw
rect 3894 5798 3950 5805
tri 3950 5798 3957 5805 sw
rect 3667 5774 3725 5798
tri 3725 5774 3749 5798 sw
tri 3767 5774 3791 5798 ne
rect 3791 5774 3841 5798
tri 3841 5774 3865 5798 sw
rect 3894 5787 3957 5798
tri 3957 5787 3968 5798 sw
tri 3894 5774 3907 5787 ne
rect 3907 5774 3968 5787
tri 3667 5756 3685 5774 ne
rect 3685 5756 3749 5774
tri 3749 5756 3767 5774 sw
tri 3791 5756 3809 5774 ne
rect 3809 5756 3865 5774
rect 3556 5755 3629 5756
tri 3629 5755 3630 5756 sw
tri 3685 5755 3686 5756 ne
rect 3686 5755 3767 5756
tri 3767 5755 3768 5756 sw
tri 3809 5755 3810 5756 ne
rect 3810 5755 3865 5756
tri 3865 5755 3884 5774 sw
tri 3907 5755 3926 5774 ne
rect 3926 5755 3968 5774
tri 3968 5755 4000 5787 sw
rect 4036 5774 4088 5839
rect 4571 5935 4703 5961
rect 4571 5883 4577 5935
rect 4629 5883 4645 5935
rect 4697 5883 4703 5935
rect 5592 5975 5593 6031
rect 5649 5975 5673 6031
rect 5729 5975 5753 6031
rect 5809 5975 5833 6031
rect 5889 5975 5913 6031
rect 5969 5975 5970 6031
rect 4571 5853 4703 5883
rect 5164 5924 5408 5933
rect 5220 5868 5258 5924
rect 5314 5868 5352 5924
tri 4703 5853 4704 5854 sw
rect 4571 5839 4704 5853
tri 4571 5829 4581 5839 ne
rect 4581 5829 4704 5839
tri 4704 5829 4728 5853 sw
tri 4581 5825 4585 5829 ne
rect 4585 5825 4728 5829
tri 4728 5825 4732 5829 sw
tri 4585 5805 4605 5825 ne
rect 4605 5805 4732 5825
tri 4732 5805 4752 5825 sw
rect 5164 5822 5408 5868
tri 4605 5783 4627 5805 ne
rect 4627 5783 4752 5805
tri 4088 5774 4097 5783 sw
tri 4627 5774 4636 5783 ne
rect 4636 5774 4752 5783
tri 4752 5774 4783 5805 sw
rect 4036 5768 4097 5774
tri 4097 5768 4103 5774 sw
tri 4636 5768 4642 5774 ne
rect 4642 5768 4783 5774
rect 4036 5761 4103 5768
tri 4036 5755 4042 5761 ne
rect 4042 5755 4103 5761
tri 4103 5755 4116 5768 sw
tri 4642 5755 4655 5768 ne
rect 4655 5755 4783 5768
tri 4783 5755 4802 5774 sw
rect 5220 5766 5258 5822
rect 5314 5766 5352 5822
rect 2805 5749 2857 5755
tri 3556 5753 3558 5755 ne
rect 3558 5753 3630 5755
tri 3630 5753 3632 5755 sw
tri 3686 5753 3688 5755 ne
rect 3688 5753 3768 5755
tri 3768 5753 3770 5755 sw
tri 3810 5753 3812 5755 ne
rect 3812 5753 3884 5755
tri 3884 5753 3886 5755 sw
tri 3926 5753 3928 5755 ne
rect 3928 5753 4000 5755
tri 4000 5753 4002 5755 sw
tri 4042 5753 4044 5755 ne
rect 4044 5753 4116 5755
tri 4116 5753 4118 5755 sw
tri 4655 5753 4657 5755 ne
rect 4657 5753 4802 5755
tri 4802 5753 4804 5755 sw
tri 3558 5749 3562 5753 ne
rect 3562 5749 3632 5753
tri 3562 5743 3568 5749 ne
rect 3568 5743 3632 5749
tri 3442 5737 3448 5743 se
rect 3448 5737 3500 5743
tri 3435 5730 3442 5737 se
rect 3442 5730 3448 5737
tri 3426 5721 3435 5730 se
rect 3435 5721 3448 5730
rect 405 5685 420 5704
tri 420 5685 439 5704 sw
rect 2473 5669 2479 5721
rect 2531 5669 2543 5721
rect 2595 5685 3448 5721
tri 3568 5733 3578 5743 ne
rect 3578 5733 3632 5743
tri 3632 5733 3652 5753 sw
tri 3688 5733 3708 5753 ne
rect 3708 5733 3770 5753
tri 3770 5733 3790 5753 sw
tri 3812 5733 3832 5753 ne
rect 3832 5745 3886 5753
tri 3886 5745 3894 5753 sw
tri 3928 5745 3936 5753 ne
rect 3936 5745 4002 5753
rect 3832 5733 3894 5745
tri 3894 5733 3906 5745 sw
tri 3936 5733 3948 5745 ne
rect 3948 5733 4002 5745
tri 4002 5733 4022 5753 sw
tri 4044 5733 4064 5753 ne
rect 4064 5733 4118 5753
tri 4118 5733 4138 5753 sw
tri 4657 5733 4677 5753 ne
rect 4677 5733 4804 5753
tri 4804 5733 4824 5753 sw
tri 3578 5730 3581 5733 ne
rect 3581 5730 3652 5733
tri 3652 5730 3655 5733 sw
tri 3708 5730 3711 5733 ne
rect 3711 5730 3790 5733
tri 3790 5730 3793 5733 sw
tri 3832 5730 3835 5733 ne
rect 3835 5730 3906 5733
rect 2595 5673 3500 5685
tri 3581 5681 3630 5730 ne
rect 3630 5681 3655 5730
tri 3655 5681 3704 5730 sw
tri 3711 5707 3734 5730 ne
rect 3734 5724 3793 5730
tri 3793 5724 3799 5730 sw
tri 3835 5724 3841 5730 ne
rect 3841 5724 3906 5730
tri 3906 5724 3915 5733 sw
tri 3948 5724 3957 5733 ne
rect 3957 5724 4022 5733
tri 4022 5724 4031 5733 sw
tri 4064 5724 4073 5733 ne
rect 4073 5724 4138 5733
tri 4138 5724 4147 5733 sw
tri 4677 5724 4686 5733 ne
rect 4686 5724 4824 5733
rect 3734 5707 3799 5724
tri 3799 5707 3816 5724 sw
tri 3841 5707 3858 5724 ne
rect 3858 5713 3915 5724
tri 3915 5713 3926 5724 sw
tri 3957 5713 3968 5724 ne
rect 3968 5713 4031 5724
tri 4031 5713 4042 5724 sw
tri 4073 5713 4084 5724 ne
rect 4084 5713 4147 5724
rect 3858 5707 3926 5713
tri 3926 5707 3932 5713 sw
tri 3968 5707 3974 5713 ne
rect 3974 5707 4042 5713
tri 4042 5707 4048 5713 sw
tri 4084 5707 4090 5713 ne
rect 4090 5707 4147 5713
tri 4147 5707 4164 5724 sw
tri 4686 5707 4703 5724 ne
rect 4703 5707 4824 5724
tri 3734 5681 3760 5707 ne
rect 3760 5682 3816 5707
tri 3816 5682 3841 5707 sw
tri 3858 5682 3883 5707 ne
rect 3883 5682 3932 5707
rect 3760 5681 3841 5682
tri 3841 5681 3842 5682 sw
tri 3883 5681 3884 5682 ne
rect 3884 5681 3932 5682
tri 3932 5681 3958 5707 sw
tri 3974 5694 3987 5707 ne
rect 3987 5694 4048 5707
tri 4048 5694 4061 5707 sw
tri 4090 5694 4103 5707 ne
rect 4103 5694 4164 5707
tri 4164 5694 4177 5707 sw
tri 4703 5694 4716 5707 ne
rect 4716 5694 4824 5707
tri 3987 5681 4000 5694 ne
rect 4000 5681 4061 5694
tri 4061 5681 4074 5694 sw
tri 4103 5681 4116 5694 ne
rect 4116 5681 4177 5694
tri 4177 5681 4190 5694 sw
tri 4716 5681 4729 5694 ne
rect 4729 5681 4824 5694
tri 4824 5681 4876 5733 sw
rect 5164 5720 5408 5766
rect 2595 5669 3448 5673
tri 3394 5621 3442 5669 ne
rect 3442 5621 3448 5669
tri 3630 5661 3650 5681 ne
rect 3650 5674 3704 5681
tri 3704 5674 3711 5681 sw
tri 3760 5674 3767 5681 ne
rect 3767 5674 3842 5681
rect 3650 5661 3711 5674
tri 3711 5661 3724 5674 sw
tri 3767 5661 3780 5674 ne
rect 3780 5661 3842 5674
tri 3842 5661 3862 5681 sw
tri 3884 5661 3904 5681 ne
rect 3904 5671 3958 5681
tri 3958 5671 3968 5681 sw
tri 4000 5671 4010 5681 ne
rect 4010 5671 4074 5681
rect 3904 5661 3968 5671
tri 3968 5661 3978 5671 sw
tri 4010 5661 4020 5671 ne
rect 4020 5661 4074 5671
tri 4074 5661 4094 5681 sw
tri 4116 5661 4136 5681 ne
rect 4136 5661 4190 5681
tri 4190 5661 4210 5681 sw
tri 4729 5661 4749 5681 ne
rect 4749 5661 4876 5681
tri 4876 5661 4896 5681 sw
rect 5220 5664 5258 5720
rect 5314 5664 5352 5720
tri 3650 5633 3678 5661 ne
rect 3678 5648 3724 5661
tri 3724 5648 3737 5661 sw
tri 3780 5648 3793 5661 ne
rect 3793 5650 3862 5661
tri 3862 5650 3873 5661 sw
tri 3904 5650 3915 5661 ne
rect 3915 5650 3978 5661
tri 3978 5650 3989 5661 sw
tri 4020 5650 4031 5661 ne
rect 4031 5650 4094 5661
tri 4094 5650 4105 5661 sw
tri 4136 5650 4147 5661 ne
rect 4147 5650 4210 5661
tri 4210 5650 4221 5661 sw
tri 4749 5650 4760 5661 ne
rect 4760 5650 4896 5661
rect 3793 5648 3873 5650
tri 3873 5648 3875 5650 sw
tri 3915 5648 3917 5650 ne
rect 3917 5648 3989 5650
rect 3678 5633 3737 5648
tri 3737 5633 3752 5648 sw
tri 3793 5633 3808 5648 ne
rect 3808 5633 3875 5648
tri 3875 5633 3890 5648 sw
tri 3917 5633 3932 5648 ne
rect 3932 5639 3989 5648
tri 3989 5639 4000 5650 sw
tri 4031 5639 4042 5650 ne
rect 4042 5639 4105 5650
tri 4105 5639 4116 5650 sw
tri 4147 5639 4158 5650 ne
rect 4158 5639 4221 5650
rect 3932 5633 4000 5639
tri 4000 5633 4006 5639 sw
tri 4042 5633 4048 5639 ne
rect 4048 5633 4116 5639
tri 4116 5633 4122 5639 sw
tri 4158 5633 4164 5639 ne
rect 4164 5633 4221 5639
tri 4221 5633 4238 5650 sw
tri 4760 5633 4777 5650 ne
rect 4777 5633 4896 5650
tri 3442 5615 3448 5621 ne
rect 3448 5615 3500 5621
tri 3678 5615 3696 5633 ne
rect 3696 5615 3752 5633
tri 3696 5607 3704 5615 ne
rect 3704 5607 3752 5615
tri 3752 5607 3778 5633 sw
tri 3808 5607 3834 5633 ne
rect 3834 5608 3890 5633
tri 3890 5608 3915 5633 sw
tri 3932 5608 3957 5633 ne
rect 3957 5608 4006 5633
rect 3834 5607 3915 5608
tri 3704 5606 3705 5607 ne
rect 3705 5606 3778 5607
tri 2897 5599 2904 5606 se
rect 2904 5470 2913 5606
rect 3049 5470 3058 5606
tri 3058 5599 3065 5606 sw
tri 3705 5599 3712 5606 ne
rect 3712 5599 3778 5606
tri 3712 5598 3713 5599 ne
rect 3713 5598 3778 5599
rect 3129 5470 3137 5598
tri 3713 5581 3730 5598 ne
rect 3730 5592 3778 5598
tri 3778 5592 3793 5607 sw
tri 3834 5592 3849 5607 ne
rect 3849 5592 3915 5607
rect 3730 5581 3793 5592
tri 3793 5581 3804 5592 sw
tri 3849 5581 3860 5592 ne
rect 3860 5581 3915 5592
tri 3915 5581 3942 5608 sw
tri 3957 5581 3984 5608 ne
rect 3984 5597 4006 5608
tri 4006 5597 4042 5633 sw
tri 4048 5620 4061 5633 ne
rect 4061 5620 4122 5633
tri 4122 5620 4135 5633 sw
tri 4164 5620 4177 5633 ne
rect 4177 5620 4238 5633
tri 4238 5620 4251 5633 sw
tri 4061 5597 4084 5620 ne
rect 4084 5607 4135 5620
tri 4135 5607 4148 5620 sw
tri 4177 5607 4190 5620 ne
rect 4190 5607 4251 5620
rect 4084 5597 4148 5607
rect 3984 5581 4042 5597
tri 4042 5581 4058 5597 sw
tri 4084 5581 4100 5597 ne
rect 4100 5581 4148 5597
tri 4148 5581 4174 5607 sw
tri 4190 5581 4216 5607 ne
rect 4216 5581 4251 5607
tri 4251 5581 4290 5620 sw
rect 4409 5581 4415 5633
rect 4467 5581 4483 5633
rect 4535 5627 4688 5633
tri 4688 5627 4694 5633 sw
tri 4777 5627 4783 5633 ne
rect 4783 5627 4896 5633
tri 4896 5627 4930 5661 sw
rect 4535 5615 4694 5627
tri 4694 5615 4706 5627 sw
tri 4783 5615 4795 5627 ne
rect 4795 5615 4930 5627
rect 4535 5609 4706 5615
tri 4706 5609 4712 5615 sw
tri 4795 5609 4801 5615 ne
rect 4801 5609 4930 5615
tri 4930 5609 4948 5627 sw
rect 5164 5618 5408 5664
rect 4535 5607 4712 5609
tri 4712 5607 4714 5609 sw
tri 4801 5607 4803 5609 ne
rect 4803 5607 4948 5609
tri 4948 5607 4950 5609 sw
rect 4535 5581 4714 5607
tri 3730 5555 3756 5581 ne
rect 3756 5566 3804 5581
tri 3804 5566 3819 5581 sw
tri 3860 5566 3875 5581 ne
rect 3875 5576 3942 5581
tri 3942 5576 3947 5581 sw
tri 3984 5576 3989 5581 ne
rect 3989 5576 4058 5581
tri 4058 5576 4063 5581 sw
tri 4100 5576 4105 5581 ne
rect 4105 5576 4174 5581
tri 4174 5576 4179 5581 sw
tri 4216 5576 4221 5581 ne
rect 4221 5576 4290 5581
tri 4290 5576 4295 5581 sw
rect 3875 5566 3947 5576
tri 3947 5566 3957 5576 sw
tri 3989 5566 3999 5576 ne
rect 3999 5566 4063 5576
rect 3756 5555 3819 5566
tri 3819 5555 3830 5566 sw
tri 3875 5555 3886 5566 ne
rect 3886 5555 3957 5566
tri 3957 5555 3968 5566 sw
tri 3999 5555 4010 5566 ne
rect 4010 5565 4063 5566
tri 4063 5565 4074 5576 sw
tri 4105 5565 4116 5576 ne
rect 4116 5565 4179 5576
tri 4179 5565 4190 5576 sw
tri 4221 5565 4232 5576 ne
rect 4232 5565 4295 5576
rect 4010 5555 4074 5565
tri 4074 5555 4084 5565 sw
tri 4116 5555 4126 5565 ne
rect 4126 5555 4190 5565
tri 4190 5555 4200 5565 sw
tri 4232 5555 4242 5565 ne
rect 4242 5555 4295 5565
tri 4295 5555 4316 5576 sw
rect 4409 5555 4714 5581
tri 3756 5549 3762 5555 ne
rect 3762 5549 3830 5555
rect 3535 5497 3541 5549
rect 3593 5497 3605 5549
rect 3657 5497 3663 5549
tri 3762 5533 3778 5549 ne
rect 3778 5510 3830 5549
tri 3830 5510 3875 5555 sw
tri 3886 5510 3931 5555 ne
rect 3931 5534 3968 5555
tri 3968 5534 3989 5555 sw
tri 4010 5534 4031 5555 ne
rect 4031 5534 4084 5555
rect 3931 5510 3989 5534
rect 3778 5503 3875 5510
tri 3875 5503 3882 5510 sw
tri 3931 5503 3938 5510 ne
rect 3938 5503 3989 5510
tri 3989 5503 4020 5534 sw
tri 4031 5503 4062 5534 ne
rect 4062 5523 4084 5534
tri 4084 5523 4116 5555 sw
tri 4126 5546 4135 5555 ne
rect 4135 5546 4200 5555
tri 4200 5546 4209 5555 sw
tri 4242 5546 4251 5555 ne
rect 4251 5546 4316 5555
tri 4316 5546 4325 5555 sw
tri 4135 5523 4158 5546 ne
rect 4158 5533 4209 5546
tri 4209 5533 4222 5546 sw
tri 4251 5533 4264 5546 ne
rect 4264 5533 4325 5546
rect 4158 5523 4222 5533
rect 4062 5503 4116 5523
tri 4116 5503 4136 5523 sw
tri 4158 5503 4178 5523 ne
rect 4178 5503 4222 5523
tri 4222 5503 4252 5533 sw
tri 4264 5503 4294 5533 ne
rect 4294 5503 4325 5533
tri 4325 5503 4368 5546 sw
rect 4409 5503 4415 5555
rect 4467 5503 4483 5555
rect 4535 5520 4714 5555
tri 4714 5520 4801 5607 sw
tri 4803 5520 4890 5607 ne
rect 4890 5599 4950 5607
tri 4950 5599 4958 5607 sw
rect 4890 5520 4958 5599
rect 4535 5503 4801 5520
rect 3535 5470 3620 5497
tri 3620 5470 3647 5497 nw
rect 3778 5484 3882 5503
tri 3882 5484 3901 5503 sw
tri 3938 5484 3957 5503 ne
rect 3957 5502 4020 5503
tri 4020 5502 4021 5503 sw
tri 4062 5502 4063 5503 ne
rect 4063 5502 4136 5503
tri 4136 5502 4137 5503 sw
tri 4178 5502 4179 5503 ne
rect 4179 5502 4252 5503
tri 4252 5502 4253 5503 sw
tri 4294 5502 4295 5503 ne
rect 4295 5502 4368 5503
tri 4368 5502 4369 5503 sw
tri 4634 5502 4635 5503 ne
rect 4635 5502 4801 5503
rect 3957 5484 4021 5502
tri 4021 5484 4039 5502 sw
tri 4063 5484 4081 5502 ne
rect 4081 5491 4137 5502
tri 4137 5491 4148 5502 sw
tri 4179 5491 4190 5502 ne
rect 4190 5491 4253 5502
tri 4253 5491 4264 5502 sw
tri 4295 5491 4306 5502 ne
rect 4306 5491 4369 5502
rect 4081 5484 4148 5491
rect 3778 5479 3901 5484
tri 3901 5479 3906 5484 sw
rect 3535 5469 3619 5470
tri 3619 5469 3620 5470 nw
tri 1259 5435 1293 5469 sw
tri 3501 5351 3535 5385 se
rect 3535 5351 3613 5469
tri 3613 5463 3619 5469 nw
tri 1426 5337 1439 5350 se
tri 1426 5299 1438 5311 ne
rect 1438 5299 1440 5311
rect 3485 5299 3491 5351
rect 3543 5299 3555 5351
rect 3607 5299 3613 5351
rect 3778 5346 3906 5479
tri 3957 5431 4010 5484 ne
rect 4010 5460 4039 5484
tri 4039 5460 4063 5484 sw
tri 4081 5460 4105 5484 ne
rect 4105 5460 4148 5484
rect 4010 5431 4063 5460
tri 4063 5431 4092 5460 sw
tri 4105 5431 4134 5460 ne
rect 4134 5449 4148 5460
tri 4148 5449 4190 5491 sw
tri 4190 5472 4209 5491 ne
rect 4209 5472 4264 5491
tri 4264 5472 4283 5491 sw
tri 4306 5472 4325 5491 ne
rect 4325 5472 4369 5491
tri 4369 5472 4399 5502 sw
tri 4635 5472 4665 5502 ne
rect 4665 5480 4801 5502
tri 4801 5480 4841 5520 sw
tri 4890 5480 4930 5520 ne
rect 4930 5480 4958 5520
tri 4958 5480 5077 5599 sw
rect 5220 5562 5258 5618
rect 5314 5562 5352 5618
rect 5592 5929 5970 5975
rect 5592 5873 5593 5929
rect 5649 5873 5673 5929
rect 5729 5873 5753 5929
rect 5809 5873 5833 5929
rect 5889 5873 5913 5929
rect 5969 5873 5970 5929
rect 13389 6021 13822 6090
rect 13389 5969 13398 6021
rect 13450 5969 13472 6021
rect 13524 5969 13545 6021
rect 13597 5969 13618 6021
rect 13670 5969 13691 6021
rect 13743 5969 13764 6021
rect 13816 5969 13822 6021
rect 13389 5949 13822 5969
tri 9416 5897 9422 5903 se
rect 9422 5897 10200 5903
tri 9402 5883 9416 5897 se
rect 9416 5883 10200 5897
tri 9396 5877 9402 5883 se
rect 9402 5877 10200 5883
rect 5592 5827 5970 5873
tri 9373 5854 9396 5877 se
rect 9396 5854 10200 5877
tri 9372 5853 9373 5854 se
rect 9373 5853 10200 5854
tri 9348 5829 9372 5853 se
rect 9372 5839 10200 5853
rect 9372 5829 9403 5839
rect 5592 5771 5593 5827
rect 5649 5771 5673 5827
rect 5729 5771 5753 5827
rect 5809 5771 5833 5827
rect 5889 5771 5913 5827
rect 5969 5771 5970 5827
tri 9344 5825 9348 5829 se
rect 9348 5825 9403 5829
tri 9324 5805 9344 5825 se
rect 9344 5805 9403 5825
tri 9293 5774 9324 5805 se
rect 9324 5783 9403 5805
rect 9459 5783 9489 5839
rect 9545 5783 9575 5839
rect 9631 5783 9661 5839
rect 9717 5783 9746 5839
rect 9802 5783 10200 5839
rect 9324 5774 10200 5783
rect 5592 5725 5970 5771
tri 9274 5755 9293 5774 se
rect 9293 5755 10200 5774
tri 9272 5753 9274 5755 se
rect 9274 5753 10200 5755
tri 9252 5733 9272 5753 se
rect 9272 5735 10200 5753
rect 9272 5733 9403 5735
rect 5592 5669 5593 5725
rect 5649 5669 5673 5725
rect 5729 5669 5753 5725
rect 5809 5669 5833 5725
rect 5889 5669 5913 5725
rect 5969 5669 5970 5725
tri 9200 5681 9252 5733 se
rect 9252 5681 9403 5733
rect 5592 5660 5970 5669
tri 9180 5661 9200 5681 se
rect 9200 5679 9403 5681
rect 9459 5679 9489 5735
rect 9545 5679 9575 5735
rect 9631 5679 9661 5735
rect 9717 5679 9746 5735
rect 9802 5679 10200 5735
rect 9200 5661 10200 5679
tri 9179 5660 9180 5661 se
rect 9180 5660 10200 5661
rect 5592 5627 5804 5660
tri 5804 5627 5837 5660 nw
tri 9172 5653 9179 5660 se
rect 9179 5653 10200 5660
tri 6184 5627 6210 5653 se
rect 6210 5631 10200 5653
rect 6210 5627 9403 5631
rect 5592 5609 5786 5627
tri 5786 5609 5804 5627 nw
tri 6166 5609 6184 5627 se
rect 6184 5609 9403 5627
rect 5592 5607 5784 5609
tri 5784 5607 5786 5609 nw
tri 6164 5607 6166 5609 se
rect 6166 5607 9403 5609
rect 5592 5599 5776 5607
tri 5776 5599 5784 5607 nw
tri 6156 5599 6164 5607 se
rect 6164 5599 9403 5607
rect 5164 5553 5408 5562
tri 5546 5553 5592 5599 se
rect 5592 5553 5657 5599
tri 5473 5480 5546 5553 se
rect 5546 5480 5657 5553
tri 5657 5480 5776 5599 nw
tri 6037 5480 6156 5599 se
rect 6156 5575 9403 5599
rect 9459 5575 9489 5631
rect 9545 5575 9575 5631
rect 9631 5575 9661 5631
rect 9717 5575 9746 5631
rect 9802 5575 10200 5631
rect 6156 5523 10200 5575
rect 10519 5523 10793 5903
rect 13389 5897 13398 5949
rect 13450 5897 13472 5949
rect 13524 5897 13545 5949
rect 13597 5897 13618 5949
rect 13670 5897 13691 5949
rect 13743 5897 13764 5949
rect 13816 5897 13822 5949
rect 13389 5877 13822 5897
rect 13389 5825 13398 5877
rect 13450 5825 13472 5877
rect 13524 5825 13545 5877
rect 13597 5825 13618 5877
rect 13670 5825 13691 5877
rect 13743 5825 13764 5877
rect 13816 5825 13822 5877
rect 13389 5805 13822 5825
rect 13389 5753 13398 5805
rect 13450 5753 13472 5805
rect 13524 5753 13545 5805
rect 13597 5753 13618 5805
rect 13670 5753 13691 5805
rect 13743 5753 13764 5805
rect 13816 5753 13822 5805
rect 13389 5733 13822 5753
rect 13389 5681 13398 5733
rect 13450 5681 13472 5733
rect 13524 5681 13545 5733
rect 13597 5681 13618 5733
rect 13670 5681 13691 5733
rect 13743 5681 13764 5733
rect 13816 5681 13822 5733
rect 13389 5661 13822 5681
rect 13389 5609 13398 5661
rect 13450 5609 13472 5661
rect 13524 5609 13545 5661
rect 13597 5609 13618 5661
rect 13670 5609 13691 5661
rect 13743 5609 13764 5661
rect 13816 5609 13822 5661
rect 13389 5608 13822 5609
rect 6156 5480 6210 5523
rect 4665 5472 4841 5480
tri 4209 5449 4232 5472 ne
rect 4232 5459 4283 5472
tri 4283 5459 4296 5472 sw
tri 4325 5459 4338 5472 ne
rect 4338 5459 4399 5472
rect 4232 5449 4296 5459
rect 4134 5431 4190 5449
tri 4190 5431 4208 5449 sw
tri 4232 5431 4250 5449 ne
rect 4250 5431 4296 5449
tri 4296 5431 4324 5459 sw
tri 4338 5431 4366 5459 ne
rect 4366 5431 4399 5459
tri 4399 5431 4440 5472 sw
tri 4665 5431 4706 5472 ne
rect 4706 5431 4841 5472
tri 4841 5431 4890 5480 sw
tri 4930 5431 4979 5480 ne
rect 4979 5431 5527 5480
tri 4010 5402 4039 5431 ne
rect 4039 5428 4092 5431
tri 4092 5428 4095 5431 sw
tri 4134 5428 4137 5431 ne
rect 4137 5428 4208 5431
tri 4208 5428 4211 5431 sw
tri 4250 5428 4253 5431 ne
rect 4253 5428 4324 5431
tri 4324 5428 4327 5431 sw
tri 4366 5428 4369 5431 ne
rect 4369 5428 4440 5431
tri 4440 5428 4443 5431 sw
tri 4706 5428 4709 5431 ne
rect 4709 5428 4890 5431
rect 4039 5402 4095 5428
tri 4095 5402 4121 5428 sw
tri 4137 5402 4163 5428 ne
rect 4163 5417 4211 5428
tri 4211 5417 4222 5428 sw
tri 4253 5417 4264 5428 ne
rect 4264 5417 4327 5428
tri 4327 5417 4338 5428 sw
tri 4369 5417 4380 5428 ne
rect 4380 5417 4443 5428
rect 4163 5402 4222 5417
tri 1438 5298 1439 5299 ne
rect 1439 5298 1440 5299
tri 1456 5294 1460 5298 ne
rect 1460 5294 1490 5298
tri 1460 5273 1481 5294 ne
rect 1481 5273 1490 5294
tri 1481 5264 1490 5273 ne
rect 1518 5294 1548 5298
tri 1548 5294 1552 5298 nw
rect 3778 5294 3784 5346
rect 3836 5294 3848 5346
rect 3900 5294 3906 5346
tri 4039 5320 4121 5402 ne
tri 4121 5386 4137 5402 sw
tri 4163 5386 4179 5402 ne
rect 4179 5386 4222 5402
rect 4121 5354 4137 5386
tri 4137 5354 4169 5386 sw
tri 4179 5354 4211 5386 ne
rect 4211 5375 4222 5386
tri 4222 5375 4264 5417 sw
tri 4264 5398 4283 5417 ne
rect 4283 5398 4338 5417
tri 4338 5398 4357 5417 sw
tri 4380 5398 4399 5417 ne
rect 4399 5398 4443 5417
tri 4443 5398 4473 5428 sw
tri 4709 5398 4739 5428 ne
rect 4739 5398 4890 5428
tri 4283 5375 4306 5398 ne
rect 4306 5385 4357 5398
tri 4357 5385 4370 5398 sw
tri 4399 5385 4412 5398 ne
rect 4412 5385 4473 5398
rect 4306 5375 4370 5385
rect 4211 5354 4264 5375
tri 4264 5354 4285 5375 sw
tri 4306 5354 4327 5375 ne
rect 4327 5354 4370 5375
tri 4370 5354 4401 5385 sw
tri 4412 5354 4443 5385 ne
rect 4443 5354 4473 5385
tri 4473 5354 4517 5398 sw
tri 4739 5354 4783 5398 ne
rect 4783 5354 4890 5398
rect 4121 5320 4169 5354
tri 4169 5320 4203 5354 sw
tri 4211 5320 4245 5354 ne
rect 4245 5343 4285 5354
tri 4285 5343 4296 5354 sw
tri 4327 5343 4338 5354 ne
rect 4338 5343 4401 5354
tri 4401 5343 4412 5354 sw
tri 4443 5343 4454 5354 ne
rect 4454 5343 4517 5354
rect 4245 5320 4296 5343
tri 4121 5294 4147 5320 ne
rect 4147 5312 4203 5320
tri 4203 5312 4211 5320 sw
tri 4245 5312 4253 5320 ne
rect 4253 5312 4296 5320
rect 4147 5294 4211 5312
tri 4211 5294 4229 5312 sw
tri 4253 5294 4271 5312 ne
rect 4271 5301 4296 5312
tri 4296 5301 4338 5343 sw
tri 4338 5324 4357 5343 ne
rect 4357 5324 4412 5343
tri 4412 5324 4431 5343 sw
tri 4454 5324 4473 5343 ne
rect 4473 5324 4517 5343
tri 4517 5324 4547 5354 sw
tri 4783 5324 4813 5354 ne
rect 4813 5350 4890 5354
tri 4890 5350 4971 5431 sw
tri 4979 5350 5060 5431 ne
rect 5060 5350 5527 5431
tri 5527 5350 5657 5480 nw
tri 6026 5469 6037 5480 se
rect 6037 5469 6210 5480
tri 6210 5469 6264 5523 nw
tri 5907 5350 6026 5469 se
rect 4813 5324 4971 5350
tri 4357 5301 4380 5324 ne
rect 4380 5311 4431 5324
tri 4431 5311 4444 5324 sw
tri 4473 5311 4486 5324 ne
rect 4486 5311 4547 5324
rect 4380 5301 4444 5311
rect 4271 5294 4338 5301
tri 4338 5294 4345 5301 sw
tri 4380 5294 4387 5301 ne
rect 4387 5294 4444 5301
tri 4444 5294 4461 5311 sw
tri 4486 5294 4503 5311 ne
rect 4503 5294 4547 5311
tri 4547 5294 4577 5324 sw
tri 4813 5294 4843 5324 ne
rect 4843 5294 4971 5324
tri 4971 5294 5027 5350 sw
tri 5851 5294 5907 5350 se
rect 5907 5294 6026 5350
rect 1518 5273 1527 5294
tri 1527 5273 1548 5294 nw
tri 4147 5273 4168 5294 ne
rect 4168 5280 4229 5294
tri 4229 5280 4243 5294 sw
tri 4271 5280 4285 5294 ne
rect 4285 5280 4345 5294
tri 4345 5280 4359 5294 sw
tri 4387 5280 4401 5294 ne
rect 4401 5280 4461 5294
tri 4461 5280 4475 5294 sw
tri 4503 5280 4517 5294 ne
rect 4517 5280 4577 5294
tri 4577 5280 4591 5294 sw
tri 4843 5280 4857 5294 ne
rect 4857 5285 5027 5294
tri 5027 5285 5036 5294 sw
tri 5842 5285 5851 5294 se
rect 5851 5285 6026 5294
tri 6026 5285 6210 5469 nw
rect 7812 5411 11206 5412
rect 7812 5355 7856 5411
rect 7912 5355 7937 5411
rect 7993 5355 8018 5411
rect 8074 5355 8099 5411
rect 8155 5355 8180 5411
rect 8236 5355 8261 5411
rect 8317 5355 8341 5411
rect 8397 5355 8421 5411
rect 8477 5355 8501 5411
rect 8557 5355 8581 5411
rect 8637 5355 8661 5411
rect 8717 5355 8741 5411
rect 8797 5355 8821 5411
rect 8877 5355 8901 5411
rect 8957 5355 8981 5411
rect 9037 5355 9061 5411
rect 9117 5355 9141 5411
rect 9197 5355 9221 5411
rect 9277 5355 9301 5411
rect 9357 5355 9381 5411
rect 9437 5355 9461 5411
rect 9517 5355 9541 5411
rect 9597 5355 9621 5411
rect 9677 5355 9701 5411
rect 9757 5355 9781 5411
rect 9837 5355 9861 5411
rect 9917 5355 9941 5411
rect 9997 5355 10021 5411
rect 10077 5355 10101 5411
rect 10157 5355 10181 5411
rect 10237 5355 10261 5411
rect 10317 5355 10341 5411
rect 10397 5355 10421 5411
rect 10477 5355 10501 5411
rect 10557 5355 10581 5411
rect 10637 5355 10661 5411
rect 10717 5355 10741 5411
rect 10797 5355 10821 5411
rect 10877 5355 10901 5411
rect 10957 5355 10981 5411
rect 11037 5355 11061 5411
rect 11117 5355 11141 5411
rect 11197 5355 11206 5411
rect 7812 5317 11206 5355
rect 4857 5280 5036 5285
rect 4168 5273 4243 5280
tri 4243 5273 4250 5280 sw
tri 4285 5273 4292 5280 ne
rect 4292 5273 4359 5280
tri 4359 5273 4366 5280 sw
tri 4401 5273 4408 5280 ne
rect 4408 5273 4475 5280
tri 4475 5273 4482 5280 sw
tri 4517 5273 4524 5280 ne
rect 4524 5273 4591 5280
tri 4591 5273 4598 5280 sw
tri 4857 5273 4864 5280 ne
rect 4864 5273 5036 5280
tri 5036 5273 5048 5285 sw
tri 5830 5273 5842 5285 se
rect 5842 5273 6014 5285
tri 6014 5273 6026 5285 nw
tri 1518 5264 1527 5273 nw
tri 4168 5264 4177 5273 ne
rect 4177 5264 4250 5273
tri 4177 5255 4186 5264 ne
rect 4186 5255 4250 5264
tri 3929 5252 3932 5255 se
tri 4186 5252 4189 5255 ne
rect 4189 5252 4250 5255
tri 4189 5247 4194 5252 ne
rect 4194 5247 4250 5252
tri 4250 5247 4276 5273 sw
tri 4292 5247 4318 5273 ne
rect 4318 5269 4366 5273
tri 4366 5269 4370 5273 sw
tri 4408 5269 4412 5273 ne
rect 4412 5269 4482 5273
tri 4482 5269 4486 5273 sw
tri 4524 5269 4528 5273 ne
rect 4528 5269 4598 5273
rect 4318 5247 4370 5269
tri 4370 5247 4392 5269 sw
tri 4412 5250 4431 5269 ne
rect 4431 5250 4486 5269
tri 4486 5250 4505 5269 sw
tri 4528 5250 4547 5269 ne
rect 4547 5250 4598 5269
tri 4598 5250 4621 5273 sw
tri 4864 5250 4887 5273 ne
rect 4887 5250 5048 5273
tri 4431 5247 4434 5250 ne
rect 4434 5247 4505 5250
tri 4505 5247 4508 5250 sw
tri 4547 5247 4550 5250 ne
rect 4550 5247 4621 5250
tri 4621 5247 4624 5250 sw
tri 4887 5247 4890 5250 ne
rect 4890 5247 5048 5250
tri 5048 5247 5074 5273 sw
tri 5804 5247 5830 5273 se
rect 5830 5247 5988 5273
tri 5988 5247 6014 5273 nw
rect 7812 5261 7856 5317
rect 7912 5261 7937 5317
rect 7993 5261 8018 5317
rect 8074 5261 8099 5317
rect 8155 5261 8180 5317
rect 8236 5261 8261 5317
rect 8317 5261 8341 5317
rect 8397 5261 8421 5317
rect 8477 5261 8501 5317
rect 8557 5261 8581 5317
rect 8637 5261 8661 5317
rect 8717 5261 8741 5317
rect 8797 5261 8821 5317
rect 8877 5261 8901 5317
rect 8957 5261 8981 5317
rect 9037 5261 9061 5317
rect 9117 5261 9141 5317
rect 9197 5261 9221 5317
rect 9277 5261 9301 5317
rect 9357 5261 9381 5317
rect 9437 5261 9461 5317
rect 9517 5261 9541 5317
rect 9597 5261 9621 5317
rect 9677 5261 9701 5317
rect 9757 5261 9781 5317
rect 9837 5261 9861 5317
rect 9917 5261 9941 5317
rect 9997 5261 10021 5317
rect 10077 5261 10101 5317
rect 10157 5261 10181 5317
rect 10237 5261 10261 5317
rect 10317 5261 10341 5317
rect 10397 5261 10421 5317
rect 10477 5261 10501 5317
rect 10557 5261 10581 5317
rect 10637 5261 10661 5317
rect 10717 5261 10741 5317
rect 10797 5261 10821 5317
rect 10877 5261 10901 5317
rect 10957 5261 10981 5317
rect 11037 5261 11061 5317
rect 11117 5261 11141 5317
rect 11197 5261 11206 5317
tri 4194 5238 4203 5247 ne
rect 4203 5238 4276 5247
tri 4276 5238 4285 5247 sw
tri 4318 5238 4327 5247 ne
rect 4327 5238 4392 5247
tri 4203 5221 4220 5238 ne
rect 4220 5221 4285 5238
tri 4285 5221 4302 5238 sw
tri 4327 5221 4344 5238 ne
rect 4344 5227 4392 5238
tri 4392 5227 4412 5247 sw
tri 4434 5227 4454 5247 ne
rect 4454 5237 4508 5247
tri 4508 5237 4518 5247 sw
tri 4550 5237 4560 5247 ne
rect 4560 5237 4624 5247
rect 4454 5227 4518 5237
rect 4344 5221 4412 5227
tri 4412 5221 4418 5227 sw
tri 4454 5221 4460 5227 ne
rect 4460 5221 4518 5227
tri 4518 5221 4534 5237 sw
tri 4560 5221 4576 5237 ne
rect 4576 5221 4624 5237
tri 4624 5221 4650 5247 sw
tri 4890 5221 4916 5247 ne
rect 4916 5221 5962 5247
tri 5962 5221 5988 5247 nw
rect 7812 5223 11206 5261
tri 4220 5206 4235 5221 ne
rect 4235 5206 4302 5221
tri 4302 5206 4317 5221 sw
tri 4344 5206 4359 5221 ne
rect 4359 5206 4418 5221
tri 4418 5206 4433 5221 sw
tri 4460 5206 4475 5221 ne
rect 4475 5206 4534 5221
tri 4534 5206 4549 5221 sw
tri 4576 5206 4591 5221 ne
rect 4591 5206 4650 5221
tri 4650 5206 4665 5221 sw
tri 4916 5206 4931 5221 ne
rect 4931 5206 5947 5221
tri 5947 5206 5962 5221 nw
tri 4235 5200 4241 5206 ne
rect 4241 5200 4317 5206
tri 3907 5199 3908 5200 ne
rect 3908 5199 3932 5200
tri -744 5165 -710 5199 nw
tri 3908 5175 3932 5199 ne
tri 4241 5175 4266 5200 ne
rect 4266 5175 4317 5200
tri 4266 5165 4276 5175 ne
rect 4276 5165 4317 5175
tri 4276 5157 4284 5165 ne
rect 4284 5164 4317 5165
tri 4317 5164 4359 5206 sw
tri 4359 5164 4401 5206 ne
rect 4401 5195 4433 5206
tri 4433 5195 4444 5206 sw
tri 4475 5195 4486 5206 ne
rect 4486 5195 4549 5206
tri 4549 5195 4560 5206 sw
tri 4591 5195 4602 5206 ne
rect 4602 5195 4665 5206
rect 4401 5176 4444 5195
tri 4444 5176 4463 5195 sw
tri 4486 5176 4505 5195 ne
rect 4505 5176 4560 5195
tri 4560 5176 4579 5195 sw
tri 4602 5176 4621 5195 ne
rect 4621 5176 4665 5195
tri 4665 5176 4695 5206 sw
tri 4931 5176 4961 5206 ne
rect 4961 5176 5895 5206
rect 4401 5164 4463 5176
rect 4284 5157 4359 5164
tri 4359 5157 4366 5164 sw
tri 4401 5157 4408 5164 ne
rect 4408 5157 4463 5164
tri 3043 5156 3044 5157 sw
tri 4284 5156 4285 5157 ne
rect 4285 5156 4366 5157
tri 4366 5156 4367 5157 sw
tri 4408 5156 4409 5157 ne
rect 4409 5156 4463 5157
tri 4285 5154 4287 5156 ne
rect 4287 5154 4367 5156
tri 4367 5154 4369 5156 sw
tri 4409 5154 4411 5156 ne
rect 4411 5154 4463 5156
tri 4463 5154 4485 5176 sw
tri 4505 5154 4527 5176 ne
rect 4527 5169 4579 5176
tri 4579 5169 4586 5176 sw
tri 4621 5169 4628 5176 ne
rect 4628 5169 4695 5176
rect 4527 5154 4586 5169
tri 4586 5154 4601 5169 sw
tri 4628 5154 4643 5169 ne
rect 4643 5154 4695 5169
tri 4695 5154 4717 5176 sw
tri 4961 5154 4983 5176 ne
rect 4983 5154 5895 5176
tri 5895 5154 5947 5206 nw
rect 7812 5167 7856 5223
rect 7912 5167 7937 5223
rect 7993 5167 8018 5223
rect 8074 5167 8099 5223
rect 8155 5167 8180 5223
rect 8236 5167 8261 5223
rect 8317 5167 8341 5223
rect 8397 5167 8421 5223
rect 8477 5167 8501 5223
rect 8557 5167 8581 5223
rect 8637 5167 8661 5223
rect 8717 5167 8741 5223
rect 8797 5167 8821 5223
rect 8877 5167 8901 5223
rect 8957 5167 8981 5223
rect 9037 5167 9061 5223
rect 9117 5167 9141 5223
rect 9197 5167 9221 5223
rect 9277 5167 9301 5223
rect 9357 5167 9381 5223
rect 9437 5167 9461 5223
rect 9517 5167 9541 5223
rect 9597 5167 9621 5223
rect 9677 5167 9701 5223
rect 9757 5167 9781 5223
rect 9837 5167 9861 5223
rect 9917 5167 9941 5223
rect 9997 5167 10021 5223
rect 10077 5167 10101 5223
rect 10157 5167 10181 5223
rect 10237 5167 10261 5223
rect 10317 5167 10341 5223
rect 10397 5167 10421 5223
rect 10477 5167 10501 5223
rect 10557 5167 10581 5223
rect 10637 5167 10661 5223
rect 10717 5167 10741 5223
rect 10797 5167 10821 5223
rect 10877 5167 10901 5223
rect 10957 5167 10981 5223
rect 11037 5167 11061 5223
rect 11117 5167 11141 5223
rect 11197 5167 11206 5223
tri 4287 5145 4296 5154 ne
rect 4296 5145 4369 5154
tri 1207 5139 1213 5145 ne
rect 1213 5139 1221 5145
tri 1213 5135 1217 5139 ne
rect 1217 5135 1221 5139
rect 1249 5139 1253 5145
tri 1253 5139 1259 5145 nw
tri 4296 5139 4302 5145 ne
rect 4302 5139 4369 5145
tri 4369 5139 4384 5154 sw
tri 4411 5139 4426 5154 ne
rect 4426 5153 4485 5154
tri 4485 5153 4486 5154 sw
tri 4527 5153 4528 5154 ne
rect 4528 5153 4601 5154
rect 4426 5139 4486 5153
tri 4486 5139 4500 5153 sw
tri 4528 5139 4542 5153 ne
rect 4542 5139 4601 5153
tri 4601 5139 4616 5154 sw
tri 4643 5139 4658 5154 ne
rect 4658 5139 4717 5154
tri 4717 5139 4732 5154 sw
tri 4983 5139 4998 5154 ne
rect 4998 5139 5880 5154
tri 5880 5139 5895 5154 nw
rect 7812 5145 11206 5167
tri 1249 5135 1253 5139 nw
tri 4302 5135 4306 5139 ne
rect 4306 5135 4384 5139
tri 1217 5131 1221 5135 ne
tri 4306 5131 4310 5135 ne
rect 4310 5132 4384 5135
tri 4384 5132 4391 5139 sw
tri 4426 5132 4433 5139 ne
rect 4433 5132 4500 5139
tri 4500 5132 4507 5139 sw
tri 4542 5132 4549 5139 ne
rect 4549 5132 4616 5139
tri 4616 5132 4623 5139 sw
tri 4658 5132 4665 5139 ne
rect 4665 5132 4732 5139
tri 4732 5132 4739 5139 sw
tri 4998 5132 5005 5139 ne
rect 5005 5132 5858 5139
rect 4310 5131 4391 5132
tri 4310 5121 4320 5131 ne
rect 4320 5121 4391 5131
tri 1407 5118 1410 5121 ne
rect 1433 5117 1455 5121
tri 1455 5117 1459 5121 nw
tri 4320 5117 4324 5121 ne
rect 4324 5117 4391 5121
tri 4391 5117 4406 5132 sw
tri 4433 5117 4448 5132 ne
rect 4448 5131 4507 5132
tri 4507 5131 4508 5132 sw
rect 4448 5117 4508 5131
tri 4549 5121 4560 5132 ne
rect 4560 5127 4623 5132
tri 4623 5127 4628 5132 sw
tri 4665 5127 4670 5132 ne
rect 4670 5127 4739 5132
rect 4560 5121 4628 5127
tri 4628 5121 4634 5127 sw
tri 4670 5121 4676 5127 ne
rect 4676 5121 4739 5127
rect 1433 5114 1452 5117
tri 1452 5114 1455 5117 nw
tri 4324 5114 4327 5117 ne
rect 4327 5114 4406 5117
tri 1433 5095 1452 5114 nw
tri 1740 5095 1759 5114 se
rect 1759 5095 2160 5114
tri 1707 5062 1740 5095 se
rect 1740 5062 2160 5095
rect 2212 5062 2224 5114
rect 2276 5062 2282 5114
tri 4327 5105 4336 5114 ne
rect 4336 5105 4406 5114
tri 3818 5095 3828 5105 ne
rect 3828 5095 3852 5105
tri 3828 5087 3836 5095 ne
rect 3836 5087 3852 5095
tri 4336 5087 4354 5105 ne
rect 4354 5099 4406 5105
tri 4406 5099 4424 5117 sw
tri 4448 5102 4463 5117 ne
rect 4354 5087 4424 5099
tri 3836 5075 3848 5087 ne
rect 3848 5075 3852 5087
tri 4354 5075 4366 5087 ne
tri 3848 5072 3851 5075 ne
rect 3851 5072 3852 5075
tri 3851 5071 3852 5072 ne
tri 1692 5047 1707 5062 se
rect 1707 5047 1766 5062
tri 1766 5047 1781 5062 nw
tri 1685 5040 1692 5047 se
rect 1692 5040 1759 5047
tri 1759 5040 1766 5047 nw
tri 1651 5006 1685 5040 se
rect 1685 5006 1725 5040
tri 1725 5006 1759 5040 nw
rect 1651 4995 1714 5006
tri 1714 4995 1725 5006 nw
tri -227 4654 -225 4656 se
tri -458 4629 -455 4632 ne
rect -455 4629 -438 4632
tri -455 4612 -438 4629 ne
rect -412 4629 -409 4632
tri -409 4629 -406 4632 nw
tri -412 4626 -409 4629 nw
rect -334 4626 -309 4629
tri -309 4626 -306 4629 nw
rect -334 4612 -323 4626
tri -323 4612 -309 4626 nw
tri -334 4601 -323 4612 nw
tri -660 4417 -631 4446 nw
tri 346 3896 362 3912 se
tri 328 3878 346 3896 se
rect 346 3878 362 3896
tri 272 3806 292 3826 ne
rect 292 3806 304 3826
tri 292 3799 299 3806 ne
rect 299 3799 304 3806
tri 299 3794 304 3799 ne
rect 356 3806 370 3826
tri 370 3806 390 3826 nw
rect 356 3799 363 3806
tri 363 3799 370 3806 nw
rect 356 3794 358 3799
tri 358 3794 363 3799 nw
tri 356 3792 358 3794 nw
rect 1651 3728 1703 4995
tri 1703 4984 1714 4995 nw
rect 1953 4841 1959 4893
rect 2011 4841 2023 4893
rect 2075 4841 2081 4893
tri 4095 4850 4100 4855 se
tri 1953 4838 1956 4841 ne
rect 1956 4838 2078 4841
tri 2078 4838 2081 4841 nw
tri 4083 4838 4095 4850 se
rect 4095 4838 4100 4850
tri 1956 4829 1965 4838 ne
rect 1965 4829 2069 4838
tri 2069 4829 2078 4838 nw
tri 1965 4821 1973 4829 ne
rect 1973 4821 2061 4829
tri 2061 4821 2069 4829 nw
rect 1973 4786 2026 4821
tri 2026 4786 2061 4821 nw
tri 1703 3728 1705 3730 sw
rect 1651 3713 1705 3728
tri 1705 3713 1720 3728 sw
rect 1651 3709 1720 3713
tri 1720 3709 1724 3713 sw
rect 1651 3708 1724 3709
tri 1724 3708 1725 3709 sw
tri 1651 3678 1681 3708 ne
rect 1681 3678 1725 3708
tri 1725 3678 1755 3708 sw
tri 1681 3673 1686 3678 ne
rect 1686 3673 1755 3678
tri 1755 3673 1760 3678 sw
tri 1686 3634 1725 3673 ne
rect 1725 3634 1760 3673
tri 1760 3634 1799 3673 sw
tri 1725 3621 1738 3634 ne
rect 1738 3621 1799 3634
tri 1799 3621 1812 3634 sw
tri 1738 3609 1750 3621 ne
rect 1750 3609 1812 3621
tri 1812 3609 1824 3621 sw
tri 1750 3560 1799 3609 ne
rect 1799 3576 1824 3609
tri 1824 3576 1857 3609 sw
rect 1799 3560 1857 3576
tri 1857 3560 1873 3576 sw
tri 1799 3557 1802 3560 ne
rect 1802 3557 1873 3560
tri 1873 3557 1876 3560 sw
tri 1802 3554 1805 3557 ne
rect 1805 3554 1876 3557
tri 1876 3554 1879 3557 sw
tri 1805 3552 1807 3554 ne
rect 1807 3552 1879 3554
tri 1879 3552 1881 3554 sw
tri 1807 3514 1845 3552 ne
rect 1845 3524 1881 3552
tri 1881 3524 1909 3552 sw
rect 1845 3514 1909 3524
tri 1845 3502 1857 3514 ne
tri 1466 3339 1490 3363 se
rect 1857 3295 1909 3514
rect 1973 3266 2025 4786
tri 2025 4785 2026 4786 nw
tri 4074 4785 4075 4786 ne
rect 4075 4785 4100 4786
tri 4075 4777 4083 4785 ne
rect 4083 4777 4100 4785
tri 4083 4760 4100 4777 ne
tri 3977 4704 3978 4705 ne
rect 3978 4704 4011 4705
tri 3978 4683 3999 4704 ne
rect 3999 4683 4011 4704
tri 3999 4674 4008 4683 ne
rect 4008 4674 4011 4683
tri 2649 4640 2683 4674 ne
tri 4008 4671 4011 4674 ne
rect 2908 4639 3054 4645
rect 2960 4635 3002 4639
rect 2908 4579 2913 4587
rect 2969 4579 2993 4635
rect 3049 4579 3054 4587
rect 2908 4573 3054 4579
rect 2960 4554 3002 4573
rect 2908 4506 2913 4521
rect 2969 4498 2993 4554
rect 3049 4506 3054 4521
rect 2960 4454 3002 4498
rect 4281 4611 4334 4617
rect 4333 4559 4334 4611
rect 4281 4547 4334 4559
rect 4333 4495 4334 4547
rect 4281 4489 4334 4495
tri 4281 4485 4285 4489 ne
rect 4285 4485 4334 4489
tri 4285 4468 4302 4485 ne
rect 2908 4448 3054 4454
tri 4152 4217 4157 4222 se
tri 4131 4196 4152 4217 se
rect 4152 4196 4157 4217
tri 4123 4188 4131 4196 se
rect 4131 4188 4157 4196
tri 2812 4077 2844 4109 sw
tri 4125 4077 4157 4109 se
rect 2812 4075 2844 4077
tri 2844 4075 2846 4077 sw
tri 4123 4075 4125 4077 se
rect 4125 4075 4157 4077
tri 4128 4013 4138 4023 ne
rect 4138 4013 4157 4023
tri 4138 3994 4157 4013 ne
rect 4302 3975 4334 4485
rect 4366 4410 4424 5087
rect 4366 4358 4369 4410
rect 4421 4358 4424 4410
rect 4366 4346 4424 4358
rect 4366 4294 4369 4346
rect 4421 4294 4424 4346
rect 4366 4288 4424 4294
tri 4334 3975 4341 3982 sw
rect 4302 3951 4341 3975
tri 4341 3951 4365 3975 sw
tri 2682 3948 2683 3949 se
tri 2649 3915 2682 3948 se
rect 2682 3915 2683 3948
tri 2711 3948 2712 3949 sw
rect 4302 3948 4365 3951
tri 4365 3948 4368 3951 sw
rect 2711 3915 2712 3948
tri 2712 3915 2745 3948 sw
tri 4142 3896 4157 3911 se
rect 4302 3896 4308 3948
rect 4360 3896 4372 3948
rect 4424 3896 4430 3948
tri 4123 3877 4142 3896 se
rect 4142 3877 4157 3896
tri 4451 3877 4463 3889 se
rect 4463 3877 4508 5117
tri 4560 5102 4579 5121 ne
rect 4579 5117 4634 5121
tri 4634 5117 4638 5121 sw
tri 4676 5117 4680 5121 ne
rect 4680 5117 4739 5121
tri 4739 5117 4754 5132 sw
tri 5005 5117 5020 5132 ne
rect 5020 5117 5858 5132
tri 5858 5117 5880 5139 nw
rect 7847 5129 11206 5145
rect 4579 5102 4638 5117
tri 4638 5102 4653 5117 sw
tri 4680 5102 4695 5117 ne
rect 4695 5102 4754 5117
tri 4754 5102 4769 5117 sw
tri 4579 5087 4594 5102 ne
rect 4594 5087 4653 5102
tri 4653 5087 4668 5102 sw
tri 4695 5087 4710 5102 ne
rect 4710 5087 4769 5102
tri 4594 5080 4601 5087 ne
rect 4601 5080 4668 5087
tri 4668 5080 4675 5087 sw
tri 4710 5080 4717 5087 ne
tri 4601 5072 4609 5080 ne
rect 4609 5075 4675 5080
tri 4675 5075 4680 5080 sw
rect 4609 5072 4680 5075
tri 4609 5053 4628 5072 ne
tri 4444 3870 4451 3877 se
rect 4451 3870 4508 3877
tri 4438 3864 4444 3870 se
rect 4444 3864 4508 3870
tri 4140 3836 4157 3853 ne
rect 4157 3836 4160 3853
rect 4264 3815 4508 3864
rect 4537 4410 4589 4416
rect 4537 4346 4589 4358
rect 4264 3806 4341 3815
tri 4341 3806 4350 3815 nw
rect 4264 3799 4334 3806
tri 4334 3799 4341 3806 nw
rect 4264 3795 4330 3799
tri 4330 3795 4334 3799 nw
tri 4172 3728 4176 3732 se
tri 4163 3719 4172 3728 se
rect 4172 3719 4176 3728
tri 4142 3678 4155 3691 ne
rect 4155 3678 4176 3691
tri 4155 3673 4160 3678 ne
rect 4160 3673 4176 3678
tri 4160 3657 4176 3673 ne
tri 2170 3621 2190 3641 se
rect 2190 3621 3939 3641
tri 3939 3621 3959 3641 sw
tri 2158 3609 2170 3621 se
rect 2170 3611 3959 3621
tri 3959 3611 3969 3621 sw
rect 2170 3609 3969 3611
tri 3969 3609 3971 3611 sw
tri 2116 3567 2158 3609 se
rect 2158 3589 3971 3609
tri 3971 3589 3991 3609 sw
rect 2158 3567 2190 3589
tri 2190 3567 2212 3589 nw
tri 3917 3567 3939 3589 ne
rect 3939 3583 3991 3589
tri 3991 3583 3997 3589 sw
rect 3939 3580 3997 3583
tri 3997 3580 4000 3583 sw
rect 3939 3571 4000 3580
tri 4000 3571 4009 3580 sw
tri 4255 3571 4264 3580 se
rect 4264 3571 4316 3795
tri 4316 3781 4330 3795 nw
tri 4395 3571 4407 3583 ne
rect 4434 3571 4435 3583
tri 4435 3571 4447 3583 nw
tri 4526 3571 4537 3582 se
rect 4537 3571 4589 4294
rect 3939 3570 4009 3571
tri 4009 3570 4010 3571 sw
tri 4254 3570 4255 3571 se
rect 4255 3570 4316 3571
tri 4434 3570 4435 3571 nw
tri 4525 3570 4526 3571 se
rect 4526 3570 4589 3571
rect 3939 3567 4010 3570
tri 4010 3567 4013 3570 sw
tri 4251 3567 4254 3570 se
rect 4254 3567 4316 3570
tri 4522 3567 4525 3570 se
rect 4525 3567 4589 3570
tri 2106 3557 2116 3567 se
rect 2116 3557 2180 3567
tri 2180 3557 2190 3567 nw
tri 3939 3557 3949 3567 ne
rect 3949 3557 4013 3567
tri 4013 3557 4023 3567 sw
tri 4241 3557 4251 3567 se
rect 4251 3557 4316 3567
tri 4512 3557 4522 3567 se
rect 4522 3560 4589 3567
rect 4522 3557 4586 3560
tri 4586 3557 4589 3560 nw
tri 2103 3554 2106 3557 se
rect 2106 3554 2177 3557
tri 2177 3554 2180 3557 nw
tri 3949 3554 3952 3557 ne
rect 3952 3554 4023 3557
tri 4023 3554 4026 3557 sw
tri 4238 3554 4241 3557 se
rect 4241 3554 4316 3557
tri 4509 3554 4512 3557 se
rect 4512 3554 4583 3557
tri 4583 3554 4586 3557 nw
tri 2101 3552 2103 3554 se
rect 2103 3552 2175 3554
tri 2175 3552 2177 3554 nw
tri 3952 3552 3954 3554 ne
rect 3954 3552 4026 3554
tri 4026 3552 4028 3554 sw
tri 4236 3552 4238 3554 se
rect 4238 3552 4316 3554
tri 4507 3552 4509 3554 se
rect 4509 3552 4581 3554
tri 4581 3552 4583 3554 nw
tri 2092 3543 2101 3552 se
rect 2101 3543 2166 3552
tri 2166 3543 2175 3552 nw
tri 3954 3543 3963 3552 ne
rect 3963 3543 4028 3552
tri 4028 3543 4037 3552 sw
tri 4227 3543 4236 3552 se
rect 4236 3543 4316 3552
tri 4498 3543 4507 3552 se
rect 4507 3543 4556 3552
rect 1857 3231 1909 3243
rect 1857 3173 1909 3179
tri 356 3020 359 3023 sw
tri 273 2989 304 3020 se
rect 356 2989 359 3020
tri 359 2989 390 3020 sw
tri -655 2986 -652 2989 sw
rect -655 2955 -652 2986
tri -652 2955 -621 2986 sw
rect -655 2889 -635 2903
tri -635 2889 -621 2903 nw
rect -655 2877 -647 2889
tri -647 2877 -635 2889 nw
tri -655 2869 -647 2877 nw
tri 2078 2671 2092 2685 se
rect 2092 2671 2144 3543
tri 2144 3521 2166 3543 nw
tri 3963 3537 3969 3543 ne
rect 3969 3537 4037 3543
tri 4037 3537 4043 3543 sw
tri 4221 3537 4227 3543 se
rect 4227 3537 4316 3543
tri 3969 3536 3970 3537 ne
rect 3970 3536 4316 3537
tri 2267 3521 2282 3536 se
rect 2282 3521 3861 3536
tri 3861 3521 3876 3536 sw
tri 3970 3521 3985 3536 ne
rect 3985 3521 4316 3536
tri 2260 3514 2267 3521 se
rect 2267 3514 3876 3521
tri 3876 3514 3883 3521 sw
tri 3985 3514 3992 3521 ne
rect 3992 3515 4316 3521
rect 3992 3514 4315 3515
tri 4315 3514 4316 3515 nw
tri 4482 3527 4498 3543 se
rect 4498 3527 4556 3543
tri 4556 3527 4581 3552 nw
rect 4482 3521 4550 3527
tri 4550 3521 4556 3527 nw
rect 4482 3514 4543 3521
tri 4543 3514 4550 3521 nw
tri 2241 3495 2260 3514 se
rect 2260 3495 3883 3514
tri 3883 3495 3902 3514 sw
tri 3992 3495 4011 3514 ne
rect 4011 3495 4288 3514
tri 2233 3487 2241 3495 se
rect 2241 3487 3902 3495
tri 3902 3487 3910 3495 sw
tri 4011 3487 4019 3495 ne
rect 4019 3487 4288 3495
tri 4288 3487 4315 3514 nw
tri 2208 3462 2233 3487 se
rect 2233 3485 3910 3487
tri 3910 3485 3912 3487 sw
tri 4019 3485 4021 3487 ne
rect 4021 3485 4286 3487
tri 4286 3485 4288 3487 nw
rect 2233 3484 3912 3485
rect 2233 3462 2282 3484
tri 2282 3462 2304 3484 nw
tri 3839 3462 3861 3484 ne
rect 3861 3462 3912 3484
tri 2191 3445 2208 3462 se
rect 2208 3445 2265 3462
tri 2265 3445 2282 3462 nw
tri 3861 3445 3878 3462 ne
rect 3878 3446 3912 3462
tri 3912 3446 3951 3485 sw
rect 3878 3445 3951 3446
rect 2191 3440 2260 3445
tri 2260 3440 2265 3445 nw
tri 3878 3440 3883 3445 ne
rect 3883 3440 3951 3445
tri 3951 3440 3957 3446 sw
tri 4170 3440 4176 3446 se
rect 4176 3440 4228 3446
rect 2191 3295 2243 3440
tri 2243 3423 2260 3440 nw
tri 3883 3423 3900 3440 ne
rect 3900 3423 3957 3440
tri 3900 3421 3902 3423 ne
rect 3902 3421 3957 3423
tri 3957 3421 3976 3440 sw
tri 4151 3421 4170 3440 se
rect 4170 3421 4176 3440
tri 3902 3412 3911 3421 ne
rect 3911 3412 4176 3421
tri 3911 3388 3935 3412 ne
rect 3935 3388 4176 3412
tri 3935 3376 3947 3388 ne
rect 3947 3376 4228 3388
tri 3947 3372 3951 3376 ne
rect 3951 3372 4176 3376
tri 3951 3369 3954 3372 ne
rect 3954 3369 4176 3372
tri 4125 3324 4170 3369 ne
rect 4170 3324 4176 3369
tri 4170 3318 4176 3324 ne
rect 4176 3318 4228 3324
rect 2191 3231 2243 3243
rect 2191 3173 2243 3179
tri 3493 3115 3506 3128 sw
tri 4163 3115 4176 3128 se
rect 3493 3094 3506 3115
tri 3506 3094 3527 3115 sw
tri 4142 3094 4163 3115 se
rect 4163 3094 4176 3115
tri 4134 3025 4151 3042 ne
rect 4151 3025 4176 3042
tri 4151 3000 4176 3025 ne
tri 4170 2941 4176 2947 se
tri 3431 2914 3458 2941 sw
tri 4143 2914 4170 2941 se
rect 4170 2914 4176 2941
tri 3186 2894 3190 2898 se
tri 3234 2894 3238 2898 sw
rect 3431 2848 3451 2862
tri 3451 2848 3465 2862 nw
tri 4133 2848 4147 2862 ne
rect 4147 2848 4176 2862
tri 3287 2842 3293 2848 ne
rect 3293 2842 3306 2848
tri 3333 2842 3339 2848 nw
rect 3431 2842 3445 2848
tri 3445 2842 3451 2848 nw
tri 4147 2842 4153 2848 ne
rect 4153 2842 4176 2848
tri 3293 2829 3306 2842 ne
rect 3431 2829 3432 2842
tri 3432 2829 3445 2842 nw
tri 4153 2829 4166 2842 ne
rect 4166 2829 4176 2842
tri 3431 2828 3432 2829 nw
tri 4166 2828 4167 2829 ne
rect 4167 2828 4176 2829
tri 4167 2825 4170 2828 ne
rect 4170 2825 4176 2828
tri 4170 2819 4176 2825 ne
rect 1627 2631 1679 2671
tri 2051 2644 2078 2671 se
rect 2078 2663 2144 2671
rect 2078 2644 2125 2663
tri 2125 2644 2144 2663 nw
tri 2047 2640 2051 2644 se
rect 2051 2640 2112 2644
tri 1679 2631 1688 2640 sw
tri 2038 2631 2047 2640 se
rect 2047 2631 2112 2640
tri 2112 2631 2125 2644 nw
rect 1627 2618 1688 2631
tri 1627 2600 1645 2618 ne
rect 1645 2611 1688 2618
tri 1688 2611 1708 2631 sw
tri 2018 2611 2038 2631 se
rect 2038 2611 2092 2631
tri 2092 2611 2112 2631 nw
rect 1645 2600 1708 2611
tri 1708 2600 1719 2611 sw
tri 2007 2600 2018 2611 se
rect 2018 2600 2081 2611
tri 2081 2600 2092 2611 nw
tri 1645 2579 1666 2600 ne
rect 1666 2579 2060 2600
tri 2060 2579 2081 2600 nw
tri 1666 2570 1675 2579 ne
rect 1675 2570 2051 2579
tri 2051 2570 2060 2579 nw
tri 1675 2566 1679 2570 ne
rect 1679 2566 2047 2570
tri 2047 2566 2051 2570 nw
tri 1679 2548 1697 2566 ne
rect 1697 2548 2029 2566
tri 2029 2548 2047 2566 nw
tri 4149 2448 4176 2475 se
tri 4135 2434 4149 2448 se
rect 4149 2434 4176 2448
tri 4095 2394 4135 2434 se
rect 4135 2394 4176 2434
tri 4157 2364 4159 2366 ne
rect 4159 2364 4176 2366
rect 2882 2347 3052 2364
tri 3052 2347 3069 2364 sw
tri 4159 2347 4176 2364 ne
rect 2882 2313 3069 2347
tri 3069 2313 3103 2347 sw
rect 2882 2312 4177 2313
tri 3030 2261 3081 2312 ne
rect 3081 2261 4177 2312
rect 4229 2261 4241 2313
rect 4293 2261 4299 2313
tri 1537 2012 1546 2021 se
tri 1513 1988 1537 2012 se
rect 1537 1988 1546 2012
tri 1512 1987 1513 1988 se
rect 1513 1987 1546 1988
tri 1598 2012 1605 2019 sw
rect 3715 2012 4215 2018
rect 1598 1988 1605 2012
tri 1605 1988 1629 2012 sw
rect 1598 1987 1629 1988
tri 1629 1987 1630 1988 sw
rect 3264 1936 3270 1988
rect 3322 1983 3388 1988
rect 3440 1936 3446 1988
rect 3264 1910 3285 1936
rect 3421 1910 3446 1936
rect 3264 1858 3270 1910
rect 3440 1858 3446 1910
rect 3767 1960 4163 2012
rect 3715 1948 4215 1960
rect 3767 1896 4163 1948
rect 3715 1890 4215 1896
rect 4482 1951 4534 3514
tri 4534 3505 4543 3514 nw
tri 4593 3435 4628 3470 se
rect 4628 3448 4680 5072
rect 4628 3435 4667 3448
tri 4667 3435 4680 3448 nw
tri 4581 3423 4593 3435 se
rect 4593 3423 4655 3435
tri 4655 3423 4667 3435 nw
tri 3264 1847 3275 1858 ne
rect 3275 1847 3285 1858
rect 3421 1847 3435 1858
tri 3435 1847 3446 1858 nw
rect 4482 1887 4534 1899
rect 4482 1829 4534 1835
tri 4562 3404 4581 3423 se
rect 4581 3404 4636 3423
tri 4636 3404 4655 3423 nw
tri 705 1496 709 1500 ne
rect 709 1496 739 1500
tri 709 1475 730 1496 ne
rect 730 1475 739 1496
rect 767 1496 788 1500
tri 788 1496 792 1500 nw
tri 767 1475 788 1496 nw
tri 730 1466 739 1475 ne
tri 2864 1361 2867 1364 ne
rect 2867 1361 2888 1364
tri 2388 1351 2398 1361 ne
rect 2436 1351 2460 1361
tri 2460 1351 2470 1361 nw
tri 2867 1351 2877 1361 ne
rect 2877 1351 2888 1361
rect 2436 1339 2448 1351
tri 2448 1339 2460 1351 nw
tri 2877 1340 2888 1351 ne
rect 2915 1361 2946 1364
tri 2946 1361 2949 1364 nw
rect 2915 1340 2925 1361
tri 2925 1340 2946 1361 nw
rect 2915 1339 2924 1340
tri 2924 1339 2925 1340 nw
tri 2436 1327 2448 1339 nw
tri 2915 1330 2924 1339 nw
tri 613 1163 634 1184 sw
tri 558 1159 562 1163 se
tri 549 1150 558 1159 se
rect 558 1150 562 1159
rect 613 1159 634 1163
tri 634 1159 638 1163 sw
rect 613 1150 638 1159
tri 638 1150 647 1159 sw
tri -267 1009 -236 1040 sw
rect -267 1006 -236 1009
tri -236 1006 -233 1009 sw
rect 846 671 852 723
rect 904 671 916 723
rect 968 671 974 723
tri -182 591 -174 599 se
tri -204 569 -182 591 se
rect -182 569 -174 591
tri -216 557 -204 569 se
rect -204 557 -174 569
tri -217 556 -216 557 se
rect -216 556 -174 557
tri -124 569 -102 591 sw
rect -124 557 -102 569
tri -102 557 -90 569 sw
rect -124 556 -90 557
tri -90 556 -89 557 sw
tri -188 503 -187 504 ne
rect -187 503 -154 504
tri -361 499 -357 503 sw
tri -187 499 -183 503 ne
rect -183 499 -154 503
tri -399 489 -389 499 se
rect -361 489 -357 499
tri -357 489 -347 499 sw
tri -183 489 -173 499 ne
rect -173 489 -154 499
tri -173 470 -154 489 ne
rect -128 473 -123 504
tri -128 470 -125 473 ne
rect -125 470 -123 473
tri -123 470 -89 504 nw
tri -125 469 -124 470 ne
tri -124 469 -123 470 nw
tri 4226 428 4245 447 se
tri 4211 413 4226 428 se
rect 4226 413 4245 428
rect 4562 386 4614 3404
tri 4614 3382 4636 3404 nw
rect 4717 2941 4769 5087
rect 7847 5073 7856 5129
rect 7912 5073 7937 5129
rect 7993 5073 8018 5129
rect 8074 5073 8099 5129
rect 8155 5073 8180 5129
rect 8236 5073 8261 5129
rect 8317 5073 8341 5129
rect 8397 5073 8421 5129
rect 8477 5073 8501 5129
rect 8557 5073 8581 5129
rect 8637 5073 8661 5129
rect 8717 5073 8741 5129
rect 8797 5073 8821 5129
rect 8877 5073 8901 5129
rect 8957 5073 8981 5129
rect 9037 5073 9061 5129
rect 9117 5073 9141 5129
rect 9197 5073 9221 5129
rect 9277 5073 9301 5129
rect 9357 5073 9381 5129
rect 9437 5073 9461 5129
rect 9517 5073 9541 5129
rect 9597 5073 9621 5129
rect 9677 5073 9701 5129
rect 9757 5073 9781 5129
rect 9837 5073 9861 5129
rect 9917 5073 9941 5129
rect 9997 5073 10021 5129
rect 10077 5073 10101 5129
rect 10157 5073 10181 5129
rect 10237 5073 10261 5129
rect 10317 5073 10341 5129
rect 10397 5073 10421 5129
rect 10477 5073 10501 5129
rect 10557 5073 10581 5129
rect 10637 5073 10661 5129
rect 10717 5073 10741 5129
rect 10797 5073 10821 5129
rect 10877 5073 10901 5129
rect 10957 5073 10981 5129
rect 11037 5073 11061 5129
rect 11117 5073 11141 5129
rect 11197 5073 11206 5129
rect 7847 5072 11206 5073
rect 13983 5273 14035 5279
rect 13983 5206 14035 5221
rect 13983 5139 14035 5154
rect 13983 5072 14035 5087
rect 4814 5047 5032 5053
rect 4814 5044 4955 5047
rect 5007 5044 5032 5047
rect 4870 4988 4894 5044
rect 4950 4995 4955 5044
rect 4950 4988 4974 4995
rect 5030 4988 5032 5044
rect 13983 5005 14035 5020
rect 4814 4975 5032 4988
rect 4814 4923 4955 4975
rect 5007 4923 5032 4975
rect 4814 4919 5032 4923
rect 4870 4863 4894 4919
rect 4950 4902 4974 4919
rect 4950 4863 4955 4902
rect 5030 4863 5032 4919
rect 4814 4850 4955 4863
rect 5007 4850 5032 4863
rect 4814 4829 5032 4850
rect 4814 4793 4955 4829
rect 5007 4793 5032 4829
rect 4870 4737 4894 4793
rect 4950 4777 4955 4793
rect 4950 4756 4974 4777
rect 4950 4737 4955 4756
rect 5030 4737 5032 4793
rect 4814 4704 4955 4737
rect 5007 4704 5032 4737
rect 4814 4683 5032 4704
rect 4814 4667 4955 4683
rect 5007 4667 5032 4683
rect 4870 4611 4894 4667
rect 4950 4631 4955 4667
rect 4950 4611 4974 4631
rect 5030 4611 5032 4667
rect 11453 4953 11985 4989
tri 11985 4953 12021 4989 sw
rect 11453 4938 12021 4953
tri 12021 4938 12036 4953 sw
rect 13983 4938 14035 4953
rect 11453 4886 12036 4938
tri 12036 4886 12088 4938 sw
rect 11453 4871 12088 4886
tri 12088 4871 12103 4886 sw
rect 13983 4871 14035 4886
rect 11453 4819 12103 4871
tri 12103 4819 12155 4871 sw
rect 11453 4803 12155 4819
tri 12155 4803 12171 4819 sw
rect 13983 4803 14035 4819
rect 11453 4751 12171 4803
tri 12171 4751 12223 4803 sw
rect 11453 4735 12223 4751
tri 12223 4735 12239 4751 sw
rect 13983 4735 14035 4751
rect 11453 4703 12239 4735
tri 12239 4703 12271 4735 sw
rect 11453 4683 13156 4703
tri 13156 4683 13176 4703 sw
rect 11453 4667 13176 4683
tri 13176 4667 13192 4683 sw
rect 13983 4667 14035 4683
rect 11453 4661 13192 4667
tri 13192 4661 13198 4667 sw
rect 11453 4650 13833 4661
tri 13135 4648 13137 4650 ne
rect 13137 4648 13833 4650
tri 13833 4648 13846 4661 sw
tri 13137 4615 13170 4648 ne
rect 13170 4615 13846 4648
tri 13846 4615 13879 4648 sw
rect 4814 4610 5032 4611
rect 4814 4558 4955 4610
rect 5007 4558 5032 4610
tri 13170 4609 13176 4615 ne
rect 13176 4609 13879 4615
tri 13811 4574 13846 4609 ne
rect 13846 4574 13879 4609
tri 13879 4574 13920 4615 sw
tri 13846 4561 13859 4574 ne
rect 13859 4561 13920 4574
tri 5513 4558 5516 4561 se
rect 5516 4558 13553 4561
tri 13553 4558 13556 4561 sw
tri 13859 4558 13862 4561 ne
rect 13862 4558 13920 4561
rect 4814 4541 5032 4558
rect 4870 4485 4894 4541
rect 4950 4537 4974 4541
rect 4950 4485 4955 4537
rect 5030 4485 5032 4541
tri 5476 4521 5513 4558 se
rect 5513 4552 13556 4558
tri 13556 4552 13562 4558 sw
tri 13862 4552 13868 4558 ne
rect 5513 4533 13562 4552
rect 5513 4521 5516 4533
tri 5516 4521 5528 4533 nw
tri 13527 4521 13539 4533 ne
rect 13539 4521 13562 4533
tri 5460 4505 5476 4521 se
rect 5476 4505 5500 4521
tri 5500 4505 5516 4521 nw
tri 13539 4505 13555 4521 ne
rect 13555 4505 13562 4521
tri 13562 4505 13609 4552 sw
rect 4814 4476 5032 4485
tri 5436 4481 5460 4505 se
rect 5460 4481 5476 4505
tri 5476 4481 5500 4505 nw
tri 5516 4481 5540 4505 se
rect 5540 4481 12584 4505
tri 5431 4476 5436 4481 se
rect 5436 4476 5465 4481
tri 5425 4470 5431 4476 se
rect 5431 4470 5465 4476
tri 5465 4470 5476 4481 nw
tri 5505 4470 5516 4481 se
rect 5516 4477 12584 4481
rect 5516 4470 5545 4477
tri 5545 4470 5552 4477 nw
tri 12558 4470 12565 4477 ne
rect 12565 4470 12584 4477
tri 12584 4470 12619 4505 sw
tri 13555 4504 13556 4505 ne
rect 13556 4504 13609 4505
tri 13609 4504 13610 4505 sw
tri 5420 4465 5425 4470 se
rect 5425 4465 5460 4470
tri 5460 4465 5465 4470 nw
tri 5500 4465 5505 4470 se
rect 5505 4465 5540 4470
tri 5540 4465 5545 4470 nw
tri 12565 4465 12570 4470 ne
rect 12570 4465 12619 4470
tri 5396 4441 5420 4465 se
rect 5420 4441 5436 4465
tri 5436 4441 5460 4465 nw
tri 5476 4441 5500 4465 se
tri 5394 4439 5396 4441 se
rect 5396 4439 5434 4441
tri 5434 4439 5436 4441 nw
tri 5474 4439 5476 4441 se
rect 5476 4439 5500 4441
rect 5075 4358 5081 4410
rect 5133 4358 5145 4410
rect 5197 4358 5203 4410
tri 5087 4328 5117 4358 ne
rect 5117 4328 5173 4358
tri 5173 4328 5203 4358 nw
tri 5117 4324 5121 4328 ne
rect 5121 3899 5173 4328
tri 5276 3951 5279 3954 ne
rect 5279 3951 5310 3954
tri 5279 3920 5310 3951 ne
tri 5173 3899 5184 3910 sw
rect 5121 3891 5184 3899
tri 5184 3891 5192 3899 sw
rect 5121 3888 5192 3891
tri 5121 3870 5139 3888 ne
rect 5139 3870 5192 3888
tri 5192 3870 5213 3891 sw
tri 5139 3858 5151 3870 ne
rect 5151 3858 5213 3870
tri 5213 3858 5225 3870 sw
tri 5151 3817 5192 3858 ne
rect 5192 3817 5225 3858
tri 5225 3817 5266 3858 sw
tri 5192 3806 5203 3817 ne
rect 5203 3806 5266 3817
tri 5203 3799 5210 3806 ne
rect 5210 3799 5266 3806
tri 5210 3795 5214 3799 ne
rect 4717 2877 4769 2889
rect 4717 2819 4769 2825
tri 5207 2382 5214 2389 se
rect 5214 2382 5266 3799
tri 5138 2313 5207 2382 se
rect 5207 2313 5266 2382
rect 5138 2261 5144 2313
rect 5196 2261 5208 2313
rect 5260 2261 5266 2313
rect 5394 1502 5422 4439
tri 5422 4427 5434 4439 nw
tri 5462 4427 5474 4439 se
rect 5474 4427 5500 4439
tri 5460 4425 5462 4427 se
rect 5462 4425 5500 4427
tri 5500 4425 5540 4465 nw
tri 12570 4451 12584 4465 ne
rect 12584 4451 12619 4465
tri 12584 4449 12586 4451 ne
rect 12586 4449 12619 4451
tri 13556 4450 13610 4504 ne
tri 13610 4450 13664 4504 sw
tri 6448 4425 6472 4449 se
rect 6472 4444 11174 4449
tri 11174 4444 11179 4449 sw
tri 12586 4444 12591 4449 ne
rect 6472 4425 11179 4444
tri 11179 4425 11198 4444 sw
tri 5450 4415 5460 4425 se
rect 5460 4415 5490 4425
tri 5490 4415 5500 4425 nw
tri 6438 4415 6448 4425 se
rect 6448 4419 11198 4425
tri 11198 4419 11204 4425 sw
rect 6448 4415 11204 4419
tri 11204 4415 11208 4419 sw
rect 5450 4410 5485 4415
tri 5485 4410 5490 4415 nw
tri 6434 4411 6438 4415 se
rect 6438 4411 11208 4415
tri 6433 4410 6434 4411 se
rect 6434 4410 6500 4411
rect 5450 3514 5478 4410
tri 5478 4403 5485 4410 nw
rect 5652 4358 5658 4410
rect 5710 4358 5722 4410
rect 5774 4403 6500 4410
tri 6500 4403 6508 4411 nw
tri 11158 4403 11166 4411 ne
rect 11166 4403 11208 4411
tri 11208 4403 11220 4415 sw
rect 5774 4383 6480 4403
tri 6480 4383 6500 4403 nw
tri 11166 4383 11186 4403 ne
rect 11186 4383 11220 4403
rect 5774 4365 6462 4383
tri 6462 4365 6480 4383 nw
tri 6575 4365 6593 4383 se
rect 6593 4370 10277 4383
tri 10277 4370 10290 4383 sw
tri 11186 4370 11199 4383 ne
rect 11199 4370 11220 4383
rect 6593 4365 10290 4370
tri 10290 4365 10295 4370 sw
tri 11199 4365 11204 4370 ne
rect 11204 4365 11220 4370
tri 11220 4365 11258 4403 sw
rect 5774 4358 6455 4365
tri 6455 4358 6462 4365 nw
tri 6568 4358 6575 4365 se
rect 6575 4358 10295 4365
tri 6559 4349 6568 4358 se
rect 6568 4349 10295 4358
tri 10295 4349 10311 4365 sw
tri 11204 4349 11220 4365 ne
tri 6543 4333 6559 4349 se
rect 6559 4347 10311 4349
tri 10311 4347 10313 4349 sw
rect 6559 4333 6593 4347
tri 6593 4333 6607 4347 nw
tri 10239 4333 10253 4347 ne
rect 10253 4333 10313 4347
tri 10313 4333 10327 4347 sw
tri 6528 4318 6543 4333 se
rect 5915 4295 6186 4318
rect 5915 4293 5924 4295
rect 5915 4241 5921 4293
rect 5915 4239 5924 4241
rect 5980 4239 6023 4295
rect 6079 4239 6121 4295
rect 6177 4293 6186 4295
rect 6180 4241 6186 4293
tri 6493 4283 6528 4318 se
rect 6528 4283 6543 4318
tri 6543 4283 6593 4333 nw
tri 10253 4296 10290 4333 ne
rect 10290 4296 10327 4333
tri 10327 4296 10364 4333 sw
tri 10290 4283 10303 4296 ne
rect 10303 4283 10364 4296
tri 6479 4269 6493 4283 se
rect 6493 4269 6529 4283
tri 6529 4269 6543 4283 nw
tri 10303 4274 10312 4283 ne
rect 6177 4239 6186 4241
rect 5915 4216 6186 4239
tri 6443 4233 6479 4269 se
rect 6479 4233 6493 4269
tri 6493 4233 6529 4269 nw
tri 6440 4230 6443 4233 se
rect 6443 4230 6490 4233
tri 6490 4230 6493 4233 nw
tri 6427 4217 6440 4230 se
rect 6440 4217 6477 4230
tri 6477 4217 6490 4230 nw
rect 10312 4217 10364 4283
tri 10364 4217 10377 4230 sw
tri 6426 4216 6427 4217 se
rect 6427 4216 6456 4217
tri 6406 4196 6426 4216 se
rect 6426 4196 6456 4216
tri 6456 4196 6477 4217 nw
rect 10312 4196 10377 4217
tri 10377 4196 10398 4217 sw
tri 6398 4188 6406 4196 se
rect 6406 4188 6448 4196
tri 6448 4188 6456 4196 nw
tri 6124 4156 6156 4188 se
rect 6156 4160 6420 4188
tri 6420 4160 6448 4188 nw
rect 6156 4156 6174 4160
tri 6174 4156 6178 4160 nw
tri 6115 4147 6124 4156 se
rect 6124 4147 6165 4156
tri 6165 4147 6174 4156 nw
tri 6112 4144 6115 4147 se
rect 6115 4144 6162 4147
tri 6162 4144 6165 4147 nw
rect 10312 4144 10318 4196
rect 10370 4144 10382 4196
rect 10434 4144 10440 4196
rect 11220 4185 11258 4365
tri 11220 4156 11249 4185 ne
rect 11249 4156 11258 4185
tri 11258 4156 11303 4201 sw
tri 11249 4147 11258 4156 ne
rect 11258 4147 11303 4156
tri 11258 4144 11261 4147 ne
rect 11261 4144 11303 4147
tri 6108 4140 6112 4144 se
rect 6112 4140 6158 4144
tri 6158 4140 6162 4144 nw
tri 9816 4140 9820 4144 ne
rect 9820 4140 9850 4144
tri 6106 4138 6108 4140 se
rect 6108 4138 6156 4140
tri 6156 4138 6158 4140 nw
rect 6877 4138 6909 4140
tri 6909 4138 6911 4140 nw
tri 9820 4138 9822 4140 ne
rect 9822 4138 9850 4140
tri 6097 4129 6106 4138 se
rect 6106 4129 6147 4138
tri 6147 4129 6156 4138 nw
rect 6877 4129 6900 4138
tri 6900 4129 6909 4138 nw
tri 9822 4129 9831 4138 ne
rect 9831 4129 9850 4138
tri 6074 4106 6097 4129 se
rect 6097 4106 6124 4129
tri 6124 4106 6147 4129 nw
tri 6877 4106 6900 4129 nw
tri 9831 4125 9835 4129 ne
rect 9835 4125 9850 4129
rect 9895 4140 9910 4144
tri 9910 4140 9914 4144 nw
tri 11261 4140 11265 4144 ne
rect 11265 4140 11303 4144
tri 11303 4140 11319 4156 sw
rect 9895 4129 9899 4140
tri 9899 4129 9910 4140 nw
tri 11265 4129 11276 4140 ne
rect 11276 4129 11319 4140
tri 11319 4129 11330 4140 sw
tri 9895 4125 9899 4129 nw
tri 11276 4125 11280 4129 ne
rect 11280 4125 11330 4129
tri 9835 4110 9850 4125 ne
tri 11280 4110 11295 4125 ne
rect 11295 4110 11330 4125
tri 11295 4106 11299 4110 ne
rect 11299 4106 11330 4110
tri 11330 4106 11353 4129 sw
tri 6070 4102 6074 4106 se
rect 6074 4102 6120 4106
tri 6120 4102 6124 4106 nw
tri 11299 4102 11303 4106 ne
rect 11303 4102 11353 4106
tri 11353 4102 11357 4106 sw
tri 5595 4077 5620 4102 se
rect 5620 4077 6095 4102
tri 6095 4077 6120 4102 nw
tri 11303 4077 11328 4102 ne
rect 11328 4077 11357 4102
tri 11357 4077 11382 4102 sw
tri 5583 4065 5595 4077 se
rect 5595 4066 6084 4077
tri 6084 4066 6095 4077 nw
tri 11328 4066 11339 4077 ne
rect 11339 4066 11382 4077
rect 5595 4065 5657 4066
tri 5657 4065 5658 4066 nw
tri 11339 4065 11340 4066 ne
rect 11340 4065 11382 4066
tri 11382 4065 11394 4077 sw
tri 5566 4048 5583 4065 se
rect 5583 4048 5640 4065
tri 5640 4048 5657 4065 nw
tri 11340 4048 11357 4065 ne
rect 11357 4048 11394 4065
tri 11394 4048 11411 4065 sw
tri 5546 4028 5566 4048 se
rect 5566 4028 5620 4048
tri 5620 4028 5640 4048 nw
tri 11357 4028 11377 4048 ne
rect 11377 4028 11411 4048
tri 5536 4018 5546 4028 se
rect 5546 4018 5610 4028
tri 5610 4018 5620 4028 nw
tri 11377 4018 11387 4028 ne
rect 11387 4018 11411 4028
rect 5536 4013 5605 4018
tri 5605 4013 5610 4018 nw
tri 11387 4013 11392 4018 ne
rect 11392 4013 11411 4018
tri 11411 4013 11446 4048 sw
rect 5536 4009 5601 4013
tri 5601 4009 5605 4013 nw
tri 11392 4009 11396 4013 ne
rect 11396 4009 11446 4013
rect 5536 4004 5596 4009
tri 5596 4004 5601 4009 nw
tri 9472 4004 9477 4009 se
tri 5478 3514 5481 3517 sw
rect 5450 3493 5481 3514
tri 5481 3493 5502 3514 sw
rect 5450 3487 5502 3493
rect 5450 3423 5502 3435
rect 5450 3365 5502 3371
tri 5533 3159 5536 3162 se
rect 5536 3159 5588 4004
tri 5588 3996 5596 4004 nw
tri 7023 3996 7031 4004 ne
rect 7031 3996 7057 4004
tri 7031 3975 7052 3996 ne
rect 7052 3975 7057 3996
tri 7052 3970 7057 3975 ne
rect 7073 3975 7079 4004
tri 7079 3975 7108 4004 nw
tri 9443 3975 9472 4004 se
rect 9472 3975 9477 4004
tri 9505 4004 9510 4009 sw
tri 11396 4004 11401 4009 ne
rect 11401 4004 11446 4009
tri 11446 4004 11455 4013 sw
rect 9505 3994 9510 4004
tri 9510 3994 9520 4004 sw
tri 11401 3994 11411 4004 ne
rect 11411 3994 11455 4004
tri 11455 3994 11465 4004 sw
rect 9505 3975 9520 3994
tri 9520 3975 9539 3994 sw
tri 11411 3975 11430 3994 ne
rect 11430 3975 11465 3994
tri 11465 3975 11484 3994 sw
rect 7073 3970 7074 3975
tri 7074 3970 7079 3975 nw
tri 11430 3974 11431 3975 ne
rect 11431 3974 11484 3975
tri 9846 3970 9850 3974 se
tri 7073 3969 7074 3970 nw
tri 9845 3969 9846 3970 se
rect 9846 3969 9850 3970
tri 9827 3951 9845 3969 se
rect 9845 3951 9850 3969
tri 9816 3940 9827 3951 se
rect 9827 3940 9850 3951
tri 9898 3973 9899 3974 sw
tri 11431 3973 11432 3974 ne
rect 11432 3973 11484 3974
rect 9898 3970 9899 3973
tri 9899 3970 9902 3973 sw
tri 10054 3970 10057 3973 sw
tri 11432 3970 11435 3973 ne
rect 11435 3970 11484 3973
tri 11484 3970 11489 3975 sw
rect 9898 3969 9902 3970
tri 9902 3969 9903 3970 sw
rect 10054 3969 10057 3970
tri 10057 3969 10058 3970 sw
tri 11435 3969 11436 3970 ne
rect 11436 3969 11489 3970
tri 11489 3969 11490 3970 sw
rect 9898 3964 9903 3969
tri 9903 3964 9908 3969 sw
rect 9898 3951 9908 3964
tri 9908 3951 9921 3964 sw
tri 9989 3951 10002 3964 se
rect 9898 3940 9921 3951
tri 9921 3940 9932 3951 sw
tri 9978 3940 9989 3951 se
rect 9989 3940 10002 3951
tri 9977 3939 9978 3940 se
rect 9978 3939 10002 3940
rect 10054 3955 10058 3969
tri 10058 3955 10072 3969 sw
tri 11436 3955 11450 3969 ne
rect 11450 3955 11490 3969
rect 10054 3951 10072 3955
tri 10072 3951 10076 3955 sw
tri 10200 3951 10204 3955 sw
tri 10904 3951 10908 3955 se
tri 11450 3951 11454 3955 ne
rect 11454 3951 11490 3955
tri 11490 3951 11508 3969 sw
rect 10054 3939 10076 3951
tri 10076 3939 10088 3951 sw
rect 10200 3940 10204 3951
tri 10204 3940 10215 3951 sw
tri 10893 3940 10904 3951 se
rect 10904 3940 10908 3951
tri 11454 3940 11465 3951 ne
rect 11465 3940 11508 3951
tri 11508 3940 11519 3951 sw
rect 10200 3921 10215 3940
tri 10215 3921 10234 3940 sw
tri 10874 3921 10893 3940 se
rect 10893 3921 10908 3940
tri 11465 3921 11484 3940 ne
rect 11484 3921 11519 3940
tri 11484 3899 11506 3921 ne
rect 11506 3899 11519 3921
tri 11519 3899 11560 3940 sw
tri 11506 3892 11513 3899 ne
rect 11513 3892 11560 3899
tri 5619 3870 5641 3892 ne
rect 5641 3870 5655 3892
tri 5641 3858 5653 3870 ne
rect 5653 3858 5655 3870
tri 5653 3856 5655 3858 ne
rect 5692 3886 5741 3892
tri 5741 3886 5747 3892 nw
tri 11513 3886 11519 3892 ne
rect 11519 3886 11560 3892
tri 11560 3886 11573 3899 sw
rect 5692 3870 5725 3886
tri 5725 3870 5741 3886 nw
tri 11519 3870 11535 3886 ne
rect 11535 3870 11573 3886
tri 11573 3870 11589 3886 sw
rect 5692 3858 5713 3870
tri 5713 3858 5725 3870 nw
tri 11535 3858 11547 3870 ne
rect 11547 3858 11589 3870
tri 11589 3858 11601 3870 sw
rect 5692 3856 5711 3858
tri 5711 3856 5713 3858 nw
tri 11547 3856 11549 3858 ne
rect 11549 3856 11601 3858
tri 5692 3837 5711 3856 nw
tri 11549 3837 11568 3856 ne
rect 11568 3837 11601 3856
tri 11568 3832 11573 3837 ne
rect 11573 3832 11601 3837
tri 11601 3832 11627 3858 sw
tri 11573 3806 11599 3832 ne
rect 11599 3806 11627 3832
tri 11627 3806 11653 3832 sw
tri 11599 3799 11606 3806 ne
rect 11606 3799 11653 3806
tri 11653 3799 11660 3806 sw
tri 11606 3780 11625 3799 ne
rect 11625 3780 11660 3799
tri 11660 3780 11679 3799 sw
tri 11625 3778 11627 3780 ne
rect 11627 3778 11679 3780
tri 11679 3778 11681 3780 sw
tri 11627 3728 11677 3778 ne
rect 11677 3728 11681 3778
tri 11681 3728 11731 3778 sw
tri 11677 3724 11681 3728 ne
rect 11681 3724 11731 3728
tri 11731 3724 11735 3728 sw
tri 11681 3713 11692 3724 ne
rect 11692 3713 11735 3724
tri 11735 3713 11746 3724 sw
tri 11692 3709 11696 3713 ne
rect 11696 3709 11746 3713
tri 11746 3709 11750 3713 sw
tri 11696 3683 11722 3709 ne
rect 11722 3683 11750 3709
tri 8050 3678 8055 3683 ne
rect 8055 3678 8084 3683
tri 8055 3673 8060 3678 ne
rect 8060 3673 8084 3678
tri 8060 3649 8084 3673 ne
rect 8111 3678 8140 3683
tri 8140 3678 8145 3683 nw
tri 11722 3678 11727 3683 ne
rect 11727 3678 11750 3683
rect 8111 3673 8135 3678
tri 8135 3673 8140 3678 nw
rect 9110 3673 10247 3678
rect 8111 3670 8132 3673
tri 8132 3670 8135 3673 nw
tri 8111 3649 8132 3670 nw
rect 9110 3621 9119 3673
rect 9171 3621 9194 3673
rect 9246 3621 9268 3673
rect 9320 3621 9342 3673
rect 9394 3626 10247 3673
rect 10299 3626 10315 3678
rect 10367 3626 10383 3678
rect 10435 3626 10451 3678
rect 10503 3626 10519 3678
rect 10571 3626 10587 3678
rect 10639 3626 10654 3678
rect 10706 3670 11373 3678
tri 11373 3670 11381 3678 sw
tri 11727 3670 11735 3678 ne
rect 11735 3670 11750 3678
tri 11750 3670 11789 3709 sw
rect 10706 3657 11381 3670
tri 11381 3657 11394 3670 sw
tri 11735 3657 11748 3670 ne
rect 11748 3657 11789 3670
tri 11789 3657 11802 3670 sw
rect 10706 3632 11394 3657
tri 11394 3632 11419 3657 sw
tri 11748 3632 11773 3657 ne
rect 11773 3632 11802 3657
tri 11802 3632 11827 3657 sw
rect 10706 3626 11419 3632
rect 9394 3621 11419 3626
rect 9110 3616 11419 3621
tri 11419 3616 11435 3632 sw
tri 11773 3616 11789 3632 ne
rect 11789 3616 11827 3632
tri 11827 3616 11843 3632 sw
rect 9110 3609 11435 3616
rect 9110 3557 9119 3609
rect 9171 3557 9194 3609
rect 9246 3557 9268 3609
rect 9320 3557 9342 3609
rect 9394 3606 11435 3609
rect 9394 3557 10247 3606
rect 9110 3554 10247 3557
rect 10299 3554 10315 3606
rect 10367 3554 10383 3606
rect 10435 3554 10451 3606
rect 10503 3554 10519 3606
rect 10571 3554 10587 3606
rect 10639 3554 10654 3606
rect 10706 3604 11435 3606
tri 11435 3604 11447 3616 sw
tri 11789 3604 11801 3616 ne
rect 11801 3604 11843 3616
tri 11843 3604 11855 3616 sw
rect 10706 3562 11447 3604
tri 11447 3562 11489 3604 sw
tri 11801 3562 11843 3604 ne
rect 11843 3562 11855 3604
tri 11855 3562 11897 3604 sw
rect 10706 3554 11489 3562
tri 11489 3554 11497 3562 sw
tri 11843 3554 11851 3562 ne
rect 11851 3554 11897 3562
tri 11259 3552 11261 3554 ne
rect 11261 3552 11497 3554
tri 11497 3552 11499 3554 sw
tri 11851 3552 11853 3554 ne
rect 11853 3552 11897 3554
tri 11261 3546 11267 3552 ne
rect 11267 3546 11499 3552
tri 11499 3546 11505 3552 sw
tri 11853 3546 11859 3552 ne
tri 11267 3514 11299 3546 ne
rect 11299 3514 11505 3546
tri 11505 3514 11537 3546 sw
tri 11299 3462 11351 3514 ne
rect 11351 3499 11537 3514
tri 11537 3499 11552 3514 sw
rect 11351 3462 11552 3499
tri 11552 3462 11589 3499 sw
rect 5826 3450 5848 3462
tri 5848 3450 5860 3462 nw
tri 11351 3450 11363 3462 ne
rect 11363 3450 11589 3462
tri 11589 3450 11601 3462 sw
tri 5826 3428 5848 3450 nw
tri 11363 3428 11385 3450 ne
rect 11385 3428 11601 3450
tri 11385 3398 11415 3428 ne
rect 11415 3398 11601 3428
tri 11601 3398 11653 3450 sw
tri 11415 3388 11425 3398 ne
rect 11425 3388 11653 3398
tri 11653 3388 11663 3398 sw
tri 11425 3336 11477 3388 ne
rect 11477 3336 11663 3388
tri 11663 3336 11715 3388 sw
tri 11477 3316 11497 3336 ne
rect 11497 3316 11715 3336
tri 11715 3316 11735 3336 sw
tri 11497 3296 11517 3316 ne
rect 11517 3305 11735 3316
tri 11735 3305 11746 3316 sw
rect 11517 3296 11746 3305
tri 11517 3291 11522 3296 ne
rect 11522 3291 11746 3296
tri 11522 3261 11552 3291 ne
tri 6509 3204 6512 3207 se
tri 6508 3203 6509 3204 se
rect 6509 3203 6512 3204
tri 6501 3196 6508 3203 se
rect 6508 3196 6512 3203
tri 6464 3159 6501 3196 se
rect 6501 3159 6512 3196
tri 6555 3159 6592 3196 sw
tri 5525 3151 5533 3159 se
rect 5533 3151 5588 3159
tri 5523 3149 5525 3151 se
rect 5525 3149 5588 3151
tri 5489 3115 5523 3149 se
rect 5523 3140 5588 3149
rect 5523 3115 5563 3140
tri 5563 3115 5588 3140 nw
tri 5462 3088 5489 3115 se
rect 5489 3088 5536 3115
tri 5536 3088 5563 3115 nw
rect 5462 1589 5514 3088
tri 5514 3066 5536 3088 nw
rect 9018 3040 10356 3049
rect 9018 2986 9095 3040
rect 9151 2986 9175 3040
rect 9231 2986 9255 3040
rect 9311 2993 10356 3040
rect 10412 2993 10453 3049
rect 10509 2993 10550 3049
rect 10606 2993 10646 3049
rect 10702 2993 10712 3049
rect 9311 2986 10712 2993
rect 9018 2934 9024 2986
rect 9076 2984 9095 2986
rect 9156 2984 9175 2986
rect 9236 2984 9255 2986
rect 9076 2942 9104 2984
rect 9156 2942 9184 2984
rect 9236 2942 9263 2984
rect 9076 2934 9095 2942
rect 9156 2934 9175 2942
rect 9236 2934 9255 2942
rect 9315 2934 9342 2986
rect 9394 2945 10712 2986
rect 9394 2934 10356 2945
rect 9018 2910 9095 2934
rect 9151 2910 9175 2934
rect 9231 2910 9255 2934
rect 9311 2910 10356 2934
tri 6402 2878 6421 2897 sw
tri 8830 2878 8849 2897 se
tri 5640 2865 5653 2878 se
rect 6402 2865 6421 2878
tri 6421 2865 6434 2878 sw
tri 8817 2865 8830 2878 se
rect 8830 2865 8849 2878
rect 6402 2863 6434 2865
tri 6434 2863 6436 2865 sw
tri 8815 2863 8817 2865 se
rect 8817 2863 8849 2865
tri 8899 2863 8921 2885 sw
rect 9018 2858 9024 2910
rect 9076 2886 9095 2910
rect 9156 2886 9175 2910
rect 9236 2886 9255 2910
rect 9076 2858 9104 2886
rect 9156 2858 9184 2886
rect 9236 2858 9263 2886
rect 9315 2858 9342 2910
rect 9394 2889 10356 2910
rect 10412 2889 10453 2945
rect 10509 2889 10550 2945
rect 10606 2889 10646 2945
rect 10702 2889 10712 2945
rect 9394 2858 10712 2889
rect 9018 2844 10712 2858
rect 9018 2834 9095 2844
rect 9151 2834 9175 2844
rect 9231 2834 9255 2844
rect 9311 2841 10712 2844
rect 9311 2834 10356 2841
tri 5684 2794 5703 2813 nw
rect 9018 2782 9024 2834
rect 9076 2788 9095 2834
rect 9156 2788 9175 2834
rect 9236 2788 9255 2834
rect 9076 2782 9104 2788
rect 9156 2782 9184 2788
rect 9236 2782 9263 2788
rect 9315 2782 9342 2834
rect 9394 2785 10356 2834
rect 10412 2785 10453 2841
rect 10509 2785 10550 2841
rect 10606 2785 10646 2841
rect 10702 2785 10712 2841
rect 9394 2782 10712 2785
rect 9018 2758 10712 2782
tri 6423 2718 6457 2752 ne
rect 9018 2706 9024 2758
rect 9076 2746 9104 2758
rect 9156 2746 9184 2758
rect 9236 2746 9263 2758
rect 9076 2706 9095 2746
rect 9156 2706 9175 2746
rect 9236 2706 9255 2746
rect 9315 2706 9342 2758
rect 9394 2737 10712 2758
rect 9394 2706 10356 2737
rect 9018 2690 9095 2706
rect 9151 2690 9175 2706
rect 9231 2690 9255 2706
rect 9311 2690 10356 2706
rect 9018 2681 10356 2690
rect 10412 2681 10453 2737
rect 10509 2681 10550 2737
rect 10606 2681 10646 2737
rect 10702 2681 10712 2737
rect 11552 2956 11746 3291
rect 11552 2904 11553 2956
rect 11605 2904 11623 2956
rect 11675 2904 11693 2956
rect 11745 2904 11746 2956
rect 11552 2891 11746 2904
rect 11552 2839 11553 2891
rect 11605 2839 11623 2891
rect 11675 2839 11693 2891
rect 11745 2839 11746 2891
rect 11552 2826 11746 2839
rect 11552 2774 11553 2826
rect 11605 2774 11623 2826
rect 11675 2774 11693 2826
rect 11745 2774 11746 2826
rect 11552 2761 11746 2774
rect 11552 2709 11553 2761
rect 11605 2709 11623 2761
rect 11675 2709 11693 2761
rect 11745 2709 11746 2761
rect 11552 2696 11746 2709
rect 11552 2644 11553 2696
rect 11605 2644 11623 2696
rect 11675 2644 11693 2696
rect 11745 2644 11746 2696
rect 11552 2631 11746 2644
rect 11552 2579 11553 2631
rect 11605 2579 11623 2631
rect 11675 2579 11693 2631
rect 11745 2579 11746 2631
rect 11552 2566 11746 2579
rect 11552 2514 11553 2566
rect 11605 2514 11623 2566
rect 11675 2514 11693 2566
rect 11745 2514 11746 2566
rect 11552 2500 11746 2514
rect 11859 2519 11897 3552
rect 12591 3514 12619 4449
tri 13610 4396 13664 4450 ne
tri 13664 4396 13718 4450 sw
tri 13664 4342 13718 4396 ne
tri 13718 4342 13772 4396 sw
tri 13718 4340 13720 4342 ne
rect 12922 4217 12928 4269
rect 12980 4217 12992 4269
rect 13044 4217 13552 4269
rect 13604 4217 13616 4269
rect 13668 4217 13674 4269
rect 12654 4129 13480 4135
rect 12654 4099 13428 4129
rect 12654 4043 12669 4099
rect 12725 4043 12759 4099
rect 12815 4043 12848 4099
rect 12904 4077 13428 4099
rect 12904 4065 13480 4077
rect 12904 4043 13428 4065
rect 12654 4013 13428 4043
rect 12654 4007 13480 4013
rect 13720 4091 13772 4342
rect 13720 4027 13772 4039
rect 13720 3969 13772 3975
rect 12933 3899 12939 3951
rect 12991 3899 13003 3951
rect 13055 3946 13220 3951
tri 13220 3946 13225 3951 sw
rect 13055 3944 13225 3946
tri 13225 3944 13227 3946 sw
rect 13055 3928 13227 3944
tri 13227 3928 13243 3944 sw
rect 13055 3922 13601 3928
rect 13055 3899 13549 3922
tri 13162 3870 13191 3899 ne
rect 13191 3870 13549 3899
tri 13191 3858 13203 3870 ne
rect 13203 3858 13601 3870
tri 13203 3806 13255 3858 ne
rect 13255 3806 13549 3858
tri 13255 3800 13261 3806 ne
rect 13261 3800 13601 3806
rect 13868 3922 13920 4558
rect 13868 3851 13920 3870
rect 13868 3780 13920 3799
rect 13983 3944 14035 4615
rect 13983 3880 14035 3892
rect 13983 3816 14035 3828
rect 13983 3758 14035 3764
rect 14063 3944 14115 8490
rect 14063 3855 14115 3892
rect 14143 8367 14195 8373
rect 14143 8300 14195 8315
rect 14143 8233 14195 8248
rect 14143 8166 14195 8181
rect 14143 8099 14195 8114
rect 14143 8032 14195 8047
rect 14143 7965 14195 7980
rect 14143 7897 14195 7913
rect 14143 7829 14195 7845
rect 14143 3946 14195 7777
rect 14143 3868 14195 3894
rect 14143 3810 14195 3816
rect 14063 3765 14115 3803
rect 13868 3722 13920 3728
rect 12933 3657 12939 3709
rect 12991 3657 13003 3709
rect 13055 3684 13227 3709
tri 13227 3684 13252 3709 sw
rect 14063 3707 14115 3713
rect 14143 3773 14195 3779
rect 14143 3709 14195 3721
tri 14132 3684 14143 3695 se
rect 13055 3657 13748 3684
tri 13205 3632 13230 3657 ne
rect 13230 3632 13748 3657
rect 13800 3632 13812 3684
rect 13864 3632 13870 3684
tri 14105 3657 14132 3684 se
rect 14132 3657 14143 3684
tri 14080 3632 14105 3657 se
rect 14105 3651 14195 3657
rect 14105 3632 14143 3651
tri 14069 3621 14080 3632 se
rect 14080 3621 14143 3632
tri 14143 3621 14173 3651 nw
tri 14052 3604 14069 3621 se
rect 14069 3604 14126 3621
tri 14126 3604 14143 3621 nw
rect 12924 3552 12930 3604
rect 12982 3552 12994 3604
rect 13046 3563 14085 3604
tri 14085 3563 14126 3604 nw
rect 14135 3563 14187 3569
rect 13046 3554 14076 3563
tri 14076 3554 14085 3563 nw
rect 13046 3552 14074 3554
tri 14074 3552 14076 3554 nw
tri 14133 3552 14135 3554 se
tri 14110 3529 14133 3552 se
rect 14133 3529 14135 3552
tri 12619 3514 12634 3529 sw
tri 14101 3520 14110 3529 se
rect 14110 3520 14135 3529
rect 13113 3514 14135 3520
rect 12591 3508 12634 3514
tri 12591 3493 12606 3508 ne
rect 12606 3493 12634 3508
tri 12606 3480 12619 3493 ne
rect 12619 3480 12634 3493
tri 12634 3480 12668 3514 sw
tri 12619 3462 12637 3480 ne
rect 12637 3462 12668 3480
tri 12668 3462 12686 3480 sw
rect 13165 3511 14135 3514
rect 13165 3499 14187 3511
rect 13165 3468 14135 3499
rect 13165 3462 13178 3468
tri 12637 3450 12649 3462 ne
rect 12649 3450 12686 3462
tri 12686 3450 12698 3462 sw
rect 13113 3450 13178 3462
tri 12649 3431 12668 3450 ne
rect 12668 3431 12698 3450
tri 12698 3431 12717 3450 sw
tri 12668 3403 12696 3431 ne
rect 12696 3403 12940 3431
tri 12910 3398 12915 3403 ne
rect 12915 3398 12940 3403
tri 12940 3398 12973 3431 sw
rect 13165 3447 13178 3450
tri 13178 3447 13199 3468 nw
tri 14108 3447 14129 3468 ne
rect 14129 3447 14135 3468
tri 13165 3434 13178 3447 nw
tri 14129 3441 14135 3447 ne
rect 14135 3441 14187 3447
tri 12915 3388 12925 3398 ne
rect 12925 3388 12973 3398
tri 12973 3388 12983 3398 sw
rect 13113 3392 13165 3398
tri 12925 3375 12938 3388 ne
rect 12938 3375 12983 3388
tri 12983 3375 12996 3388 sw
tri 12938 3373 12940 3375 ne
rect 12940 3373 12996 3375
tri 12940 3336 12977 3373 ne
rect 12977 3336 12996 3373
tri 12996 3336 13035 3375 sw
rect 14067 3336 14073 3388
rect 14125 3336 14137 3388
rect 14189 3336 14195 3388
tri 12977 3317 12996 3336 ne
rect 12996 3317 13035 3336
tri 13035 3317 13054 3336 sw
tri 14133 3317 14152 3336 ne
rect 14152 3317 14195 3336
tri 12996 3296 13017 3317 ne
rect 13017 3296 13054 3317
tri 13054 3296 13075 3317 sw
tri 14152 3302 14167 3317 ne
rect 13849 3296 13953 3302
tri 13017 3294 13019 3296 ne
rect 13019 3294 13075 3296
rect 12064 3292 12888 3294
tri 12888 3292 12890 3294 sw
tri 13019 3292 13021 3294 ne
rect 13021 3292 13075 3294
tri 13075 3292 13079 3296 sw
rect 12064 3291 12913 3292
rect 12064 3239 12100 3291
rect 12152 3239 12169 3291
rect 12221 3239 12238 3291
rect 12290 3239 12307 3291
rect 12359 3239 12376 3291
rect 12428 3239 12445 3291
rect 12497 3239 12514 3291
rect 12566 3239 12583 3291
rect 12635 3239 12651 3291
rect 12703 3239 12719 3291
rect 12771 3239 12787 3291
rect 12839 3239 12855 3291
rect 12907 3259 12913 3291
tri 12913 3259 12946 3292 sw
tri 13021 3259 13054 3292 ne
rect 13054 3267 13079 3292
tri 13079 3267 13104 3292 sw
tri 13843 3267 13849 3273 se
rect 13849 3267 13875 3296
rect 13054 3259 13104 3267
tri 13104 3259 13112 3267 sw
tri 13835 3259 13843 3267 se
rect 13843 3259 13875 3267
rect 12907 3244 12946 3259
tri 12946 3244 12961 3259 sw
tri 13054 3244 13069 3259 ne
rect 13069 3244 13112 3259
tri 13112 3244 13127 3259 sw
tri 13820 3244 13835 3259 se
rect 13835 3244 13875 3259
rect 13927 3244 13953 3296
rect 12907 3239 12961 3244
rect 12064 3209 12961 3239
tri 12961 3209 12996 3244 sw
tri 13069 3209 13104 3244 ne
rect 13104 3209 13127 3244
rect 12064 3204 12996 3209
tri 12996 3204 13001 3209 sw
tri 13104 3204 13109 3209 ne
rect 13109 3204 13127 3209
tri 13127 3204 13167 3244 sw
tri 13780 3204 13820 3244 se
rect 13820 3204 13953 3244
rect 12064 3203 13001 3204
rect 12064 3151 12100 3203
rect 12152 3151 12169 3203
rect 12221 3151 12238 3203
rect 12290 3151 12307 3203
rect 12359 3151 12376 3203
rect 12428 3151 12445 3203
rect 12497 3151 12514 3203
rect 12566 3151 12583 3203
rect 12635 3151 12651 3203
rect 12703 3151 12719 3203
rect 12771 3151 12787 3203
rect 12839 3151 12855 3203
rect 12907 3201 13001 3203
tri 13001 3201 13004 3204 sw
tri 13109 3201 13112 3204 ne
rect 13112 3201 13167 3204
tri 13167 3201 13170 3204 sw
tri 13777 3201 13780 3204 se
rect 13780 3201 13875 3204
rect 12907 3151 13004 3201
rect 12064 3149 13004 3151
tri 13004 3149 13056 3201 sw
tri 13112 3149 13164 3201 ne
rect 13164 3149 13443 3201
rect 13495 3149 13507 3201
rect 13559 3149 13565 3201
tri 13728 3152 13777 3201 se
rect 13777 3152 13875 3201
rect 13927 3152 13953 3204
tri 13725 3149 13728 3152 se
rect 13728 3149 13953 3152
rect 12064 3124 13056 3149
tri 13056 3124 13081 3149 sw
tri 13700 3124 13725 3149 se
rect 13725 3124 13953 3149
rect 12064 3115 13081 3124
rect 12064 3063 12100 3115
rect 12152 3063 12169 3115
rect 12221 3063 12238 3115
rect 12290 3063 12307 3115
rect 12359 3063 12376 3115
rect 12428 3063 12445 3115
rect 12497 3063 12514 3115
rect 12566 3063 12583 3115
rect 12635 3063 12651 3115
rect 12703 3063 12719 3115
rect 12771 3063 12787 3115
rect 12839 3063 12855 3115
rect 12907 3112 13081 3115
tri 13081 3112 13093 3124 sw
tri 13648 3112 13660 3124 se
rect 13660 3112 13953 3124
rect 12907 3101 13093 3112
tri 13093 3101 13104 3112 sw
tri 13637 3101 13648 3112 se
rect 13648 3101 13875 3112
rect 12907 3063 13875 3101
rect 12064 3060 13875 3063
rect 13927 3060 13953 3112
rect 14011 3152 14017 3204
rect 14069 3152 14081 3204
rect 14133 3152 14139 3204
rect 12064 3017 13953 3060
tri 13984 3077 14011 3104 se
rect 14011 3077 14056 3152
tri 14056 3118 14090 3152 nw
rect 13984 3069 14056 3077
rect 13984 3059 14046 3069
tri 14046 3059 14056 3069 nw
rect 12064 2995 13681 3017
tri 13681 2995 13703 3017 nw
rect 12064 2977 13039 2995
tri 13039 2977 13057 2995 nw
rect 12064 2975 13035 2977
rect 12064 2919 12073 2975
rect 12129 2919 12198 2975
rect 12254 2919 12323 2975
rect 12379 2919 12448 2975
rect 12504 2919 12573 2975
rect 12629 2919 12698 2975
rect 12754 2919 12823 2975
rect 12879 2973 13035 2975
tri 13035 2973 13039 2977 nw
rect 12879 2919 12888 2973
rect 12064 2869 12888 2919
rect 12064 2813 12073 2869
rect 12129 2813 12198 2869
rect 12254 2813 12323 2869
rect 12379 2813 12448 2869
rect 12504 2813 12573 2869
rect 12629 2813 12698 2869
rect 12754 2813 12823 2869
rect 12879 2813 12888 2869
tri 12888 2826 13035 2973 nw
tri 13928 2826 13984 2882 se
rect 13984 2826 14030 3059
tri 14030 3043 14046 3059 nw
tri 14151 3043 14167 3059 se
rect 14167 3043 14195 3317
tri 14133 3025 14151 3043 se
rect 14151 3025 14195 3043
rect 14067 2973 14073 3025
rect 14125 2973 14137 3025
rect 14189 2973 14195 3025
rect 12064 2763 12888 2813
rect 12064 2707 12073 2763
rect 12129 2707 12198 2763
rect 12254 2707 12323 2763
rect 12379 2707 12448 2763
rect 12504 2707 12573 2763
rect 12629 2707 12698 2763
rect 12754 2707 12823 2763
rect 12879 2707 12888 2763
tri 13902 2800 13928 2826 se
rect 13928 2800 14030 2826
rect 12064 2657 12888 2707
rect 12960 2700 12969 2756
rect 13025 2700 13049 2756
rect 13105 2748 13579 2756
tri 13579 2748 13587 2756 sw
rect 13902 2748 13908 2800
rect 13960 2748 13972 2800
rect 14024 2748 14030 2800
rect 13105 2700 13587 2748
rect 12064 2601 12073 2657
rect 12129 2601 12198 2657
rect 12254 2601 12323 2657
rect 12379 2601 12448 2657
rect 12504 2601 12573 2657
rect 12629 2601 12698 2657
rect 12754 2601 12823 2657
rect 12879 2601 12888 2657
tri 13493 2622 13571 2700 ne
rect 13571 2622 13587 2700
tri 13587 2622 13713 2748 sw
tri 13571 2614 13579 2622 ne
rect 13579 2614 13722 2622
rect 12064 2551 12888 2601
tri 13579 2570 13623 2614 ne
rect 13623 2570 13722 2614
rect 13774 2570 13786 2622
rect 13838 2570 13850 2622
rect 13902 2570 13915 2622
rect 13967 2570 13973 2622
tri 11859 2506 11872 2519 ne
rect 11872 2506 11897 2519
tri 11897 2506 11926 2535 sw
tri 8912 2481 8921 2490 ne
rect 8921 2481 8946 2490
tri 8921 2456 8946 2481 ne
rect 8974 2481 8999 2490
tri 8999 2481 9008 2490 nw
tri 8974 2456 8999 2481 nw
rect 11552 2448 11553 2500
rect 11605 2448 11623 2500
rect 11675 2448 11693 2500
rect 11745 2448 11746 2500
tri 11872 2481 11897 2506 ne
rect 11897 2481 11926 2506
tri 11897 2452 11926 2481 ne
tri 11926 2463 11969 2506 sw
rect 12064 2495 12073 2551
rect 12129 2495 12198 2551
rect 12254 2495 12323 2551
rect 12379 2495 12448 2551
rect 12504 2495 12573 2551
rect 12629 2495 12698 2551
rect 12754 2495 12823 2551
rect 12879 2495 12888 2551
rect 12064 2493 12888 2495
rect 11926 2452 11969 2463
tri 11969 2452 11980 2463 sw
rect 13105 2458 13463 2463
rect 11552 2434 11746 2448
tri 9222 2398 9227 2403 sw
rect 9222 2382 9227 2398
tri 9227 2382 9243 2398 sw
rect 11552 2382 11553 2434
rect 11605 2382 11623 2434
rect 11675 2382 11693 2434
rect 11745 2382 11746 2434
tri 11926 2398 11980 2452 ne
tri 11980 2398 12034 2452 sw
rect 13105 2402 13114 2458
rect 13170 2402 13194 2458
rect 13250 2402 13463 2458
rect 13105 2398 13463 2402
rect 9222 2379 9243 2382
tri 9243 2379 9246 2382 sw
rect 11552 2376 11746 2382
tri 11980 2376 12002 2398 ne
rect 12002 2382 12034 2398
tri 12034 2382 12050 2398 sw
tri 13402 2382 13418 2398 ne
rect 13418 2382 13463 2398
tri 13463 2382 13544 2463 sw
rect 12002 2376 12050 2382
tri 12002 2351 12027 2376 ne
rect 12027 2351 12050 2376
tri 9662 2344 9669 2351 ne
rect 9669 2344 9696 2351
tri 12027 2344 12034 2351 ne
rect 12034 2344 12050 2351
tri 12050 2344 12088 2382 sw
tri 13418 2344 13456 2382 ne
rect 13456 2344 13544 2382
tri 9669 2323 9690 2344 ne
rect 9690 2323 9696 2344
rect 7595 2300 7862 2323
tri 9426 2317 9432 2323 se
rect 9432 2317 9645 2323
tri 9690 2317 9696 2323 ne
tri 12034 2317 12061 2344 ne
rect 12061 2337 13337 2344
tri 13337 2337 13344 2344 sw
tri 13456 2337 13463 2344 ne
rect 13463 2337 13544 2344
rect 12061 2317 13344 2337
tri 9422 2313 9426 2317 se
rect 9426 2313 9645 2317
tri 9415 2306 9422 2313 se
rect 9422 2306 9496 2313
tri 9409 2300 9415 2306 se
rect 9415 2300 9496 2306
rect 7595 2248 7601 2300
rect 7653 2299 7703 2300
rect 7755 2299 7804 2300
rect 7595 2243 7609 2248
rect 7665 2243 7701 2299
rect 7757 2243 7792 2299
rect 7856 2248 7862 2300
tri 9399 2290 9409 2300 se
rect 9409 2290 9496 2300
tri 9393 2284 9399 2290 se
rect 9399 2284 9496 2290
rect 9090 2278 9496 2284
rect 7848 2243 7862 2248
tri 8927 2246 8946 2265 se
rect 7595 2225 7862 2243
tri 8907 2226 8927 2246 se
rect 8927 2226 8946 2246
tri 8906 2225 8907 2226 se
rect 8907 2225 8946 2226
tri 8899 2218 8906 2225 se
rect 8906 2218 8946 2225
tri 8974 2246 8980 2252 sw
rect 8974 2226 8980 2246
tri 8980 2226 9000 2246 sw
rect 9090 2226 9091 2278
rect 9143 2275 9159 2278
rect 9211 2275 9227 2278
rect 9279 2275 9496 2278
rect 9151 2226 9159 2275
rect 9311 2261 9496 2275
rect 9548 2261 9582 2313
rect 9634 2261 9645 2313
tri 12061 2306 12072 2317 ne
rect 12072 2306 13344 2317
tri 13321 2300 13327 2306 ne
rect 13327 2300 13344 2306
tri 13344 2300 13381 2337 sw
tri 13463 2300 13500 2337 ne
rect 13500 2300 13544 2337
tri 13327 2290 13337 2300 ne
rect 13337 2290 13381 2300
rect 9311 2249 9645 2261
rect 8974 2218 9000 2226
tri 9000 2218 9008 2226 sw
rect 9090 2219 9095 2226
rect 9151 2219 9175 2226
rect 9231 2219 9255 2226
rect 9311 2219 9496 2249
rect 9090 2197 9496 2219
rect 9548 2197 9582 2249
rect 9634 2197 9645 2249
tri 13337 2246 13381 2290 ne
tri 13381 2256 13425 2300 sw
tri 13500 2256 13544 2300 ne
tri 13544 2256 13670 2382 sw
rect 13381 2246 13425 2256
tri 13425 2246 13435 2256 sw
tri 13544 2246 13554 2256 ne
rect 13554 2246 13670 2256
rect 9090 2193 9645 2197
rect 9090 2141 9091 2193
rect 9151 2141 9159 2193
rect 9090 2137 9095 2141
rect 9151 2137 9175 2141
rect 9231 2137 9255 2141
rect 9311 2137 9645 2193
tri 13381 2192 13435 2246 ne
tri 13435 2192 13489 2246 sw
tri 13554 2192 13608 2246 ne
rect 13608 2192 13670 2246
tri 13435 2159 13468 2192 ne
rect 13468 2159 13489 2192
rect 9090 2128 9645 2137
tri 9724 2138 9745 2159 sw
tri 13468 2138 13489 2159 ne
tri 13489 2138 13543 2192 sw
tri 13608 2138 13662 2192 ne
rect 13662 2138 13670 2192
tri 9692 2128 9697 2133 se
rect 9090 2125 9514 2128
tri 9514 2125 9517 2128 nw
tri 9689 2125 9692 2128 se
rect 9692 2125 9697 2128
rect 9724 2125 9745 2138
tri 9745 2125 9758 2138 sw
tri 13489 2125 13502 2138 ne
rect 13502 2130 13543 2138
tri 13543 2130 13551 2138 sw
tri 13662 2130 13670 2138 ne
tri 13670 2130 13796 2256 sw
rect 13502 2125 13551 2130
rect 9090 2110 9490 2125
rect 9090 2107 9095 2110
rect 9151 2107 9175 2110
rect 9231 2107 9255 2110
tri 5703 2055 5723 2075 sw
rect 9090 2055 9091 2107
rect 9151 2055 9159 2107
rect 9311 2101 9490 2110
tri 9490 2101 9514 2125 nw
tri 13502 2101 13526 2125 ne
rect 13526 2107 13551 2125
tri 13551 2107 13574 2130 sw
tri 13670 2107 13693 2130 ne
rect 13693 2107 13796 2130
rect 13526 2101 13597 2107
rect 9311 2084 9473 2101
tri 9473 2084 9490 2101 nw
tri 13526 2084 13543 2101 ne
rect 13543 2084 13545 2101
rect 9311 2082 9471 2084
tri 9471 2082 9473 2084 nw
tri 13543 2082 13545 2084 ne
rect 5703 2052 5723 2055
tri 5723 2052 5726 2055 sw
rect 9090 2054 9095 2055
rect 9151 2054 9175 2055
rect 9231 2054 9255 2055
rect 9311 2054 9441 2082
rect 9090 2052 9441 2054
tri 9441 2052 9471 2082 nw
rect 5703 2051 5726 2052
tri 5726 2051 5727 2052 sw
rect 9090 2051 9440 2052
tri 9440 2051 9441 2052 nw
rect 5703 2049 5727 2051
tri 5727 2049 5729 2051 sw
rect 9090 2049 9438 2051
tri 9438 2049 9440 2051 nw
tri 13693 2094 13706 2107 ne
rect 5703 2045 5729 2049
tri 5729 2045 5733 2049 sw
tri 9090 2045 9094 2049 ne
rect 9094 2046 9435 2049
tri 9435 2046 9438 2049 nw
rect 9094 2045 9311 2046
tri 9311 2045 9312 2046 nw
rect 5703 2041 5733 2045
tri 5733 2041 5737 2045 sw
rect 13545 2037 13597 2049
tri 5872 1985 5876 1989 ne
rect 5876 1985 5906 1989
tri 5876 1955 5906 1985 ne
rect 13545 1979 13597 1985
tri 5726 1830 5732 1836 ne
rect 5732 1830 5752 1836
tri 5732 1810 5752 1830 ne
rect 5802 1830 5830 1836
tri 5830 1830 5836 1836 nw
rect 5802 1810 5810 1830
tri 5810 1810 5830 1830 nw
tri 8600 1810 8620 1830 ne
rect 8620 1810 8634 1830
tri 5802 1802 5810 1810 nw
tri 8620 1802 8628 1810 ne
rect 8628 1802 8634 1810
tri 8628 1796 8634 1802 ne
tri 7744 1755 7778 1789 ne
rect 12709 1687 12764 1702
rect 12709 1681 12768 1687
tri 12722 1635 12768 1681 ne
tri 5514 1589 5543 1618 sw
rect 5462 1537 5468 1589
rect 5520 1537 5532 1589
rect 5584 1537 5590 1589
tri 5422 1502 5446 1526 sw
rect 5394 1496 5446 1502
tri 7830 1505 7851 1526 sw
rect 7830 1492 7851 1505
tri 7851 1492 7864 1505 sw
tri 8686 1499 8692 1505 sw
rect 8686 1471 8692 1499
tri 8692 1471 8720 1499 sw
tri 8769 1471 8797 1499 se
tri 10924 1471 10950 1497 se
rect 10950 1471 12172 1497
tri 12172 1471 12198 1497 sw
rect 5394 1430 5446 1444
tri 10872 1419 10924 1471 se
rect 10924 1419 12198 1471
tri 12198 1419 12250 1471 sw
tri 8763 1385 8797 1419 ne
tri 10838 1385 10872 1419 se
rect 10872 1385 12250 1419
tri 12250 1385 12284 1419 sw
rect 5394 1372 5446 1378
tri 10825 1372 10838 1385 se
rect 10838 1372 12284 1385
tri 12284 1372 12297 1385 sw
tri 10817 1364 10825 1372 se
rect 10825 1364 12297 1372
tri 12297 1364 12305 1372 sw
tri 10814 1361 10817 1364 se
rect 10817 1361 12305 1364
tri 12305 1361 12308 1364 sw
tri 10792 1339 10814 1361 se
rect 10814 1348 12308 1361
rect 10814 1339 11153 1348
tri 11153 1339 11162 1348 nw
tri 12089 1339 12098 1348 ne
rect 12098 1339 12308 1348
tri 12308 1339 12330 1361 sw
rect 7595 1296 7604 1300
rect 7660 1296 7701 1300
rect 7757 1296 7797 1300
rect 7853 1296 7862 1300
rect 7595 1244 7601 1296
rect 7660 1244 7669 1296
rect 7789 1244 7797 1296
rect 7856 1244 7862 1296
rect 9771 1287 9777 1339
rect 9829 1287 9842 1339
rect 9771 1275 9842 1287
rect 9771 1223 9777 1275
rect 9829 1223 9842 1275
rect 9771 1211 9842 1223
rect 9771 1159 9777 1211
rect 9829 1159 9842 1211
rect 10086 1338 11152 1339
tri 11152 1338 11153 1339 nw
tri 12098 1338 12099 1339 ne
rect 12099 1338 12717 1339
rect 10086 1286 11100 1338
tri 11100 1286 11152 1338 nw
tri 12099 1286 12151 1338 ne
rect 12151 1286 12509 1338
rect 12561 1286 12584 1338
rect 12636 1286 12659 1338
rect 12711 1286 12717 1338
rect 10086 1270 11084 1286
tri 11084 1270 11100 1286 nw
tri 12151 1270 12167 1286 ne
rect 12167 1270 12717 1286
rect 10086 1218 11032 1270
tri 11032 1218 11084 1270 nw
tri 12167 1265 12172 1270 ne
rect 12172 1265 12509 1270
tri 12172 1218 12219 1265 ne
rect 12219 1218 12509 1265
rect 12561 1218 12584 1270
rect 12636 1218 12659 1270
rect 12711 1218 12717 1270
rect 10086 1202 11016 1218
tri 11016 1202 11032 1218 nw
tri 12219 1202 12235 1218 ne
rect 12235 1202 12717 1218
rect 10086 1159 10973 1202
tri 10973 1159 11016 1202 nw
tri 12235 1159 12278 1202 ne
rect 12278 1159 12509 1202
tri 12278 1150 12287 1159 ne
rect 12287 1150 12509 1159
rect 12561 1150 12584 1202
rect 12636 1150 12659 1202
rect 12711 1150 12717 1202
tri 12287 1134 12303 1150 ne
rect 12303 1134 12717 1150
tri 12303 1087 12350 1134 ne
rect 12350 1087 12509 1134
tri 5901 1082 5906 1087 se
tri 12350 1082 12355 1087 ne
rect 12355 1082 12509 1087
rect 12561 1082 12584 1134
rect 12636 1082 12659 1134
rect 12711 1082 12717 1134
rect 13021 1239 13333 1245
rect 13073 1187 13281 1239
rect 13021 1175 13333 1187
rect 13073 1123 13281 1175
rect 13021 1117 13333 1123
rect 13706 1173 13796 2107
rect 13706 1121 13725 1173
rect 13777 1121 13796 1173
tri 5900 1081 5901 1082 se
rect 5901 1081 5906 1082
tri 5880 1061 5900 1081 se
rect 5900 1061 5906 1081
tri 12748 1061 12768 1081 se
tri 5872 1053 5880 1061 se
rect 5880 1053 5906 1061
tri 12740 1053 12748 1061 se
rect 12748 1053 12768 1061
tri 12734 1047 12740 1053 se
rect 12740 1047 12768 1053
rect 13706 1061 13796 1121
rect 13706 1009 13725 1061
rect 13777 1009 13796 1061
tri 5872 967 5906 1001 ne
rect 13706 948 13796 1009
rect 13706 896 13725 948
rect 13777 896 13796 948
rect 6974 835 6999 844
tri 6999 835 7008 844 nw
rect 13706 835 13796 896
tri 6974 810 6999 835 nw
tri 6810 783 6814 787 ne
rect 6814 783 6844 787
tri 6814 753 6844 783 ne
rect 6865 783 6897 787
tri 6897 783 6901 787 nw
rect 13706 783 13725 835
rect 13777 783 13796 835
rect 6865 753 6867 783
tri 6867 753 6897 783 nw
tri 6865 751 6867 753 nw
tri 6587 722 6612 747 ne
rect 6612 722 6621 747
tri 6612 713 6621 722 ne
rect 13706 722 13796 783
tri 7150 692 7163 705 sw
rect 7150 686 7163 692
tri 7163 686 7169 692 sw
tri 7554 686 7560 692 se
rect 7150 685 7169 686
tri 7169 685 7170 686 sw
rect 13706 670 13725 722
rect 13777 670 13796 722
tri 7547 640 7560 653 ne
rect 11304 621 11356 627
rect 7132 591 7147 598
tri 7147 591 7154 598 nw
tri 7132 576 7147 591 nw
rect 11304 557 11356 569
rect 13706 609 13796 670
rect 13706 557 13725 609
rect 13777 557 13796 609
rect 13706 521 13796 557
tri 10036 428 10064 456 sw
tri 10846 428 10873 455 sw
tri 9974 390 10012 428 se
rect 10036 390 10064 428
tri 10064 390 10102 428 sw
rect 10846 421 10873 428
tri 10873 421 10880 428 sw
tri 4401 361 4407 367 se
tri -399 351 -389 361 ne
rect -361 351 -357 361
tri -357 351 -347 361 nw
tri 4392 352 4401 361 se
rect 4401 352 4407 361
tri 4391 351 4392 352 se
rect 4392 351 4407 352
tri -361 347 -357 351 nw
tri 4387 347 4391 351 se
rect 4391 347 4407 351
tri 4378 338 4387 347 se
rect 4387 338 4407 347
tri 4374 334 4378 338 se
rect 4378 334 4407 338
tri 4373 333 4374 334 se
rect 4374 333 4407 334
tri 8515 378 8527 390 se
rect 8527 378 8528 390
tri 11116 361 11123 368 se
tri 11107 352 11116 361 se
rect 11116 352 11123 361
tri 8513 347 8518 352 ne
rect 8518 347 8527 352
tri 8518 338 8527 347 ne
tri 11093 338 11107 352 se
rect 11107 338 11123 352
tri 11089 334 11093 338 se
rect 11093 334 11123 338
rect 4562 322 4614 334
tri 3766 277 3800 311 se
tri 3823 277 3857 311 sw
tri 7636 277 7649 290 ne
rect 7649 277 7662 290
rect 4562 264 4614 270
tri 7649 266 7660 277 ne
rect 7660 266 7662 277
rect 9598 257 9604 309
rect 9656 257 9668 309
rect 9720 257 10369 309
rect 10360 253 10369 257
rect 10425 253 10449 309
rect 10505 253 10514 309
tri 10636 262 10638 264 ne
rect 10638 262 10670 264
tri 10638 253 10647 262 ne
rect 10647 253 10670 262
tri 10647 251 10649 253 ne
rect 10649 251 10670 253
tri 10649 242 10658 251 ne
rect 10658 242 10670 251
tri 10658 230 10670 242 ne
tri 10722 242 10731 251 sw
rect 10722 230 10731 242
tri 10731 230 10743 242 sw
rect 10722 217 10743 230
tri 10743 217 10756 230 sw
rect 7595 -43 7602 9
rect 7595 -47 7604 -43
rect 7660 -47 7701 9
rect 7757 -47 7797 9
rect 7855 -43 7862 9
rect 7853 -47 7862 -43
rect 7595 -55 7862 -47
rect 7595 -107 7602 -55
rect 7654 -71 7703 -55
rect 7755 -71 7803 -55
rect 7595 -127 7604 -107
rect 7660 -127 7701 -71
rect 7757 -127 7797 -71
rect 7855 -107 7862 -55
rect 7853 -127 7862 -107
tri 11223 -127 11304 -46 se
rect 11304 -102 11356 505
tri 11196 -154 11223 -127 se
rect 11223 -154 11304 -127
tri 11304 -154 11356 -102 nw
rect 12966 267 13439 314
rect 12966 211 12970 267
rect 13026 211 13066 267
rect 13122 211 13162 267
rect 13218 211 13258 267
rect 13314 262 13439 267
rect 13491 262 13508 314
rect 13560 262 13577 314
rect 13629 262 13646 314
rect 13698 262 13714 314
rect 13766 262 13782 314
rect 13834 262 13850 314
rect 13902 262 13918 314
rect 13970 262 14008 314
rect 13314 242 14008 262
rect 13314 211 13439 242
rect 12966 190 13439 211
rect 13491 190 13508 242
rect 13560 190 13577 242
rect 13629 190 13646 242
rect 13698 190 13714 242
rect 13766 190 13782 242
rect 13834 190 13850 242
rect 13902 190 13918 242
rect 13970 190 14008 242
rect 12966 183 14008 190
rect 12966 127 12970 183
rect 13026 127 13066 183
rect 13122 127 13162 183
rect 13218 127 13258 183
rect 13314 170 14008 183
rect 13314 127 13439 170
rect 12966 118 13439 127
rect 13491 118 13508 170
rect 13560 118 13577 170
rect 13629 118 13646 170
rect 13698 118 13714 170
rect 13766 118 13782 170
rect 13834 118 13850 170
rect 13902 118 13918 170
rect 13970 118 14008 170
rect 12966 99 14008 118
rect 12966 43 12970 99
rect 13026 43 13066 99
rect 13122 43 13162 99
rect 13218 43 13258 99
rect 13314 43 14008 99
rect 12966 15 14008 43
rect 12966 -41 12970 15
rect 13026 -41 13066 15
rect 13122 -41 13162 15
rect 13218 -41 13258 15
rect 13314 -41 14008 15
rect 12966 -69 14008 -41
rect 12966 -125 12970 -69
rect 13026 -125 13066 -69
rect 13122 -125 13162 -69
rect 13218 -125 13258 -69
rect 13314 -125 14008 -69
rect 12966 -154 14008 -125
tri 11189 -161 11196 -154 se
rect 11196 -161 11297 -154
tri 11297 -161 11304 -154 nw
tri 8880 -219 8938 -161 se
rect 8938 -213 11245 -161
tri 11245 -213 11297 -161 nw
rect 12966 -210 12970 -154
rect 13026 -210 13066 -154
rect 13122 -210 13162 -154
rect 13218 -210 13258 -154
rect 13314 -210 14008 -154
rect 8938 -219 8954 -213
tri 8954 -219 8960 -213 nw
rect 12966 -219 14008 -210
tri 8864 -235 8880 -219 se
rect 8880 -235 8938 -219
tri 8938 -235 8954 -219 nw
tri 8861 -238 8864 -235 se
rect 8864 -238 8935 -235
tri 8935 -238 8938 -235 nw
rect 8861 -399 8913 -238
tri 8913 -260 8935 -238 nw
tri 8913 -399 8928 -384 sw
tri 464 -403 468 -399 sw
tri 426 -413 436 -403 se
rect 464 -413 468 -403
tri 468 -413 478 -403 sw
rect 8861 -406 8928 -399
tri 8928 -406 8935 -399 sw
tri 8861 -413 8868 -406 ne
rect 8868 -413 8935 -406
tri 8868 -426 8881 -413 ne
rect 8881 -426 8935 -413
tri -176 -448 -154 -426 se
tri 8881 -448 8903 -426 ne
rect 8903 -448 8935 -426
tri 8903 -480 8935 -448 ne
tri 8935 -480 9009 -406 sw
tri 8935 -502 8957 -480 ne
tri 8883 -2183 8957 -2109 se
rect 8957 -2131 9009 -480
tri 8957 -2183 9009 -2131 nw
tri 8809 -2257 8883 -2183 se
tri 8883 -2257 8957 -2183 nw
tri 8711 -2355 8809 -2257 se
rect 8809 -2355 8839 -2257
tri 8839 -2301 8883 -2257 nw
rect 8711 -2381 8839 -2355
rect 8711 -2433 8717 -2381
rect 8769 -2433 8781 -2381
rect 8833 -2433 8839 -2381
rect 14822 -10026 14874 -8127
rect 14822 -10090 14874 -10078
rect 14822 -10148 14874 -10142
<< via2 >>
rect 1129 8813 1185 8869
rect 1129 8733 1185 8789
rect 1295 8543 1340 8593
rect 1340 8543 1351 8593
rect 1377 8543 1404 8593
rect 1404 8543 1416 8593
rect 1416 8543 1433 8593
rect 1459 8543 1468 8593
rect 1468 8543 1480 8593
rect 1480 8543 1515 8593
rect 1541 8543 1544 8593
rect 1544 8543 1596 8593
rect 1596 8543 1597 8593
rect 1295 8537 1351 8543
rect 1377 8537 1433 8543
rect 1459 8537 1515 8543
rect 1541 8537 1597 8543
rect 1295 8453 1351 8509
rect 1377 8453 1433 8509
rect 1459 8453 1515 8509
rect 1541 8453 1597 8509
rect 1295 8369 1351 8425
rect 1377 8369 1433 8425
rect 1459 8369 1515 8425
rect 1541 8369 1597 8425
rect 1295 8324 1351 8341
rect 1377 8324 1433 8341
rect 1459 8324 1515 8341
rect 1541 8324 1597 8341
rect 1295 8285 1340 8324
rect 1340 8285 1351 8324
rect 1377 8285 1404 8324
rect 1404 8285 1416 8324
rect 1416 8285 1433 8324
rect 1459 8285 1468 8324
rect 1468 8285 1480 8324
rect 1480 8285 1515 8324
rect 1541 8285 1544 8324
rect 1544 8285 1596 8324
rect 1596 8285 1597 8324
rect 1295 8201 1351 8257
rect 1377 8201 1433 8257
rect 1459 8201 1515 8257
rect 1541 8201 1597 8257
rect 1295 8117 1351 8173
rect 1377 8117 1433 8173
rect 1459 8117 1515 8173
rect 1541 8117 1597 8173
rect 4814 8127 4870 8183
rect 4894 8127 4950 8183
rect 4974 8134 5007 8183
rect 5007 8134 5030 8183
rect 4974 8127 5030 8134
rect 1295 8033 1351 8089
rect 1377 8033 1433 8089
rect 1459 8033 1515 8089
rect 1541 8033 1597 8089
rect 1295 7964 1340 8005
rect 1340 7964 1351 8005
rect 1377 7964 1404 8005
rect 1404 7964 1416 8005
rect 1416 7964 1433 8005
rect 1459 7964 1468 8005
rect 1468 7964 1480 8005
rect 1480 7964 1515 8005
rect 1541 7964 1544 8005
rect 1544 7964 1596 8005
rect 1596 7964 1597 8005
rect 1295 7949 1351 7964
rect 1377 7949 1433 7964
rect 1459 7949 1515 7964
rect 1541 7949 1597 7964
rect 4814 8004 4870 8060
rect 4894 8004 4950 8060
rect 4974 8058 5007 8060
rect 5007 8058 5030 8060
rect 4974 8034 5030 8058
rect 4974 8004 5007 8034
rect 5007 8004 5030 8034
rect 1295 7865 1351 7921
rect 1377 7865 1433 7921
rect 1459 7865 1515 7921
rect 1541 7865 1597 7921
rect 1295 7781 1351 7837
rect 1377 7781 1433 7837
rect 1459 7781 1515 7837
rect 1541 7781 1597 7837
rect 1295 7701 1351 7753
rect 1377 7701 1433 7753
rect 1459 7701 1515 7753
rect 1541 7701 1597 7753
rect 1295 7697 1340 7701
rect 1340 7697 1351 7701
rect 1377 7697 1404 7701
rect 1404 7697 1416 7701
rect 1416 7697 1433 7701
rect 1459 7697 1468 7701
rect 1468 7697 1480 7701
rect 1480 7697 1515 7701
rect 1541 7697 1544 7701
rect 1544 7697 1596 7701
rect 1596 7697 1597 7701
rect 4814 7881 4870 7937
rect 4894 7881 4950 7937
rect 4974 7906 5007 7937
rect 5007 7906 5030 7937
rect 4974 7882 5030 7906
rect 4974 7881 5007 7882
rect 5007 7881 5030 7882
rect 4814 7757 4870 7813
rect 4894 7757 4950 7813
rect 4974 7806 5030 7813
rect 4974 7757 5007 7806
rect 5007 7757 5030 7806
rect 6479 7781 6535 7837
rect 6561 7781 6617 7837
rect 6643 7781 6699 7837
rect 6725 7781 6781 7837
rect 6807 7781 6863 7837
rect 6888 7781 6944 7837
rect 6969 7781 7025 7837
rect 7050 7781 7106 7837
rect 7131 7781 7187 7837
rect 7212 7781 7268 7837
rect 7293 7781 7349 7837
rect 7374 7781 7430 7837
rect 7455 7781 7511 7837
rect 7536 7781 7592 7837
rect 7617 7781 7673 7837
rect 7698 7781 7754 7837
rect 7779 7781 7835 7837
rect 7860 7781 7916 7837
rect 7941 7781 7997 7837
rect 8022 7781 8078 7837
rect 8103 7781 8159 7837
rect 8184 7781 8240 7837
rect 8265 7781 8321 7837
rect 8346 7781 8402 7837
rect 8427 7781 8483 7837
rect 8508 7781 8564 7837
rect 8589 7781 8645 7837
rect 8670 7781 8726 7837
rect 8751 7781 8807 7837
rect 8832 7781 8888 7837
rect 8913 7781 8969 7837
rect 8994 7781 9050 7837
rect 9075 7781 9131 7837
rect 9156 7781 9212 7837
rect 9237 7781 9293 7837
rect 9318 7781 9374 7837
rect 9399 7781 9455 7837
rect 9480 7781 9536 7837
rect 9561 7781 9617 7837
rect 9642 7781 9698 7837
rect 1295 7649 1340 7669
rect 1340 7649 1351 7669
rect 1377 7649 1404 7669
rect 1404 7649 1416 7669
rect 1416 7649 1433 7669
rect 1459 7649 1468 7669
rect 1468 7649 1480 7669
rect 1480 7649 1515 7669
rect 1541 7649 1544 7669
rect 1544 7649 1596 7669
rect 1596 7649 1597 7669
rect 1295 7613 1351 7649
rect 1377 7613 1433 7649
rect 1459 7613 1515 7649
rect 1541 7613 1597 7649
rect 1295 7529 1351 7585
rect 1377 7529 1433 7585
rect 1459 7529 1515 7585
rect 1541 7529 1597 7585
rect 6479 7687 6535 7743
rect 6561 7687 6617 7743
rect 6643 7687 6699 7743
rect 6725 7687 6781 7743
rect 6807 7687 6863 7743
rect 6888 7687 6944 7743
rect 6969 7687 7025 7743
rect 7050 7687 7106 7743
rect 7131 7687 7187 7743
rect 7212 7687 7268 7743
rect 7293 7687 7349 7743
rect 7374 7687 7430 7743
rect 7455 7687 7511 7743
rect 7536 7687 7592 7743
rect 7617 7687 7673 7743
rect 7698 7687 7754 7743
rect 7779 7687 7835 7743
rect 7860 7687 7916 7743
rect 7941 7687 7997 7743
rect 8022 7687 8078 7743
rect 8103 7687 8159 7743
rect 8184 7687 8240 7743
rect 8265 7687 8321 7743
rect 8346 7687 8402 7743
rect 8427 7687 8483 7743
rect 8508 7687 8564 7743
rect 8589 7687 8645 7743
rect 8670 7687 8726 7743
rect 8751 7687 8807 7743
rect 8832 7687 8888 7743
rect 8913 7687 8969 7743
rect 8994 7687 9050 7743
rect 9075 7687 9131 7743
rect 9156 7687 9212 7743
rect 9237 7687 9293 7743
rect 9318 7687 9374 7743
rect 9399 7687 9455 7743
rect 9480 7687 9536 7743
rect 9561 7687 9617 7743
rect 9642 7687 9698 7743
rect 6479 7593 6535 7649
rect 6561 7593 6617 7649
rect 6643 7593 6699 7649
rect 6725 7593 6781 7649
rect 6807 7593 6863 7649
rect 6888 7593 6944 7649
rect 6969 7593 7025 7649
rect 7050 7593 7106 7649
rect 7131 7593 7187 7649
rect 7212 7593 7268 7649
rect 7293 7593 7349 7649
rect 7374 7593 7430 7649
rect 7455 7593 7511 7649
rect 7536 7593 7592 7649
rect 7617 7593 7673 7649
rect 7698 7593 7754 7649
rect 7779 7593 7835 7649
rect 7860 7593 7916 7649
rect 7941 7593 7997 7649
rect 8022 7593 8078 7649
rect 8103 7593 8159 7649
rect 8184 7593 8240 7649
rect 8265 7593 8321 7649
rect 8346 7593 8402 7649
rect 8427 7593 8483 7649
rect 8508 7593 8564 7649
rect 8589 7593 8645 7649
rect 8670 7593 8726 7649
rect 8751 7593 8807 7649
rect 8832 7593 8888 7649
rect 8913 7593 8969 7649
rect 8994 7593 9050 7649
rect 9075 7593 9131 7649
rect 9156 7593 9212 7649
rect 9237 7593 9293 7649
rect 9318 7593 9374 7649
rect 9399 7593 9455 7649
rect 9480 7593 9536 7649
rect 9561 7593 9617 7649
rect 9642 7593 9698 7649
rect 1295 7445 1351 7501
rect 1377 7445 1433 7501
rect 1459 7445 1515 7501
rect 1541 7445 1597 7501
rect 6479 7499 6535 7555
rect 6561 7499 6617 7555
rect 6643 7499 6699 7555
rect 6725 7499 6781 7555
rect 6807 7499 6863 7555
rect 6888 7499 6944 7555
rect 6969 7499 7025 7555
rect 7050 7499 7106 7555
rect 7131 7499 7187 7555
rect 7212 7499 7268 7555
rect 7293 7499 7349 7555
rect 7374 7499 7430 7555
rect 7455 7499 7511 7555
rect 7536 7499 7592 7555
rect 7617 7499 7673 7555
rect 7698 7499 7754 7555
rect 7779 7499 7835 7555
rect 7860 7499 7916 7555
rect 7941 7499 7997 7555
rect 8022 7499 8078 7555
rect 8103 7499 8159 7555
rect 8184 7499 8240 7555
rect 8265 7499 8321 7555
rect 8346 7499 8402 7555
rect 8427 7499 8483 7555
rect 8508 7499 8564 7555
rect 8589 7499 8645 7555
rect 8670 7499 8726 7555
rect 8751 7499 8807 7555
rect 8832 7499 8888 7555
rect 8913 7499 8969 7555
rect 8994 7499 9050 7555
rect 9075 7499 9131 7555
rect 9156 7499 9212 7555
rect 9237 7499 9293 7555
rect 9318 7499 9374 7555
rect 9399 7499 9455 7555
rect 9480 7499 9536 7555
rect 9561 7499 9617 7555
rect 9642 7499 9698 7555
rect 1295 7389 1351 7417
rect 1377 7389 1433 7417
rect 1459 7389 1515 7417
rect 1541 7389 1597 7417
rect 1295 7361 1340 7389
rect 1340 7361 1351 7389
rect 1377 7361 1404 7389
rect 1404 7361 1416 7389
rect 1416 7361 1433 7389
rect 1459 7361 1468 7389
rect 1468 7361 1480 7389
rect 1480 7361 1515 7389
rect 1541 7361 1544 7389
rect 1544 7361 1596 7389
rect 1596 7361 1597 7389
rect 1295 7321 1351 7333
rect 1377 7321 1433 7333
rect 1459 7321 1515 7333
rect 1541 7321 1597 7333
rect 1295 7277 1336 7321
rect 1336 7277 1349 7321
rect 1349 7277 1351 7321
rect 1377 7277 1401 7321
rect 1401 7277 1414 7321
rect 1414 7277 1433 7321
rect 1459 7277 1466 7321
rect 1466 7277 1479 7321
rect 1479 7277 1515 7321
rect 1541 7277 1544 7321
rect 1544 7277 1596 7321
rect 1596 7277 1597 7321
rect 5164 7365 5220 7421
rect 5258 7365 5314 7421
rect 5352 7365 5408 7421
rect 1003 6989 1059 7045
rect 5164 7263 5220 7319
rect 5258 7263 5314 7319
rect 5352 7263 5408 7319
rect 8856 7305 8912 7361
rect 8947 7305 9003 7361
rect 9038 7305 9094 7361
rect 9129 7305 9185 7361
rect 9219 7305 9275 7361
rect 5164 7161 5220 7217
rect 5258 7161 5314 7217
rect 5352 7161 5408 7217
rect 5164 7059 5220 7115
rect 5258 7059 5314 7115
rect 5352 7059 5408 7115
rect 1003 6909 1059 6965
rect 5593 7218 5649 7274
rect 5673 7218 5729 7274
rect 5753 7218 5809 7274
rect 5833 7218 5889 7274
rect 5913 7218 5969 7274
rect 5593 7130 5649 7186
rect 5673 7130 5729 7186
rect 5753 7130 5809 7186
rect 5833 7130 5889 7186
rect 5913 7130 5969 7186
rect 8856 7169 8912 7225
rect 8947 7169 9003 7225
rect 9038 7169 9094 7225
rect 9129 7169 9185 7225
rect 9219 7169 9275 7225
rect 9403 7357 9459 7413
rect 9490 7357 9546 7413
rect 9577 7357 9633 7413
rect 9664 7357 9720 7413
rect 9750 7357 9806 7413
rect 9403 7265 9459 7321
rect 9490 7265 9546 7321
rect 9577 7265 9633 7321
rect 9664 7265 9720 7321
rect 9750 7265 9806 7321
rect 9403 7173 9459 7229
rect 9490 7173 9546 7229
rect 9577 7173 9633 7229
rect 9664 7173 9720 7229
rect 9750 7173 9806 7229
rect 5593 7041 5649 7097
rect 5673 7041 5729 7097
rect 5753 7041 5809 7097
rect 5833 7041 5889 7097
rect 5913 7041 5969 7097
rect 9403 7081 9459 7137
rect 9490 7081 9546 7137
rect 9577 7081 9633 7137
rect 9664 7081 9720 7137
rect 9750 7081 9806 7137
rect 5593 6952 5649 7008
rect 5673 6952 5729 7008
rect 5753 6952 5809 7008
rect 5833 6952 5889 7008
rect 5913 6952 5969 7008
rect 1801 6700 1857 6702
rect 1905 6700 1961 6702
rect 2008 6700 2064 6702
rect 2111 6700 2167 6702
rect 1801 6648 1837 6700
rect 1837 6648 1857 6700
rect 1905 6648 1957 6700
rect 1957 6648 1961 6700
rect 2008 6648 2025 6700
rect 2025 6648 2040 6700
rect 2040 6648 2064 6700
rect 2111 6648 2159 6700
rect 2159 6648 2167 6700
rect 1801 6646 1857 6648
rect 1905 6646 1961 6648
rect 2008 6646 2064 6648
rect 2111 6646 2167 6648
rect 2987 6499 3030 6546
rect 3030 6499 3043 6546
rect 3074 6499 3102 6546
rect 3102 6499 3122 6546
rect 3122 6499 3130 6546
rect 3161 6499 3174 6546
rect 3174 6499 3194 6546
rect 3194 6499 3217 6546
rect 3247 6499 3266 6546
rect 3266 6499 3303 6546
rect 2987 6490 3043 6499
rect 3074 6490 3130 6499
rect 3161 6490 3217 6499
rect 3247 6490 3303 6499
rect 2987 6427 3030 6456
rect 3030 6427 3043 6456
rect 3074 6427 3102 6456
rect 3102 6427 3122 6456
rect 3122 6427 3130 6456
rect 3161 6427 3174 6456
rect 3174 6427 3194 6456
rect 3194 6427 3217 6456
rect 3247 6427 3266 6456
rect 3266 6427 3303 6456
rect 2987 6407 3043 6427
rect 3074 6407 3130 6427
rect 3161 6407 3217 6427
rect 3247 6407 3303 6427
rect 2987 6400 3030 6407
rect 3030 6400 3043 6407
rect 3074 6400 3102 6407
rect 3102 6400 3122 6407
rect 3122 6400 3130 6407
rect 3161 6400 3174 6407
rect 3174 6400 3194 6407
rect 3194 6400 3217 6407
rect 3247 6400 3266 6407
rect 3266 6400 3303 6407
rect 2987 6355 3030 6366
rect 3030 6355 3043 6366
rect 3074 6355 3102 6366
rect 3102 6355 3122 6366
rect 3122 6355 3130 6366
rect 3161 6355 3174 6366
rect 3174 6355 3194 6366
rect 3194 6355 3217 6366
rect 3247 6355 3266 6366
rect 3266 6355 3303 6366
rect 2987 6335 3043 6355
rect 3074 6335 3130 6355
rect 3161 6335 3217 6355
rect 3247 6335 3303 6355
rect 2987 6310 3030 6335
rect 3030 6310 3043 6335
rect 3074 6310 3102 6335
rect 3102 6310 3122 6335
rect 3122 6310 3130 6335
rect 3161 6310 3174 6335
rect 3174 6310 3194 6335
rect 3194 6310 3217 6335
rect 3247 6310 3266 6335
rect 3266 6310 3303 6335
rect 2987 6263 3043 6276
rect 3074 6263 3130 6276
rect 3161 6263 3217 6276
rect 3247 6263 3303 6276
rect 2987 6220 3030 6263
rect 3030 6220 3043 6263
rect 3074 6220 3102 6263
rect 3102 6220 3122 6263
rect 3122 6220 3130 6263
rect 3161 6220 3174 6263
rect 3174 6220 3194 6263
rect 3194 6220 3217 6263
rect 3247 6220 3266 6263
rect 3266 6220 3303 6263
rect 8856 6619 8912 6675
rect 8947 6619 9003 6675
rect 9038 6619 9094 6675
rect 9129 6619 9185 6675
rect 9219 6619 9275 6675
rect 8856 6539 8912 6595
rect 8947 6539 9003 6595
rect 9038 6539 9094 6595
rect 9129 6539 9185 6595
rect 9219 6539 9275 6595
rect 8856 6459 8912 6515
rect 8947 6459 9003 6515
rect 9038 6459 9094 6515
rect 9129 6459 9185 6515
rect 9219 6459 9275 6515
rect 8856 6379 8912 6435
rect 8947 6379 9003 6435
rect 9038 6379 9094 6435
rect 9129 6379 9185 6435
rect 9219 6379 9275 6435
rect 5593 5975 5649 6031
rect 5673 5975 5729 6031
rect 5753 5975 5809 6031
rect 5833 5975 5889 6031
rect 5913 5975 5969 6031
rect 5164 5868 5220 5924
rect 5258 5868 5314 5924
rect 5352 5868 5408 5924
rect 5164 5766 5220 5822
rect 5258 5766 5314 5822
rect 5352 5766 5408 5822
rect 5164 5664 5220 5720
rect 5258 5664 5314 5720
rect 5352 5664 5408 5720
rect 2913 5470 3049 5606
rect 5164 5562 5220 5618
rect 5258 5562 5314 5618
rect 5352 5562 5408 5618
rect 5593 5873 5649 5929
rect 5673 5873 5729 5929
rect 5753 5873 5809 5929
rect 5833 5873 5889 5929
rect 5913 5873 5969 5929
rect 5593 5771 5649 5827
rect 5673 5771 5729 5827
rect 5753 5771 5809 5827
rect 5833 5771 5889 5827
rect 5913 5771 5969 5827
rect 9403 5783 9459 5839
rect 9489 5783 9545 5839
rect 9575 5783 9631 5839
rect 9661 5783 9717 5839
rect 9746 5783 9802 5839
rect 5593 5669 5649 5725
rect 5673 5669 5729 5725
rect 5753 5669 5809 5725
rect 5833 5669 5889 5725
rect 5913 5669 5969 5725
rect 9403 5679 9459 5735
rect 9489 5679 9545 5735
rect 9575 5679 9631 5735
rect 9661 5679 9717 5735
rect 9746 5679 9802 5735
rect 9403 5575 9459 5631
rect 9489 5575 9545 5631
rect 9575 5575 9631 5631
rect 9661 5575 9717 5631
rect 9746 5575 9802 5631
rect 7856 5355 7912 5411
rect 7937 5355 7993 5411
rect 8018 5355 8074 5411
rect 8099 5355 8155 5411
rect 8180 5355 8236 5411
rect 8261 5355 8317 5411
rect 8341 5355 8397 5411
rect 8421 5355 8477 5411
rect 8501 5355 8557 5411
rect 8581 5355 8637 5411
rect 8661 5355 8717 5411
rect 8741 5355 8797 5411
rect 8821 5355 8877 5411
rect 8901 5355 8957 5411
rect 8981 5355 9037 5411
rect 9061 5355 9117 5411
rect 9141 5355 9197 5411
rect 9221 5355 9277 5411
rect 9301 5355 9357 5411
rect 9381 5355 9437 5411
rect 9461 5355 9517 5411
rect 9541 5355 9597 5411
rect 9621 5355 9677 5411
rect 9701 5355 9757 5411
rect 9781 5355 9837 5411
rect 9861 5355 9917 5411
rect 9941 5355 9997 5411
rect 10021 5355 10077 5411
rect 10101 5355 10157 5411
rect 10181 5355 10237 5411
rect 10261 5355 10317 5411
rect 10341 5355 10397 5411
rect 10421 5355 10477 5411
rect 10501 5355 10557 5411
rect 10581 5355 10637 5411
rect 10661 5355 10717 5411
rect 10741 5355 10797 5411
rect 10821 5355 10877 5411
rect 10901 5355 10957 5411
rect 10981 5355 11037 5411
rect 11061 5355 11117 5411
rect 11141 5355 11197 5411
rect 7856 5261 7912 5317
rect 7937 5261 7993 5317
rect 8018 5261 8074 5317
rect 8099 5261 8155 5317
rect 8180 5261 8236 5317
rect 8261 5261 8317 5317
rect 8341 5261 8397 5317
rect 8421 5261 8477 5317
rect 8501 5261 8557 5317
rect 8581 5261 8637 5317
rect 8661 5261 8717 5317
rect 8741 5261 8797 5317
rect 8821 5261 8877 5317
rect 8901 5261 8957 5317
rect 8981 5261 9037 5317
rect 9061 5261 9117 5317
rect 9141 5261 9197 5317
rect 9221 5261 9277 5317
rect 9301 5261 9357 5317
rect 9381 5261 9437 5317
rect 9461 5261 9517 5317
rect 9541 5261 9597 5317
rect 9621 5261 9677 5317
rect 9701 5261 9757 5317
rect 9781 5261 9837 5317
rect 9861 5261 9917 5317
rect 9941 5261 9997 5317
rect 10021 5261 10077 5317
rect 10101 5261 10157 5317
rect 10181 5261 10237 5317
rect 10261 5261 10317 5317
rect 10341 5261 10397 5317
rect 10421 5261 10477 5317
rect 10501 5261 10557 5317
rect 10581 5261 10637 5317
rect 10661 5261 10717 5317
rect 10741 5261 10797 5317
rect 10821 5261 10877 5317
rect 10901 5261 10957 5317
rect 10981 5261 11037 5317
rect 11061 5261 11117 5317
rect 11141 5261 11197 5317
rect 7856 5167 7912 5223
rect 7937 5167 7993 5223
rect 8018 5167 8074 5223
rect 8099 5167 8155 5223
rect 8180 5167 8236 5223
rect 8261 5167 8317 5223
rect 8341 5167 8397 5223
rect 8421 5167 8477 5223
rect 8501 5167 8557 5223
rect 8581 5167 8637 5223
rect 8661 5167 8717 5223
rect 8741 5167 8797 5223
rect 8821 5167 8877 5223
rect 8901 5167 8957 5223
rect 8981 5167 9037 5223
rect 9061 5167 9117 5223
rect 9141 5167 9197 5223
rect 9221 5167 9277 5223
rect 9301 5167 9357 5223
rect 9381 5167 9437 5223
rect 9461 5167 9517 5223
rect 9541 5167 9597 5223
rect 9621 5167 9677 5223
rect 9701 5167 9757 5223
rect 9781 5167 9837 5223
rect 9861 5167 9917 5223
rect 9941 5167 9997 5223
rect 10021 5167 10077 5223
rect 10101 5167 10157 5223
rect 10181 5167 10237 5223
rect 10261 5167 10317 5223
rect 10341 5167 10397 5223
rect 10421 5167 10477 5223
rect 10501 5167 10557 5223
rect 10581 5167 10637 5223
rect 10661 5167 10717 5223
rect 10741 5167 10797 5223
rect 10821 5167 10877 5223
rect 10901 5167 10957 5223
rect 10981 5167 11037 5223
rect 11061 5167 11117 5223
rect 11141 5167 11197 5223
rect 2913 4587 2960 4635
rect 2960 4587 2969 4635
rect 2913 4579 2969 4587
rect 2993 4587 3002 4635
rect 3002 4587 3049 4635
rect 2993 4579 3049 4587
rect 2913 4521 2960 4554
rect 2960 4521 2969 4554
rect 2913 4506 2969 4521
rect 2913 4498 2960 4506
rect 2960 4498 2969 4506
rect 2993 4521 3002 4554
rect 3002 4521 3049 4554
rect 2993 4506 3049 4521
rect 2993 4498 3002 4506
rect 3002 4498 3049 4506
rect 3285 1936 3322 1983
rect 3322 1936 3388 1983
rect 3388 1936 3421 1983
rect 3285 1910 3421 1936
rect 3285 1858 3322 1910
rect 3322 1858 3388 1910
rect 3388 1858 3421 1910
rect 3285 1847 3421 1858
rect 7856 5073 7912 5129
rect 7937 5073 7993 5129
rect 8018 5073 8074 5129
rect 8099 5073 8155 5129
rect 8180 5073 8236 5129
rect 8261 5073 8317 5129
rect 8341 5073 8397 5129
rect 8421 5073 8477 5129
rect 8501 5073 8557 5129
rect 8581 5073 8637 5129
rect 8661 5073 8717 5129
rect 8741 5073 8797 5129
rect 8821 5073 8877 5129
rect 8901 5073 8957 5129
rect 8981 5073 9037 5129
rect 9061 5073 9117 5129
rect 9141 5073 9197 5129
rect 9221 5073 9277 5129
rect 9301 5073 9357 5129
rect 9381 5073 9437 5129
rect 9461 5073 9517 5129
rect 9541 5073 9597 5129
rect 9621 5073 9677 5129
rect 9701 5073 9757 5129
rect 9781 5073 9837 5129
rect 9861 5073 9917 5129
rect 9941 5073 9997 5129
rect 10021 5073 10077 5129
rect 10101 5073 10157 5129
rect 10181 5073 10237 5129
rect 10261 5073 10317 5129
rect 10341 5073 10397 5129
rect 10421 5073 10477 5129
rect 10501 5073 10557 5129
rect 10581 5073 10637 5129
rect 10661 5073 10717 5129
rect 10741 5073 10797 5129
rect 10821 5073 10877 5129
rect 10901 5073 10957 5129
rect 10981 5073 11037 5129
rect 11061 5073 11117 5129
rect 11141 5073 11197 5129
rect 4814 4988 4870 5044
rect 4894 4988 4950 5044
rect 4974 4995 5007 5044
rect 5007 4995 5030 5044
rect 4974 4988 5030 4995
rect 4814 4863 4870 4919
rect 4894 4863 4950 4919
rect 4974 4902 5030 4919
rect 4974 4863 5007 4902
rect 5007 4863 5030 4902
rect 4814 4737 4870 4793
rect 4894 4737 4950 4793
rect 4974 4777 5007 4793
rect 5007 4777 5030 4793
rect 4974 4756 5030 4777
rect 4974 4737 5007 4756
rect 5007 4737 5030 4756
rect 4814 4611 4870 4667
rect 4894 4611 4950 4667
rect 4974 4631 5007 4667
rect 5007 4631 5030 4667
rect 4974 4611 5030 4631
rect 4814 4485 4870 4541
rect 4894 4485 4950 4541
rect 4974 4537 5030 4541
rect 4974 4485 5007 4537
rect 5007 4485 5030 4537
rect 5924 4293 5980 4295
rect 5924 4241 5973 4293
rect 5973 4241 5980 4293
rect 5924 4239 5980 4241
rect 6023 4293 6079 4295
rect 6023 4241 6025 4293
rect 6025 4241 6077 4293
rect 6077 4241 6079 4293
rect 6023 4239 6079 4241
rect 6121 4293 6177 4295
rect 6121 4241 6128 4293
rect 6128 4241 6177 4293
rect 6121 4239 6177 4241
rect 9095 2986 9151 3040
rect 9175 2986 9231 3040
rect 9255 2986 9311 3040
rect 10356 2993 10412 3049
rect 10453 2993 10509 3049
rect 10550 2993 10606 3049
rect 10646 2993 10702 3049
rect 9095 2984 9104 2986
rect 9104 2984 9151 2986
rect 9175 2984 9184 2986
rect 9184 2984 9231 2986
rect 9255 2984 9263 2986
rect 9263 2984 9311 2986
rect 9095 2934 9104 2942
rect 9104 2934 9151 2942
rect 9175 2934 9184 2942
rect 9184 2934 9231 2942
rect 9255 2934 9263 2942
rect 9263 2934 9311 2942
rect 9095 2910 9151 2934
rect 9175 2910 9231 2934
rect 9255 2910 9311 2934
rect 9095 2886 9104 2910
rect 9104 2886 9151 2910
rect 9175 2886 9184 2910
rect 9184 2886 9231 2910
rect 9255 2886 9263 2910
rect 9263 2886 9311 2910
rect 10356 2889 10412 2945
rect 10453 2889 10509 2945
rect 10550 2889 10606 2945
rect 10646 2889 10702 2945
rect 9095 2834 9151 2844
rect 9175 2834 9231 2844
rect 9255 2834 9311 2844
rect 9095 2788 9104 2834
rect 9104 2788 9151 2834
rect 9175 2788 9184 2834
rect 9184 2788 9231 2834
rect 9255 2788 9263 2834
rect 9263 2788 9311 2834
rect 10356 2785 10412 2841
rect 10453 2785 10509 2841
rect 10550 2785 10606 2841
rect 10646 2785 10702 2841
rect 9095 2706 9104 2746
rect 9104 2706 9151 2746
rect 9175 2706 9184 2746
rect 9184 2706 9231 2746
rect 9255 2706 9263 2746
rect 9263 2706 9311 2746
rect 9095 2690 9151 2706
rect 9175 2690 9231 2706
rect 9255 2690 9311 2706
rect 10356 2681 10412 2737
rect 10453 2681 10509 2737
rect 10550 2681 10606 2737
rect 10646 2681 10702 2737
rect 12669 4043 12725 4099
rect 12759 4043 12815 4099
rect 12848 4043 12904 4099
rect 12073 2919 12129 2975
rect 12198 2919 12254 2975
rect 12323 2919 12379 2975
rect 12448 2919 12504 2975
rect 12573 2919 12629 2975
rect 12698 2919 12754 2975
rect 12823 2919 12879 2975
rect 12073 2813 12129 2869
rect 12198 2813 12254 2869
rect 12323 2813 12379 2869
rect 12448 2813 12504 2869
rect 12573 2813 12629 2869
rect 12698 2813 12754 2869
rect 12823 2813 12879 2869
rect 12073 2707 12129 2763
rect 12198 2707 12254 2763
rect 12323 2707 12379 2763
rect 12448 2707 12504 2763
rect 12573 2707 12629 2763
rect 12698 2707 12754 2763
rect 12823 2707 12879 2763
rect 12969 2700 13025 2756
rect 13049 2700 13105 2756
rect 12073 2601 12129 2657
rect 12198 2601 12254 2657
rect 12323 2601 12379 2657
rect 12448 2601 12504 2657
rect 12573 2601 12629 2657
rect 12698 2601 12754 2657
rect 12823 2601 12879 2657
rect 12073 2495 12129 2551
rect 12198 2495 12254 2551
rect 12323 2495 12379 2551
rect 12448 2495 12504 2551
rect 12573 2495 12629 2551
rect 12698 2495 12754 2551
rect 12823 2495 12879 2551
rect 13114 2402 13170 2458
rect 13194 2402 13250 2458
rect 7609 2248 7653 2299
rect 7653 2248 7665 2299
rect 7609 2243 7665 2248
rect 7701 2248 7703 2299
rect 7703 2248 7755 2299
rect 7755 2248 7757 2299
rect 7701 2243 7757 2248
rect 7792 2248 7804 2299
rect 7804 2248 7848 2299
rect 7792 2243 7848 2248
rect 9095 2226 9143 2275
rect 9143 2226 9151 2275
rect 9175 2226 9211 2275
rect 9211 2226 9227 2275
rect 9227 2226 9231 2275
rect 9255 2226 9279 2275
rect 9279 2226 9311 2275
rect 9095 2219 9151 2226
rect 9175 2219 9231 2226
rect 9255 2219 9311 2226
rect 9095 2141 9143 2193
rect 9143 2141 9151 2193
rect 9175 2141 9211 2193
rect 9211 2141 9227 2193
rect 9227 2141 9231 2193
rect 9255 2141 9279 2193
rect 9279 2141 9311 2193
rect 9095 2137 9151 2141
rect 9175 2137 9231 2141
rect 9255 2137 9311 2141
rect 9095 2107 9151 2110
rect 9175 2107 9231 2110
rect 9255 2107 9311 2110
rect 9095 2055 9143 2107
rect 9143 2055 9151 2107
rect 9175 2055 9211 2107
rect 9211 2055 9227 2107
rect 9227 2055 9231 2107
rect 9255 2055 9279 2107
rect 9279 2055 9311 2107
rect 9095 2054 9151 2055
rect 9175 2054 9231 2055
rect 9255 2054 9311 2055
rect 7604 1296 7660 1300
rect 7701 1296 7757 1300
rect 7797 1296 7853 1300
rect 7604 1244 7653 1296
rect 7653 1244 7660 1296
rect 7701 1244 7721 1296
rect 7721 1244 7737 1296
rect 7737 1244 7757 1296
rect 7797 1244 7804 1296
rect 7804 1244 7853 1296
rect 10369 253 10425 309
rect 10449 253 10505 309
rect 7604 -43 7654 9
rect 7654 -43 7660 9
rect 7604 -47 7660 -43
rect 7701 -43 7703 9
rect 7703 -43 7755 9
rect 7755 -43 7757 9
rect 7701 -47 7757 -43
rect 7797 -43 7803 9
rect 7803 -43 7853 9
rect 7797 -47 7853 -43
rect 7604 -107 7654 -71
rect 7654 -107 7660 -71
rect 7604 -127 7660 -107
rect 7701 -107 7703 -71
rect 7703 -107 7755 -71
rect 7755 -107 7757 -71
rect 7701 -127 7757 -107
rect 7797 -107 7803 -71
rect 7803 -107 7853 -71
rect 7797 -127 7853 -107
rect 12970 211 13026 267
rect 13066 211 13122 267
rect 13162 211 13218 267
rect 13258 211 13314 267
rect 12970 127 13026 183
rect 13066 127 13122 183
rect 13162 127 13218 183
rect 13258 127 13314 183
rect 12970 43 13026 99
rect 13066 43 13122 99
rect 13162 43 13218 99
rect 13258 43 13314 99
rect 12970 -41 13026 15
rect 13066 -41 13122 15
rect 13162 -41 13218 15
rect 13258 -41 13314 15
rect 12970 -125 13026 -69
rect 13066 -125 13122 -69
rect 13162 -125 13218 -69
rect 13258 -125 13314 -69
rect 12970 -210 13026 -154
rect 13066 -210 13122 -154
rect 13162 -210 13218 -154
rect 13258 -210 13314 -154
<< metal3 >>
rect 2972 9884 3324 9892
rect 2972 9820 2974 9884
rect 3038 9820 3068 9884
rect 3132 9820 3162 9884
rect 3226 9820 3256 9884
rect 3320 9820 3324 9884
rect 2972 9792 3324 9820
rect 2972 9728 2974 9792
rect 3038 9728 3068 9792
rect 3132 9728 3162 9792
rect 3226 9728 3256 9792
rect 3320 9728 3324 9792
rect 2972 9700 3324 9728
rect 2972 9636 2974 9700
rect 3038 9636 3068 9700
rect 3132 9636 3162 9700
rect 3226 9636 3256 9700
rect 3320 9636 3324 9700
rect 2972 9608 3324 9636
rect 2972 9544 2974 9608
rect 3038 9544 3068 9608
rect 3132 9544 3162 9608
rect 3226 9544 3256 9608
rect 3320 9544 3324 9608
rect 2972 9516 3324 9544
rect 2972 9452 2974 9516
rect 3038 9452 3068 9516
rect 3132 9452 3162 9516
rect 3226 9452 3256 9516
rect 3320 9452 3324 9516
rect 2972 9423 3324 9452
rect 2972 9359 2974 9423
rect 3038 9359 3068 9423
rect 3132 9359 3162 9423
rect 3226 9359 3256 9423
rect 3320 9359 3324 9423
rect 1124 8869 1190 8874
rect 1124 8813 1129 8869
rect 1185 8813 1190 8869
rect 1124 8789 1190 8813
rect 1124 8733 1129 8789
rect 1185 8733 1190 8789
rect 998 7045 1064 7050
rect 998 6989 1003 7045
rect 1059 6989 1064 7045
rect 998 6965 1064 6989
rect 998 6909 1003 6965
rect 1059 6909 1064 6965
tri 908 3636 998 3726 se
rect 998 3636 1064 6909
rect 908 3572 914 3636
rect 978 3572 994 3636
rect 1058 3572 1064 3636
tri 1087 2495 1124 2532 se
rect 1124 2495 1190 8733
rect 1287 8593 1664 8620
rect 1287 8537 1295 8593
rect 1351 8537 1377 8593
rect 1433 8537 1459 8593
rect 1515 8537 1541 8593
rect 1597 8537 1664 8593
rect 1287 8509 1664 8537
rect 1287 8453 1295 8509
rect 1351 8453 1377 8509
rect 1433 8453 1459 8509
rect 1515 8453 1541 8509
rect 1597 8453 1664 8509
rect 1287 8425 1664 8453
rect 1287 8369 1295 8425
rect 1351 8369 1377 8425
rect 1433 8369 1459 8425
rect 1515 8369 1541 8425
rect 1597 8369 1664 8425
rect 1287 8341 1664 8369
rect 1287 8285 1295 8341
rect 1351 8285 1377 8341
rect 1433 8285 1459 8341
rect 1515 8285 1541 8341
rect 1597 8285 1664 8341
rect 1287 8257 1664 8285
rect 1287 8201 1295 8257
rect 1351 8201 1377 8257
rect 1433 8201 1459 8257
rect 1515 8201 1541 8257
rect 1597 8201 1664 8257
rect 1287 8173 1664 8201
rect 1287 8117 1295 8173
rect 1351 8117 1377 8173
rect 1433 8117 1459 8173
rect 1515 8117 1541 8173
rect 1597 8117 1664 8173
rect 1287 8089 1664 8117
rect 1287 8033 1295 8089
rect 1351 8033 1377 8089
rect 1433 8033 1459 8089
rect 1515 8033 1541 8089
rect 1597 8033 1664 8089
rect 1287 8005 1664 8033
rect 1287 7949 1295 8005
rect 1351 7949 1377 8005
rect 1433 7949 1459 8005
rect 1515 7949 1541 8005
rect 1597 7949 1664 8005
rect 1287 7921 1664 7949
rect 1287 7865 1295 7921
rect 1351 7865 1377 7921
rect 1433 7865 1459 7921
rect 1515 7865 1541 7921
rect 1597 7865 1664 7921
rect 1287 7837 1664 7865
rect 1287 7781 1295 7837
rect 1351 7781 1377 7837
rect 1433 7781 1459 7837
rect 1515 7781 1541 7837
rect 1597 7781 1664 7837
rect 1287 7753 1664 7781
rect 1287 7697 1295 7753
rect 1351 7697 1377 7753
rect 1433 7697 1459 7753
rect 1515 7697 1541 7753
rect 1597 7697 1664 7753
rect 1287 7669 1664 7697
rect 1287 7613 1295 7669
rect 1351 7613 1377 7669
rect 1433 7613 1459 7669
rect 1515 7613 1541 7669
rect 1597 7613 1664 7669
rect 1287 7585 1664 7613
rect 1287 7529 1295 7585
rect 1351 7529 1377 7585
rect 1433 7529 1459 7585
rect 1515 7529 1541 7585
rect 1597 7529 1664 7585
rect 1287 7501 1664 7529
rect 1287 7445 1295 7501
rect 1351 7445 1377 7501
rect 1433 7445 1459 7501
rect 1515 7445 1541 7501
rect 1597 7445 1664 7501
rect 1287 7417 1664 7445
rect 1287 7361 1295 7417
rect 1351 7361 1377 7417
rect 1433 7361 1459 7417
rect 1515 7361 1541 7417
rect 1597 7361 1664 7417
rect 1287 7333 1664 7361
rect 1287 7277 1295 7333
rect 1351 7277 1377 7333
rect 1433 7277 1459 7333
rect 1515 7277 1541 7333
rect 1597 7277 1664 7333
rect 1287 3443 1664 7277
rect 1796 6702 2172 6707
rect 1796 6646 1801 6702
rect 1857 6646 1905 6702
rect 1961 6646 2008 6702
rect 2064 6646 2111 6702
rect 2167 6646 2172 6702
rect 1796 6641 2172 6646
rect 2972 6546 3324 9359
rect 2972 6490 2987 6546
rect 3043 6490 3074 6546
rect 3130 6490 3161 6546
rect 3217 6490 3247 6546
rect 3303 6490 3324 6546
rect 2972 6456 3324 6490
rect 2972 6400 2987 6456
rect 3043 6400 3074 6456
rect 3130 6400 3161 6456
rect 3217 6400 3247 6456
rect 3303 6400 3324 6456
rect 2972 6366 3324 6400
rect 2972 6310 2987 6366
rect 3043 6310 3074 6366
rect 3130 6310 3161 6366
rect 3217 6310 3247 6366
rect 3303 6310 3324 6366
rect 2972 6276 3324 6310
rect 2972 6220 2987 6276
rect 3043 6220 3074 6276
rect 3130 6220 3161 6276
rect 3217 6220 3247 6276
rect 3303 6220 3324 6276
rect 2972 6208 3324 6220
rect 4640 8183 5039 8197
rect 4640 8127 4814 8183
rect 4870 8127 4894 8183
rect 4950 8127 4974 8183
rect 5030 8127 5039 8183
rect 4640 8060 5039 8127
rect 4640 8004 4814 8060
rect 4870 8004 4894 8060
rect 4950 8004 4974 8060
rect 5030 8004 5039 8060
rect 4640 7937 5039 8004
rect 4640 7881 4814 7937
rect 4870 7881 4894 7937
rect 4950 7881 4974 7937
rect 5030 7881 5039 7937
rect 4640 7813 5039 7881
rect 4640 7757 4814 7813
rect 4870 7757 4894 7813
rect 4950 7757 4974 7813
rect 5030 7757 5039 7813
rect 2908 5606 3054 5611
rect 2908 5470 2913 5606
rect 3049 5470 3054 5606
rect 2908 4635 3054 5470
rect 2908 4579 2913 4635
rect 2969 4579 2993 4635
rect 3049 4579 3054 4635
rect 2908 4554 3054 4579
rect 2908 4498 2913 4554
rect 2969 4498 2993 4554
rect 3049 4498 3054 4554
rect 2908 4493 3054 4498
rect 4640 5044 5039 7757
rect 6474 7837 9703 7843
rect 6474 7781 6479 7837
rect 6535 7781 6561 7837
rect 6617 7781 6643 7837
rect 6699 7781 6725 7837
rect 6781 7781 6807 7837
rect 6863 7781 6888 7837
rect 6944 7781 6969 7837
rect 7025 7781 7050 7837
rect 7106 7781 7131 7837
rect 7187 7781 7212 7837
rect 7268 7781 7293 7837
rect 7349 7781 7374 7837
rect 7430 7781 7455 7837
rect 7511 7781 7536 7837
rect 7592 7781 7617 7837
rect 7673 7781 7698 7837
rect 7754 7781 7779 7837
rect 7835 7781 7860 7837
rect 7916 7781 7941 7837
rect 7997 7781 8022 7837
rect 8078 7781 8103 7837
rect 8159 7781 8184 7837
rect 8240 7781 8265 7837
rect 8321 7781 8346 7837
rect 8402 7781 8427 7837
rect 8483 7781 8508 7837
rect 8564 7781 8589 7837
rect 8645 7781 8670 7837
rect 8726 7781 8751 7837
rect 8807 7781 8832 7837
rect 8888 7781 8913 7837
rect 8969 7781 8994 7837
rect 9050 7781 9075 7837
rect 9131 7781 9156 7837
rect 9212 7781 9237 7837
rect 9293 7781 9318 7837
rect 9374 7781 9399 7837
rect 9455 7781 9480 7837
rect 9536 7781 9561 7837
rect 9617 7781 9642 7837
rect 9698 7781 9703 7837
rect 6474 7743 9703 7781
rect 6474 7687 6479 7743
rect 6535 7687 6561 7743
rect 6617 7687 6643 7743
rect 6699 7687 6725 7743
rect 6781 7687 6807 7743
rect 6863 7687 6888 7743
rect 6944 7687 6969 7743
rect 7025 7687 7050 7743
rect 7106 7687 7131 7743
rect 7187 7687 7212 7743
rect 7268 7687 7293 7743
rect 7349 7687 7374 7743
rect 7430 7687 7455 7743
rect 7511 7687 7536 7743
rect 7592 7687 7617 7743
rect 7673 7687 7698 7743
rect 7754 7687 7779 7743
rect 7835 7687 7860 7743
rect 7916 7687 7941 7743
rect 7997 7687 8022 7743
rect 8078 7687 8103 7743
rect 8159 7687 8184 7743
rect 8240 7687 8265 7743
rect 8321 7687 8346 7743
rect 8402 7687 8427 7743
rect 8483 7687 8508 7743
rect 8564 7687 8589 7743
rect 8645 7687 8670 7743
rect 8726 7687 8751 7743
rect 8807 7687 8832 7743
rect 8888 7687 8913 7743
rect 8969 7687 8994 7743
rect 9050 7687 9075 7743
rect 9131 7687 9156 7743
rect 9212 7687 9237 7743
rect 9293 7687 9318 7743
rect 9374 7687 9399 7743
rect 9455 7687 9480 7743
rect 9536 7687 9561 7743
rect 9617 7687 9642 7743
rect 9698 7687 9703 7743
rect 6474 7649 9703 7687
rect 6474 7593 6479 7649
rect 6535 7593 6561 7649
rect 6617 7593 6643 7649
rect 6699 7593 6725 7649
rect 6781 7593 6807 7649
rect 6863 7593 6888 7649
rect 6944 7593 6969 7649
rect 7025 7593 7050 7649
rect 7106 7593 7131 7649
rect 7187 7593 7212 7649
rect 7268 7593 7293 7649
rect 7349 7593 7374 7649
rect 7430 7593 7455 7649
rect 7511 7593 7536 7649
rect 7592 7593 7617 7649
rect 7673 7593 7698 7649
rect 7754 7593 7779 7649
rect 7835 7593 7860 7649
rect 7916 7593 7941 7649
rect 7997 7593 8022 7649
rect 8078 7593 8103 7649
rect 8159 7593 8184 7649
rect 8240 7593 8265 7649
rect 8321 7593 8346 7649
rect 8402 7593 8427 7649
rect 8483 7593 8508 7649
rect 8564 7593 8589 7649
rect 8645 7593 8670 7649
rect 8726 7593 8751 7649
rect 8807 7593 8832 7649
rect 8888 7593 8913 7649
rect 8969 7593 8994 7649
rect 9050 7593 9075 7649
rect 9131 7593 9156 7649
rect 9212 7593 9237 7649
rect 9293 7593 9318 7649
rect 9374 7593 9399 7649
rect 9455 7593 9480 7649
rect 9536 7593 9561 7649
rect 9617 7593 9642 7649
rect 9698 7593 9703 7649
rect 6474 7555 9703 7593
rect 6474 7499 6479 7555
rect 6535 7499 6561 7555
rect 6617 7499 6643 7555
rect 6699 7499 6725 7555
rect 6781 7499 6807 7555
rect 6863 7499 6888 7555
rect 6944 7499 6969 7555
rect 7025 7499 7050 7555
rect 7106 7499 7131 7555
rect 7187 7499 7212 7555
rect 7268 7499 7293 7555
rect 7349 7499 7374 7555
rect 7430 7499 7455 7555
rect 7511 7499 7536 7555
rect 7592 7499 7617 7555
rect 7673 7499 7698 7555
rect 7754 7499 7779 7555
rect 7835 7499 7860 7555
rect 7916 7499 7941 7555
rect 7997 7499 8022 7555
rect 8078 7499 8103 7555
rect 8159 7499 8184 7555
rect 8240 7499 8265 7555
rect 8321 7499 8346 7555
rect 8402 7499 8427 7555
rect 8483 7499 8508 7555
rect 8564 7499 8589 7555
rect 8645 7499 8670 7555
rect 8726 7499 8751 7555
rect 8807 7499 8832 7555
rect 8888 7499 8913 7555
rect 8969 7499 8994 7555
rect 9050 7499 9075 7555
rect 9131 7499 9156 7555
rect 9212 7499 9237 7555
rect 9293 7499 9318 7555
rect 9374 7499 9399 7555
rect 9455 7499 9480 7555
rect 9536 7499 9561 7555
rect 9617 7499 9642 7555
rect 9698 7499 9703 7555
rect 6474 7493 9703 7499
rect 6474 7426 7059 7493
tri 7059 7426 7126 7493 nw
rect 5159 7421 5413 7426
rect 5159 7365 5164 7421
rect 5220 7365 5258 7421
rect 5314 7365 5352 7421
rect 5408 7365 5413 7421
rect 5159 7319 5413 7365
rect 5159 7263 5164 7319
rect 5220 7263 5258 7319
rect 5314 7263 5352 7319
rect 5408 7263 5413 7319
rect 6474 7420 7053 7426
tri 7053 7420 7059 7426 nw
rect 6474 7413 7046 7420
tri 7046 7413 7053 7420 nw
rect 9394 7413 9821 7420
rect 6474 7366 6999 7413
tri 6999 7366 7046 7413 nw
rect 6474 7361 6994 7366
tri 6994 7361 6999 7366 nw
rect 8847 7361 9284 7366
rect 5159 7217 5413 7263
rect 5159 7161 5164 7217
rect 5220 7161 5258 7217
rect 5314 7161 5352 7217
rect 5408 7161 5413 7217
rect 5159 7115 5413 7161
rect 5159 7059 5164 7115
rect 5220 7059 5258 7115
rect 5314 7059 5352 7115
rect 5408 7059 5413 7115
rect 5159 5924 5413 7059
rect 5159 5868 5164 5924
rect 5220 5868 5258 5924
rect 5314 5868 5352 5924
rect 5408 5868 5413 5924
rect 5159 5822 5413 5868
rect 5159 5766 5164 5822
rect 5220 5766 5258 5822
rect 5314 5766 5352 5822
rect 5408 5766 5413 5822
rect 5159 5720 5413 5766
rect 5159 5664 5164 5720
rect 5220 5664 5258 5720
rect 5314 5664 5352 5720
rect 5408 5664 5413 5720
rect 5159 5618 5413 5664
rect 5587 7274 5975 7279
rect 5587 7218 5593 7274
rect 5649 7218 5673 7274
rect 5729 7218 5753 7274
rect 5809 7218 5833 7274
rect 5889 7218 5913 7274
rect 5969 7218 5975 7274
rect 5587 7186 5975 7218
rect 5587 7130 5593 7186
rect 5649 7130 5673 7186
rect 5729 7130 5753 7186
rect 5809 7130 5833 7186
rect 5889 7130 5913 7186
rect 5969 7130 5975 7186
rect 5587 7097 5975 7130
rect 5587 7041 5593 7097
rect 5649 7041 5673 7097
rect 5729 7041 5753 7097
rect 5809 7041 5833 7097
rect 5889 7041 5913 7097
rect 5969 7041 5975 7097
rect 5587 7008 5975 7041
rect 5587 6952 5593 7008
rect 5649 6952 5673 7008
rect 5729 6952 5753 7008
rect 5809 6952 5833 7008
rect 5889 6952 5913 7008
rect 5969 6952 5975 7008
rect 5587 6031 5975 6952
rect 5587 5975 5593 6031
rect 5649 5975 5673 6031
rect 5729 5975 5753 6031
rect 5809 5975 5833 6031
rect 5889 5975 5913 6031
rect 5969 5975 5975 6031
rect 5587 5929 5975 5975
rect 5587 5873 5593 5929
rect 5649 5873 5673 5929
rect 5729 5873 5753 5929
rect 5809 5873 5833 5929
rect 5889 5873 5913 5929
rect 5969 5873 5975 5929
rect 5587 5827 5975 5873
rect 5587 5771 5593 5827
rect 5649 5771 5673 5827
rect 5729 5771 5753 5827
rect 5809 5771 5833 5827
rect 5889 5771 5913 5827
rect 5969 5771 5975 5827
rect 5587 5725 5975 5771
rect 5587 5669 5593 5725
rect 5649 5669 5673 5725
rect 5729 5669 5753 5725
rect 5809 5669 5833 5725
rect 5889 5669 5913 5725
rect 5969 5669 5975 5725
rect 5587 5660 5975 5669
tri 6285 6779 6474 6968 se
rect 6474 6783 6951 7361
tri 6951 7318 6994 7361 nw
rect 6474 6779 6947 6783
tri 6947 6779 6951 6783 nw
rect 8847 7305 8856 7361
rect 8912 7305 8947 7361
rect 9003 7305 9038 7361
rect 9094 7305 9129 7361
rect 9185 7305 9219 7361
rect 9275 7305 9284 7361
rect 8847 7225 9284 7305
rect 8847 7169 8856 7225
rect 8912 7169 8947 7225
rect 9003 7169 9038 7225
rect 9094 7169 9129 7225
rect 9185 7169 9219 7225
rect 9275 7169 9284 7225
rect 6285 6675 6843 6779
tri 6843 6675 6947 6779 nw
rect 8847 6675 9284 7169
rect 6285 6619 6787 6675
tri 6787 6619 6843 6675 nw
rect 8847 6619 8856 6675
rect 8912 6619 8947 6675
rect 9003 6619 9038 6675
rect 9094 6619 9129 6675
rect 9185 6619 9219 6675
rect 9275 6619 9284 6675
rect 6285 6595 6763 6619
tri 6763 6595 6787 6619 nw
rect 8847 6595 9284 6619
rect 5159 5562 5164 5618
rect 5220 5562 5258 5618
rect 5314 5562 5352 5618
rect 5408 5562 5413 5618
rect 5159 5557 5413 5562
rect 4640 4988 4814 5044
rect 4870 4988 4894 5044
rect 4950 4988 4974 5044
rect 5030 4988 5039 5044
rect 4640 4919 5039 4988
rect 4640 4863 4814 4919
rect 4870 4863 4894 4919
rect 4950 4863 4974 4919
rect 5030 4863 5039 4919
rect 4640 4793 5039 4863
rect 4640 4737 4814 4793
rect 4870 4737 4894 4793
rect 4950 4737 4974 4793
rect 5030 4737 5039 4793
rect 4640 4667 5039 4737
rect 4640 4611 4814 4667
rect 4870 4611 4894 4667
rect 4950 4611 4974 4667
rect 5030 4611 5039 4667
rect 4640 4541 5039 4611
rect 1287 3379 1291 3443
rect 1355 3379 1393 3443
rect 1457 3379 1495 3443
rect 1559 3379 1597 3443
rect 1661 3379 1664 3443
rect 1287 3363 1664 3379
rect 1287 3299 1291 3363
rect 1355 3299 1393 3363
rect 1457 3299 1495 3363
rect 1559 3299 1597 3363
rect 1661 3299 1664 3363
rect 1287 3283 1664 3299
rect 1287 3219 1291 3283
rect 1355 3219 1393 3283
rect 1457 3219 1495 3283
rect 1559 3219 1597 3283
rect 1661 3219 1664 3283
rect 4640 4485 4814 4541
rect 4870 4485 4894 4541
rect 4950 4485 4974 4541
rect 5030 4485 5039 4541
rect 4640 3280 5039 4485
rect 5915 4295 6182 4318
rect 5915 4239 5924 4295
rect 5980 4239 6023 4295
rect 6079 4239 6121 4295
rect 6177 4239 6182 4295
rect 5915 3655 6182 4239
rect 1287 3202 1664 3219
rect 1287 3138 1291 3202
rect 1355 3138 1393 3202
rect 1457 3138 1495 3202
rect 1559 3138 1597 3202
rect 1661 3138 1664 3202
rect 1287 3121 1664 3138
rect 1287 3057 1291 3121
rect 1355 3057 1393 3121
rect 1457 3057 1495 3121
rect 1559 3057 1597 3121
rect 1661 3057 1664 3121
rect 1287 3040 1664 3057
rect 1287 2976 1291 3040
rect 1355 2976 1393 3040
rect 1457 2976 1495 3040
rect 1559 2976 1597 3040
rect 1661 2976 1664 3040
rect 1287 2959 1664 2976
rect 1287 2895 1291 2959
rect 1355 2895 1393 2959
rect 1457 2895 1495 2959
rect 1559 2895 1597 2959
rect 1661 2895 1664 2959
rect 1287 2878 1664 2895
rect 1287 2814 1291 2878
rect 1355 2814 1393 2878
rect 1457 2814 1495 2878
rect 1559 2814 1597 2878
rect 1661 2814 1664 2878
rect 1287 2797 1664 2814
rect 1287 2733 1291 2797
rect 1355 2733 1393 2797
rect 1457 2733 1495 2797
rect 1559 2733 1597 2797
rect 1661 2733 1664 2797
rect 1287 2716 1664 2733
rect 1287 2652 1291 2716
rect 1355 2652 1393 2716
rect 1457 2652 1495 2716
rect 1559 2652 1597 2716
rect 1661 2652 1664 2716
rect 1287 2635 1664 2652
rect 1287 2571 1291 2635
rect 1355 2571 1393 2635
rect 1457 2571 1495 2635
rect 1559 2571 1597 2635
rect 1661 2571 1664 2635
rect 1287 2563 1664 2571
tri 1059 2467 1087 2495 se
rect 1087 2467 1190 2495
tri 1054 2462 1059 2467 se
rect 1059 2462 1190 2467
tri 1190 2462 1195 2467 sw
rect 1039 2398 1045 2462
rect 1109 2398 1125 2462
rect 1189 2398 1195 2462
rect 3264 1983 3446 1988
rect 3264 1847 3285 1983
rect 3421 1847 3446 1983
rect 3264 1304 3446 1847
rect 6285 960 6754 6595
tri 6754 6586 6763 6595 nw
rect 8847 6539 8856 6595
rect 8912 6539 8947 6595
rect 9003 6539 9038 6595
rect 9094 6539 9129 6595
rect 9185 6539 9219 6595
rect 9275 6539 9284 6595
rect 8847 6515 9284 6539
rect 8847 6459 8856 6515
rect 8912 6459 8947 6515
rect 9003 6459 9038 6515
rect 9094 6459 9129 6515
rect 9185 6459 9219 6515
rect 9275 6459 9284 6515
rect 8847 6435 9284 6459
rect 8847 6379 8856 6435
rect 8912 6379 8947 6435
rect 9003 6379 9038 6435
rect 9094 6379 9129 6435
rect 9185 6379 9219 6435
rect 9275 6379 9284 6435
rect 8847 6374 9284 6379
rect 9394 7357 9403 7413
rect 9459 7357 9490 7413
rect 9546 7357 9577 7413
rect 9633 7357 9664 7413
rect 9720 7357 9750 7413
rect 9806 7357 9821 7413
rect 9394 7321 9821 7357
rect 9394 7265 9403 7321
rect 9459 7265 9490 7321
rect 9546 7265 9577 7321
rect 9633 7265 9664 7321
rect 9720 7265 9750 7321
rect 9806 7265 9821 7321
rect 9394 7229 9821 7265
rect 9394 7173 9403 7229
rect 9459 7173 9490 7229
rect 9546 7173 9577 7229
rect 9633 7173 9664 7229
rect 9720 7173 9750 7229
rect 9806 7173 9821 7229
rect 9394 7137 9821 7173
rect 9394 7081 9403 7137
rect 9459 7081 9490 7137
rect 9546 7081 9577 7137
rect 9633 7081 9664 7137
rect 9720 7081 9750 7137
rect 9806 7081 9821 7137
rect 9394 5839 9821 7081
rect 9394 5783 9403 5839
rect 9459 5783 9489 5839
rect 9545 5783 9575 5839
rect 9631 5783 9661 5839
rect 9717 5783 9746 5839
rect 9802 5783 9821 5839
rect 9394 5735 9821 5783
rect 9394 5679 9403 5735
rect 9459 5679 9489 5735
rect 9545 5679 9575 5735
rect 9631 5679 9661 5735
rect 9717 5679 9746 5735
rect 9802 5679 9821 5735
rect 9394 5631 9821 5679
rect 9394 5575 9403 5631
rect 9459 5575 9489 5631
rect 9545 5575 9575 5631
rect 9631 5575 9661 5631
rect 9717 5575 9746 5631
rect 9802 5575 9821 5631
rect 9394 5569 9821 5575
rect 7851 5411 11202 5417
rect 7851 5355 7856 5411
rect 7912 5355 7937 5411
rect 7993 5355 8018 5411
rect 8074 5355 8099 5411
rect 8155 5355 8180 5411
rect 8236 5355 8261 5411
rect 8317 5355 8341 5411
rect 8397 5355 8421 5411
rect 8477 5355 8501 5411
rect 8557 5355 8581 5411
rect 8637 5355 8661 5411
rect 8717 5355 8741 5411
rect 8797 5355 8821 5411
rect 8877 5355 8901 5411
rect 8957 5355 8981 5411
rect 9037 5355 9061 5411
rect 9117 5355 9141 5411
rect 9197 5355 9221 5411
rect 9277 5355 9301 5411
rect 9357 5355 9381 5411
rect 9437 5355 9461 5411
rect 9517 5355 9541 5411
rect 9597 5355 9621 5411
rect 9677 5355 9701 5411
rect 9757 5355 9781 5411
rect 9837 5355 9861 5411
rect 9917 5355 9941 5411
rect 9997 5355 10021 5411
rect 10077 5355 10101 5411
rect 10157 5355 10181 5411
rect 10237 5355 10261 5411
rect 10317 5355 10341 5411
rect 10397 5355 10421 5411
rect 10477 5355 10501 5411
rect 10557 5355 10581 5411
rect 10637 5355 10661 5411
rect 10717 5355 10741 5411
rect 10797 5355 10821 5411
rect 10877 5355 10901 5411
rect 10957 5355 10981 5411
rect 11037 5355 11061 5411
rect 11117 5355 11141 5411
rect 11197 5355 11202 5411
rect 7851 5317 11202 5355
rect 7851 5261 7856 5317
rect 7912 5261 7937 5317
rect 7993 5261 8018 5317
rect 8074 5261 8099 5317
rect 8155 5261 8180 5317
rect 8236 5261 8261 5317
rect 8317 5261 8341 5317
rect 8397 5261 8421 5317
rect 8477 5261 8501 5317
rect 8557 5261 8581 5317
rect 8637 5261 8661 5317
rect 8717 5261 8741 5317
rect 8797 5261 8821 5317
rect 8877 5261 8901 5317
rect 8957 5261 8981 5317
rect 9037 5261 9061 5317
rect 9117 5261 9141 5317
rect 9197 5261 9221 5317
rect 9277 5261 9301 5317
rect 9357 5261 9381 5317
rect 9437 5261 9461 5317
rect 9517 5261 9541 5317
rect 9597 5261 9621 5317
rect 9677 5261 9701 5317
rect 9757 5261 9781 5317
rect 9837 5261 9861 5317
rect 9917 5261 9941 5317
rect 9997 5261 10021 5317
rect 10077 5261 10101 5317
rect 10157 5261 10181 5317
rect 10237 5261 10261 5317
rect 10317 5261 10341 5317
rect 10397 5261 10421 5317
rect 10477 5261 10501 5317
rect 10557 5261 10581 5317
rect 10637 5261 10661 5317
rect 10717 5261 10741 5317
rect 10797 5261 10821 5317
rect 10877 5261 10901 5317
rect 10957 5261 10981 5317
rect 11037 5261 11061 5317
rect 11117 5261 11141 5317
rect 11197 5261 11202 5317
rect 7851 5223 11202 5261
rect 7851 5167 7856 5223
rect 7912 5167 7937 5223
rect 7993 5167 8018 5223
rect 8074 5167 8099 5223
rect 8155 5167 8180 5223
rect 8236 5167 8261 5223
rect 8317 5167 8341 5223
rect 8397 5167 8421 5223
rect 8477 5167 8501 5223
rect 8557 5167 8581 5223
rect 8637 5167 8661 5223
rect 8717 5167 8741 5223
rect 8797 5167 8821 5223
rect 8877 5167 8901 5223
rect 8957 5167 8981 5223
rect 9037 5167 9061 5223
rect 9117 5167 9141 5223
rect 9197 5167 9221 5223
rect 9277 5167 9301 5223
rect 9357 5167 9381 5223
rect 9437 5167 9461 5223
rect 9517 5167 9541 5223
rect 9597 5167 9621 5223
rect 9677 5167 9701 5223
rect 9757 5167 9781 5223
rect 9837 5167 9861 5223
rect 9917 5167 9941 5223
rect 9997 5167 10021 5223
rect 10077 5167 10101 5223
rect 10157 5167 10181 5223
rect 10237 5167 10261 5223
rect 10317 5167 10341 5223
rect 10397 5167 10421 5223
rect 10477 5167 10501 5223
rect 10557 5167 10581 5223
rect 10637 5167 10661 5223
rect 10717 5167 10741 5223
rect 10797 5167 10821 5223
rect 10877 5167 10901 5223
rect 10957 5167 10981 5223
rect 11037 5167 11061 5223
rect 11117 5167 11141 5223
rect 11197 5167 11202 5223
rect 7851 5129 11202 5167
rect 7851 5073 7856 5129
rect 7912 5073 7937 5129
rect 7993 5073 8018 5129
rect 8074 5073 8099 5129
rect 8155 5073 8180 5129
rect 8236 5073 8261 5129
rect 8317 5073 8341 5129
rect 8397 5073 8421 5129
rect 8477 5073 8501 5129
rect 8557 5073 8581 5129
rect 8637 5073 8661 5129
rect 8717 5073 8741 5129
rect 8797 5073 8821 5129
rect 8877 5073 8901 5129
rect 8957 5073 8981 5129
rect 9037 5073 9061 5129
rect 9117 5073 9141 5129
rect 9197 5073 9221 5129
rect 9277 5073 9301 5129
rect 9357 5073 9381 5129
rect 9437 5073 9461 5129
rect 9517 5073 9541 5129
rect 9597 5073 9621 5129
rect 9677 5073 9701 5129
rect 9757 5073 9781 5129
rect 9837 5073 9861 5129
rect 9917 5073 9941 5129
rect 9997 5073 10021 5129
rect 10077 5073 10101 5129
rect 10157 5073 10181 5129
rect 10237 5073 10261 5129
rect 10317 5073 10341 5129
rect 10397 5073 10421 5129
rect 10477 5073 10501 5129
rect 10557 5073 10581 5129
rect 10637 5073 10661 5129
rect 10717 5073 10741 5129
rect 10797 5073 10821 5129
rect 10877 5073 10901 5129
rect 10957 5073 10981 5129
rect 11037 5073 11061 5129
rect 11117 5073 11141 5129
rect 11197 5073 11202 5129
rect 7851 5067 11202 5073
tri 9271 4912 9426 5067 ne
rect 9426 4912 9914 5067
tri 9914 4912 10069 5067 nw
rect 9090 3040 9316 3049
rect 9090 2984 9095 3040
rect 9151 2984 9175 3040
rect 9231 2984 9255 3040
rect 9311 2984 9316 3040
rect 9090 2942 9316 2984
rect 9090 2886 9095 2942
rect 9151 2886 9175 2942
rect 9231 2886 9255 2942
rect 9311 2886 9316 2942
rect 9090 2844 9316 2886
rect 9090 2788 9095 2844
rect 9151 2788 9175 2844
rect 9231 2788 9255 2844
rect 9311 2788 9316 2844
rect 9090 2746 9316 2788
rect 9090 2690 9095 2746
rect 9151 2690 9175 2746
rect 9231 2690 9255 2746
rect 9311 2690 9316 2746
rect 6285 896 6288 960
rect 6352 896 6368 960
rect 6432 896 6448 960
rect 6512 896 6528 960
rect 6592 896 6608 960
rect 6672 896 6688 960
rect 6752 896 6754 960
rect 6285 872 6754 896
rect 6285 808 6288 872
rect 6352 808 6368 872
rect 6432 808 6448 872
rect 6512 808 6528 872
rect 6592 808 6608 872
rect 6672 808 6688 872
rect 6752 808 6754 872
rect 6285 784 6754 808
rect 6285 720 6288 784
rect 6352 720 6368 784
rect 6432 720 6448 784
rect 6512 720 6528 784
rect 6592 720 6608 784
rect 6672 720 6688 784
rect 6752 720 6754 784
rect 6285 696 6754 720
rect 6285 632 6288 696
rect 6352 632 6368 696
rect 6432 632 6448 696
rect 6512 632 6528 696
rect 6592 632 6608 696
rect 6672 632 6688 696
rect 6752 632 6754 696
rect 6285 608 6754 632
rect 6285 544 6288 608
rect 6352 544 6368 608
rect 6432 544 6448 608
rect 6512 544 6528 608
rect 6592 544 6608 608
rect 6672 544 6688 608
rect 6752 544 6754 608
rect 6285 519 6754 544
rect 6285 455 6288 519
rect 6352 455 6368 519
rect 6432 455 6448 519
rect 6512 455 6528 519
rect 6592 455 6608 519
rect 6672 455 6688 519
rect 6752 455 6754 519
rect 6285 430 6754 455
rect 6285 366 6288 430
rect 6352 366 6368 430
rect 6432 366 6448 430
rect 6512 366 6528 430
rect 6592 366 6608 430
rect 6672 366 6688 430
rect 6752 366 6754 430
rect 6285 360 6754 366
rect 7595 2299 7862 2323
rect 7595 2243 7609 2299
rect 7665 2243 7701 2299
rect 7757 2243 7792 2299
rect 7848 2243 7862 2299
rect 7595 1300 7862 2243
rect 9090 2275 9316 2690
rect 9090 2219 9095 2275
rect 9151 2219 9175 2275
rect 9231 2219 9255 2275
rect 9311 2219 9316 2275
rect 9090 2193 9316 2219
rect 9090 2137 9095 2193
rect 9151 2137 9175 2193
rect 9231 2137 9255 2193
rect 9311 2137 9316 2193
rect 9090 2110 9316 2137
rect 9090 2054 9095 2110
rect 9151 2054 9175 2110
rect 9231 2054 9255 2110
rect 9311 2054 9316 2110
rect 9090 2049 9316 2054
rect 7595 1244 7604 1300
rect 7660 1244 7701 1300
rect 7757 1244 7797 1300
rect 7853 1244 7862 1300
rect 7595 9 7862 1244
rect 7595 -47 7604 9
rect 7660 -47 7701 9
rect 7757 -47 7797 9
rect 7853 -47 7862 9
rect 7595 -71 7862 -47
rect 7595 -127 7604 -71
rect 7660 -127 7701 -71
rect 7757 -127 7797 -71
rect 7853 -127 7862 -71
rect 7595 -132 7862 -127
rect 9426 8 9895 4912
tri 9895 4893 9914 4912 nw
tri 12601 4135 13014 4548 se
rect 13014 4396 13308 5783
rect 13014 4135 13016 4396
tri 12570 4104 12601 4135 se
rect 12601 4104 13016 4135
tri 13016 4104 13308 4396 nw
rect 12068 4099 12919 4104
rect 12068 4043 12669 4099
rect 12725 4043 12759 4099
rect 12815 4043 12848 4099
rect 12904 4043 12919 4099
rect 12068 4007 12919 4043
tri 12919 4007 13016 4104 nw
rect 9426 -56 9429 8
rect 9493 -56 9509 8
rect 9573 -56 9589 8
rect 9653 -56 9669 8
rect 9733 -56 9749 8
rect 9813 -56 9829 8
rect 9893 -56 9895 8
rect 9426 -80 9895 -56
rect 9426 -144 9429 -80
rect 9493 -144 9509 -80
rect 9573 -144 9589 -80
rect 9653 -144 9669 -80
rect 9733 -144 9749 -80
rect 9813 -144 9829 -80
rect 9893 -144 9895 -80
rect 9426 -168 9895 -144
rect 9426 -232 9429 -168
rect 9493 -232 9509 -168
rect 9573 -232 9589 -168
rect 9653 -232 9669 -168
rect 9733 -232 9749 -168
rect 9813 -232 9829 -168
rect 9893 -232 9895 -168
rect 9426 -256 9895 -232
rect 9426 -320 9429 -256
rect 9493 -320 9509 -256
rect 9573 -320 9589 -256
rect 9653 -320 9669 -256
rect 9733 -320 9749 -256
rect 9813 -320 9829 -256
rect 9893 -320 9895 -256
rect 9426 -344 9895 -320
rect 9426 -408 9429 -344
rect 9493 -408 9509 -344
rect 9573 -408 9589 -344
rect 9653 -408 9669 -344
rect 9733 -408 9749 -344
rect 9813 -408 9829 -344
rect 9893 -408 9895 -344
rect 9426 -433 9895 -408
rect 9426 -497 9429 -433
rect 9493 -497 9509 -433
rect 9573 -497 9589 -433
rect 9653 -497 9669 -433
rect 9733 -497 9749 -433
rect 9813 -497 9829 -433
rect 9893 -497 9895 -433
rect 9426 -522 9895 -497
rect 9426 -586 9429 -522
rect 9493 -586 9509 -522
rect 9573 -586 9589 -522
rect 9653 -586 9669 -522
rect 9733 -586 9749 -522
rect 9813 -586 9829 -522
rect 9893 -586 9895 -522
rect 9426 -592 9895 -586
rect 10347 3049 10711 3059
rect 10347 2993 10356 3049
rect 10412 2993 10453 3049
rect 10509 2993 10550 3049
rect 10606 2993 10646 3049
rect 10702 2993 10711 3049
rect 10347 2945 10711 2993
rect 10347 2889 10356 2945
rect 10412 2889 10453 2945
rect 10509 2889 10550 2945
rect 10606 2889 10646 2945
rect 10702 2889 10711 2945
rect 10347 2841 10711 2889
rect 10347 2785 10356 2841
rect 10412 2785 10453 2841
rect 10509 2785 10550 2841
rect 10606 2785 10646 2841
rect 10702 2785 10711 2841
rect 10347 2737 10711 2785
rect 10347 2681 10356 2737
rect 10412 2681 10453 2737
rect 10509 2681 10550 2737
rect 10606 2681 10646 2737
rect 10702 2681 10711 2737
rect 10347 309 10711 2681
rect 12068 2975 12884 4007
tri 12884 3972 12919 4007 nw
rect 12068 2919 12073 2975
rect 12129 2919 12198 2975
rect 12254 2919 12323 2975
rect 12379 2919 12448 2975
rect 12504 2919 12573 2975
rect 12629 2919 12698 2975
rect 12754 2919 12823 2975
rect 12879 2919 12884 2975
rect 12068 2869 12884 2919
rect 12068 2813 12073 2869
rect 12129 2813 12198 2869
rect 12254 2813 12323 2869
rect 12379 2813 12448 2869
rect 12504 2813 12573 2869
rect 12629 2813 12698 2869
rect 12754 2813 12823 2869
rect 12879 2813 12884 2869
rect 12068 2763 12884 2813
rect 12068 2707 12073 2763
rect 12129 2707 12198 2763
rect 12254 2707 12323 2763
rect 12379 2707 12448 2763
rect 12504 2707 12573 2763
rect 12629 2707 12698 2763
rect 12754 2707 12823 2763
rect 12879 2707 12884 2763
rect 12068 2657 12884 2707
rect 12964 3572 12970 3636
rect 13034 3572 13050 3636
rect 13114 3572 13120 3636
rect 12964 2756 13120 3572
rect 12964 2700 12969 2756
rect 13025 2700 13049 2756
rect 13105 2700 13120 2756
rect 12964 2695 13120 2700
rect 12068 2601 12073 2657
rect 12129 2601 12198 2657
rect 12254 2601 12323 2657
rect 12379 2601 12448 2657
rect 12504 2601 12573 2657
rect 12629 2601 12698 2657
rect 12754 2601 12823 2657
rect 12879 2601 12884 2657
rect 12068 2551 12884 2601
rect 12068 2495 12073 2551
rect 12129 2495 12198 2551
rect 12254 2495 12323 2551
rect 12379 2495 12448 2551
rect 12504 2495 12573 2551
rect 12629 2495 12698 2551
rect 12754 2495 12823 2551
rect 12879 2495 12884 2551
rect 12068 1047 12884 2495
rect 13109 2462 13268 2463
rect 13109 2458 13118 2462
rect 13182 2458 13198 2462
rect 13109 2402 13114 2458
rect 13182 2402 13194 2458
rect 13109 2398 13118 2402
rect 13182 2398 13198 2402
rect 13262 2398 13268 2462
rect 13109 2397 13268 2398
rect 12965 2255 13320 2273
rect 12965 2191 12969 2255
rect 13033 2191 13063 2255
rect 13127 2191 13157 2255
rect 13221 2191 13251 2255
rect 13315 2191 13320 2255
rect 12965 2167 13320 2191
rect 12965 2103 12969 2167
rect 13033 2103 13063 2167
rect 13127 2103 13157 2167
rect 13221 2103 13251 2167
rect 13315 2103 13320 2167
rect 12965 2079 13320 2103
rect 12965 2015 12969 2079
rect 13033 2015 13063 2079
rect 13127 2015 13157 2079
rect 13221 2015 13251 2079
rect 13315 2015 13320 2079
rect 12965 1991 13320 2015
rect 12965 1927 12969 1991
rect 13033 1927 13063 1991
rect 13127 1927 13157 1991
rect 13221 1927 13251 1991
rect 13315 1927 13320 1991
rect 12965 1903 13320 1927
rect 12965 1839 12969 1903
rect 13033 1839 13063 1903
rect 13127 1839 13157 1903
rect 13221 1839 13251 1903
rect 13315 1839 13320 1903
rect 12965 1814 13320 1839
rect 12965 1750 12969 1814
rect 13033 1750 13063 1814
rect 13127 1750 13157 1814
rect 13221 1750 13251 1814
rect 13315 1750 13320 1814
rect 12965 1725 13320 1750
rect 12965 1661 12969 1725
rect 13033 1661 13063 1725
rect 13127 1661 13157 1725
rect 13221 1661 13251 1725
rect 13315 1661 13320 1725
rect 12965 1636 13320 1661
rect 12965 1572 12969 1636
rect 13033 1572 13063 1636
rect 13127 1572 13157 1636
rect 13221 1572 13251 1636
rect 13315 1572 13320 1636
rect 12965 1547 13320 1572
rect 12965 1483 12969 1547
rect 13033 1483 13063 1547
rect 13127 1483 13157 1547
rect 13221 1483 13251 1547
rect 13315 1483 13320 1547
rect 12965 1458 13320 1483
rect 12965 1394 12969 1458
rect 13033 1394 13063 1458
rect 13127 1394 13157 1458
rect 13221 1394 13251 1458
rect 13315 1394 13320 1458
rect 10347 253 10369 309
rect 10425 253 10449 309
rect 10505 253 10711 309
tri 10341 -7548 10347 -7542 se
rect 10347 -8480 10711 253
rect 12965 267 13320 1394
rect 12965 211 12970 267
rect 13026 211 13066 267
rect 13122 211 13162 267
rect 13218 211 13258 267
rect 13314 211 13320 267
rect 12965 183 13320 211
rect 12965 127 12970 183
rect 13026 127 13066 183
rect 13122 127 13162 183
rect 13218 127 13258 183
rect 13314 127 13320 183
rect 12965 99 13320 127
rect 12965 43 12970 99
rect 13026 43 13066 99
rect 13122 43 13162 99
rect 13218 43 13258 99
rect 13314 43 13320 99
rect 12965 15 13320 43
rect 12965 -41 12970 15
rect 13026 -41 13066 15
rect 13122 -41 13162 15
rect 13218 -41 13258 15
rect 13314 -41 13320 15
rect 12965 -69 13320 -41
rect 12965 -125 12970 -69
rect 13026 -125 13066 -69
rect 13122 -125 13162 -69
rect 13218 -125 13258 -69
rect 13314 -125 13320 -69
rect 12965 -154 13320 -125
rect 12965 -210 12970 -154
rect 13026 -210 13066 -154
rect 13122 -210 13162 -154
rect 13218 -210 13258 -154
rect 13314 -210 13320 -154
rect 12965 -219 13320 -210
rect 14175 -10153 14185 -10087
<< via3 >>
rect 2974 9820 3038 9884
rect 3068 9820 3132 9884
rect 3162 9820 3226 9884
rect 3256 9820 3320 9884
rect 2974 9728 3038 9792
rect 3068 9728 3132 9792
rect 3162 9728 3226 9792
rect 3256 9728 3320 9792
rect 2974 9636 3038 9700
rect 3068 9636 3132 9700
rect 3162 9636 3226 9700
rect 3256 9636 3320 9700
rect 2974 9544 3038 9608
rect 3068 9544 3132 9608
rect 3162 9544 3226 9608
rect 3256 9544 3320 9608
rect 2974 9452 3038 9516
rect 3068 9452 3132 9516
rect 3162 9452 3226 9516
rect 3256 9452 3320 9516
rect 2974 9359 3038 9423
rect 3068 9359 3132 9423
rect 3162 9359 3226 9423
rect 3256 9359 3320 9423
rect 914 3572 978 3636
rect 994 3572 1058 3636
rect 1291 3379 1355 3443
rect 1393 3379 1457 3443
rect 1495 3379 1559 3443
rect 1597 3379 1661 3443
rect 1291 3299 1355 3363
rect 1393 3299 1457 3363
rect 1495 3299 1559 3363
rect 1597 3299 1661 3363
rect 1291 3219 1355 3283
rect 1393 3219 1457 3283
rect 1495 3219 1559 3283
rect 1597 3219 1661 3283
rect 1291 3138 1355 3202
rect 1393 3138 1457 3202
rect 1495 3138 1559 3202
rect 1597 3138 1661 3202
rect 1291 3057 1355 3121
rect 1393 3057 1457 3121
rect 1495 3057 1559 3121
rect 1597 3057 1661 3121
rect 1291 2976 1355 3040
rect 1393 2976 1457 3040
rect 1495 2976 1559 3040
rect 1597 2976 1661 3040
rect 1291 2895 1355 2959
rect 1393 2895 1457 2959
rect 1495 2895 1559 2959
rect 1597 2895 1661 2959
rect 1291 2814 1355 2878
rect 1393 2814 1457 2878
rect 1495 2814 1559 2878
rect 1597 2814 1661 2878
rect 1291 2733 1355 2797
rect 1393 2733 1457 2797
rect 1495 2733 1559 2797
rect 1597 2733 1661 2797
rect 1291 2652 1355 2716
rect 1393 2652 1457 2716
rect 1495 2652 1559 2716
rect 1597 2652 1661 2716
rect 1291 2571 1355 2635
rect 1393 2571 1457 2635
rect 1495 2571 1559 2635
rect 1597 2571 1661 2635
rect 1045 2398 1109 2462
rect 1125 2398 1189 2462
rect 6288 896 6352 960
rect 6368 896 6432 960
rect 6448 896 6512 960
rect 6528 896 6592 960
rect 6608 896 6672 960
rect 6688 896 6752 960
rect 6288 808 6352 872
rect 6368 808 6432 872
rect 6448 808 6512 872
rect 6528 808 6592 872
rect 6608 808 6672 872
rect 6688 808 6752 872
rect 6288 720 6352 784
rect 6368 720 6432 784
rect 6448 720 6512 784
rect 6528 720 6592 784
rect 6608 720 6672 784
rect 6688 720 6752 784
rect 6288 632 6352 696
rect 6368 632 6432 696
rect 6448 632 6512 696
rect 6528 632 6592 696
rect 6608 632 6672 696
rect 6688 632 6752 696
rect 6288 544 6352 608
rect 6368 544 6432 608
rect 6448 544 6512 608
rect 6528 544 6592 608
rect 6608 544 6672 608
rect 6688 544 6752 608
rect 6288 455 6352 519
rect 6368 455 6432 519
rect 6448 455 6512 519
rect 6528 455 6592 519
rect 6608 455 6672 519
rect 6688 455 6752 519
rect 6288 366 6352 430
rect 6368 366 6432 430
rect 6448 366 6512 430
rect 6528 366 6592 430
rect 6608 366 6672 430
rect 6688 366 6752 430
rect 9429 -56 9493 8
rect 9509 -56 9573 8
rect 9589 -56 9653 8
rect 9669 -56 9733 8
rect 9749 -56 9813 8
rect 9829 -56 9893 8
rect 9429 -144 9493 -80
rect 9509 -144 9573 -80
rect 9589 -144 9653 -80
rect 9669 -144 9733 -80
rect 9749 -144 9813 -80
rect 9829 -144 9893 -80
rect 9429 -232 9493 -168
rect 9509 -232 9573 -168
rect 9589 -232 9653 -168
rect 9669 -232 9733 -168
rect 9749 -232 9813 -168
rect 9829 -232 9893 -168
rect 9429 -320 9493 -256
rect 9509 -320 9573 -256
rect 9589 -320 9653 -256
rect 9669 -320 9733 -256
rect 9749 -320 9813 -256
rect 9829 -320 9893 -256
rect 9429 -408 9493 -344
rect 9509 -408 9573 -344
rect 9589 -408 9653 -344
rect 9669 -408 9733 -344
rect 9749 -408 9813 -344
rect 9829 -408 9893 -344
rect 9429 -497 9493 -433
rect 9509 -497 9573 -433
rect 9589 -497 9653 -433
rect 9669 -497 9733 -433
rect 9749 -497 9813 -433
rect 9829 -497 9893 -433
rect 9429 -586 9493 -522
rect 9509 -586 9573 -522
rect 9589 -586 9653 -522
rect 9669 -586 9733 -522
rect 9749 -586 9813 -522
rect 9829 -586 9893 -522
rect 12970 3572 13034 3636
rect 13050 3572 13114 3636
rect 13118 2458 13182 2462
rect 13198 2458 13262 2462
rect 13118 2402 13170 2458
rect 13170 2402 13182 2458
rect 13198 2402 13250 2458
rect 13250 2402 13262 2458
rect 13118 2398 13182 2402
rect 13198 2398 13262 2402
rect 12969 2191 13033 2255
rect 13063 2191 13127 2255
rect 13157 2191 13221 2255
rect 13251 2191 13315 2255
rect 12969 2103 13033 2167
rect 13063 2103 13127 2167
rect 13157 2103 13221 2167
rect 13251 2103 13315 2167
rect 12969 2015 13033 2079
rect 13063 2015 13127 2079
rect 13157 2015 13221 2079
rect 13251 2015 13315 2079
rect 12969 1927 13033 1991
rect 13063 1927 13127 1991
rect 13157 1927 13221 1991
rect 13251 1927 13315 1991
rect 12969 1839 13033 1903
rect 13063 1839 13127 1903
rect 13157 1839 13221 1903
rect 13251 1839 13315 1903
rect 12969 1750 13033 1814
rect 13063 1750 13127 1814
rect 13157 1750 13221 1814
rect 13251 1750 13315 1814
rect 12969 1661 13033 1725
rect 13063 1661 13127 1725
rect 13157 1661 13221 1725
rect 13251 1661 13315 1725
rect 12969 1572 13033 1636
rect 13063 1572 13127 1636
rect 13157 1572 13221 1636
rect 13251 1572 13315 1636
rect 12969 1483 13033 1547
rect 13063 1483 13127 1547
rect 13157 1483 13221 1547
rect 13251 1483 13315 1547
rect 12969 1394 13033 1458
rect 13063 1394 13127 1458
rect 13157 1394 13221 1458
rect 13251 1394 13315 1458
<< metal4 >>
rect 2971 9884 3323 9885
rect 2971 9820 2974 9884
rect 3038 9820 3068 9884
rect 3132 9820 3162 9884
rect 3226 9820 3256 9884
rect 3320 9820 3323 9884
rect 2971 9798 3323 9820
rect 2971 9792 8650 9798
rect 2971 9728 2974 9792
rect 3038 9728 3068 9792
rect 3132 9728 3162 9792
rect 3226 9728 3256 9792
rect 3320 9728 8650 9792
rect 2971 9700 8650 9728
rect 2971 9636 2974 9700
rect 3038 9636 3068 9700
rect 3132 9636 3162 9700
rect 3226 9636 3256 9700
rect 3320 9636 8650 9700
rect 2971 9608 8650 9636
rect 2971 9544 2974 9608
rect 3038 9544 3068 9608
rect 3132 9544 3162 9608
rect 3226 9544 3256 9608
rect 3320 9544 8650 9608
rect 2971 9516 8650 9544
rect 2971 9452 2974 9516
rect 3038 9452 3068 9516
rect 3132 9452 3162 9516
rect 3226 9452 3256 9516
rect 3320 9452 8650 9516
rect 2971 9446 8650 9452
rect 2971 9423 3323 9446
rect 2971 9359 2974 9423
rect 3038 9359 3068 9423
rect 3132 9359 3162 9423
rect 3226 9359 3256 9423
rect 3320 9359 3323 9423
rect 2971 9358 3323 9359
rect 913 3636 13115 3637
rect 913 3572 914 3636
rect 978 3572 994 3636
rect 1058 3572 12970 3636
rect 13034 3572 13050 3636
rect 13114 3572 13115 3636
rect 913 3571 13115 3572
rect 1288 3443 1664 3444
rect 1288 3379 1291 3443
rect 1355 3379 1393 3443
rect 1457 3379 1495 3443
rect 1559 3379 1597 3443
rect 1661 3379 1664 3443
rect 1288 3363 1664 3379
rect 1288 3299 1291 3363
rect 1355 3299 1393 3363
rect 1457 3299 1495 3363
rect 1559 3299 1597 3363
rect 1661 3299 1664 3363
rect 1288 3283 1664 3299
rect 1288 3219 1291 3283
rect 1355 3219 1393 3283
rect 1457 3219 1495 3283
rect 1559 3219 1597 3283
rect 1661 3219 1664 3283
rect 1288 3202 1664 3219
rect 1288 3138 1291 3202
rect 1355 3138 1393 3202
rect 1457 3138 1495 3202
rect 1559 3138 1597 3202
rect 1661 3138 1664 3202
rect 1288 3121 1664 3138
rect 1288 3057 1291 3121
rect 1355 3057 1393 3121
rect 1457 3057 1495 3121
rect 1559 3057 1597 3121
rect 1661 3057 1664 3121
rect 1288 3040 1664 3057
rect 1288 2976 1291 3040
rect 1355 2976 1393 3040
rect 1457 2976 1495 3040
rect 1559 2976 1597 3040
rect 1661 2976 1664 3040
rect 1288 2959 1664 2976
rect 1288 2895 1291 2959
rect 1355 2895 1393 2959
rect 1457 2895 1495 2959
rect 1559 2895 1597 2959
rect 1661 2895 1664 2959
rect 1288 2878 1664 2895
rect 1288 2814 1291 2878
rect 1355 2814 1393 2878
rect 1457 2814 1495 2878
rect 1559 2814 1597 2878
rect 1661 2814 1664 2878
rect 1288 2797 1664 2814
rect 1288 2733 1291 2797
rect 1355 2733 1393 2797
rect 1457 2733 1495 2797
rect 1559 2733 1597 2797
rect 1661 2733 1664 2797
rect 1288 2716 1664 2733
rect 1288 2652 1291 2716
rect 1355 2652 1393 2716
rect 1457 2652 1495 2716
rect 1559 2652 1597 2716
rect 1661 2652 1664 2716
rect 1288 2635 1664 2652
rect 1288 2571 1291 2635
rect 1355 2571 1393 2635
rect 1457 2571 1495 2635
rect 1559 2571 1597 2635
rect 1661 2571 1664 2635
rect 1288 2570 1664 2571
rect 1044 2462 13269 2463
rect 1044 2398 1045 2462
rect 1109 2398 1125 2462
rect 1189 2398 13118 2462
rect 13182 2398 13198 2462
rect 13262 2398 13269 2462
rect 1044 2397 13269 2398
rect 12966 2255 13318 2256
rect 12966 2191 12969 2255
rect 13033 2191 13063 2255
rect 13127 2191 13157 2255
rect 13221 2191 13251 2255
rect 13315 2191 13318 2255
rect 12966 2167 13318 2191
rect 12966 2103 12969 2167
rect 13033 2103 13063 2167
rect 13127 2103 13157 2167
rect 13221 2103 13251 2167
rect 13315 2103 13318 2167
rect 12966 2079 13318 2103
rect 12966 2015 12969 2079
rect 13033 2015 13063 2079
rect 13127 2015 13157 2079
rect 13221 2015 13251 2079
rect 13315 2015 13318 2079
rect 12966 1991 13318 2015
rect 12966 1927 12969 1991
rect 13033 1927 13063 1991
rect 13127 1927 13157 1991
rect 13221 1927 13251 1991
rect 13315 1927 13318 1991
rect 12966 1903 13318 1927
rect 12966 1839 12969 1903
rect 13033 1839 13063 1903
rect 13127 1839 13157 1903
rect 13221 1839 13251 1903
rect 13315 1839 13318 1903
rect 12966 1814 13318 1839
rect 12966 1750 12969 1814
rect 13033 1750 13063 1814
rect 13127 1750 13157 1814
rect 13221 1750 13251 1814
rect 13315 1750 13318 1814
rect 12966 1725 13318 1750
rect 12966 1661 12969 1725
rect 13033 1661 13063 1725
rect 13127 1661 13157 1725
rect 13221 1661 13251 1725
rect 13315 1661 13318 1725
rect 12966 1636 13318 1661
rect 12966 1572 12969 1636
rect 13033 1572 13063 1636
rect 13127 1572 13157 1636
rect 13221 1572 13251 1636
rect 13315 1572 13318 1636
rect 12966 1547 13318 1572
rect 12966 1483 12969 1547
rect 13033 1483 13063 1547
rect 13127 1483 13157 1547
rect 13221 1483 13251 1547
rect 13315 1483 13318 1547
rect 12966 1458 13318 1483
rect 12966 1394 12969 1458
rect 13033 1394 13063 1458
rect 13127 1394 13157 1458
rect 13221 1394 13251 1458
rect 13315 1394 13318 1458
rect 12966 1393 13318 1394
rect 6285 960 6755 961
rect 6285 896 6288 960
rect 6352 896 6368 960
rect 6432 896 6448 960
rect 6512 896 6528 960
rect 6592 896 6608 960
rect 6672 896 6688 960
rect 6752 896 6755 960
rect 6285 872 6755 896
rect 6285 808 6288 872
rect 6352 808 6368 872
rect 6432 808 6448 872
rect 6512 808 6528 872
rect 6592 808 6608 872
rect 6672 808 6688 872
rect 6752 808 6755 872
rect 6285 784 6755 808
rect 6285 720 6288 784
rect 6352 720 6368 784
rect 6432 720 6448 784
rect 6512 720 6528 784
rect 6592 720 6608 784
rect 6672 720 6688 784
rect 6752 720 6755 784
rect 6285 696 6755 720
rect 6285 632 6288 696
rect 6352 632 6368 696
rect 6432 632 6448 696
rect 6512 632 6528 696
rect 6592 632 6608 696
rect 6672 632 6688 696
rect 6752 632 6755 696
rect 6285 608 6755 632
rect 6285 544 6288 608
rect 6352 544 6368 608
rect 6432 544 6448 608
rect 6512 544 6528 608
rect 6592 544 6608 608
rect 6672 544 6688 608
rect 6752 544 6755 608
rect 6285 519 6755 544
rect 6285 455 6288 519
rect 6352 455 6368 519
rect 6432 455 6448 519
rect 6512 455 6528 519
rect 6592 455 6608 519
rect 6672 455 6688 519
rect 6752 455 6755 519
rect 6285 430 6755 455
rect 6285 366 6288 430
rect 6352 366 6368 430
rect 6432 366 6448 430
rect 6512 366 6528 430
rect 6592 366 6608 430
rect 6672 366 6688 430
rect 6752 366 6755 430
rect 6285 365 6755 366
rect 9426 8 9896 9
rect 9426 -56 9429 8
rect 9493 -56 9509 8
rect 9573 -56 9589 8
rect 9653 -56 9669 8
rect 9733 -56 9749 8
rect 9813 -56 9829 8
rect 9893 -56 9896 8
rect 9426 -80 9896 -56
rect 9426 -144 9429 -80
rect 9493 -144 9509 -80
rect 9573 -144 9589 -80
rect 9653 -144 9669 -80
rect 9733 -144 9749 -80
rect 9813 -144 9829 -80
rect 9893 -144 9896 -80
rect 9426 -168 9896 -144
rect 9426 -232 9429 -168
rect 9493 -232 9509 -168
rect 9573 -232 9589 -168
rect 9653 -232 9669 -168
rect 9733 -232 9749 -168
rect 9813 -232 9829 -168
rect 9893 -232 9896 -168
rect 9426 -256 9896 -232
rect 9426 -320 9429 -256
rect 9493 -320 9509 -256
rect 9573 -320 9589 -256
rect 9653 -320 9669 -256
rect 9733 -320 9749 -256
rect 9813 -320 9829 -256
rect 9893 -320 9896 -256
rect 9426 -344 9896 -320
rect 9426 -408 9429 -344
rect 9493 -408 9509 -344
rect 9573 -408 9589 -344
rect 9653 -408 9669 -344
rect 9733 -408 9749 -344
rect 9813 -408 9829 -344
rect 9893 -408 9896 -344
rect 9426 -433 9896 -408
rect 9426 -497 9429 -433
rect 9493 -497 9509 -433
rect 9573 -497 9589 -433
rect 9653 -497 9669 -433
rect 9733 -497 9749 -433
rect 9813 -497 9829 -433
rect 9893 -497 9896 -433
rect 9426 -522 9896 -497
rect 9426 -586 9429 -522
rect 9493 -586 9509 -522
rect 9573 -586 9589 -522
rect 9653 -586 9669 -522
rect 9733 -586 9749 -522
rect 9813 -586 9829 -522
rect 9893 -586 9896 -522
rect 9426 -587 9896 -586
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_0
timestamp 1627201311
transform 1 0 3419 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_1
timestamp 1627201311
transform 1 0 2619 0 -1 6379
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_2
timestamp 1627201311
transform 1 0 2619 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_3
timestamp 1627201311
transform 1 0 3419 0 -1 6379
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_4
timestamp 1627201311
transform -1 0 8708 0 1 9409
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_5
timestamp 1627201311
transform 1 0 8626 0 1 9409
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_6
timestamp 1627201311
transform 0 1 12464 1 0 3136
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_7
timestamp 1627201311
transform 0 -1 12368 1 0 3136
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_8
timestamp 1627201311
transform 0 1 12464 -1 0 3218
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_9
timestamp 1627201311
transform 0 -1 11869 1 0 3136
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_10
timestamp 1627201311
transform -1 0 1901 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_11
timestamp 1627201311
transform -1 0 2701 0 -1 6879
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_12
timestamp 1627201311
transform -1 0 2701 0 -1 6379
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_13
timestamp 1627201311
transform -1 0 1901 0 -1 6379
box 0 0 882 404
use sky130_fd_pr__nfet_01v8__example_55959141808594  sky130_fd_pr__nfet_01v8__example_55959141808594_0
timestamp 1627201311
transform 0 -1 14630 -1 0 2528
box -28 0 2156 471
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_0
timestamp 1627201311
transform 1 0 13603 0 1 3415
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_1
timestamp 1627201311
transform 1 0 14151 0 1 3415
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_2
timestamp 1627201311
transform 1 0 14423 0 1 3415
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_55959141808593  sky130_fd_pr__nfet_01v8__example_55959141808593_3
timestamp 1627201311
transform 1 0 13875 0 1 3415
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_0
timestamp 1627201311
transform 1 0 14424 0 1 3035
box -28 0 128 29
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_1
timestamp 1627201311
transform 1 0 13880 0 1 3035
box -28 0 128 29
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_2
timestamp 1627201311
transform 1 0 13608 0 1 3035
box -28 0 128 29
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_3
timestamp 1627201311
transform 1 0 14152 0 1 3035
box -28 0 128 29
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_4
timestamp 1627201311
transform 1 0 13608 0 -1 3321
box -28 0 128 29
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_5
timestamp 1627201311
transform 1 0 14152 0 -1 3321
box -28 0 128 29
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_6
timestamp 1627201311
transform 1 0 14424 0 -1 3321
box -28 0 128 29
use sky130_fd_pr__nfet_01v8__example_55959141808592  sky130_fd_pr__nfet_01v8__example_55959141808592_7
timestamp 1627201311
transform 1 0 13880 0 -1 3321
box -28 0 128 29
use sky130_fd_pr__pfet_01v8__example_55959141808591  sky130_fd_pr__pfet_01v8__example_55959141808591_0
timestamp 1627201311
transform 0 1 1282 -1 0 8427
box -28 0 1064 1491
use sky130_fd_io__gpiov2_amux_ctl_logic  sky130_fd_io__gpiov2_amux_ctl_logic_0
timestamp 1627201311
transform 1 0 -26998 0 1 6306
box 25855 -16459 42060 1976
use sky130_fd_io__amux_switch_1v2b  sky130_fd_io__amux_switch_1v2b_0
timestamp 1627201311
transform 1 0 4755 0 -1 8802
box -50 -73 10379 2429
use sky130_fd_io__amux_switch_1v2b  sky130_fd_io__amux_switch_1v2b_1
timestamp 1627201311
transform 1 0 4755 0 1 4180
box -50 -73 10379 2429
<< labels >>
flabel metal4 s 8389 9734 8389 9734 0 FreeSans 440 0 0 0 PAD
port 1 nsew
flabel locali s 2651 6421 2651 6421 0 FreeSans 440 0 0 0 PAD
port 1 nsew
flabel locali s 8640 9507 8736 9716 3 FreeSans 520 0 0 0 PAD
port 1 nsew
flabel metal2 s 7812 5145 9070 5412 3 FreeSans 520 0 0 0 AMUXBUS_B
port 2 nsew
flabel metal2 s 7824 7592 8467 7821 3 FreeSans 520 0 0 0 AMUXBUS_A
port 3 nsew
flabel metal1 s 1166 8058 1194 8086 3 FreeSans 520 0 0 0 VDDIO_Q
port 4 nsew
flabel metal1 s 11819 3200 11819 3200 0 FreeSans 440 0 0 0 VSSA
port 5 nsew
flabel metal1 s 13265 -8570 13293 -8542 3 FreeSans 520 0 0 0 VCCD
port 6 nsew
flabel metal1 s 8575 8695 8603 8723 3 FreeSans 520 0 0 0 VDDA
port 7 nsew
flabel metal1 s 4964 8043 4992 8071 3 FreeSans 520 0 0 0 VDDIO_Q
port 4 nsew
flabel metal1 s 14310 1324 14562 1760 3 FreeSans 520 0 0 0 VSSIO_Q
port 8 nsew
flabel metal1 s 8762 2572 8790 2600 3 FreeSans 520 0 0 0 OUT
port 9 nsew
flabel metal1 s 13634 -7974 13662 -7946 3 FreeSans 520 180 0 0 HLD_I_H_N
port 10 nsew
flabel metal1 s 14429 -7926 14457 -7898 3 FreeSans 520 180 0 0 HLD_I_H
port 11 nsew
flabel metal1 s 2154 1374 2182 1402 3 FreeSans 520 0 0 0 ENABLE_VSWITCH_H
port 12 nsew
flabel metal1 s 434 5213 462 5241 3 FreeSans 520 0 0 0 ENABLE_VDDA_H
port 13 nsew
flabel metal1 s 5210 3259 5238 3287 3 FreeSans 520 0 0 0 ANALOG_SEL
port 14 nsew
flabel metal1 s 8762 3259 8790 3287 3 FreeSans 520 0 0 0 ANALOG_POL
port 15 nsew
flabel metal1 s 6754 2593 6782 2621 3 FreeSans 520 0 0 0 ANALOG_EN
port 16 nsew
flabel metal1 s 13244 -8912 13272 -8884 3 FreeSans 520 0 0 0 ANALOG_EN
port 16 nsew
flabel metal1 s 328 2480 356 2508 3 FreeSans 520 0 0 0 VSWITCH
port 17 nsew
flabel metal1 s 14072 -8266 14100 -8238 3 FreeSans 280 0 0 0 VSSD
port 18 nsew
flabel metal1 s 13347 -9239 13375 -9211 3 FreeSans 280 180 0 0 VSSD
port 18 nsew
flabel metal1 s -76 -954 -48 -926 3 FreeSans 520 0 0 0 VSSD
port 18 nsew
flabel metal1 s 5825 1210 5853 1238 3 FreeSans 520 0 0 0 VSSD
port 18 nsew
flabel metal1 s 13361 -9225 13361 -9225 3 FreeSans 520 0 0 0 VSSD
port 18 nsew
flabel metal1 s -768 5488 -740 5516 3 FreeSans 520 0 0 0 VSSA
port 5 nsew
flabel metal1 s -225 1614 -197 1642 3 FreeSans 520 0 0 0 VSSA
port 5 nsew
flabel metal1 s 1940 1748 1968 1776 3 FreeSans 520 0 0 0 VSSA
port 5 nsew
flabel metal1 s 470 4570 498 4598 3 FreeSans 520 0 0 0 VSSA
port 5 nsew
flabel metal1 s -228 5437 -200 5465 3 FreeSans 520 0 0 0 VSSA
port 5 nsew
flabel metal1 s 1365 5487 1393 5515 3 FreeSans 520 0 0 0 VSSA
port 5 nsew
flabel metal1 s 1789 4559 1817 4587 3 FreeSans 520 0 0 0 VSSA
port 5 nsew
flabel metal1 s 1789 3124 1817 3152 3 FreeSans 520 0 0 0 VSSA
port 5 nsew
flabel metal1 s -214 5451 -214 5451 3 FreeSans 520 0 0 0 VSSA
port 5 nsew
flabel metal1 s 13260 -7040 13288 -7012 3 FreeSans 520 180 0 0 VDDIO_Q
port 4 nsew
flabel metal1 s 9628 838 9656 866 3 FreeSans 520 0 0 0 VDDIO_Q
port 4 nsew
flabel metal1 s -702 7906 -674 7934 3 FreeSans 520 0 0 0 VDDA
port 7 nsew
flabel metal1 s 6886 2928 6914 2956 3 FreeSans 520 0 0 0 VCCD
port 6 nsew
flabel comment s 14051 274 14051 274 0 FreeSans 440 0 0 0 CONDIODE
flabel comment s -796 3405 -796 3405 0 FreeSans 440 90 0 0 CONDIODE
flabel comment s 14233 4211 14233 4211 0 FreeSans 440 0 0 0 CONDIODE
flabel comment s -276 1601 -276 1601 0 FreeSans 440 90 0 0 CONDIODE
flabel comment s 3163 2234 3163 2234 0 FreeSans 440 0 0 0 CONDIODE
flabel comment s 14263 2739 14263 2739 0 FreeSans 440 0 0 0 CONDIODE
flabel comment s 13455 4177 13455 4177 0 FreeSans 440 0 0 0 NMIDA_VCCD
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 25932566
string GDS_START 25415808
<< end >>
