magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 1 49 724 157
rect 0 0 768 49
<< scnmos >>
rect 80 47 110 131
rect 285 47 315 131
rect 357 47 387 131
rect 429 47 459 131
rect 515 47 545 131
rect 615 47 645 131
<< scpmoshvt >>
rect 129 481 159 609
rect 229 481 259 609
rect 315 481 345 609
rect 469 481 499 609
rect 555 481 585 609
rect 627 481 657 609
<< ndiff >>
rect 27 106 80 131
rect 27 72 35 106
rect 69 72 80 106
rect 27 47 80 72
rect 110 106 163 131
rect 110 72 121 106
rect 155 72 163 106
rect 110 47 163 72
rect 232 106 285 131
rect 232 72 240 106
rect 274 72 285 106
rect 232 47 285 72
rect 315 47 357 131
rect 387 47 429 131
rect 459 106 515 131
rect 459 72 470 106
rect 504 72 515 106
rect 459 47 515 72
rect 545 99 615 131
rect 545 65 563 99
rect 597 65 615 99
rect 545 47 615 65
rect 645 106 698 131
rect 645 72 656 106
rect 690 72 698 106
rect 645 47 698 72
<< pdiff >>
rect 76 597 129 609
rect 76 563 84 597
rect 118 563 129 597
rect 76 527 129 563
rect 76 493 84 527
rect 118 493 129 527
rect 76 481 129 493
rect 159 597 229 609
rect 159 563 177 597
rect 211 563 229 597
rect 159 527 229 563
rect 159 493 177 527
rect 211 493 229 527
rect 159 481 229 493
rect 259 599 315 609
rect 259 565 270 599
rect 304 565 315 599
rect 259 527 315 565
rect 259 493 270 527
rect 304 493 315 527
rect 259 481 315 493
rect 345 597 469 609
rect 345 563 356 597
rect 390 563 424 597
rect 458 563 469 597
rect 345 527 469 563
rect 345 493 356 527
rect 390 493 424 527
rect 458 493 469 527
rect 345 481 469 493
rect 499 599 555 609
rect 499 565 510 599
rect 544 565 555 599
rect 499 527 555 565
rect 499 493 510 527
rect 544 493 555 527
rect 499 481 555 493
rect 585 481 627 609
rect 657 597 710 609
rect 657 563 668 597
rect 702 563 710 597
rect 657 527 710 563
rect 657 493 668 527
rect 702 493 710 527
rect 657 481 710 493
<< ndiffc >>
rect 35 72 69 106
rect 121 72 155 106
rect 240 72 274 106
rect 470 72 504 106
rect 563 65 597 99
rect 656 72 690 106
<< pdiffc >>
rect 84 563 118 597
rect 84 493 118 527
rect 177 563 211 597
rect 177 493 211 527
rect 270 565 304 599
rect 270 493 304 527
rect 356 563 390 597
rect 424 563 458 597
rect 356 493 390 527
rect 424 493 458 527
rect 510 565 544 599
rect 510 493 544 527
rect 668 563 702 597
rect 668 493 702 527
<< poly >>
rect 129 609 159 635
rect 229 609 259 635
rect 315 609 345 635
rect 469 609 499 635
rect 555 609 585 635
rect 627 609 657 635
rect 129 443 159 481
rect 80 427 159 443
rect 80 393 109 427
rect 143 393 159 427
rect 80 359 159 393
rect 80 325 109 359
rect 143 325 159 359
rect 229 350 259 481
rect 315 365 345 481
rect 469 373 499 481
rect 80 309 159 325
rect 207 334 273 350
rect 80 131 110 309
rect 207 300 223 334
rect 257 300 273 334
rect 207 266 273 300
rect 207 232 223 266
rect 257 232 273 266
rect 207 216 273 232
rect 315 349 387 365
rect 315 315 337 349
rect 371 315 387 349
rect 315 281 387 315
rect 315 247 337 281
rect 371 247 387 281
rect 315 231 387 247
rect 243 183 273 216
rect 243 153 315 183
rect 285 131 315 153
rect 357 131 387 231
rect 429 357 501 373
rect 555 365 585 481
rect 627 443 657 481
rect 627 413 693 443
rect 429 323 451 357
rect 485 323 501 357
rect 429 289 501 323
rect 429 255 451 289
rect 485 255 501 289
rect 429 239 501 255
rect 543 349 609 365
rect 543 315 559 349
rect 593 315 609 349
rect 543 281 609 315
rect 543 247 559 281
rect 593 247 609 281
rect 429 131 459 239
rect 543 231 609 247
rect 663 325 693 413
rect 663 309 743 325
rect 663 275 693 309
rect 727 275 743 309
rect 663 241 743 275
rect 543 183 573 231
rect 663 207 693 241
rect 727 207 743 241
rect 663 191 743 207
rect 663 183 693 191
rect 515 153 573 183
rect 615 153 693 183
rect 515 131 545 153
rect 615 131 645 153
rect 80 21 110 47
rect 285 21 315 47
rect 357 21 387 47
rect 429 21 459 47
rect 515 21 545 47
rect 615 21 645 47
<< polycont >>
rect 109 393 143 427
rect 109 325 143 359
rect 223 300 257 334
rect 223 232 257 266
rect 337 315 371 349
rect 337 247 371 281
rect 451 323 485 357
rect 451 255 485 289
rect 559 315 593 349
rect 559 247 593 281
rect 693 275 727 309
rect 693 207 727 241
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 17 597 134 613
rect 17 563 84 597
rect 118 563 134 597
rect 17 527 134 563
rect 17 493 84 527
rect 118 493 134 527
rect 17 477 134 493
rect 168 597 227 649
rect 168 563 177 597
rect 211 563 227 597
rect 168 527 227 563
rect 168 493 177 527
rect 211 493 227 527
rect 168 477 227 493
rect 261 599 314 615
rect 261 565 270 599
rect 304 565 314 599
rect 261 527 314 565
rect 261 493 270 527
rect 304 493 314 527
rect 17 106 71 477
rect 261 443 314 493
rect 348 597 468 649
rect 348 563 356 597
rect 390 563 424 597
rect 458 563 468 597
rect 348 527 468 563
rect 348 493 356 527
rect 390 493 424 527
rect 458 493 468 527
rect 348 477 468 493
rect 502 599 560 615
rect 502 565 510 599
rect 544 565 560 599
rect 502 527 560 565
rect 502 493 510 527
rect 544 493 560 527
rect 502 443 560 493
rect 652 597 718 649
rect 652 563 668 597
rect 702 563 718 597
rect 652 527 718 563
rect 652 493 668 527
rect 702 493 718 527
rect 652 477 718 493
rect 105 427 560 443
rect 105 393 109 427
rect 143 407 560 427
rect 143 393 159 407
rect 105 359 159 393
rect 105 325 109 359
rect 143 325 159 359
rect 105 182 159 325
rect 207 334 272 373
rect 207 300 223 334
rect 257 300 272 334
rect 207 266 272 300
rect 207 232 223 266
rect 257 232 272 266
rect 207 216 272 232
rect 309 349 371 373
rect 309 315 337 349
rect 309 281 371 315
rect 309 247 337 281
rect 105 148 275 182
rect 17 72 35 106
rect 69 72 71 106
rect 17 53 71 72
rect 105 106 171 114
rect 105 72 121 106
rect 155 72 171 106
rect 105 17 171 72
rect 224 106 275 148
rect 224 72 240 106
rect 274 72 275 106
rect 309 75 371 247
rect 405 357 502 373
rect 405 323 451 357
rect 485 323 502 357
rect 405 289 502 323
rect 405 255 451 289
rect 485 255 502 289
rect 405 228 502 255
rect 543 349 643 365
rect 543 315 559 349
rect 593 315 643 349
rect 543 281 643 315
rect 543 247 559 281
rect 593 247 643 281
rect 543 228 643 247
rect 677 309 751 440
rect 677 275 693 309
rect 727 275 751 309
rect 677 241 751 275
rect 677 207 693 241
rect 727 207 751 241
rect 454 139 706 173
rect 454 106 513 139
rect 224 56 275 72
rect 454 72 470 106
rect 504 72 513 106
rect 650 106 706 139
rect 454 56 513 72
rect 547 99 613 105
rect 547 65 563 99
rect 597 65 613 99
rect 547 17 613 65
rect 650 72 656 106
rect 690 72 706 106
rect 650 56 706 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2111a_0
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4258612
string GDS_START 4249726
<< end >>
