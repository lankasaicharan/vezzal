magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4466 1975
<< nwell >>
rect -38 415 3206 704
rect -38 331 2264 415
rect 2518 331 3206 415
rect 2518 321 2874 331
<< pwell >>
rect 2354 241 2476 329
rect 2866 241 3164 247
rect 13 216 585 229
rect 13 211 865 216
rect 2354 211 3164 241
rect 13 157 1117 211
rect 1765 201 3164 211
rect 1379 157 3164 201
rect 13 49 3164 157
rect 0 0 3168 49
<< scnmos >>
rect 96 119 126 203
rect 174 119 204 203
rect 260 119 290 203
rect 332 119 362 203
rect 472 119 502 203
rect 725 106 755 190
rect 950 101 980 185
rect 1202 47 1232 131
rect 1288 47 1318 131
rect 1360 47 1390 131
rect 1462 47 1492 175
rect 1548 47 1578 175
rect 1650 47 1680 175
rect 1850 57 1880 185
rect 1934 57 1964 185
rect 2036 101 2066 185
rect 2114 101 2144 185
rect 2249 57 2279 185
rect 2335 57 2365 185
rect 2455 57 2485 185
rect 2649 131 2679 215
rect 2751 47 2781 215
rect 2949 137 2979 221
rect 3051 53 3081 221
<< scpmoshvt >>
rect 84 481 114 609
rect 194 481 224 609
rect 272 481 302 609
rect 358 481 388 609
rect 572 481 602 609
rect 770 474 800 602
rect 968 457 998 585
rect 1186 457 1216 541
rect 1272 457 1302 541
rect 1350 457 1380 541
rect 1468 373 1498 541
rect 1554 373 1584 541
rect 1650 373 1680 541
rect 1736 373 1766 541
rect 1831 431 1861 599
rect 1933 515 1963 599
rect 2064 515 2094 599
rect 2263 451 2293 619
rect 2365 451 2395 619
rect 2449 451 2479 619
rect 2649 357 2679 485
rect 2751 357 2781 609
rect 2949 367 2979 495
rect 3051 367 3081 619
<< ndiff >>
rect 39 178 96 203
rect 39 144 51 178
rect 85 144 96 178
rect 39 119 96 144
rect 126 119 174 203
rect 204 178 260 203
rect 204 144 215 178
rect 249 144 260 178
rect 204 119 260 144
rect 290 119 332 203
rect 362 174 472 203
rect 362 140 373 174
rect 407 140 472 174
rect 362 119 472 140
rect 502 182 559 203
rect 502 148 513 182
rect 547 148 559 182
rect 502 119 559 148
rect 641 165 725 190
rect 641 131 653 165
rect 687 131 725 165
rect 641 106 725 131
rect 755 175 839 190
rect 755 141 793 175
rect 827 141 839 175
rect 755 106 839 141
rect 893 173 950 185
rect 893 139 905 173
rect 939 139 950 173
rect 893 101 950 139
rect 980 114 1091 185
rect 2380 291 2450 303
rect 2380 257 2404 291
rect 2438 257 2450 291
rect 2380 245 2450 257
rect 2380 185 2440 245
rect 1405 131 1462 175
rect 980 101 1045 114
rect 995 80 1045 101
rect 1079 80 1091 114
rect 995 68 1091 80
rect 1145 111 1202 131
rect 1145 77 1157 111
rect 1191 77 1202 111
rect 1145 47 1202 77
rect 1232 111 1288 131
rect 1232 77 1243 111
rect 1277 77 1288 111
rect 1232 47 1288 77
rect 1318 47 1360 131
rect 1390 123 1462 131
rect 1390 89 1417 123
rect 1451 89 1462 123
rect 1390 47 1462 89
rect 1492 128 1548 175
rect 1492 94 1503 128
rect 1537 94 1548 128
rect 1492 47 1548 94
rect 1578 163 1650 175
rect 1578 129 1605 163
rect 1639 129 1650 163
rect 1578 47 1650 129
rect 1680 93 1737 175
rect 1680 59 1691 93
rect 1725 59 1737 93
rect 1680 47 1737 59
rect 1791 111 1850 185
rect 1791 77 1803 111
rect 1837 77 1850 111
rect 1791 57 1850 77
rect 1880 57 1934 185
rect 1964 173 2036 185
rect 1964 139 1975 173
rect 2009 139 2036 173
rect 1964 101 2036 139
rect 2066 101 2114 185
rect 2144 125 2249 185
rect 2144 101 2188 125
rect 1964 57 2021 101
rect 2176 91 2188 101
rect 2222 91 2249 125
rect 2176 57 2249 91
rect 2279 108 2335 185
rect 2279 74 2290 108
rect 2324 74 2335 108
rect 2279 57 2335 74
rect 2365 57 2455 185
rect 2485 108 2538 185
rect 2592 180 2649 215
rect 2592 146 2604 180
rect 2638 146 2649 180
rect 2592 131 2649 146
rect 2679 184 2751 215
rect 2679 150 2706 184
rect 2740 150 2751 184
rect 2679 131 2751 150
rect 2485 74 2496 108
rect 2530 74 2538 108
rect 2485 57 2538 74
rect 2694 93 2751 131
rect 2694 59 2706 93
rect 2740 59 2751 93
rect 2694 47 2751 59
rect 2781 199 2838 215
rect 2781 165 2792 199
rect 2826 165 2838 199
rect 2781 103 2838 165
rect 2892 196 2949 221
rect 2892 162 2904 196
rect 2938 162 2949 196
rect 2892 137 2949 162
rect 2979 209 3051 221
rect 2979 175 3006 209
rect 3040 175 3051 209
rect 2979 137 3051 175
rect 2781 69 2792 103
rect 2826 69 2838 103
rect 2781 47 2838 69
rect 2994 99 3051 137
rect 2994 65 3006 99
rect 3040 65 3051 99
rect 2994 53 3051 65
rect 3081 209 3138 221
rect 3081 175 3092 209
rect 3126 175 3138 209
rect 3081 103 3138 175
rect 3081 69 3092 103
rect 3126 69 3138 103
rect 3081 53 3138 69
<< pdiff >>
rect 27 597 84 609
rect 27 563 39 597
rect 73 563 84 597
rect 27 527 84 563
rect 27 493 39 527
rect 73 493 84 527
rect 27 481 84 493
rect 114 565 194 609
rect 114 531 141 565
rect 175 531 194 565
rect 114 481 194 531
rect 224 481 272 609
rect 302 527 358 609
rect 302 493 313 527
rect 347 493 358 527
rect 302 481 358 493
rect 388 597 461 609
rect 388 563 415 597
rect 449 563 461 597
rect 388 527 461 563
rect 388 493 415 527
rect 449 493 461 527
rect 388 481 461 493
rect 515 597 572 609
rect 515 563 527 597
rect 561 563 572 597
rect 515 527 572 563
rect 515 493 527 527
rect 561 493 572 527
rect 515 481 572 493
rect 602 597 659 609
rect 602 563 613 597
rect 647 563 659 597
rect 602 527 659 563
rect 602 493 613 527
rect 647 493 659 527
rect 602 481 659 493
rect 713 590 770 602
rect 713 556 725 590
rect 759 556 770 590
rect 713 520 770 556
rect 713 486 725 520
rect 759 486 770 520
rect 713 474 770 486
rect 800 590 857 602
rect 800 556 811 590
rect 845 556 857 590
rect 800 520 857 556
rect 800 486 811 520
rect 845 486 857 520
rect 800 474 857 486
rect 911 573 968 585
rect 911 539 923 573
rect 957 539 968 573
rect 911 503 968 539
rect 911 469 923 503
rect 957 469 968 503
rect 911 457 968 469
rect 998 573 1071 585
rect 998 539 1025 573
rect 1059 539 1071 573
rect 2206 599 2263 619
rect 1395 586 1453 598
rect 1395 552 1407 586
rect 1441 552 1453 586
rect 1395 541 1453 552
rect 1781 541 1831 599
rect 998 503 1071 539
rect 998 469 1025 503
rect 1059 469 1071 503
rect 998 457 1071 469
rect 1129 516 1186 541
rect 1129 482 1141 516
rect 1175 482 1186 516
rect 1129 457 1186 482
rect 1216 516 1272 541
rect 1216 482 1227 516
rect 1261 482 1272 516
rect 1216 457 1272 482
rect 1302 457 1350 541
rect 1380 457 1468 541
rect 1395 373 1468 457
rect 1498 529 1554 541
rect 1498 495 1509 529
rect 1543 495 1554 529
rect 1498 442 1554 495
rect 1498 408 1509 442
rect 1543 408 1554 442
rect 1498 373 1554 408
rect 1584 373 1650 541
rect 1680 520 1736 541
rect 1680 486 1691 520
rect 1725 486 1736 520
rect 1680 373 1736 486
rect 1766 431 1831 541
rect 1861 578 1933 599
rect 1861 544 1872 578
rect 1906 544 1933 578
rect 1861 515 1933 544
rect 1963 515 2064 599
rect 2094 596 2263 599
rect 2094 562 2218 596
rect 2252 562 2263 596
rect 2094 515 2263 562
rect 1861 431 1918 515
rect 1766 373 1816 431
rect 2206 451 2263 515
rect 2293 597 2365 619
rect 2293 563 2320 597
rect 2354 563 2365 597
rect 2293 516 2365 563
rect 2293 482 2320 516
rect 2354 482 2365 516
rect 2293 451 2365 482
rect 2395 451 2449 619
rect 2479 596 2536 619
rect 2479 562 2490 596
rect 2524 562 2536 596
rect 2479 451 2536 562
rect 2694 591 2751 609
rect 2694 557 2706 591
rect 2740 557 2751 591
rect 2694 485 2751 557
rect 2592 416 2649 485
rect 2592 382 2604 416
rect 2638 382 2649 416
rect 2592 357 2649 382
rect 2679 357 2751 485
rect 2781 597 2838 609
rect 2781 563 2792 597
rect 2826 563 2838 597
rect 2781 500 2838 563
rect 2994 607 3051 619
rect 2994 573 3006 607
rect 3040 573 3051 607
rect 2781 466 2792 500
rect 2826 466 2838 500
rect 2994 510 3051 573
rect 2994 495 3006 510
rect 2781 403 2838 466
rect 2781 369 2792 403
rect 2826 369 2838 403
rect 2781 357 2838 369
rect 2892 483 2949 495
rect 2892 449 2904 483
rect 2938 449 2949 483
rect 2892 413 2949 449
rect 2892 379 2904 413
rect 2938 379 2949 413
rect 2892 367 2949 379
rect 2979 476 3006 495
rect 3040 476 3051 510
rect 2979 413 3051 476
rect 2979 379 3006 413
rect 3040 379 3051 413
rect 2979 367 3051 379
rect 3081 597 3138 619
rect 3081 563 3092 597
rect 3126 563 3138 597
rect 3081 505 3138 563
rect 3081 471 3092 505
rect 3126 471 3138 505
rect 3081 413 3138 471
rect 3081 379 3092 413
rect 3126 379 3138 413
rect 3081 367 3138 379
<< ndiffc >>
rect 51 144 85 178
rect 215 144 249 178
rect 373 140 407 174
rect 513 148 547 182
rect 653 131 687 165
rect 793 141 827 175
rect 905 139 939 173
rect 2404 257 2438 291
rect 1045 80 1079 114
rect 1157 77 1191 111
rect 1243 77 1277 111
rect 1417 89 1451 123
rect 1503 94 1537 128
rect 1605 129 1639 163
rect 1691 59 1725 93
rect 1803 77 1837 111
rect 1975 139 2009 173
rect 2188 91 2222 125
rect 2290 74 2324 108
rect 2604 146 2638 180
rect 2706 150 2740 184
rect 2496 74 2530 108
rect 2706 59 2740 93
rect 2792 165 2826 199
rect 2904 162 2938 196
rect 3006 175 3040 209
rect 2792 69 2826 103
rect 3006 65 3040 99
rect 3092 175 3126 209
rect 3092 69 3126 103
<< pdiffc >>
rect 39 563 73 597
rect 39 493 73 527
rect 141 531 175 565
rect 313 493 347 527
rect 415 563 449 597
rect 415 493 449 527
rect 527 563 561 597
rect 527 493 561 527
rect 613 563 647 597
rect 613 493 647 527
rect 725 556 759 590
rect 725 486 759 520
rect 811 556 845 590
rect 811 486 845 520
rect 923 539 957 573
rect 923 469 957 503
rect 1025 539 1059 573
rect 1407 552 1441 586
rect 1025 469 1059 503
rect 1141 482 1175 516
rect 1227 482 1261 516
rect 1509 495 1543 529
rect 1509 408 1543 442
rect 1691 486 1725 520
rect 1872 544 1906 578
rect 2218 562 2252 596
rect 2320 563 2354 597
rect 2320 482 2354 516
rect 2490 562 2524 596
rect 2706 557 2740 591
rect 2604 382 2638 416
rect 2792 563 2826 597
rect 3006 573 3040 607
rect 2792 466 2826 500
rect 2792 369 2826 403
rect 2904 449 2938 483
rect 2904 379 2938 413
rect 3006 476 3040 510
rect 3006 379 3040 413
rect 3092 563 3126 597
rect 3092 471 3126 505
rect 3092 379 3126 413
<< poly >>
rect 84 609 114 635
rect 194 609 224 635
rect 272 609 302 635
rect 358 609 388 635
rect 572 609 602 635
rect 770 602 800 628
rect 968 615 1861 645
rect 84 454 114 481
rect 80 424 114 454
rect 194 449 224 481
rect 80 377 110 424
rect 44 361 110 377
rect 188 419 224 449
rect 188 376 218 419
rect 44 327 60 361
rect 94 327 110 361
rect 44 293 110 327
rect 152 360 218 376
rect 272 371 302 481
rect 358 449 388 481
rect 572 449 602 481
rect 968 585 998 615
rect 358 419 430 449
rect 572 419 609 449
rect 770 434 800 474
rect 1186 541 1216 567
rect 1272 541 1302 615
rect 1831 599 1861 615
rect 1933 599 1963 625
rect 2064 599 2094 625
rect 2263 619 2293 645
rect 2365 619 2395 645
rect 2449 619 2479 645
rect 1350 541 1380 567
rect 1468 541 1498 567
rect 1554 541 1584 567
rect 1650 541 1680 567
rect 1736 541 1766 567
rect 400 371 430 419
rect 152 326 168 360
rect 202 326 218 360
rect 152 310 218 326
rect 260 355 358 371
rect 260 321 308 355
rect 342 321 358 355
rect 44 259 60 293
rect 94 262 110 293
rect 94 259 126 262
rect 44 232 126 259
rect 96 203 126 232
rect 174 203 204 310
rect 260 305 358 321
rect 400 355 531 371
rect 400 321 481 355
rect 515 321 531 355
rect 400 305 531 321
rect 260 203 290 305
rect 400 248 430 305
rect 579 248 609 419
rect 689 418 800 434
rect 689 384 705 418
rect 739 404 800 418
rect 739 384 755 404
rect 689 350 755 384
rect 689 316 705 350
rect 739 316 755 350
rect 689 300 755 316
rect 332 218 430 248
rect 472 218 609 248
rect 332 203 362 218
rect 472 203 502 218
rect 725 190 755 300
rect 803 330 869 346
rect 803 296 819 330
rect 853 296 869 330
rect 803 262 869 296
rect 803 228 819 262
rect 853 235 869 262
rect 968 235 998 457
rect 1046 401 1112 417
rect 1046 367 1062 401
rect 1096 367 1112 401
rect 1046 333 1112 367
rect 1046 299 1062 333
rect 1096 313 1112 333
rect 1186 313 1216 457
rect 1272 431 1302 457
rect 1350 356 1380 457
rect 1933 491 1963 515
rect 1933 467 2016 491
rect 1933 461 1966 467
rect 1950 433 1966 461
rect 2000 433 2016 467
rect 2064 483 2094 515
rect 2064 467 2174 483
rect 2064 453 2124 467
rect 1831 413 1861 431
rect 1950 417 2016 433
rect 2108 433 2124 453
rect 2158 433 2174 467
rect 2751 609 2781 635
rect 3051 619 3081 645
rect 2649 485 2679 511
rect 1831 383 1908 413
rect 1096 299 1216 313
rect 1046 283 1216 299
rect 1297 340 1380 356
rect 1468 341 1498 373
rect 1297 306 1313 340
rect 1347 320 1380 340
rect 1432 325 1498 341
rect 1554 339 1584 373
rect 1347 306 1390 320
rect 1297 290 1390 306
rect 1186 248 1216 283
rect 1186 242 1304 248
rect 853 228 1136 235
rect 803 205 1136 228
rect 1186 218 1318 242
rect 1274 212 1318 218
rect 96 93 126 119
rect 174 51 204 119
rect 260 93 290 119
rect 332 93 362 119
rect 472 51 502 119
rect 950 185 980 205
rect 725 80 755 106
rect 1106 176 1136 205
rect 1106 146 1232 176
rect 1202 131 1232 146
rect 1288 131 1318 212
rect 1360 131 1390 290
rect 1432 291 1448 325
rect 1482 291 1498 325
rect 1432 275 1498 291
rect 1540 323 1606 339
rect 1540 289 1556 323
rect 1590 289 1606 323
rect 1462 175 1492 275
rect 1540 255 1606 289
rect 1540 221 1556 255
rect 1590 221 1606 255
rect 1540 205 1606 221
rect 1650 263 1680 373
rect 1736 335 1766 373
rect 1878 369 1908 383
rect 2108 399 2174 433
rect 2263 419 2293 451
rect 1878 339 2066 369
rect 2108 365 2124 399
rect 2158 365 2174 399
rect 2108 349 2174 365
rect 2216 403 2293 419
rect 2365 409 2395 451
rect 2216 369 2232 403
rect 2266 389 2293 403
rect 2335 393 2401 409
rect 2266 369 2282 389
rect 2216 353 2282 369
rect 2335 359 2351 393
rect 2385 359 2401 393
rect 1736 305 1836 335
rect 1806 291 1836 305
rect 1806 275 1880 291
rect 1650 247 1764 263
rect 1650 213 1714 247
rect 1748 213 1764 247
rect 1806 241 1822 275
rect 1856 241 1880 275
rect 1806 225 1880 241
rect 1922 275 1988 291
rect 1922 241 1938 275
rect 1972 241 1988 275
rect 1922 225 1988 241
rect 1548 175 1578 205
rect 1650 197 1764 213
rect 1650 175 1680 197
rect 1850 185 1880 225
rect 1934 185 1964 225
rect 2036 185 2066 339
rect 2114 185 2144 349
rect 2249 185 2279 353
rect 2335 341 2401 359
rect 2449 387 2479 451
rect 2449 371 2560 387
rect 2449 357 2510 371
rect 2335 185 2365 341
rect 2494 337 2510 357
rect 2544 337 2560 371
rect 2949 495 2979 521
rect 2494 303 2560 337
rect 2649 303 2679 357
rect 2751 317 2781 357
rect 2494 269 2510 303
rect 2544 269 2560 303
rect 2494 253 2560 269
rect 2613 287 2679 303
rect 2613 253 2629 287
rect 2663 253 2679 287
rect 2494 230 2524 253
rect 2613 237 2679 253
rect 2727 301 2793 317
rect 2727 267 2743 301
rect 2777 281 2793 301
rect 2949 281 2979 367
rect 3051 327 3081 367
rect 2777 267 2979 281
rect 2727 251 2979 267
rect 3021 311 3087 327
rect 3021 277 3037 311
rect 3071 277 3087 311
rect 3021 261 3087 277
rect 2455 200 2524 230
rect 2649 215 2679 237
rect 2751 215 2781 251
rect 2949 221 2979 251
rect 3051 221 3081 261
rect 2455 185 2485 200
rect 950 75 980 101
rect 174 21 502 51
rect 2036 75 2066 101
rect 2114 75 2144 101
rect 2649 105 2679 131
rect 1202 21 1232 47
rect 1288 21 1318 47
rect 1360 21 1390 47
rect 1462 21 1492 47
rect 1548 21 1578 47
rect 1650 21 1680 47
rect 1850 31 1880 57
rect 1934 31 1964 57
rect 2249 31 2279 57
rect 2335 31 2365 57
rect 2455 31 2485 57
rect 2949 111 2979 137
rect 2751 21 2781 47
rect 3051 27 3081 53
<< polycont >>
rect 60 327 94 361
rect 168 326 202 360
rect 308 321 342 355
rect 60 259 94 293
rect 481 321 515 355
rect 705 384 739 418
rect 705 316 739 350
rect 819 296 853 330
rect 819 228 853 262
rect 1062 367 1096 401
rect 1062 299 1096 333
rect 1966 433 2000 467
rect 2124 433 2158 467
rect 1313 306 1347 340
rect 1448 291 1482 325
rect 1556 289 1590 323
rect 1556 221 1590 255
rect 2124 365 2158 399
rect 2232 369 2266 403
rect 2351 359 2385 393
rect 1714 213 1748 247
rect 1822 241 1856 275
rect 1938 241 1972 275
rect 2510 337 2544 371
rect 2510 269 2544 303
rect 2629 253 2663 287
rect 2743 267 2777 301
rect 3037 277 3071 311
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 23 597 89 613
rect 23 563 39 597
rect 73 563 89 597
rect 23 527 89 563
rect 23 493 39 527
rect 73 493 89 527
rect 23 447 89 493
rect 125 565 191 649
rect 125 531 141 565
rect 175 531 191 565
rect 125 483 191 531
rect 227 597 465 613
rect 227 579 415 597
rect 227 447 261 579
rect 399 563 415 579
rect 449 563 465 597
rect 23 413 261 447
rect 297 527 363 543
rect 297 493 313 527
rect 347 493 363 527
rect 297 441 363 493
rect 399 527 465 563
rect 399 493 415 527
rect 449 493 465 527
rect 399 477 465 493
rect 511 597 561 649
rect 511 563 527 597
rect 511 527 561 563
rect 511 493 527 527
rect 511 477 561 493
rect 597 597 663 613
rect 597 563 613 597
rect 647 563 663 597
rect 597 527 663 563
rect 597 493 613 527
rect 647 493 663 527
rect 597 477 663 493
rect 709 590 775 649
rect 709 556 725 590
rect 759 556 775 590
rect 709 520 775 556
rect 709 486 725 520
rect 759 486 775 520
rect 297 407 429 441
rect 25 361 110 377
rect 25 327 60 361
rect 94 327 110 361
rect 25 293 110 327
rect 152 360 257 376
rect 152 326 168 360
rect 202 326 257 360
rect 152 310 257 326
rect 293 355 359 371
rect 293 321 308 355
rect 342 321 359 355
rect 293 305 359 321
rect 25 259 60 293
rect 94 259 110 293
rect 395 269 429 407
rect 597 371 631 477
rect 709 470 775 486
rect 811 590 869 606
rect 845 556 869 590
rect 811 520 869 556
rect 845 486 869 520
rect 465 355 631 371
rect 465 321 481 355
rect 515 337 631 355
rect 689 418 755 434
rect 689 384 705 418
rect 739 384 755 418
rect 689 350 755 384
rect 515 321 547 337
rect 465 305 547 321
rect 25 243 110 259
rect 199 235 477 269
rect 35 178 101 207
rect 35 144 51 178
rect 85 144 101 178
rect 35 17 101 144
rect 199 178 265 235
rect 199 144 215 178
rect 249 144 265 178
rect 199 115 265 144
rect 357 174 407 199
rect 357 140 373 174
rect 357 17 407 140
rect 443 87 477 235
rect 513 182 547 305
rect 689 316 705 350
rect 739 316 755 350
rect 811 346 869 486
rect 689 300 755 316
rect 793 330 869 346
rect 793 296 819 330
rect 853 296 869 330
rect 513 123 547 148
rect 583 230 757 264
rect 583 87 617 230
rect 443 53 617 87
rect 653 165 687 194
rect 653 17 687 131
rect 723 87 757 230
rect 793 262 869 296
rect 793 228 819 262
rect 853 228 869 262
rect 793 175 869 228
rect 827 141 869 175
rect 793 123 869 141
rect 905 573 973 589
rect 905 539 923 573
rect 957 539 973 573
rect 905 503 973 539
rect 905 469 923 503
rect 957 469 973 503
rect 905 417 973 469
rect 1009 573 1075 649
rect 1009 539 1025 573
rect 1059 539 1075 573
rect 1391 586 1457 649
rect 1391 552 1407 586
rect 1441 552 1457 586
rect 1009 503 1075 539
rect 1009 469 1025 503
rect 1059 469 1075 503
rect 1009 453 1075 469
rect 1125 516 1191 545
rect 1125 482 1141 516
rect 1175 482 1191 516
rect 1125 453 1191 482
rect 905 401 1112 417
rect 905 383 1062 401
rect 905 173 939 383
rect 1009 367 1062 383
rect 1096 367 1112 401
rect 1009 333 1112 367
rect 1009 299 1062 333
rect 1096 299 1112 333
rect 1009 283 1112 299
rect 1009 282 1043 283
rect 985 276 1043 282
rect 985 242 991 276
rect 1025 242 1043 276
rect 985 236 1043 242
rect 1157 200 1191 453
rect 905 123 939 139
rect 975 166 1191 200
rect 975 87 1009 166
rect 723 53 1009 87
rect 1045 114 1095 130
rect 1079 80 1095 114
rect 1045 17 1095 80
rect 1141 111 1191 166
rect 1141 77 1157 111
rect 1141 53 1191 77
rect 1227 516 1261 545
rect 1391 536 1457 552
rect 1493 529 1559 545
rect 1493 500 1509 529
rect 1227 239 1261 482
rect 1297 495 1509 500
rect 1543 495 1559 529
rect 1297 466 1559 495
rect 1297 354 1331 466
rect 1493 442 1559 466
rect 1675 520 1741 649
rect 1675 486 1691 520
rect 1725 486 1741 520
rect 1856 578 1922 603
rect 1856 544 1872 578
rect 1906 553 1922 578
rect 2202 596 2268 649
rect 2202 562 2218 596
rect 2252 562 2268 596
rect 1906 544 2079 553
rect 1856 519 2079 544
rect 2202 536 2268 562
rect 2304 597 2370 613
rect 2304 563 2320 597
rect 2354 563 2370 597
rect 1675 462 1741 486
rect 1922 467 2009 483
rect 1369 424 1433 430
rect 1369 390 1375 424
rect 1409 390 1433 424
rect 1493 408 1509 442
rect 1543 426 1559 442
rect 1922 433 1966 467
rect 2000 433 2009 467
rect 1543 408 1872 426
rect 1493 392 1872 408
rect 1399 356 1433 390
rect 1297 340 1363 354
rect 1297 306 1313 340
rect 1347 306 1363 340
rect 1297 290 1363 306
rect 1399 325 1505 356
rect 1399 291 1448 325
rect 1482 291 1505 325
rect 1399 275 1505 291
rect 1541 323 1599 339
rect 1541 289 1556 323
rect 1590 289 1599 323
rect 1541 255 1599 289
rect 1541 239 1556 255
rect 1227 221 1556 239
rect 1590 221 1599 255
rect 1227 205 1599 221
rect 1227 111 1293 205
rect 1227 77 1243 111
rect 1277 77 1293 111
rect 1227 53 1293 77
rect 1401 123 1451 169
rect 1401 89 1417 123
rect 1401 17 1451 89
rect 1487 128 1553 169
rect 1635 163 1669 392
rect 1806 275 1872 392
rect 1589 129 1605 163
rect 1639 129 1669 163
rect 1705 247 1764 263
rect 1705 213 1714 247
rect 1748 213 1764 247
rect 1806 241 1822 275
rect 1856 241 1872 275
rect 1806 225 1872 241
rect 1922 417 2009 433
rect 1922 276 1991 417
rect 2045 304 2079 519
rect 2304 516 2370 563
rect 2474 596 2540 649
rect 2474 562 2490 596
rect 2524 562 2540 596
rect 2474 536 2540 562
rect 2690 591 2756 649
rect 2690 557 2706 591
rect 2740 557 2756 591
rect 2690 536 2756 557
rect 2792 597 2863 613
rect 2826 563 2863 597
rect 2304 500 2320 516
rect 2115 482 2320 500
rect 2354 500 2370 516
rect 2792 500 2863 563
rect 2354 482 2756 500
rect 2115 467 2756 482
rect 2115 433 2124 467
rect 2158 466 2756 467
rect 2158 433 2174 466
rect 2115 399 2174 433
rect 2115 365 2124 399
rect 2158 365 2174 399
rect 2115 349 2174 365
rect 2216 424 2282 430
rect 2216 403 2239 424
rect 2216 369 2232 403
rect 2273 390 2282 424
rect 2266 369 2282 390
rect 2216 353 2282 369
rect 2318 393 2394 409
rect 2318 359 2351 393
rect 2385 359 2394 393
rect 2318 343 2394 359
rect 2318 304 2352 343
rect 2430 307 2464 466
rect 2588 416 2654 430
rect 2588 387 2604 416
rect 1922 275 1951 276
rect 1922 241 1938 275
rect 1985 242 1991 276
rect 1972 241 1991 242
rect 1922 225 1991 241
rect 2027 270 2352 304
rect 2388 291 2464 307
rect 1705 189 1764 213
rect 2027 189 2061 270
rect 2388 257 2404 291
rect 2438 257 2464 291
rect 2388 241 2464 257
rect 2500 382 2604 387
rect 2638 382 2654 416
rect 2500 371 2654 382
rect 2500 337 2510 371
rect 2544 353 2654 371
rect 2544 337 2560 353
rect 2500 303 2560 337
rect 2722 317 2756 466
rect 2826 466 2863 500
rect 2990 607 3040 649
rect 2990 573 3006 607
rect 2990 510 3040 573
rect 2792 403 2863 466
rect 2826 369 2863 403
rect 2792 353 2863 369
rect 2500 269 2510 303
rect 2544 269 2560 303
rect 1705 155 1923 189
rect 1487 94 1503 128
rect 1537 94 1553 128
rect 1487 93 1553 94
rect 1787 111 1853 119
rect 1487 59 1691 93
rect 1725 59 1741 93
rect 1487 53 1741 59
rect 1787 77 1803 111
rect 1837 77 1853 111
rect 1787 17 1853 77
rect 1889 87 1923 155
rect 1959 173 2061 189
rect 1959 139 1975 173
rect 2009 139 2061 173
rect 1959 123 2061 139
rect 2097 200 2352 234
rect 2500 200 2560 269
rect 2613 287 2679 303
rect 2613 253 2629 287
rect 2663 253 2679 287
rect 2613 236 2679 253
rect 2722 301 2793 317
rect 2722 267 2743 301
rect 2777 267 2793 301
rect 2722 251 2793 267
rect 2829 215 2863 353
rect 2097 87 2131 200
rect 2318 180 2654 200
rect 2318 166 2604 180
rect 1889 53 2131 87
rect 2172 125 2238 164
rect 2638 146 2654 180
rect 2172 91 2188 125
rect 2222 91 2238 125
rect 2172 17 2238 91
rect 2274 108 2340 130
rect 2274 74 2290 108
rect 2324 87 2340 108
rect 2480 108 2530 130
rect 2604 127 2654 146
rect 2690 184 2740 200
rect 2690 150 2706 184
rect 2480 87 2496 108
rect 2324 74 2496 87
rect 2274 53 2530 74
rect 2690 93 2740 150
rect 2690 59 2706 93
rect 2690 17 2740 59
rect 2776 199 2863 215
rect 2776 165 2792 199
rect 2826 165 2863 199
rect 2776 103 2863 165
rect 2904 483 2954 499
rect 2938 449 2954 483
rect 2904 413 2954 449
rect 2938 379 2954 413
rect 2904 327 2954 379
rect 2990 476 3006 510
rect 2990 413 3040 476
rect 2990 379 3006 413
rect 2990 363 3040 379
rect 3076 597 3150 613
rect 3076 563 3092 597
rect 3126 563 3150 597
rect 3076 505 3150 563
rect 3076 471 3092 505
rect 3126 471 3150 505
rect 3076 413 3150 471
rect 3076 379 3092 413
rect 3126 379 3150 413
rect 3076 363 3150 379
rect 2904 311 3080 327
rect 2904 277 3037 311
rect 3071 277 3080 311
rect 2904 261 3080 277
rect 2904 196 2954 261
rect 3116 225 3150 363
rect 2938 162 2954 196
rect 2904 133 2954 162
rect 2990 209 3040 225
rect 2990 175 3006 209
rect 2776 69 2792 103
rect 2826 69 2863 103
rect 2776 53 2863 69
rect 2990 99 3040 175
rect 2990 65 3006 99
rect 2990 17 3040 65
rect 3076 209 3150 225
rect 3076 175 3092 209
rect 3126 175 3150 209
rect 3076 103 3150 175
rect 3076 69 3092 103
rect 3126 69 3150 103
rect 3076 53 3150 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 991 242 1025 276
rect 1375 390 1409 424
rect 2239 403 2273 424
rect 2239 390 2266 403
rect 2266 390 2273 403
rect 1951 275 1985 276
rect 1951 242 1972 275
rect 1972 242 1985 275
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
<< metal1 >>
rect 0 683 3168 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3168 683
rect 0 617 3168 649
rect 1363 424 1421 430
rect 1363 390 1375 424
rect 1409 421 1421 424
rect 2227 424 2285 430
rect 2227 421 2239 424
rect 1409 393 2239 421
rect 1409 390 1421 393
rect 1363 384 1421 390
rect 2227 390 2239 393
rect 2273 390 2285 424
rect 2227 384 2285 390
rect 979 276 1037 282
rect 979 242 991 276
rect 1025 273 1037 276
rect 1939 276 1997 282
rect 1939 273 1951 276
rect 1025 245 1951 273
rect 1025 242 1037 245
rect 979 236 1037 242
rect 1939 242 1951 245
rect 1985 242 1997 276
rect 1939 236 1997 242
rect 0 17 3168 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3168 17
rect 0 -49 3168 -17
<< labels >>
flabel pwell s 0 0 3168 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 3168 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfbbp_1
flabel metal1 s 0 617 3168 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 3168 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 3103 94 3137 128 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 3103 168 3137 202 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2815 390 2849 424 0 FreeSans 340 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 2815 464 2849 498 0 FreeSans 340 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 2815 538 2849 572 0 FreeSans 340 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 2623 242 2657 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 SET_B
port 6 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3168 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 7004052
string GDS_START 6981462
<< end >>
