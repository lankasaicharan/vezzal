magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 4426 1852
<< nwell >>
rect -38 261 3166 582
<< pwell >>
rect 1 21 3111 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 183 47 213 177
rect 267 47 297 177
rect 371 47 401 177
rect 455 47 485 177
rect 559 47 589 177
rect 643 47 673 177
rect 747 47 777 177
rect 831 47 861 177
rect 935 47 965 177
rect 1019 47 1049 177
rect 1123 47 1153 177
rect 1207 47 1237 177
rect 1311 47 1341 177
rect 1395 47 1425 177
rect 1499 47 1529 177
rect 1583 47 1613 177
rect 1677 47 1707 177
rect 1771 47 1801 177
rect 1875 47 1905 177
rect 1959 47 1989 177
rect 2063 47 2093 177
rect 2147 47 2177 177
rect 2241 47 2271 177
rect 2335 47 2365 177
rect 2439 47 2469 177
rect 2523 47 2553 177
rect 2627 47 2657 177
rect 2711 47 2741 177
rect 2815 47 2845 177
rect 2899 47 2929 177
rect 3003 47 3033 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
rect 1115 297 1151 497
rect 1209 297 1245 497
rect 1303 297 1339 497
rect 1397 297 1433 497
rect 1491 297 1527 497
rect 1585 297 1621 497
rect 1679 297 1715 497
rect 1773 297 1809 497
rect 1867 297 1903 497
rect 1961 297 1997 497
rect 2055 297 2091 497
rect 2149 297 2185 497
rect 2243 297 2279 497
rect 2337 297 2373 497
rect 2431 297 2467 497
rect 2525 297 2561 497
rect 2619 297 2655 497
rect 2713 297 2749 497
rect 2807 297 2843 497
rect 2901 297 2937 497
rect 2995 297 3031 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 93 183 177
rect 109 59 129 93
rect 163 59 183 93
rect 109 47 183 59
rect 213 161 267 177
rect 213 127 223 161
rect 257 127 267 161
rect 213 93 267 127
rect 213 59 223 93
rect 257 59 267 93
rect 213 47 267 59
rect 297 93 371 177
rect 297 59 317 93
rect 351 59 371 93
rect 297 47 371 59
rect 401 161 455 177
rect 401 127 411 161
rect 445 127 455 161
rect 401 93 455 127
rect 401 59 411 93
rect 445 59 455 93
rect 401 47 455 59
rect 485 93 559 177
rect 485 59 505 93
rect 539 59 559 93
rect 485 47 559 59
rect 589 161 643 177
rect 589 127 599 161
rect 633 127 643 161
rect 589 93 643 127
rect 589 59 599 93
rect 633 59 643 93
rect 589 47 643 59
rect 673 93 747 177
rect 673 59 693 93
rect 727 59 747 93
rect 673 47 747 59
rect 777 161 831 177
rect 777 127 787 161
rect 821 127 831 161
rect 777 93 831 127
rect 777 59 787 93
rect 821 59 831 93
rect 777 47 831 59
rect 861 93 935 177
rect 861 59 881 93
rect 915 59 935 93
rect 861 47 935 59
rect 965 161 1019 177
rect 965 127 975 161
rect 1009 127 1019 161
rect 965 93 1019 127
rect 965 59 975 93
rect 1009 59 1019 93
rect 965 47 1019 59
rect 1049 93 1123 177
rect 1049 59 1069 93
rect 1103 59 1123 93
rect 1049 47 1123 59
rect 1153 161 1207 177
rect 1153 127 1163 161
rect 1197 127 1207 161
rect 1153 93 1207 127
rect 1153 59 1163 93
rect 1197 59 1207 93
rect 1153 47 1207 59
rect 1237 93 1311 177
rect 1237 59 1257 93
rect 1291 59 1311 93
rect 1237 47 1311 59
rect 1341 161 1395 177
rect 1341 127 1351 161
rect 1385 127 1395 161
rect 1341 93 1395 127
rect 1341 59 1351 93
rect 1385 59 1395 93
rect 1341 47 1395 59
rect 1425 93 1499 177
rect 1425 59 1445 93
rect 1479 59 1499 93
rect 1425 47 1499 59
rect 1529 161 1583 177
rect 1529 127 1539 161
rect 1573 127 1583 161
rect 1529 93 1583 127
rect 1529 59 1539 93
rect 1573 59 1583 93
rect 1529 47 1583 59
rect 1613 161 1677 177
rect 1613 127 1633 161
rect 1667 127 1677 161
rect 1613 47 1677 127
rect 1707 93 1771 177
rect 1707 59 1727 93
rect 1761 59 1771 93
rect 1707 47 1771 59
rect 1801 161 1875 177
rect 1801 127 1821 161
rect 1855 127 1875 161
rect 1801 47 1875 127
rect 1905 93 1959 177
rect 1905 59 1915 93
rect 1949 59 1959 93
rect 1905 47 1959 59
rect 1989 161 2063 177
rect 1989 127 2009 161
rect 2043 127 2063 161
rect 1989 47 2063 127
rect 2093 93 2147 177
rect 2093 59 2103 93
rect 2137 59 2147 93
rect 2093 47 2147 59
rect 2177 161 2241 177
rect 2177 127 2197 161
rect 2231 127 2241 161
rect 2177 47 2241 127
rect 2271 93 2335 177
rect 2271 59 2291 93
rect 2325 59 2335 93
rect 2271 47 2335 59
rect 2365 161 2439 177
rect 2365 127 2385 161
rect 2419 127 2439 161
rect 2365 47 2439 127
rect 2469 93 2523 177
rect 2469 59 2479 93
rect 2513 59 2523 93
rect 2469 47 2523 59
rect 2553 161 2627 177
rect 2553 127 2573 161
rect 2607 127 2627 161
rect 2553 47 2627 127
rect 2657 93 2711 177
rect 2657 59 2667 93
rect 2701 59 2711 93
rect 2657 47 2711 59
rect 2741 161 2815 177
rect 2741 127 2761 161
rect 2795 127 2815 161
rect 2741 47 2815 127
rect 2845 93 2899 177
rect 2845 59 2855 93
rect 2889 59 2899 93
rect 2845 47 2899 59
rect 2929 161 3003 177
rect 2929 127 2949 161
rect 2983 127 3003 161
rect 2929 47 3003 127
rect 3033 161 3085 177
rect 3033 127 3043 161
rect 3077 127 3085 161
rect 3033 93 3085 127
rect 3033 59 3043 93
rect 3077 59 3085 93
rect 3033 47 3085 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 417 81 451
rect 27 383 35 417
rect 69 383 81 417
rect 27 349 81 383
rect 27 315 35 349
rect 69 315 81 349
rect 27 297 81 315
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 349 175 383
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 417 269 451
rect 211 383 223 417
rect 257 383 269 417
rect 211 297 269 383
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 349 363 383
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 417 457 451
rect 399 383 411 417
rect 445 383 457 417
rect 399 297 457 383
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 349 551 383
rect 493 315 505 349
rect 539 315 551 349
rect 493 297 551 315
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 417 645 451
rect 587 383 599 417
rect 633 383 645 417
rect 587 297 645 383
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 349 739 383
rect 681 315 693 349
rect 727 315 739 349
rect 681 297 739 315
rect 775 485 833 497
rect 775 451 787 485
rect 821 451 833 485
rect 775 417 833 451
rect 775 383 787 417
rect 821 383 833 417
rect 775 297 833 383
rect 869 485 927 497
rect 869 451 881 485
rect 915 451 927 485
rect 869 417 927 451
rect 869 383 881 417
rect 915 383 927 417
rect 869 349 927 383
rect 869 315 881 349
rect 915 315 927 349
rect 869 297 927 315
rect 963 485 1021 497
rect 963 451 975 485
rect 1009 451 1021 485
rect 963 417 1021 451
rect 963 383 975 417
rect 1009 383 1021 417
rect 963 297 1021 383
rect 1057 485 1115 497
rect 1057 451 1069 485
rect 1103 451 1115 485
rect 1057 417 1115 451
rect 1057 383 1069 417
rect 1103 383 1115 417
rect 1057 349 1115 383
rect 1057 315 1069 349
rect 1103 315 1115 349
rect 1057 297 1115 315
rect 1151 485 1209 497
rect 1151 451 1163 485
rect 1197 451 1209 485
rect 1151 417 1209 451
rect 1151 383 1163 417
rect 1197 383 1209 417
rect 1151 297 1209 383
rect 1245 485 1303 497
rect 1245 451 1257 485
rect 1291 451 1303 485
rect 1245 417 1303 451
rect 1245 383 1257 417
rect 1291 383 1303 417
rect 1245 349 1303 383
rect 1245 315 1257 349
rect 1291 315 1303 349
rect 1245 297 1303 315
rect 1339 485 1397 497
rect 1339 451 1351 485
rect 1385 451 1397 485
rect 1339 417 1397 451
rect 1339 383 1351 417
rect 1385 383 1397 417
rect 1339 297 1397 383
rect 1433 485 1491 497
rect 1433 451 1445 485
rect 1479 451 1491 485
rect 1433 417 1491 451
rect 1433 383 1445 417
rect 1479 383 1491 417
rect 1433 349 1491 383
rect 1433 315 1445 349
rect 1479 315 1491 349
rect 1433 297 1491 315
rect 1527 485 1585 497
rect 1527 451 1539 485
rect 1573 451 1585 485
rect 1527 417 1585 451
rect 1527 383 1539 417
rect 1573 383 1585 417
rect 1527 297 1585 383
rect 1621 485 1679 497
rect 1621 451 1633 485
rect 1667 451 1679 485
rect 1621 417 1679 451
rect 1621 383 1633 417
rect 1667 383 1679 417
rect 1621 349 1679 383
rect 1621 315 1633 349
rect 1667 315 1679 349
rect 1621 297 1679 315
rect 1715 485 1773 497
rect 1715 451 1727 485
rect 1761 451 1773 485
rect 1715 417 1773 451
rect 1715 383 1727 417
rect 1761 383 1773 417
rect 1715 297 1773 383
rect 1809 485 1867 497
rect 1809 451 1821 485
rect 1855 451 1867 485
rect 1809 417 1867 451
rect 1809 383 1821 417
rect 1855 383 1867 417
rect 1809 349 1867 383
rect 1809 315 1821 349
rect 1855 315 1867 349
rect 1809 297 1867 315
rect 1903 485 1961 497
rect 1903 451 1915 485
rect 1949 451 1961 485
rect 1903 417 1961 451
rect 1903 383 1915 417
rect 1949 383 1961 417
rect 1903 297 1961 383
rect 1997 485 2055 497
rect 1997 451 2009 485
rect 2043 451 2055 485
rect 1997 417 2055 451
rect 1997 383 2009 417
rect 2043 383 2055 417
rect 1997 349 2055 383
rect 1997 315 2009 349
rect 2043 315 2055 349
rect 1997 297 2055 315
rect 2091 485 2149 497
rect 2091 451 2103 485
rect 2137 451 2149 485
rect 2091 417 2149 451
rect 2091 383 2103 417
rect 2137 383 2149 417
rect 2091 297 2149 383
rect 2185 485 2243 497
rect 2185 451 2197 485
rect 2231 451 2243 485
rect 2185 417 2243 451
rect 2185 383 2197 417
rect 2231 383 2243 417
rect 2185 349 2243 383
rect 2185 315 2197 349
rect 2231 315 2243 349
rect 2185 297 2243 315
rect 2279 485 2337 497
rect 2279 451 2291 485
rect 2325 451 2337 485
rect 2279 417 2337 451
rect 2279 383 2291 417
rect 2325 383 2337 417
rect 2279 297 2337 383
rect 2373 485 2431 497
rect 2373 451 2385 485
rect 2419 451 2431 485
rect 2373 417 2431 451
rect 2373 383 2385 417
rect 2419 383 2431 417
rect 2373 349 2431 383
rect 2373 315 2385 349
rect 2419 315 2431 349
rect 2373 297 2431 315
rect 2467 485 2525 497
rect 2467 451 2479 485
rect 2513 451 2525 485
rect 2467 417 2525 451
rect 2467 383 2479 417
rect 2513 383 2525 417
rect 2467 297 2525 383
rect 2561 485 2619 497
rect 2561 451 2573 485
rect 2607 451 2619 485
rect 2561 417 2619 451
rect 2561 383 2573 417
rect 2607 383 2619 417
rect 2561 349 2619 383
rect 2561 315 2573 349
rect 2607 315 2619 349
rect 2561 297 2619 315
rect 2655 485 2713 497
rect 2655 451 2667 485
rect 2701 451 2713 485
rect 2655 417 2713 451
rect 2655 383 2667 417
rect 2701 383 2713 417
rect 2655 297 2713 383
rect 2749 485 2807 497
rect 2749 451 2761 485
rect 2795 451 2807 485
rect 2749 417 2807 451
rect 2749 383 2761 417
rect 2795 383 2807 417
rect 2749 349 2807 383
rect 2749 315 2761 349
rect 2795 315 2807 349
rect 2749 297 2807 315
rect 2843 485 2901 497
rect 2843 451 2855 485
rect 2889 451 2901 485
rect 2843 417 2901 451
rect 2843 383 2855 417
rect 2889 383 2901 417
rect 2843 297 2901 383
rect 2937 485 2995 497
rect 2937 451 2949 485
rect 2983 451 2995 485
rect 2937 417 2995 451
rect 2937 383 2949 417
rect 2983 383 2995 417
rect 2937 349 2995 383
rect 2937 315 2949 349
rect 2983 315 2995 349
rect 2937 297 2995 315
rect 3031 485 3085 497
rect 3031 451 3043 485
rect 3077 451 3085 485
rect 3031 417 3085 451
rect 3031 383 3043 417
rect 3077 383 3085 417
rect 3031 349 3085 383
rect 3031 315 3043 349
rect 3077 315 3085 349
rect 3031 297 3085 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 129 59 163 93
rect 223 127 257 161
rect 223 59 257 93
rect 317 59 351 93
rect 411 127 445 161
rect 411 59 445 93
rect 505 59 539 93
rect 599 127 633 161
rect 599 59 633 93
rect 693 59 727 93
rect 787 127 821 161
rect 787 59 821 93
rect 881 59 915 93
rect 975 127 1009 161
rect 975 59 1009 93
rect 1069 59 1103 93
rect 1163 127 1197 161
rect 1163 59 1197 93
rect 1257 59 1291 93
rect 1351 127 1385 161
rect 1351 59 1385 93
rect 1445 59 1479 93
rect 1539 127 1573 161
rect 1539 59 1573 93
rect 1633 127 1667 161
rect 1727 59 1761 93
rect 1821 127 1855 161
rect 1915 59 1949 93
rect 2009 127 2043 161
rect 2103 59 2137 93
rect 2197 127 2231 161
rect 2291 59 2325 93
rect 2385 127 2419 161
rect 2479 59 2513 93
rect 2573 127 2607 161
rect 2667 59 2701 93
rect 2761 127 2795 161
rect 2855 59 2889 93
rect 2949 127 2983 161
rect 3043 127 3077 161
rect 3043 59 3077 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 129 451 163 485
rect 129 383 163 417
rect 129 315 163 349
rect 223 451 257 485
rect 223 383 257 417
rect 317 451 351 485
rect 317 383 351 417
rect 317 315 351 349
rect 411 451 445 485
rect 411 383 445 417
rect 505 451 539 485
rect 505 383 539 417
rect 505 315 539 349
rect 599 451 633 485
rect 599 383 633 417
rect 693 451 727 485
rect 693 383 727 417
rect 693 315 727 349
rect 787 451 821 485
rect 787 383 821 417
rect 881 451 915 485
rect 881 383 915 417
rect 881 315 915 349
rect 975 451 1009 485
rect 975 383 1009 417
rect 1069 451 1103 485
rect 1069 383 1103 417
rect 1069 315 1103 349
rect 1163 451 1197 485
rect 1163 383 1197 417
rect 1257 451 1291 485
rect 1257 383 1291 417
rect 1257 315 1291 349
rect 1351 451 1385 485
rect 1351 383 1385 417
rect 1445 451 1479 485
rect 1445 383 1479 417
rect 1445 315 1479 349
rect 1539 451 1573 485
rect 1539 383 1573 417
rect 1633 451 1667 485
rect 1633 383 1667 417
rect 1633 315 1667 349
rect 1727 451 1761 485
rect 1727 383 1761 417
rect 1821 451 1855 485
rect 1821 383 1855 417
rect 1821 315 1855 349
rect 1915 451 1949 485
rect 1915 383 1949 417
rect 2009 451 2043 485
rect 2009 383 2043 417
rect 2009 315 2043 349
rect 2103 451 2137 485
rect 2103 383 2137 417
rect 2197 451 2231 485
rect 2197 383 2231 417
rect 2197 315 2231 349
rect 2291 451 2325 485
rect 2291 383 2325 417
rect 2385 451 2419 485
rect 2385 383 2419 417
rect 2385 315 2419 349
rect 2479 451 2513 485
rect 2479 383 2513 417
rect 2573 451 2607 485
rect 2573 383 2607 417
rect 2573 315 2607 349
rect 2667 451 2701 485
rect 2667 383 2701 417
rect 2761 451 2795 485
rect 2761 383 2795 417
rect 2761 315 2795 349
rect 2855 451 2889 485
rect 2855 383 2889 417
rect 2949 451 2983 485
rect 2949 383 2983 417
rect 2949 315 2983 349
rect 3043 451 3077 485
rect 3043 383 3077 417
rect 3043 315 3077 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 1115 497 1151 523
rect 1209 497 1245 523
rect 1303 497 1339 523
rect 1397 497 1433 523
rect 1491 497 1527 523
rect 1585 497 1621 523
rect 1679 497 1715 523
rect 1773 497 1809 523
rect 1867 497 1903 523
rect 1961 497 1997 523
rect 2055 497 2091 523
rect 2149 497 2185 523
rect 2243 497 2279 523
rect 2337 497 2373 523
rect 2431 497 2467 523
rect 2525 497 2561 523
rect 2619 497 2655 523
rect 2713 497 2749 523
rect 2807 497 2843 523
rect 2901 497 2937 523
rect 2995 497 3031 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 1115 282 1151 297
rect 1209 282 1245 297
rect 1303 282 1339 297
rect 1397 282 1433 297
rect 1491 282 1527 297
rect 1585 282 1621 297
rect 1679 282 1715 297
rect 1773 282 1809 297
rect 1867 282 1903 297
rect 1961 282 1997 297
rect 2055 282 2091 297
rect 2149 282 2185 297
rect 2243 282 2279 297
rect 2337 282 2373 297
rect 2431 282 2467 297
rect 2525 282 2561 297
rect 2619 282 2655 297
rect 2713 282 2749 297
rect 2807 282 2843 297
rect 2901 282 2937 297
rect 2995 282 3031 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 831 265 871 282
rect 925 265 965 282
rect 1019 265 1059 282
rect 1113 265 1153 282
rect 1207 265 1247 282
rect 1301 265 1341 282
rect 1395 265 1435 282
rect 1489 265 1529 282
rect 79 249 1529 265
rect 79 215 95 249
rect 129 215 163 249
rect 197 215 231 249
rect 265 215 299 249
rect 333 215 367 249
rect 401 215 435 249
rect 469 215 503 249
rect 537 215 571 249
rect 605 215 639 249
rect 673 215 707 249
rect 741 215 775 249
rect 809 215 843 249
rect 877 215 911 249
rect 945 215 979 249
rect 1013 215 1047 249
rect 1081 215 1115 249
rect 1149 215 1183 249
rect 1217 215 1251 249
rect 1285 215 1319 249
rect 1353 215 1387 249
rect 1421 215 1455 249
rect 1489 215 1529 249
rect 79 199 1529 215
rect 79 177 109 199
rect 183 177 213 199
rect 267 177 297 199
rect 371 177 401 199
rect 455 177 485 199
rect 559 177 589 199
rect 643 177 673 199
rect 747 177 777 199
rect 831 177 861 199
rect 935 177 965 199
rect 1019 177 1049 199
rect 1123 177 1153 199
rect 1207 177 1237 199
rect 1311 177 1341 199
rect 1395 177 1425 199
rect 1499 177 1529 199
rect 1583 265 1623 282
rect 1677 265 1717 282
rect 1771 265 1811 282
rect 1865 265 1905 282
rect 1959 265 1999 282
rect 2053 265 2093 282
rect 2147 265 2187 282
rect 2241 265 2281 282
rect 2335 265 2375 282
rect 2429 265 2469 282
rect 2523 265 2563 282
rect 2617 265 2657 282
rect 2711 265 2751 282
rect 2805 265 2845 282
rect 2899 265 2939 282
rect 2993 265 3033 282
rect 1583 249 3033 265
rect 1583 215 1717 249
rect 1751 215 1785 249
rect 1819 215 1853 249
rect 1887 215 1921 249
rect 1955 215 1989 249
rect 2023 215 2057 249
rect 2091 215 2125 249
rect 2159 215 2193 249
rect 2227 215 2261 249
rect 2295 215 2329 249
rect 2363 215 2397 249
rect 2431 215 2465 249
rect 2499 215 2533 249
rect 2567 215 2601 249
rect 2635 215 2669 249
rect 2703 215 2737 249
rect 2771 215 2805 249
rect 2839 215 3033 249
rect 1583 199 3033 215
rect 1583 177 1613 199
rect 1677 177 1707 199
rect 1771 177 1801 199
rect 1875 177 1905 199
rect 1959 177 1989 199
rect 2063 177 2093 199
rect 2147 177 2177 199
rect 2241 177 2271 199
rect 2335 177 2365 199
rect 2439 177 2469 199
rect 2523 177 2553 199
rect 2627 177 2657 199
rect 2711 177 2741 199
rect 2815 177 2845 199
rect 2899 177 2929 199
rect 3003 177 3033 199
rect 79 21 109 47
rect 183 21 213 47
rect 267 21 297 47
rect 371 21 401 47
rect 455 21 485 47
rect 559 21 589 47
rect 643 21 673 47
rect 747 21 777 47
rect 831 21 861 47
rect 935 21 965 47
rect 1019 21 1049 47
rect 1123 21 1153 47
rect 1207 21 1237 47
rect 1311 21 1341 47
rect 1395 21 1425 47
rect 1499 21 1529 47
rect 1583 21 1613 47
rect 1677 21 1707 47
rect 1771 21 1801 47
rect 1875 21 1905 47
rect 1959 21 1989 47
rect 2063 21 2093 47
rect 2147 21 2177 47
rect 2241 21 2271 47
rect 2335 21 2365 47
rect 2439 21 2469 47
rect 2523 21 2553 47
rect 2627 21 2657 47
rect 2711 21 2741 47
rect 2815 21 2845 47
rect 2899 21 2929 47
rect 3003 21 3033 47
<< polycont >>
rect 95 215 129 249
rect 163 215 197 249
rect 231 215 265 249
rect 299 215 333 249
rect 367 215 401 249
rect 435 215 469 249
rect 503 215 537 249
rect 571 215 605 249
rect 639 215 673 249
rect 707 215 741 249
rect 775 215 809 249
rect 843 215 877 249
rect 911 215 945 249
rect 979 215 1013 249
rect 1047 215 1081 249
rect 1115 215 1149 249
rect 1183 215 1217 249
rect 1251 215 1285 249
rect 1319 215 1353 249
rect 1387 215 1421 249
rect 1455 215 1489 249
rect 1717 215 1751 249
rect 1785 215 1819 249
rect 1853 215 1887 249
rect 1921 215 1955 249
rect 1989 215 2023 249
rect 2057 215 2091 249
rect 2125 215 2159 249
rect 2193 215 2227 249
rect 2261 215 2295 249
rect 2329 215 2363 249
rect 2397 215 2431 249
rect 2465 215 2499 249
rect 2533 215 2567 249
rect 2601 215 2635 249
rect 2669 215 2703 249
rect 2737 215 2771 249
rect 2805 215 2839 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3128 561
rect 25 485 79 527
rect 25 451 35 485
rect 69 451 79 485
rect 25 417 79 451
rect 25 383 35 417
rect 69 383 79 417
rect 25 349 79 383
rect 25 315 35 349
rect 69 315 79 349
rect 25 299 79 315
rect 113 485 179 493
rect 113 451 129 485
rect 163 451 179 485
rect 113 417 179 451
rect 113 383 129 417
rect 163 383 179 417
rect 113 349 179 383
rect 213 485 267 527
rect 213 451 223 485
rect 257 451 267 485
rect 213 417 267 451
rect 213 383 223 417
rect 257 383 267 417
rect 213 367 267 383
rect 301 485 367 493
rect 301 451 317 485
rect 351 451 367 485
rect 301 417 367 451
rect 301 383 317 417
rect 351 383 367 417
rect 113 315 129 349
rect 163 333 179 349
rect 301 349 367 383
rect 401 485 455 527
rect 401 451 411 485
rect 445 451 455 485
rect 401 417 455 451
rect 401 383 411 417
rect 445 383 455 417
rect 401 367 455 383
rect 489 485 555 493
rect 489 451 505 485
rect 539 451 555 485
rect 489 417 555 451
rect 489 383 505 417
rect 539 383 555 417
rect 301 333 317 349
rect 163 315 317 333
rect 351 333 367 349
rect 489 349 555 383
rect 589 485 643 527
rect 589 451 599 485
rect 633 451 643 485
rect 589 417 643 451
rect 589 383 599 417
rect 633 383 643 417
rect 589 367 643 383
rect 677 485 743 493
rect 677 451 693 485
rect 727 451 743 485
rect 677 417 743 451
rect 677 383 693 417
rect 727 383 743 417
rect 489 333 505 349
rect 351 315 505 333
rect 539 333 555 349
rect 677 349 743 383
rect 777 485 831 527
rect 777 451 787 485
rect 821 451 831 485
rect 777 417 831 451
rect 777 383 787 417
rect 821 383 831 417
rect 777 367 831 383
rect 865 485 931 493
rect 865 451 881 485
rect 915 451 931 485
rect 865 417 931 451
rect 865 383 881 417
rect 915 383 931 417
rect 677 333 693 349
rect 539 315 693 333
rect 727 333 743 349
rect 865 349 931 383
rect 965 485 1019 527
rect 965 451 975 485
rect 1009 451 1019 485
rect 965 417 1019 451
rect 965 383 975 417
rect 1009 383 1019 417
rect 965 367 1019 383
rect 1053 485 1119 493
rect 1053 451 1069 485
rect 1103 451 1119 485
rect 1053 417 1119 451
rect 1053 383 1069 417
rect 1103 383 1119 417
rect 865 333 881 349
rect 727 315 881 333
rect 915 333 931 349
rect 1053 349 1119 383
rect 1153 485 1207 527
rect 1153 451 1163 485
rect 1197 451 1207 485
rect 1153 417 1207 451
rect 1153 383 1163 417
rect 1197 383 1207 417
rect 1153 367 1207 383
rect 1241 485 1307 493
rect 1241 451 1257 485
rect 1291 451 1307 485
rect 1241 417 1307 451
rect 1241 383 1257 417
rect 1291 383 1307 417
rect 1053 333 1069 349
rect 915 315 1069 333
rect 1103 333 1119 349
rect 1241 349 1307 383
rect 1341 485 1395 527
rect 1341 451 1351 485
rect 1385 451 1395 485
rect 1341 417 1395 451
rect 1341 383 1351 417
rect 1385 383 1395 417
rect 1341 367 1395 383
rect 1429 485 1495 493
rect 1429 451 1445 485
rect 1479 451 1495 485
rect 1429 417 1495 451
rect 1429 383 1445 417
rect 1479 383 1495 417
rect 1241 333 1257 349
rect 1103 315 1257 333
rect 1291 333 1307 349
rect 1429 349 1495 383
rect 1529 485 1583 527
rect 1529 451 1539 485
rect 1573 451 1583 485
rect 1529 417 1583 451
rect 1529 383 1539 417
rect 1573 383 1583 417
rect 1529 367 1583 383
rect 1617 485 1683 493
rect 1617 451 1633 485
rect 1667 451 1683 485
rect 1617 417 1683 451
rect 1617 383 1633 417
rect 1667 383 1683 417
rect 1429 333 1445 349
rect 1291 315 1445 333
rect 1479 333 1495 349
rect 1617 349 1683 383
rect 1717 485 1771 527
rect 1717 451 1727 485
rect 1761 451 1771 485
rect 1717 417 1771 451
rect 1717 383 1727 417
rect 1761 383 1771 417
rect 1717 367 1771 383
rect 1805 485 1871 493
rect 1805 451 1821 485
rect 1855 451 1871 485
rect 1805 417 1871 451
rect 1805 383 1821 417
rect 1855 383 1871 417
rect 1617 333 1633 349
rect 1479 315 1633 333
rect 1667 333 1683 349
rect 1805 349 1871 383
rect 1905 485 1959 527
rect 1905 451 1915 485
rect 1949 451 1959 485
rect 1905 417 1959 451
rect 1905 383 1915 417
rect 1949 383 1959 417
rect 1905 367 1959 383
rect 1993 485 2059 493
rect 1993 451 2009 485
rect 2043 451 2059 485
rect 1993 417 2059 451
rect 1993 383 2009 417
rect 2043 383 2059 417
rect 1805 333 1821 349
rect 1667 315 1821 333
rect 1855 333 1871 349
rect 1993 349 2059 383
rect 2093 485 2147 527
rect 2093 451 2103 485
rect 2137 451 2147 485
rect 2093 417 2147 451
rect 2093 383 2103 417
rect 2137 383 2147 417
rect 2093 367 2147 383
rect 2181 485 2247 493
rect 2181 451 2197 485
rect 2231 451 2247 485
rect 2181 417 2247 451
rect 2181 383 2197 417
rect 2231 383 2247 417
rect 1993 333 2009 349
rect 1855 315 2009 333
rect 2043 333 2059 349
rect 2181 349 2247 383
rect 2281 485 2335 527
rect 2281 451 2291 485
rect 2325 451 2335 485
rect 2281 417 2335 451
rect 2281 383 2291 417
rect 2325 383 2335 417
rect 2281 367 2335 383
rect 2369 485 2435 493
rect 2369 451 2385 485
rect 2419 451 2435 485
rect 2369 417 2435 451
rect 2369 383 2385 417
rect 2419 383 2435 417
rect 2181 333 2197 349
rect 2043 315 2197 333
rect 2231 333 2247 349
rect 2369 349 2435 383
rect 2469 485 2523 527
rect 2469 451 2479 485
rect 2513 451 2523 485
rect 2469 417 2523 451
rect 2469 383 2479 417
rect 2513 383 2523 417
rect 2469 367 2523 383
rect 2557 485 2623 493
rect 2557 451 2573 485
rect 2607 451 2623 485
rect 2557 417 2623 451
rect 2557 383 2573 417
rect 2607 383 2623 417
rect 2369 333 2385 349
rect 2231 315 2385 333
rect 2419 333 2435 349
rect 2557 349 2623 383
rect 2657 485 2711 527
rect 2657 451 2667 485
rect 2701 451 2711 485
rect 2657 417 2711 451
rect 2657 383 2667 417
rect 2701 383 2711 417
rect 2657 367 2711 383
rect 2745 485 2811 493
rect 2745 451 2761 485
rect 2795 451 2811 485
rect 2745 417 2811 451
rect 2745 383 2761 417
rect 2795 383 2811 417
rect 2557 333 2573 349
rect 2419 315 2573 333
rect 2607 333 2623 349
rect 2745 349 2811 383
rect 2845 485 2899 527
rect 2845 451 2855 485
rect 2889 451 2899 485
rect 2845 417 2899 451
rect 2845 383 2855 417
rect 2889 383 2899 417
rect 2845 367 2899 383
rect 2933 485 2999 493
rect 2933 451 2949 485
rect 2983 451 2999 485
rect 2933 417 2999 451
rect 2933 383 2949 417
rect 2983 383 2999 417
rect 2745 333 2761 349
rect 2607 315 2761 333
rect 2795 333 2811 349
rect 2933 349 2999 383
rect 2933 333 2949 349
rect 2795 315 2949 333
rect 2983 315 2999 349
rect 113 299 2999 315
rect 3033 485 3087 527
rect 3033 451 3043 485
rect 3077 451 3087 485
rect 3033 417 3087 451
rect 3033 383 3043 417
rect 3077 383 3087 417
rect 3033 349 3087 383
rect 3033 315 3043 349
rect 3077 315 3087 349
rect 3033 299 3087 315
rect 79 249 1505 265
rect 79 215 95 249
rect 129 215 163 249
rect 197 215 231 249
rect 265 215 299 249
rect 333 215 367 249
rect 401 215 435 249
rect 469 215 503 249
rect 537 215 571 249
rect 605 215 639 249
rect 673 215 707 249
rect 741 215 775 249
rect 809 215 843 249
rect 877 215 911 249
rect 945 215 979 249
rect 1013 215 1047 249
rect 1081 215 1115 249
rect 1149 215 1183 249
rect 1217 215 1251 249
rect 1285 215 1319 249
rect 1353 215 1387 249
rect 1421 215 1455 249
rect 1489 215 1505 249
rect 79 211 1505 215
rect 1585 211 1667 299
rect 2945 265 2999 299
rect 1701 249 2855 265
rect 1701 215 1717 249
rect 1751 215 1785 249
rect 1819 215 1853 249
rect 1887 215 1921 249
rect 1955 215 1989 249
rect 2023 215 2057 249
rect 2091 215 2125 249
rect 2159 215 2193 249
rect 2227 215 2261 249
rect 2295 215 2329 249
rect 2363 215 2397 249
rect 2431 215 2465 249
rect 2499 215 2533 249
rect 2567 215 2601 249
rect 2635 215 2669 249
rect 2703 215 2737 249
rect 2771 215 2805 249
rect 2839 215 2855 249
rect 1701 211 2855 215
rect 2945 211 3023 265
rect 1607 177 1667 211
rect 2945 177 2999 211
rect 19 161 1573 177
rect 19 127 35 161
rect 69 143 223 161
rect 69 127 85 143
rect 19 93 85 127
rect 207 127 223 143
rect 257 143 411 161
rect 257 127 273 143
rect 19 59 35 93
rect 69 59 85 93
rect 19 51 85 59
rect 119 93 173 109
rect 119 59 129 93
rect 163 59 173 93
rect 119 17 173 59
rect 207 93 273 127
rect 395 127 411 143
rect 445 143 599 161
rect 445 127 461 143
rect 207 59 223 93
rect 257 59 273 93
rect 207 51 273 59
rect 307 93 361 109
rect 307 59 317 93
rect 351 59 361 93
rect 307 17 361 59
rect 395 93 461 127
rect 583 127 599 143
rect 633 143 787 161
rect 633 127 649 143
rect 395 59 411 93
rect 445 59 461 93
rect 395 51 461 59
rect 495 93 549 109
rect 495 59 505 93
rect 539 59 549 93
rect 495 17 549 59
rect 583 93 649 127
rect 771 127 787 143
rect 821 143 975 161
rect 821 127 837 143
rect 583 59 599 93
rect 633 59 649 93
rect 583 51 649 59
rect 683 93 737 109
rect 683 59 693 93
rect 727 59 737 93
rect 683 17 737 59
rect 771 93 837 127
rect 959 127 975 143
rect 1009 143 1163 161
rect 1009 127 1025 143
rect 771 59 787 93
rect 821 59 837 93
rect 771 51 837 59
rect 871 93 925 109
rect 871 59 881 93
rect 915 59 925 93
rect 871 17 925 59
rect 959 93 1025 127
rect 1147 127 1163 143
rect 1197 143 1351 161
rect 1197 127 1213 143
rect 959 59 975 93
rect 1009 59 1025 93
rect 959 51 1025 59
rect 1059 93 1113 109
rect 1059 59 1069 93
rect 1103 59 1113 93
rect 1059 17 1113 59
rect 1147 93 1213 127
rect 1335 127 1351 143
rect 1385 143 1539 161
rect 1385 127 1401 143
rect 1147 59 1163 93
rect 1197 59 1213 93
rect 1147 51 1213 59
rect 1247 93 1301 109
rect 1247 59 1257 93
rect 1291 59 1301 93
rect 1247 17 1301 59
rect 1335 93 1401 127
rect 1523 127 1539 143
rect 1607 161 2999 177
rect 1607 127 1633 161
rect 1667 127 1821 161
rect 1855 127 2009 161
rect 2043 127 2197 161
rect 2231 127 2385 161
rect 2419 127 2573 161
rect 2607 127 2761 161
rect 2795 127 2949 161
rect 2983 127 2999 161
rect 3043 161 3093 177
rect 3077 127 3093 161
rect 1335 59 1351 93
rect 1385 59 1401 93
rect 1335 51 1401 59
rect 1435 93 1489 109
rect 1435 59 1445 93
rect 1479 59 1489 93
rect 1435 17 1489 59
rect 1523 93 1573 127
rect 3043 93 3093 127
rect 1523 59 1539 93
rect 1573 59 1727 93
rect 1761 59 1915 93
rect 1949 59 2103 93
rect 2137 59 2291 93
rect 2325 59 2479 93
rect 2513 59 2667 93
rect 2701 59 2855 93
rect 2889 59 3043 93
rect 3077 59 3093 93
rect 1523 51 3093 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3128 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 3065 527 3099 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
rect 3065 -17 3099 17
<< metal1 >>
rect 0 561 3128 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3128 561
rect 0 496 3128 527
rect 0 17 3128 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3128 17
rect 0 -48 3128 -17
<< labels >>
flabel locali s 1593 221 1627 255 0 FreeSans 250 0 0 0 Y
port 7 nsew signal output
flabel locali s 2237 221 2271 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 765 221 799 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand2_16
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 3128 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 3516752
string GDS_START 3495032
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
