magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 43 49 575 243
rect 0 0 576 49
<< scnmos >>
rect 122 49 152 217
rect 208 49 238 217
rect 294 49 324 217
rect 380 49 410 217
rect 466 49 496 217
<< scpmoshvt >>
rect 122 367 152 619
rect 208 367 238 619
rect 294 367 324 619
rect 380 367 410 619
rect 466 367 496 619
<< ndiff >>
rect 69 181 122 217
rect 69 147 77 181
rect 111 147 122 181
rect 69 95 122 147
rect 69 61 77 95
rect 111 61 122 95
rect 69 49 122 61
rect 152 205 208 217
rect 152 171 163 205
rect 197 171 208 205
rect 152 101 208 171
rect 152 67 163 101
rect 197 67 208 101
rect 152 49 208 67
rect 238 181 294 217
rect 238 147 249 181
rect 283 147 294 181
rect 238 95 294 147
rect 238 61 249 95
rect 283 61 294 95
rect 238 49 294 61
rect 324 205 380 217
rect 324 171 335 205
rect 369 171 380 205
rect 324 101 380 171
rect 324 67 335 101
rect 369 67 380 101
rect 324 49 380 67
rect 410 130 466 217
rect 410 96 421 130
rect 455 96 466 130
rect 410 49 466 96
rect 496 190 549 217
rect 496 156 507 190
rect 541 156 549 190
rect 496 101 549 156
rect 496 67 507 101
rect 541 67 549 101
rect 496 49 549 67
<< pdiff >>
rect 65 611 122 619
rect 65 577 77 611
rect 111 577 122 611
rect 65 533 122 577
rect 65 499 77 533
rect 111 499 122 533
rect 65 457 122 499
rect 65 423 77 457
rect 111 423 122 457
rect 65 367 122 423
rect 152 599 208 619
rect 152 565 163 599
rect 197 565 208 599
rect 152 506 208 565
rect 152 472 163 506
rect 197 472 208 506
rect 152 413 208 472
rect 152 379 163 413
rect 197 379 208 413
rect 152 367 208 379
rect 238 611 294 619
rect 238 577 249 611
rect 283 577 294 611
rect 238 533 294 577
rect 238 499 249 533
rect 283 499 294 533
rect 238 457 294 499
rect 238 423 249 457
rect 283 423 294 457
rect 238 367 294 423
rect 324 599 380 619
rect 324 565 335 599
rect 369 565 380 599
rect 324 506 380 565
rect 324 472 335 506
rect 369 472 380 506
rect 324 413 380 472
rect 324 379 335 413
rect 369 379 380 413
rect 324 367 380 379
rect 410 607 466 619
rect 410 573 421 607
rect 455 573 466 607
rect 410 531 466 573
rect 410 497 421 531
rect 455 497 466 531
rect 410 453 466 497
rect 410 419 421 453
rect 455 419 466 453
rect 410 367 466 419
rect 496 599 549 619
rect 496 565 507 599
rect 541 565 549 599
rect 496 506 549 565
rect 496 472 507 506
rect 541 472 549 506
rect 496 413 549 472
rect 496 379 507 413
rect 541 379 549 413
rect 496 367 549 379
<< ndiffc >>
rect 77 147 111 181
rect 77 61 111 95
rect 163 171 197 205
rect 163 67 197 101
rect 249 147 283 181
rect 249 61 283 95
rect 335 171 369 205
rect 335 67 369 101
rect 421 96 455 130
rect 507 156 541 190
rect 507 67 541 101
<< pdiffc >>
rect 77 577 111 611
rect 77 499 111 533
rect 77 423 111 457
rect 163 565 197 599
rect 163 472 197 506
rect 163 379 197 413
rect 249 577 283 611
rect 249 499 283 533
rect 249 423 283 457
rect 335 565 369 599
rect 335 472 369 506
rect 335 379 369 413
rect 421 573 455 607
rect 421 497 455 531
rect 421 419 455 453
rect 507 565 541 599
rect 507 472 541 506
rect 507 379 541 413
<< poly >>
rect 122 619 152 645
rect 208 619 238 645
rect 294 619 324 645
rect 380 619 410 645
rect 466 619 496 645
rect 122 335 152 367
rect 208 335 238 367
rect 294 335 324 367
rect 380 335 410 367
rect 122 319 410 335
rect 122 285 156 319
rect 190 285 224 319
rect 258 285 292 319
rect 326 285 360 319
rect 394 285 410 319
rect 122 269 410 285
rect 122 217 152 269
rect 208 217 238 269
rect 294 217 324 269
rect 380 217 410 269
rect 466 308 496 367
rect 466 292 532 308
rect 466 258 482 292
rect 516 258 532 292
rect 466 242 532 258
rect 466 217 496 242
rect 122 23 152 49
rect 208 23 238 49
rect 294 23 324 49
rect 380 23 410 49
rect 466 23 496 49
<< polycont >>
rect 156 285 190 319
rect 224 285 258 319
rect 292 285 326 319
rect 360 285 394 319
rect 482 258 516 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 61 611 127 649
rect 61 577 77 611
rect 111 577 127 611
rect 61 533 127 577
rect 61 499 77 533
rect 111 499 127 533
rect 61 457 127 499
rect 61 423 77 457
rect 111 423 127 457
rect 161 599 199 615
rect 161 565 163 599
rect 197 565 199 599
rect 161 506 199 565
rect 161 472 163 506
rect 197 472 199 506
rect 161 413 199 472
rect 233 611 299 649
rect 233 577 249 611
rect 283 577 299 611
rect 233 533 299 577
rect 233 499 249 533
rect 283 499 299 533
rect 233 457 299 499
rect 233 423 249 457
rect 283 423 299 457
rect 333 599 371 615
rect 333 565 335 599
rect 369 565 371 599
rect 333 506 371 565
rect 333 472 335 506
rect 369 472 371 506
rect 161 389 163 413
rect 19 379 163 389
rect 197 389 199 413
rect 333 413 371 472
rect 405 607 471 649
rect 405 573 421 607
rect 455 573 471 607
rect 405 531 471 573
rect 405 497 421 531
rect 455 497 471 531
rect 405 453 471 497
rect 405 419 421 453
rect 455 419 471 453
rect 505 599 557 615
rect 505 565 507 599
rect 541 565 557 599
rect 505 506 557 565
rect 505 472 507 506
rect 541 472 557 506
rect 333 389 335 413
rect 197 379 335 389
rect 369 379 371 413
rect 505 413 557 472
rect 505 385 507 413
rect 19 355 371 379
rect 405 379 507 385
rect 541 379 557 413
rect 19 249 102 355
rect 405 351 557 379
rect 405 321 444 351
rect 140 319 444 321
rect 140 285 156 319
rect 190 285 224 319
rect 258 285 292 319
rect 326 285 360 319
rect 394 285 444 319
rect 140 283 444 285
rect 19 215 371 249
rect 161 205 199 215
rect 61 147 77 181
rect 111 147 127 181
rect 61 95 127 147
rect 61 61 77 95
rect 111 61 127 95
rect 61 17 127 61
rect 161 171 163 205
rect 197 171 199 205
rect 333 205 371 215
rect 161 101 199 171
rect 161 67 163 101
rect 197 67 199 101
rect 161 51 199 67
rect 233 147 249 181
rect 283 147 299 181
rect 233 95 299 147
rect 233 61 249 95
rect 283 61 299 95
rect 233 17 299 61
rect 333 171 335 205
rect 369 171 371 205
rect 405 206 444 283
rect 478 292 557 308
rect 478 258 482 292
rect 516 258 557 292
rect 478 240 557 258
rect 405 190 557 206
rect 405 172 507 190
rect 333 101 371 171
rect 505 156 507 172
rect 541 156 557 190
rect 333 67 335 101
rect 369 67 371 101
rect 333 51 371 67
rect 405 130 471 138
rect 405 96 421 130
rect 455 96 471 130
rect 405 17 471 96
rect 505 101 557 156
rect 505 67 507 101
rect 541 67 557 101
rect 505 51 557 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 buf_4
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5101886
string GDS_START 5096136
<< end >>
