magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2586 1852
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 1 21 1265 203
rect 29 -17 63 21
<< scnmos >>
rect 82 47 112 177
rect 186 47 216 177
rect 280 47 310 177
rect 374 47 404 177
rect 572 47 602 177
rect 656 47 686 177
rect 750 47 780 177
rect 865 47 895 177
rect 1053 47 1083 177
rect 1157 47 1187 177
<< scpmoshvt >>
rect 84 297 120 497
rect 178 297 214 497
rect 272 297 308 497
rect 366 297 402 497
rect 564 297 600 497
rect 658 297 694 497
rect 752 297 788 497
rect 857 297 893 497
rect 1055 297 1091 497
rect 1149 297 1185 497
<< ndiff >>
rect 27 95 82 177
rect 27 61 38 95
rect 72 61 82 95
rect 27 47 82 61
rect 112 163 186 177
rect 112 129 132 163
rect 166 129 186 163
rect 112 95 186 129
rect 112 61 132 95
rect 166 61 186 95
rect 112 47 186 61
rect 216 95 280 177
rect 216 61 226 95
rect 260 61 280 95
rect 216 47 280 61
rect 310 163 374 177
rect 310 129 320 163
rect 354 129 374 163
rect 310 95 374 129
rect 310 61 320 95
rect 354 61 374 95
rect 310 47 374 61
rect 404 95 456 177
rect 404 61 414 95
rect 448 61 456 95
rect 404 47 456 61
rect 510 163 572 177
rect 510 129 518 163
rect 552 129 572 163
rect 510 95 572 129
rect 510 61 518 95
rect 552 61 572 95
rect 510 47 572 61
rect 602 95 656 177
rect 602 61 612 95
rect 646 61 656 95
rect 602 47 656 61
rect 686 125 750 177
rect 686 91 706 125
rect 740 91 750 125
rect 686 47 750 91
rect 780 163 865 177
rect 780 129 811 163
rect 845 129 865 163
rect 780 47 865 129
rect 895 95 947 177
rect 895 61 905 95
rect 939 61 947 95
rect 895 47 947 61
rect 1001 95 1053 177
rect 1001 61 1009 95
rect 1043 61 1053 95
rect 1001 47 1053 61
rect 1083 163 1157 177
rect 1083 129 1103 163
rect 1137 129 1157 163
rect 1083 47 1157 129
rect 1187 95 1239 177
rect 1187 61 1197 95
rect 1231 61 1239 95
rect 1187 47 1239 61
<< pdiff >>
rect 27 477 84 497
rect 27 443 38 477
rect 72 443 84 477
rect 27 297 84 443
rect 120 477 178 497
rect 120 443 132 477
rect 166 443 178 477
rect 120 297 178 443
rect 214 477 272 497
rect 214 443 226 477
rect 260 443 272 477
rect 214 297 272 443
rect 308 409 366 497
rect 308 375 320 409
rect 354 375 366 409
rect 308 297 366 375
rect 402 477 456 497
rect 402 443 414 477
rect 448 443 456 477
rect 402 297 456 443
rect 510 477 564 497
rect 510 443 518 477
rect 552 443 564 477
rect 510 409 564 443
rect 510 375 518 409
rect 552 375 564 409
rect 510 297 564 375
rect 600 477 658 497
rect 600 443 612 477
rect 646 443 658 477
rect 600 297 658 443
rect 694 477 752 497
rect 694 443 706 477
rect 740 443 752 477
rect 694 409 752 443
rect 694 375 706 409
rect 740 375 752 409
rect 694 297 752 375
rect 788 477 857 497
rect 788 443 811 477
rect 845 443 857 477
rect 788 297 857 443
rect 893 477 947 497
rect 893 443 905 477
rect 939 443 947 477
rect 893 409 947 443
rect 893 375 905 409
rect 939 375 947 409
rect 893 297 947 375
rect 1001 477 1055 497
rect 1001 443 1009 477
rect 1043 443 1055 477
rect 1001 409 1055 443
rect 1001 375 1009 409
rect 1043 375 1055 409
rect 1001 297 1055 375
rect 1091 409 1149 497
rect 1091 375 1103 409
rect 1137 375 1149 409
rect 1091 341 1149 375
rect 1091 307 1103 341
rect 1137 307 1149 341
rect 1091 297 1149 307
rect 1185 477 1243 497
rect 1185 443 1197 477
rect 1231 443 1243 477
rect 1185 409 1243 443
rect 1185 375 1197 409
rect 1231 375 1243 409
rect 1185 297 1243 375
<< ndiffc >>
rect 38 61 72 95
rect 132 129 166 163
rect 132 61 166 95
rect 226 61 260 95
rect 320 129 354 163
rect 320 61 354 95
rect 414 61 448 95
rect 518 129 552 163
rect 518 61 552 95
rect 612 61 646 95
rect 706 91 740 125
rect 811 129 845 163
rect 905 61 939 95
rect 1009 61 1043 95
rect 1103 129 1137 163
rect 1197 61 1231 95
<< pdiffc >>
rect 38 443 72 477
rect 132 443 166 477
rect 226 443 260 477
rect 320 375 354 409
rect 414 443 448 477
rect 518 443 552 477
rect 518 375 552 409
rect 612 443 646 477
rect 706 443 740 477
rect 706 375 740 409
rect 811 443 845 477
rect 905 443 939 477
rect 905 375 939 409
rect 1009 443 1043 477
rect 1009 375 1043 409
rect 1103 375 1137 409
rect 1103 307 1137 341
rect 1197 443 1231 477
rect 1197 375 1231 409
<< poly >>
rect 84 497 120 523
rect 178 497 214 523
rect 272 497 308 523
rect 366 497 402 523
rect 564 497 600 523
rect 658 497 694 523
rect 752 497 788 523
rect 857 497 893 523
rect 1055 497 1091 523
rect 1149 497 1185 523
rect 84 282 120 297
rect 178 282 214 297
rect 272 282 308 297
rect 366 282 402 297
rect 564 282 600 297
rect 658 282 694 297
rect 752 282 788 297
rect 857 282 893 297
rect 1055 282 1091 297
rect 1149 282 1185 297
rect 82 265 122 282
rect 176 265 216 282
rect 270 265 310 282
rect 364 265 404 282
rect 562 265 602 282
rect 656 265 696 282
rect 750 265 790 282
rect 855 265 895 282
rect 82 249 216 265
rect 82 215 135 249
rect 169 215 216 249
rect 82 199 216 215
rect 268 249 404 265
rect 268 215 278 249
rect 312 215 404 249
rect 268 199 404 215
rect 558 249 700 265
rect 558 215 568 249
rect 602 215 646 249
rect 680 215 700 249
rect 558 199 700 215
rect 750 249 895 265
rect 750 215 760 249
rect 794 215 838 249
rect 872 215 895 249
rect 750 199 895 215
rect 82 177 112 199
rect 186 177 216 199
rect 280 177 310 199
rect 374 177 404 199
rect 572 177 602 199
rect 656 177 686 199
rect 750 177 780 199
rect 865 177 895 199
rect 1053 265 1093 282
rect 1147 265 1187 282
rect 1053 249 1187 265
rect 1053 215 1095 249
rect 1129 215 1187 249
rect 1053 199 1187 215
rect 1053 177 1083 199
rect 1157 177 1187 199
rect 82 21 112 47
rect 186 21 216 47
rect 280 21 310 47
rect 374 21 404 47
rect 572 21 602 47
rect 656 21 686 47
rect 750 21 780 47
rect 865 21 895 47
rect 1053 21 1083 47
rect 1157 21 1187 47
<< polycont >>
rect 135 215 169 249
rect 278 215 312 249
rect 568 215 602 249
rect 646 215 680 249
rect 760 215 794 249
rect 838 215 872 249
rect 1095 215 1129 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 24 477 80 493
rect 24 459 38 477
rect 24 427 29 459
rect 72 443 80 477
rect 63 427 80 443
rect 124 477 174 527
rect 124 443 132 477
rect 166 443 174 477
rect 124 427 174 443
rect 218 477 456 493
rect 218 443 226 477
rect 260 459 414 477
rect 218 427 233 443
rect 267 427 268 459
rect 406 443 414 459
rect 448 443 456 477
rect 406 427 456 443
rect 497 477 560 493
rect 497 443 518 477
rect 552 443 560 477
rect 497 425 560 443
rect 604 477 654 527
rect 604 443 612 477
rect 646 443 654 477
rect 604 427 654 443
rect 698 477 748 493
rect 698 443 706 477
rect 740 443 748 477
rect 312 409 362 425
rect 312 391 320 409
rect 24 375 320 391
rect 354 391 362 409
rect 518 409 560 425
rect 354 375 484 391
rect 24 357 484 375
rect 552 391 560 409
rect 698 409 748 443
rect 792 477 853 527
rect 792 443 811 477
rect 845 443 853 477
rect 792 427 853 443
rect 897 477 1239 493
rect 897 443 905 477
rect 939 443 1009 477
rect 1043 459 1197 477
rect 1043 443 1051 459
rect 698 391 706 409
rect 552 375 706 391
rect 740 391 748 409
rect 897 409 1051 443
rect 1189 443 1197 459
rect 1231 443 1239 477
rect 897 391 905 409
rect 740 375 905 391
rect 939 375 1009 409
rect 1043 375 1051 409
rect 518 357 1051 375
rect 1095 409 1145 425
rect 1095 375 1103 409
rect 1137 375 1145 409
rect 24 181 58 357
rect 450 323 484 357
rect 1095 341 1145 375
rect 1189 409 1239 443
rect 1189 375 1197 409
rect 1231 375 1239 409
rect 1189 359 1239 375
rect 151 289 416 323
rect 450 289 1037 323
rect 151 255 185 289
rect 372 255 416 289
rect 109 249 185 255
rect 109 215 135 249
rect 169 215 185 249
rect 229 221 233 255
rect 267 249 338 255
rect 267 221 278 249
rect 229 215 278 221
rect 312 215 338 249
rect 372 249 706 255
rect 372 215 568 249
rect 602 215 646 249
rect 680 215 706 249
rect 744 249 765 255
rect 799 249 898 255
rect 744 215 760 249
rect 799 221 838 249
rect 794 215 838 221
rect 872 215 898 249
rect 1003 249 1037 289
rect 1095 307 1103 341
rect 1137 325 1145 341
rect 1137 307 1270 325
rect 1095 283 1270 307
rect 1003 215 1095 249
rect 1129 215 1145 249
rect 1197 181 1270 283
rect 24 163 370 181
rect 24 145 132 163
rect 106 129 132 145
rect 166 145 320 163
rect 166 129 182 145
rect 38 95 72 111
rect 38 17 72 61
rect 106 95 182 129
rect 294 129 320 145
rect 354 129 370 163
rect 106 61 132 95
rect 166 61 182 95
rect 106 51 182 61
rect 226 95 260 111
rect 226 17 260 61
rect 294 95 370 129
rect 502 163 740 181
rect 502 129 518 163
rect 552 145 740 163
rect 552 129 568 145
rect 294 61 320 95
rect 354 61 370 95
rect 294 51 370 61
rect 414 95 448 111
rect 414 17 448 61
rect 502 95 568 129
rect 680 125 740 145
rect 795 163 1270 181
rect 795 129 811 163
rect 845 145 1103 163
rect 845 129 861 145
rect 1077 129 1103 145
rect 1137 145 1270 163
rect 1137 129 1153 145
rect 502 61 518 95
rect 552 61 568 95
rect 502 51 568 61
rect 612 95 646 111
rect 612 17 646 61
rect 680 91 706 125
rect 1009 95 1043 111
rect 740 91 905 95
rect 680 61 905 91
rect 939 61 956 95
rect 680 51 956 61
rect 1009 17 1043 61
rect 1197 95 1231 111
rect 1197 17 1231 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 443 38 459
rect 38 443 63 459
rect 29 425 63 443
rect 233 443 260 459
rect 260 443 267 459
rect 233 425 267 443
rect 233 221 267 255
rect 765 249 799 255
rect 765 221 794 249
rect 794 221 799 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 17 459 75 465
rect 17 425 29 459
rect 63 456 75 459
rect 221 459 279 465
rect 221 456 233 459
rect 63 428 233 456
rect 63 425 75 428
rect 17 419 75 425
rect 221 425 233 428
rect 267 425 279 459
rect 221 419 279 425
rect 221 255 279 261
rect 221 221 233 255
rect 267 252 279 255
rect 753 255 811 261
rect 753 252 765 255
rect 267 224 765 252
rect 267 221 279 224
rect 221 215 279 221
rect 753 221 765 224
rect 799 221 811 255
rect 753 215 811 221
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel metal1 s 765 221 799 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1225 289 1259 323 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel locali s 213 289 247 323 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 xor2_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1288 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 42966
string GDS_START 33408
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
