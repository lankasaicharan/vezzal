magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3698 1975
<< nwell >>
rect -38 331 2438 704
rect 1011 280 1440 331
<< pwell >>
rect 1 157 1522 207
rect 2203 165 2399 249
rect 2094 157 2399 165
rect 1 49 2399 157
rect 0 0 2400 49
<< scnmos >>
rect 84 97 114 181
rect 156 97 186 181
rect 250 97 280 181
rect 336 97 366 181
rect 408 97 438 181
rect 540 97 570 181
rect 612 97 642 181
rect 684 97 714 181
rect 816 97 846 181
rect 1039 97 1069 181
rect 1117 97 1147 181
rect 1189 97 1219 181
rect 1314 97 1344 181
rect 1386 97 1416 181
rect 1681 47 1711 131
rect 1799 47 1829 131
rect 1887 47 1917 131
rect 1959 47 1989 131
rect 2177 55 2207 139
rect 2286 55 2316 223
<< scpmoshvt >>
rect 84 487 114 615
rect 184 487 214 615
rect 307 487 337 615
rect 393 487 423 615
rect 465 487 495 615
rect 812 387 842 515
rect 1033 466 1063 594
rect 1165 466 1195 594
rect 1274 394 1324 594
rect 1515 419 1565 619
rect 1607 419 1657 619
rect 1715 419 1765 619
rect 1807 419 1857 619
rect 1959 419 2009 619
rect 2177 367 2207 495
rect 2286 367 2316 619
<< ndiff >>
rect 27 154 84 181
rect 27 120 39 154
rect 73 120 84 154
rect 27 97 84 120
rect 114 97 156 181
rect 186 148 250 181
rect 186 114 205 148
rect 239 114 250 148
rect 186 97 250 114
rect 280 148 336 181
rect 280 114 291 148
rect 325 114 336 148
rect 280 97 336 114
rect 366 97 408 181
rect 438 169 540 181
rect 438 135 472 169
rect 506 135 540 169
rect 438 97 540 135
rect 570 97 612 181
rect 642 97 684 181
rect 714 97 816 181
rect 846 156 903 181
rect 846 122 857 156
rect 891 122 903 156
rect 846 97 903 122
rect 982 160 1039 181
rect 982 126 994 160
rect 1028 126 1039 160
rect 982 97 1039 126
rect 1069 97 1117 181
rect 1147 97 1189 181
rect 1219 110 1314 181
rect 1219 97 1246 110
rect 736 71 794 97
rect 1234 76 1246 97
rect 1280 97 1314 110
rect 1344 97 1386 181
rect 1416 169 1496 181
rect 1416 135 1450 169
rect 1484 135 1496 169
rect 1416 97 1496 135
rect 2229 177 2286 223
rect 2229 143 2241 177
rect 2275 143 2286 177
rect 2229 139 2286 143
rect 1280 76 1292 97
rect 736 37 748 71
rect 782 37 794 71
rect 1234 64 1292 76
rect 1624 110 1681 131
rect 1624 76 1636 110
rect 1670 76 1681 110
rect 1624 47 1681 76
rect 1711 73 1799 131
rect 1711 47 1738 73
rect 736 27 794 37
rect 1726 39 1738 47
rect 1772 47 1799 73
rect 1829 110 1887 131
rect 1829 76 1841 110
rect 1875 76 1887 110
rect 1829 47 1887 76
rect 1917 47 1959 131
rect 1989 110 2046 131
rect 1989 76 2000 110
rect 2034 76 2046 110
rect 1989 47 2046 76
rect 2120 114 2177 139
rect 2120 80 2132 114
rect 2166 80 2177 114
rect 2120 55 2177 80
rect 2207 101 2286 139
rect 2207 67 2241 101
rect 2275 67 2286 101
rect 2207 55 2286 67
rect 2316 211 2373 223
rect 2316 177 2327 211
rect 2361 177 2373 211
rect 2316 101 2373 177
rect 2316 67 2327 101
rect 2361 67 2373 101
rect 2316 55 2373 67
rect 1772 39 1784 47
rect 1726 27 1784 39
<< pdiff >>
rect 864 629 922 639
rect 27 603 84 615
rect 27 569 39 603
rect 73 569 84 603
rect 27 487 84 569
rect 114 567 184 615
rect 114 533 139 567
rect 173 533 184 567
rect 114 487 184 533
rect 214 603 307 615
rect 214 569 248 603
rect 282 569 307 603
rect 214 535 307 569
rect 214 501 248 535
rect 282 501 307 535
rect 214 487 307 501
rect 337 566 393 615
rect 337 532 348 566
rect 382 532 393 566
rect 337 487 393 532
rect 423 487 465 615
rect 495 566 552 615
rect 495 532 506 566
rect 540 532 552 566
rect 864 595 876 629
rect 910 595 922 629
rect 495 487 552 532
rect 864 515 922 595
rect 732 425 812 515
rect 732 391 744 425
rect 778 391 812 425
rect 732 387 812 391
rect 842 387 922 515
rect 976 582 1033 594
rect 976 548 988 582
rect 1022 548 1033 582
rect 976 466 1033 548
rect 1063 466 1165 594
rect 1195 582 1274 594
rect 1195 548 1229 582
rect 1263 548 1274 582
rect 1195 466 1274 548
rect 732 380 790 387
rect 1085 362 1143 466
rect 1085 328 1097 362
rect 1131 328 1143 362
rect 1085 316 1143 328
rect 1217 394 1274 466
rect 1324 394 1404 594
rect 1458 498 1515 619
rect 1458 464 1470 498
rect 1504 464 1515 498
rect 1458 419 1515 464
rect 1565 419 1607 619
rect 1657 590 1715 619
rect 1657 556 1670 590
rect 1704 556 1715 590
rect 1657 419 1715 556
rect 1765 419 1807 619
rect 1857 599 1959 619
rect 1857 565 1891 599
rect 1925 565 1959 599
rect 1857 514 1959 565
rect 1857 480 1891 514
rect 1925 480 1959 514
rect 1857 419 1959 480
rect 2009 590 2066 619
rect 2009 556 2020 590
rect 2054 556 2066 590
rect 2009 419 2066 556
rect 2229 607 2286 619
rect 2229 573 2241 607
rect 2275 573 2286 607
rect 2229 510 2286 573
rect 2229 495 2241 510
rect 2120 482 2177 495
rect 2120 448 2132 482
rect 2166 448 2177 482
rect 1346 362 1404 394
rect 1346 328 1358 362
rect 1392 328 1404 362
rect 1346 316 1404 328
rect 2120 413 2177 448
rect 2120 379 2132 413
rect 2166 379 2177 413
rect 2120 367 2177 379
rect 2207 476 2241 495
rect 2275 476 2286 510
rect 2207 413 2286 476
rect 2207 379 2241 413
rect 2275 379 2286 413
rect 2207 367 2286 379
rect 2316 599 2373 619
rect 2316 565 2327 599
rect 2361 565 2373 599
rect 2316 506 2373 565
rect 2316 472 2327 506
rect 2361 472 2373 506
rect 2316 413 2373 472
rect 2316 379 2327 413
rect 2361 379 2373 413
rect 2316 367 2373 379
<< ndiffc >>
rect 39 120 73 154
rect 205 114 239 148
rect 291 114 325 148
rect 472 135 506 169
rect 857 122 891 156
rect 994 126 1028 160
rect 1246 76 1280 110
rect 1450 135 1484 169
rect 2241 143 2275 177
rect 748 37 782 71
rect 1636 76 1670 110
rect 1738 39 1772 73
rect 1841 76 1875 110
rect 2000 76 2034 110
rect 2132 80 2166 114
rect 2241 67 2275 101
rect 2327 177 2361 211
rect 2327 67 2361 101
<< pdiffc >>
rect 39 569 73 603
rect 139 533 173 567
rect 248 569 282 603
rect 248 501 282 535
rect 348 532 382 566
rect 506 532 540 566
rect 876 595 910 629
rect 744 391 778 425
rect 988 548 1022 582
rect 1229 548 1263 582
rect 1097 328 1131 362
rect 1470 464 1504 498
rect 1670 556 1704 590
rect 1891 565 1925 599
rect 1891 480 1925 514
rect 2020 556 2054 590
rect 2241 573 2275 607
rect 2132 448 2166 482
rect 1358 328 1392 362
rect 2132 379 2166 413
rect 2241 476 2275 510
rect 2241 379 2275 413
rect 2327 565 2361 599
rect 2327 472 2361 506
rect 2327 379 2361 413
<< poly >>
rect 84 615 114 641
rect 184 615 214 641
rect 307 615 337 641
rect 393 615 423 641
rect 465 615 495 641
rect 812 515 842 541
rect 1033 594 1063 620
rect 1165 594 1195 620
rect 1274 594 1324 620
rect 1515 619 1565 645
rect 1607 619 1657 645
rect 1715 619 1765 645
rect 1807 619 1857 645
rect 1959 619 2009 645
rect 2286 619 2316 645
rect 84 282 114 487
rect 184 451 214 487
rect 184 435 255 451
rect 184 415 205 435
rect 21 266 114 282
rect 21 232 37 266
rect 71 232 114 266
rect 21 216 114 232
rect 84 181 114 216
rect 156 401 205 415
rect 239 401 255 435
rect 156 385 255 401
rect 156 181 186 385
rect 307 337 337 487
rect 228 321 337 337
rect 393 365 423 487
rect 465 365 495 487
rect 812 365 842 387
rect 393 339 941 365
rect 393 335 891 339
rect 228 287 244 321
rect 278 307 337 321
rect 278 287 294 307
rect 228 253 294 287
rect 228 219 244 253
rect 278 219 294 253
rect 400 269 466 285
rect 400 249 416 269
rect 228 203 294 219
rect 336 235 416 249
rect 450 235 466 269
rect 336 219 466 235
rect 250 181 280 203
rect 336 181 366 219
rect 408 181 438 219
rect 540 181 570 335
rect 816 305 891 335
rect 925 305 941 339
rect 612 277 714 293
rect 612 243 628 277
rect 662 243 714 277
rect 612 227 714 243
rect 612 181 642 227
rect 684 181 714 227
rect 816 271 941 305
rect 1033 284 1063 466
rect 1165 294 1195 466
rect 2177 495 2207 521
rect 1274 294 1324 394
rect 816 237 891 271
rect 925 237 941 271
rect 816 221 941 237
rect 1009 268 1075 284
rect 1009 234 1025 268
rect 1059 234 1075 268
rect 1165 278 1344 294
rect 1165 258 1264 278
rect 816 181 846 221
rect 1009 218 1075 234
rect 1117 244 1264 258
rect 1298 258 1344 278
rect 1298 244 1416 258
rect 1117 228 1416 244
rect 1039 181 1069 218
rect 1117 181 1147 228
rect 1189 181 1219 228
rect 1314 181 1344 228
rect 1386 181 1416 228
rect 84 71 114 97
rect 156 71 186 97
rect 250 71 280 97
rect 336 71 366 97
rect 408 71 438 97
rect 540 71 570 97
rect 612 71 642 97
rect 684 71 714 97
rect 816 71 846 97
rect 1039 71 1069 97
rect 1117 71 1147 97
rect 1189 71 1219 97
rect 1515 117 1565 419
rect 1607 387 1657 419
rect 1607 371 1673 387
rect 1607 337 1623 371
rect 1657 337 1673 371
rect 1607 321 1673 337
rect 1715 261 1765 419
rect 1677 231 1765 261
rect 1807 387 1857 419
rect 1807 371 1911 387
rect 1807 337 1861 371
rect 1895 337 1911 371
rect 1807 321 1911 337
rect 1677 218 1745 231
rect 1677 184 1693 218
rect 1727 184 1745 218
rect 1677 168 1745 184
rect 1807 183 1837 321
rect 1959 273 2009 419
rect 1681 131 1711 168
rect 1799 153 1837 183
rect 1887 267 2009 273
rect 2177 267 2207 367
rect 2286 329 2316 367
rect 1887 257 2207 267
rect 2249 313 2316 329
rect 2249 279 2265 313
rect 2299 279 2316 313
rect 2249 263 2316 279
rect 1887 223 1903 257
rect 1937 237 2207 257
rect 1937 223 1989 237
rect 1887 207 1989 223
rect 1799 131 1829 153
rect 1887 131 1917 207
rect 1959 131 1989 207
rect 2177 139 2207 237
rect 2286 223 2316 263
rect 1515 101 1584 117
rect 1314 71 1344 97
rect 1386 71 1416 97
rect 1515 67 1534 101
rect 1568 67 1584 101
rect 1515 51 1584 67
rect 1681 21 1711 47
rect 1799 21 1829 47
rect 1887 21 1917 47
rect 1959 21 1989 47
rect 2177 29 2207 55
rect 2286 29 2316 55
<< polycont >>
rect 37 232 71 266
rect 205 401 239 435
rect 244 287 278 321
rect 244 219 278 253
rect 416 235 450 269
rect 891 305 925 339
rect 628 243 662 277
rect 891 237 925 271
rect 1025 234 1059 268
rect 1264 244 1298 278
rect 1623 337 1657 371
rect 1861 337 1895 371
rect 1693 184 1727 218
rect 2265 279 2299 313
rect 1903 223 1937 257
rect 1534 67 1568 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 23 603 89 649
rect 23 569 39 603
rect 73 569 89 603
rect 23 553 89 569
rect 123 567 189 615
rect 123 533 139 567
rect 173 533 189 567
rect 123 519 189 533
rect 121 485 189 519
rect 232 603 298 649
rect 860 629 926 649
rect 232 569 248 603
rect 282 569 298 603
rect 232 535 298 569
rect 232 501 248 535
rect 282 501 298 535
rect 232 485 298 501
rect 332 566 398 615
rect 332 532 348 566
rect 382 532 398 566
rect 121 350 155 485
rect 332 483 398 532
rect 490 566 556 615
rect 860 595 876 629
rect 910 595 926 629
rect 490 532 506 566
rect 540 532 556 566
rect 988 582 1127 598
rect 490 483 556 532
rect 189 435 263 451
rect 189 401 205 435
rect 239 424 263 435
rect 189 390 223 401
rect 257 390 263 424
rect 189 384 263 390
rect 121 321 294 350
rect 121 316 244 321
rect 21 266 87 282
rect 21 232 37 266
rect 71 232 87 266
rect 21 216 87 232
rect 121 182 155 316
rect 228 287 244 316
rect 278 287 294 321
rect 228 253 294 287
rect 228 219 244 253
rect 278 219 294 253
rect 228 203 294 219
rect 23 154 155 182
rect 332 169 366 483
rect 23 120 39 154
rect 73 148 155 154
rect 189 148 239 169
rect 73 120 89 148
rect 23 93 89 120
rect 189 114 205 148
rect 189 17 239 114
rect 275 148 366 169
rect 275 114 291 148
rect 325 114 366 148
rect 275 93 366 114
rect 400 269 466 285
rect 400 235 416 269
rect 450 235 466 269
rect 400 219 466 235
rect 400 85 434 219
rect 500 207 556 483
rect 592 527 954 561
rect 1022 581 1127 582
rect 1022 548 1087 581
rect 988 547 1087 548
rect 1121 547 1127 581
rect 988 532 1127 547
rect 1177 582 1279 598
rect 1177 581 1229 582
rect 1177 547 1183 581
rect 1217 548 1229 581
rect 1263 548 1279 582
rect 1217 547 1279 548
rect 1177 532 1279 547
rect 1313 581 1620 615
rect 592 289 626 527
rect 920 498 954 527
rect 1313 498 1347 581
rect 660 459 886 493
rect 920 464 1347 498
rect 1454 498 1552 547
rect 1454 464 1470 498
rect 1504 464 1552 498
rect 660 357 694 459
rect 852 430 886 459
rect 1454 430 1552 464
rect 728 391 744 425
rect 778 391 814 425
rect 852 396 1552 430
rect 660 323 746 357
rect 592 277 678 289
rect 592 243 628 277
rect 662 243 678 277
rect 592 241 678 243
rect 712 207 746 323
rect 500 185 746 207
rect 472 173 746 185
rect 780 185 814 391
rect 875 339 1097 362
rect 875 305 891 339
rect 925 328 1097 339
rect 1131 328 1147 362
rect 1342 328 1358 362
rect 1392 328 1408 362
rect 925 305 975 328
rect 875 271 975 305
rect 875 237 891 271
rect 925 237 975 271
rect 875 221 975 237
rect 472 169 534 173
rect 506 135 534 169
rect 780 156 907 185
rect 780 139 857 156
rect 472 119 534 135
rect 568 122 857 139
rect 891 122 907 156
rect 568 105 907 122
rect 941 184 975 221
rect 1009 268 1127 284
rect 1009 234 1025 268
rect 1059 234 1127 268
rect 1009 218 1127 234
rect 1177 278 1319 294
rect 1177 244 1264 278
rect 1298 244 1319 278
rect 1177 228 1319 244
rect 1374 262 1408 328
rect 1518 295 1552 396
rect 1586 498 1620 581
rect 1654 590 1720 615
rect 1654 581 1670 590
rect 1654 547 1663 581
rect 1704 556 1720 590
rect 1697 547 1720 556
rect 1654 532 1720 547
rect 1875 599 1941 615
rect 1875 565 1891 599
rect 1925 565 1941 599
rect 1875 514 1941 565
rect 2004 590 2087 615
rect 2004 556 2020 590
rect 2054 581 2087 590
rect 2004 547 2047 556
rect 2081 547 2087 581
rect 2004 532 2087 547
rect 2225 607 2275 649
rect 2225 573 2241 607
rect 1875 498 1891 514
rect 1586 480 1891 498
rect 1925 498 1941 514
rect 2225 510 2275 573
rect 1925 480 2059 498
rect 1586 464 2059 480
rect 1586 387 1620 464
rect 1845 424 1991 430
rect 1845 390 1855 424
rect 1889 390 1991 424
rect 1586 371 1673 387
rect 1586 337 1623 371
rect 1657 337 1673 371
rect 1586 329 1673 337
rect 1845 371 1991 390
rect 1845 337 1861 371
rect 1895 337 1991 371
rect 1845 310 1991 337
rect 1518 273 1811 295
rect 1374 228 1484 262
rect 1518 261 1953 273
rect 1434 227 1484 228
rect 1777 257 1953 261
rect 1434 218 1743 227
rect 941 160 1044 184
rect 941 126 994 160
rect 1028 126 1044 160
rect 941 119 1044 126
rect 1161 160 1400 194
rect 568 85 602 105
rect 400 51 602 85
rect 841 85 907 105
rect 1161 85 1195 160
rect 732 37 748 71
rect 782 37 798 71
rect 841 51 1195 85
rect 1230 110 1296 126
rect 1230 76 1246 110
rect 1280 76 1296 110
rect 732 17 798 37
rect 1230 17 1296 76
rect 1366 85 1400 160
rect 1434 184 1693 218
rect 1727 184 1743 218
rect 1777 223 1903 257
rect 1937 223 1953 257
rect 1777 207 1953 223
rect 1434 175 1743 184
rect 1434 169 1484 175
rect 1434 135 1450 169
rect 1434 119 1484 135
rect 1518 101 1584 117
rect 1518 85 1534 101
rect 1366 67 1534 85
rect 1568 67 1584 101
rect 1366 51 1584 67
rect 1636 110 1891 141
rect 2025 135 2059 464
rect 1670 107 1841 110
rect 1670 76 1686 107
rect 1636 51 1686 76
rect 1825 76 1841 107
rect 1875 76 1891 110
rect 1722 39 1738 73
rect 1772 39 1788 73
rect 1825 51 1891 76
rect 1984 110 2059 135
rect 1984 76 2000 110
rect 2034 76 2059 110
rect 1984 51 2059 76
rect 2116 482 2182 498
rect 2116 448 2132 482
rect 2166 448 2182 482
rect 2116 413 2182 448
rect 2116 379 2132 413
rect 2166 379 2182 413
rect 2116 329 2182 379
rect 2225 476 2241 510
rect 2225 413 2275 476
rect 2225 379 2241 413
rect 2225 363 2275 379
rect 2311 599 2383 615
rect 2311 565 2327 599
rect 2361 565 2383 599
rect 2311 506 2383 565
rect 2311 472 2327 506
rect 2361 472 2383 506
rect 2311 413 2383 472
rect 2311 379 2327 413
rect 2361 379 2383 413
rect 2311 363 2383 379
rect 2116 313 2315 329
rect 2116 279 2265 313
rect 2299 279 2315 313
rect 2116 263 2315 279
rect 2116 114 2182 263
rect 2349 227 2383 363
rect 2311 211 2383 227
rect 2116 80 2132 114
rect 2166 80 2182 114
rect 2116 51 2182 80
rect 2225 177 2275 193
rect 2225 143 2241 177
rect 2225 101 2275 143
rect 2225 67 2241 101
rect 1722 17 1788 39
rect 2225 17 2275 67
rect 2311 177 2327 211
rect 2361 177 2383 211
rect 2311 101 2383 177
rect 2311 67 2327 101
rect 2361 67 2383 101
rect 2311 51 2383 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 223 401 239 424
rect 239 401 257 424
rect 223 390 257 401
rect 1087 547 1121 581
rect 1183 547 1217 581
rect 1663 556 1670 581
rect 1670 556 1697 581
rect 1663 547 1697 556
rect 2047 556 2054 581
rect 2054 556 2081 581
rect 2047 547 2081 556
rect 1855 390 1889 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
<< metal1 >>
rect 0 683 2400 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2400 683
rect 0 617 2400 649
rect 14 581 2386 589
rect 14 547 1087 581
rect 1121 547 1183 581
rect 1217 547 1663 581
rect 1697 547 2047 581
rect 2081 547 2386 581
rect 14 535 2386 547
rect 211 424 269 430
rect 211 390 223 424
rect 257 421 269 424
rect 1843 424 1901 430
rect 1843 421 1855 424
rect 257 393 1855 421
rect 257 390 269 393
rect 211 384 269 390
rect 1843 390 1855 393
rect 1889 390 1901 424
rect 1843 384 1901 390
rect 0 17 2400 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2400 17
rect 0 -49 2400 -17
<< labels >>
flabel pwell s 0 0 2400 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2400 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 srdlrtp_1
flabel metal1 s 14 535 2386 589 0 FreeSans 200 0 0 0 KAPWR
port 5 nsew power bidirectional
flabel metal1 s 1855 390 1889 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel metal1 s 0 617 2400 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2400 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 2335 94 2369 128 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 2335 168 2369 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 SLEEP_B
port 4 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 SLEEP_B
port 4 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2400 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5377920
string GDS_START 5361896
<< end >>
