magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 4850 1975
<< nwell >>
rect -38 332 3590 704
<< pwell >>
rect 658 191 954 248
rect 658 184 1452 191
rect 1768 184 2264 228
rect 2848 184 3551 248
rect 1 49 3551 184
rect 0 0 3552 49
<< scpmos >>
rect 90 464 120 592
rect 190 464 220 592
rect 274 464 304 592
rect 388 464 418 592
rect 472 464 502 592
rect 678 368 708 592
rect 844 368 874 592
rect 1071 463 1101 547
rect 1171 463 1201 547
rect 1255 463 1285 547
rect 1472 463 1502 547
rect 1582 463 1612 547
rect 1858 424 1888 592
rect 1948 424 1978 592
rect 2038 424 2068 592
rect 2128 424 2158 592
rect 2337 455 2367 539
rect 2545 508 2575 592
rect 2635 508 2665 592
rect 2837 494 2867 578
rect 2944 368 2974 592
rect 3034 368 3064 592
rect 3236 368 3266 568
rect 3346 368 3376 592
rect 3436 368 3466 592
<< nmoslvt >>
rect 84 74 114 158
rect 199 74 229 158
rect 277 74 307 158
rect 465 74 495 158
rect 543 74 573 158
rect 741 74 771 222
rect 841 74 871 222
rect 1039 81 1069 165
rect 1244 81 1274 165
rect 1322 81 1352 165
rect 1537 74 1567 158
rect 1615 74 1645 158
rect 1861 74 1891 202
rect 1951 74 1981 202
rect 2037 74 2067 202
rect 2137 74 2167 202
rect 2471 74 2501 158
rect 2549 74 2579 158
rect 2627 74 2657 158
rect 2729 74 2759 158
rect 2941 74 2971 222
rect 3031 74 3061 222
rect 3239 94 3269 222
rect 3352 74 3382 222
rect 3438 74 3468 222
<< ndiff >>
rect 684 186 741 222
rect 27 133 84 158
rect 27 99 39 133
rect 73 99 84 133
rect 27 74 84 99
rect 114 120 199 158
rect 114 86 146 120
rect 180 86 199 120
rect 114 74 199 86
rect 229 74 277 158
rect 307 130 465 158
rect 307 96 414 130
rect 448 96 465 130
rect 307 74 465 96
rect 495 74 543 158
rect 573 130 630 158
rect 573 96 584 130
rect 618 96 630 130
rect 573 74 630 96
rect 684 152 696 186
rect 730 152 741 186
rect 684 118 741 152
rect 684 84 696 118
rect 730 84 741 118
rect 684 74 741 84
rect 771 186 841 222
rect 771 152 782 186
rect 816 152 841 186
rect 771 118 841 152
rect 771 84 782 118
rect 816 84 841 118
rect 771 74 841 84
rect 871 186 928 222
rect 871 152 882 186
rect 916 152 928 186
rect 871 118 928 152
rect 871 84 882 118
rect 916 84 928 118
rect 871 74 928 84
rect 982 153 1039 165
rect 982 119 994 153
rect 1028 119 1039 153
rect 982 81 1039 119
rect 1069 144 1244 165
rect 1069 110 1180 144
rect 1214 110 1244 144
rect 1069 81 1244 110
rect 1274 81 1322 165
rect 1352 124 1426 165
rect 1794 190 1861 202
rect 1352 90 1363 124
rect 1397 90 1426 124
rect 1352 81 1426 90
rect 1480 133 1537 158
rect 1480 99 1492 133
rect 1526 99 1537 133
rect 1480 74 1537 99
rect 1567 74 1615 158
rect 1645 120 1735 158
rect 1645 86 1656 120
rect 1690 86 1735 120
rect 1645 74 1735 86
rect 1794 156 1806 190
rect 1840 156 1861 190
rect 1794 120 1861 156
rect 1794 86 1806 120
rect 1840 86 1861 120
rect 1794 74 1861 86
rect 1891 135 1951 202
rect 1891 101 1906 135
rect 1940 101 1951 135
rect 1891 74 1951 101
rect 1981 190 2037 202
rect 1981 156 1992 190
rect 2026 156 2037 190
rect 1981 120 2037 156
rect 1981 86 1992 120
rect 2026 86 2037 120
rect 1981 74 2037 86
rect 2067 179 2137 202
rect 2067 145 2092 179
rect 2126 145 2137 179
rect 2067 74 2137 145
rect 2167 121 2238 202
rect 2167 87 2192 121
rect 2226 87 2238 121
rect 2167 74 2238 87
rect 2292 130 2471 158
rect 2292 96 2304 130
rect 2338 96 2426 130
rect 2460 96 2471 130
rect 2292 74 2471 96
rect 2501 74 2549 158
rect 2579 74 2627 158
rect 2657 131 2729 158
rect 2657 97 2668 131
rect 2702 97 2729 131
rect 2657 74 2729 97
rect 2759 133 2816 158
rect 2759 99 2770 133
rect 2804 99 2816 133
rect 2759 74 2816 99
rect 2874 142 2941 222
rect 2874 108 2886 142
rect 2920 108 2941 142
rect 2874 74 2941 108
rect 2971 210 3031 222
rect 2971 176 2986 210
rect 3020 176 3031 210
rect 2971 120 3031 176
rect 2971 86 2986 120
rect 3020 86 3031 120
rect 2971 74 3031 86
rect 3061 210 3127 222
rect 3061 176 3081 210
rect 3115 176 3127 210
rect 3061 120 3127 176
rect 3061 86 3081 120
rect 3115 86 3127 120
rect 3182 210 3239 222
rect 3182 176 3194 210
rect 3228 176 3239 210
rect 3182 140 3239 176
rect 3182 106 3194 140
rect 3228 106 3239 140
rect 3182 94 3239 106
rect 3269 210 3352 222
rect 3269 176 3307 210
rect 3341 176 3352 210
rect 3269 120 3352 176
rect 3269 94 3307 120
rect 3061 74 3127 86
rect 3295 86 3307 94
rect 3341 86 3352 120
rect 3295 74 3352 86
rect 3382 210 3438 222
rect 3382 176 3393 210
rect 3427 176 3438 210
rect 3382 120 3438 176
rect 3382 86 3393 120
rect 3427 86 3438 120
rect 3382 74 3438 86
rect 3468 210 3525 222
rect 3468 176 3479 210
rect 3513 176 3525 210
rect 3468 120 3525 176
rect 3468 86 3479 120
rect 3513 86 3525 120
rect 3468 74 3525 86
<< pdiff >>
rect 31 580 90 592
rect 31 546 43 580
rect 77 546 90 580
rect 31 510 90 546
rect 31 476 43 510
rect 77 476 90 510
rect 31 464 90 476
rect 120 580 190 592
rect 120 546 143 580
rect 177 546 190 580
rect 120 512 190 546
rect 120 478 143 512
rect 177 478 190 512
rect 120 464 190 478
rect 220 464 274 592
rect 304 580 388 592
rect 304 546 329 580
rect 363 546 388 580
rect 304 510 388 546
rect 304 476 329 510
rect 363 476 388 510
rect 304 464 388 476
rect 418 464 472 592
rect 502 580 565 592
rect 502 546 517 580
rect 551 546 565 580
rect 502 464 565 546
rect 619 421 678 592
rect 619 387 631 421
rect 665 387 678 421
rect 619 368 678 387
rect 708 580 844 592
rect 708 546 721 580
rect 755 546 794 580
rect 828 546 844 580
rect 708 368 844 546
rect 874 562 940 592
rect 874 528 894 562
rect 928 528 940 562
rect 874 368 940 528
rect 1012 520 1071 547
rect 1012 486 1024 520
rect 1058 486 1071 520
rect 1012 463 1071 486
rect 1101 520 1171 547
rect 1101 486 1124 520
rect 1158 486 1171 520
rect 1101 463 1171 486
rect 1201 463 1255 547
rect 1285 535 1472 547
rect 1285 501 1322 535
rect 1356 501 1472 535
rect 1285 463 1472 501
rect 1502 520 1582 547
rect 1502 486 1515 520
rect 1549 486 1582 520
rect 1502 463 1582 486
rect 1612 531 1729 547
rect 1612 497 1683 531
rect 1717 497 1729 531
rect 1612 463 1729 497
rect 1789 580 1858 592
rect 1789 546 1801 580
rect 1835 546 1858 580
rect 1789 476 1858 546
rect 1789 442 1801 476
rect 1835 442 1858 476
rect 1789 424 1858 442
rect 1888 562 1948 592
rect 1888 528 1901 562
rect 1935 528 1948 562
rect 1888 424 1948 528
rect 1978 580 2038 592
rect 1978 546 1991 580
rect 2025 546 2038 580
rect 1978 470 2038 546
rect 1978 436 1991 470
rect 2025 436 2038 470
rect 1978 424 2038 436
rect 2068 509 2128 592
rect 2068 475 2081 509
rect 2115 475 2128 509
rect 2068 424 2128 475
rect 2158 580 2217 592
rect 2158 546 2171 580
rect 2205 546 2217 580
rect 2158 510 2217 546
rect 2158 476 2171 510
rect 2205 476 2217 510
rect 2158 424 2217 476
rect 2277 527 2337 539
rect 2277 493 2289 527
rect 2323 493 2337 527
rect 2277 455 2337 493
rect 2367 514 2426 539
rect 2367 480 2380 514
rect 2414 480 2426 514
rect 2367 455 2426 480
rect 2486 567 2545 592
rect 2486 533 2498 567
rect 2532 533 2545 567
rect 2486 508 2545 533
rect 2575 567 2635 592
rect 2575 533 2588 567
rect 2622 533 2635 567
rect 2575 508 2635 533
rect 2665 567 2724 592
rect 2885 580 2944 592
rect 2885 578 2897 580
rect 2665 533 2678 567
rect 2712 533 2724 567
rect 2665 508 2724 533
rect 2778 556 2837 578
rect 2778 522 2790 556
rect 2824 522 2837 556
rect 2778 494 2837 522
rect 2867 546 2897 578
rect 2931 546 2944 580
rect 2867 497 2944 546
rect 2867 494 2897 497
rect 2885 463 2897 494
rect 2931 463 2944 497
rect 2885 414 2944 463
rect 2885 380 2897 414
rect 2931 380 2944 414
rect 2885 368 2944 380
rect 2974 580 3034 592
rect 2974 546 2987 580
rect 3021 546 3034 580
rect 2974 497 3034 546
rect 2974 463 2987 497
rect 3021 463 3034 497
rect 2974 414 3034 463
rect 2974 380 2987 414
rect 3021 380 3034 414
rect 2974 368 3034 380
rect 3064 580 3123 592
rect 3064 546 3077 580
rect 3111 546 3123 580
rect 3287 580 3346 592
rect 3287 568 3299 580
rect 3064 497 3123 546
rect 3064 463 3077 497
rect 3111 463 3123 497
rect 3064 414 3123 463
rect 3064 380 3077 414
rect 3111 380 3123 414
rect 3064 368 3123 380
rect 3177 556 3236 568
rect 3177 522 3189 556
rect 3223 522 3236 556
rect 3177 485 3236 522
rect 3177 451 3189 485
rect 3223 451 3236 485
rect 3177 414 3236 451
rect 3177 380 3189 414
rect 3223 380 3236 414
rect 3177 368 3236 380
rect 3266 546 3299 568
rect 3333 546 3346 580
rect 3266 497 3346 546
rect 3266 463 3299 497
rect 3333 463 3346 497
rect 3266 414 3346 463
rect 3266 380 3299 414
rect 3333 380 3346 414
rect 3266 368 3346 380
rect 3376 580 3436 592
rect 3376 546 3389 580
rect 3423 546 3436 580
rect 3376 497 3436 546
rect 3376 463 3389 497
rect 3423 463 3436 497
rect 3376 414 3436 463
rect 3376 380 3389 414
rect 3423 380 3436 414
rect 3376 368 3436 380
rect 3466 580 3525 592
rect 3466 546 3479 580
rect 3513 546 3525 580
rect 3466 497 3525 546
rect 3466 463 3479 497
rect 3513 463 3525 497
rect 3466 414 3525 463
rect 3466 380 3479 414
rect 3513 380 3525 414
rect 3466 368 3525 380
<< ndiffc >>
rect 39 99 73 133
rect 146 86 180 120
rect 414 96 448 130
rect 584 96 618 130
rect 696 152 730 186
rect 696 84 730 118
rect 782 152 816 186
rect 782 84 816 118
rect 882 152 916 186
rect 882 84 916 118
rect 994 119 1028 153
rect 1180 110 1214 144
rect 1363 90 1397 124
rect 1492 99 1526 133
rect 1656 86 1690 120
rect 1806 156 1840 190
rect 1806 86 1840 120
rect 1906 101 1940 135
rect 1992 156 2026 190
rect 1992 86 2026 120
rect 2092 145 2126 179
rect 2192 87 2226 121
rect 2304 96 2338 130
rect 2426 96 2460 130
rect 2668 97 2702 131
rect 2770 99 2804 133
rect 2886 108 2920 142
rect 2986 176 3020 210
rect 2986 86 3020 120
rect 3081 176 3115 210
rect 3081 86 3115 120
rect 3194 176 3228 210
rect 3194 106 3228 140
rect 3307 176 3341 210
rect 3307 86 3341 120
rect 3393 176 3427 210
rect 3393 86 3427 120
rect 3479 176 3513 210
rect 3479 86 3513 120
<< pdiffc >>
rect 43 546 77 580
rect 43 476 77 510
rect 143 546 177 580
rect 143 478 177 512
rect 329 546 363 580
rect 329 476 363 510
rect 517 546 551 580
rect 631 387 665 421
rect 721 546 755 580
rect 794 546 828 580
rect 894 528 928 562
rect 1024 486 1058 520
rect 1124 486 1158 520
rect 1322 501 1356 535
rect 1515 486 1549 520
rect 1683 497 1717 531
rect 1801 546 1835 580
rect 1801 442 1835 476
rect 1901 528 1935 562
rect 1991 546 2025 580
rect 1991 436 2025 470
rect 2081 475 2115 509
rect 2171 546 2205 580
rect 2171 476 2205 510
rect 2289 493 2323 527
rect 2380 480 2414 514
rect 2498 533 2532 567
rect 2588 533 2622 567
rect 2678 533 2712 567
rect 2790 522 2824 556
rect 2897 546 2931 580
rect 2897 463 2931 497
rect 2897 380 2931 414
rect 2987 546 3021 580
rect 2987 463 3021 497
rect 2987 380 3021 414
rect 3077 546 3111 580
rect 3077 463 3111 497
rect 3077 380 3111 414
rect 3189 522 3223 556
rect 3189 451 3223 485
rect 3189 380 3223 414
rect 3299 546 3333 580
rect 3299 463 3333 497
rect 3299 380 3333 414
rect 3389 546 3423 580
rect 3389 463 3423 497
rect 3389 380 3423 414
rect 3479 546 3513 580
rect 3479 463 3513 497
rect 3479 380 3513 414
<< poly >>
rect 90 592 120 618
rect 190 592 220 618
rect 274 592 304 618
rect 388 592 418 618
rect 472 592 502 618
rect 678 592 708 618
rect 844 592 874 618
rect 955 615 1774 645
rect 90 449 120 464
rect 190 449 220 464
rect 274 449 304 464
rect 388 449 418 464
rect 472 449 502 464
rect 87 360 123 449
rect 187 360 223 449
rect 83 344 223 360
rect 83 310 99 344
rect 133 310 167 344
rect 201 330 223 344
rect 201 310 217 330
rect 83 294 217 310
rect 271 294 307 449
rect 385 428 421 449
rect 355 412 421 428
rect 355 378 371 412
rect 405 378 421 412
rect 355 362 421 378
rect 469 392 505 449
rect 469 362 573 392
rect 543 324 573 362
rect 678 353 708 368
rect 844 353 874 368
rect 84 158 114 294
rect 277 246 307 294
rect 393 298 495 314
rect 393 264 409 298
rect 443 264 495 298
rect 163 230 229 246
rect 163 196 179 230
rect 213 196 229 230
rect 163 180 229 196
rect 199 158 229 180
rect 277 230 343 246
rect 277 196 293 230
rect 327 196 343 230
rect 277 180 343 196
rect 393 230 495 264
rect 393 196 409 230
rect 443 196 495 230
rect 393 180 495 196
rect 277 158 307 180
rect 465 158 495 180
rect 543 308 627 324
rect 543 274 577 308
rect 611 274 627 308
rect 543 240 627 274
rect 675 310 711 353
rect 841 336 877 353
rect 955 336 985 615
rect 1071 547 1101 573
rect 1168 562 1204 615
rect 1171 547 1201 562
rect 1255 547 1285 573
rect 1472 547 1502 573
rect 1582 547 1612 573
rect 1071 448 1101 463
rect 1068 392 1104 448
rect 1171 437 1201 463
rect 1255 448 1285 463
rect 1472 448 1502 463
rect 1582 448 1612 463
rect 1252 406 1288 448
rect 841 320 985 336
rect 675 294 799 310
rect 675 260 749 294
rect 783 260 799 294
rect 675 244 799 260
rect 841 286 894 320
rect 928 286 985 320
rect 841 270 985 286
rect 543 206 577 240
rect 611 206 627 240
rect 741 222 771 244
rect 841 222 871 270
rect 543 190 627 206
rect 543 158 573 190
rect 955 210 985 270
rect 1046 376 1112 392
rect 1252 390 1393 406
rect 1252 376 1343 390
rect 1046 342 1062 376
rect 1096 342 1112 376
rect 1046 308 1112 342
rect 1327 356 1343 376
rect 1377 356 1393 390
rect 1327 340 1393 356
rect 1046 274 1062 308
rect 1096 288 1112 308
rect 1204 312 1274 328
rect 1204 288 1220 312
rect 1096 278 1220 288
rect 1254 278 1274 312
rect 1096 274 1274 278
rect 1046 258 1274 274
rect 1204 244 1274 258
rect 1204 210 1220 244
rect 1254 210 1274 244
rect 1363 253 1393 340
rect 1469 310 1505 448
rect 1579 376 1615 448
rect 1744 392 1774 615
rect 1858 592 1888 618
rect 1948 592 1978 618
rect 2038 592 2068 618
rect 2128 592 2158 618
rect 2232 613 2471 643
rect 1858 409 1888 424
rect 1948 409 1978 424
rect 2038 409 2068 424
rect 2128 409 2158 424
rect 2232 409 2262 613
rect 2337 539 2367 565
rect 2337 440 2367 455
rect 1744 376 1813 392
rect 1579 360 1645 376
rect 1579 326 1595 360
rect 1629 326 1645 360
rect 1744 342 1763 376
rect 1797 342 1813 376
rect 1744 326 1813 342
rect 1579 310 1645 326
rect 1471 308 1505 310
rect 1471 292 1537 308
rect 1471 258 1487 292
rect 1521 262 1537 292
rect 1521 258 1567 262
rect 1363 237 1429 253
rect 1363 217 1379 237
rect 955 180 1069 210
rect 1204 194 1274 210
rect 1039 165 1069 180
rect 1244 165 1274 194
rect 1322 203 1379 217
rect 1413 203 1429 237
rect 1471 232 1567 258
rect 1322 187 1429 203
rect 1322 165 1352 187
rect 1537 158 1567 232
rect 1615 158 1645 310
rect 1855 277 1891 409
rect 1945 277 1981 409
rect 2035 379 2262 409
rect 2334 324 2370 440
rect 1855 247 1981 277
rect 2076 294 2370 324
rect 2076 290 2278 294
rect 2076 270 2092 290
rect 1706 230 1891 247
rect 1706 196 1722 230
rect 1756 217 1891 230
rect 1756 196 1772 217
rect 1861 202 1891 217
rect 1951 202 1981 247
rect 2037 256 2092 270
rect 2126 256 2160 290
rect 2194 256 2228 290
rect 2262 256 2278 290
rect 2037 240 2278 256
rect 2441 246 2471 613
rect 2545 592 2575 618
rect 2635 592 2665 618
rect 2837 578 2867 604
rect 2944 592 2974 618
rect 3034 592 3064 618
rect 2545 493 2575 508
rect 2635 493 2665 508
rect 2542 392 2578 493
rect 2632 394 2668 493
rect 2837 479 2867 494
rect 2834 462 2870 479
rect 2729 446 2870 462
rect 2729 412 2745 446
rect 2779 432 2870 446
rect 2779 412 2795 432
rect 2513 376 2579 392
rect 2513 342 2529 376
rect 2563 342 2579 376
rect 2513 308 2579 342
rect 2513 274 2529 308
rect 2563 274 2579 308
rect 2513 258 2579 274
rect 2621 378 2687 394
rect 2621 344 2637 378
rect 2671 344 2687 378
rect 2621 310 2687 344
rect 2621 276 2637 310
rect 2671 276 2687 310
rect 2621 260 2687 276
rect 2729 378 2795 412
rect 2729 344 2745 378
rect 2779 344 2795 378
rect 3236 568 3266 594
rect 3346 592 3376 618
rect 3436 592 3466 618
rect 2944 353 2974 368
rect 3034 353 3064 368
rect 3236 353 3266 368
rect 3346 353 3376 368
rect 3436 353 3466 368
rect 2729 310 2795 344
rect 2729 276 2745 310
rect 2779 290 2795 310
rect 2941 290 2977 353
rect 3031 290 3067 353
rect 3233 290 3269 353
rect 3343 326 3379 353
rect 3433 326 3469 353
rect 2779 276 3269 290
rect 2729 260 3269 276
rect 3311 310 3469 326
rect 3311 276 3327 310
rect 3361 290 3469 310
rect 3361 276 3468 290
rect 3311 260 3468 276
rect 2037 202 2067 240
rect 2137 202 2167 240
rect 2344 230 2471 246
rect 1706 180 1772 196
rect 84 48 114 74
rect 199 48 229 74
rect 277 48 307 74
rect 465 48 495 74
rect 543 48 573 74
rect 741 48 771 74
rect 841 48 871 74
rect 1039 55 1069 81
rect 1244 55 1274 81
rect 1322 55 1352 81
rect 2344 196 2360 230
rect 2394 210 2471 230
rect 2394 196 2501 210
rect 2344 180 2501 196
rect 2471 158 2501 180
rect 2549 158 2579 258
rect 2627 158 2657 260
rect 2729 158 2759 260
rect 2941 222 2971 260
rect 3031 222 3061 260
rect 3239 222 3269 260
rect 3352 222 3382 260
rect 3438 222 3468 260
rect 1537 48 1567 74
rect 1615 48 1645 74
rect 1861 48 1891 74
rect 1951 48 1981 74
rect 2037 48 2067 74
rect 2137 48 2167 74
rect 2471 48 2501 74
rect 2549 48 2579 74
rect 2627 48 2657 74
rect 2729 48 2759 74
rect 2941 48 2971 74
rect 3031 48 3061 74
rect 3239 68 3269 94
rect 3352 48 3382 74
rect 3438 48 3468 74
<< polycont >>
rect 99 310 133 344
rect 167 310 201 344
rect 371 378 405 412
rect 409 264 443 298
rect 179 196 213 230
rect 293 196 327 230
rect 409 196 443 230
rect 577 274 611 308
rect 749 260 783 294
rect 894 286 928 320
rect 577 206 611 240
rect 1062 342 1096 376
rect 1343 356 1377 390
rect 1062 274 1096 308
rect 1220 278 1254 312
rect 1220 210 1254 244
rect 1595 326 1629 360
rect 1763 342 1797 376
rect 1487 258 1521 292
rect 1379 203 1413 237
rect 1722 196 1756 230
rect 2092 256 2126 290
rect 2160 256 2194 290
rect 2228 256 2262 290
rect 2745 412 2779 446
rect 2529 342 2563 376
rect 2529 274 2563 308
rect 2637 344 2671 378
rect 2637 276 2671 310
rect 2745 344 2779 378
rect 2745 276 2779 310
rect 3327 276 3361 310
rect 2360 196 2394 230
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3552 683
rect 17 580 93 596
rect 17 546 43 580
rect 77 546 93 580
rect 17 510 93 546
rect 17 476 43 510
rect 77 476 93 510
rect 17 428 93 476
rect 127 580 193 649
rect 127 546 143 580
rect 177 546 193 580
rect 127 512 193 546
rect 127 478 143 512
rect 177 478 193 512
rect 127 462 193 478
rect 301 580 391 596
rect 301 546 329 580
rect 363 546 391 580
rect 301 510 391 546
rect 499 580 569 649
rect 499 546 517 580
rect 551 546 569 580
rect 499 530 569 546
rect 705 580 844 649
rect 705 546 721 580
rect 755 546 794 580
rect 828 546 844 580
rect 705 530 844 546
rect 878 581 1248 615
rect 878 562 944 581
rect 301 476 329 510
rect 363 496 391 510
rect 878 528 894 562
rect 928 528 944 562
rect 363 476 777 496
rect 878 494 944 528
rect 978 520 1074 547
rect 301 462 777 476
rect 17 412 421 428
rect 17 394 371 412
rect 17 246 51 394
rect 355 378 371 394
rect 405 378 421 412
rect 355 362 421 378
rect 85 344 217 360
rect 85 310 99 344
rect 133 310 167 344
rect 201 314 217 344
rect 201 310 459 314
rect 85 298 459 310
rect 85 280 409 298
rect 393 264 409 280
rect 443 264 459 298
rect 17 230 229 246
rect 17 196 179 230
rect 213 196 229 230
rect 17 180 229 196
rect 277 230 359 246
rect 277 196 293 230
rect 327 196 359 230
rect 17 133 89 180
rect 17 99 39 133
rect 73 99 89 133
rect 17 70 89 99
rect 123 120 204 136
rect 123 86 146 120
rect 180 86 204 120
rect 277 88 359 196
rect 393 230 459 264
rect 393 196 409 230
rect 443 196 459 230
rect 393 180 459 196
rect 493 146 527 462
rect 743 460 777 462
rect 978 486 1024 520
rect 1058 486 1074 520
rect 978 460 1074 486
rect 615 421 709 428
rect 743 426 1074 460
rect 1108 520 1180 547
rect 1108 486 1124 520
rect 1158 486 1180 520
rect 1108 459 1180 486
rect 615 387 631 421
rect 665 392 709 421
rect 665 387 944 392
rect 615 358 944 387
rect 561 308 641 324
rect 561 274 577 308
rect 611 274 641 308
rect 561 240 641 274
rect 561 206 577 240
rect 611 206 641 240
rect 561 190 641 206
rect 675 202 709 358
rect 878 320 944 358
rect 743 294 839 310
rect 743 260 749 294
rect 783 260 839 294
rect 878 286 894 320
rect 928 286 944 320
rect 878 270 944 286
rect 743 236 839 260
rect 675 186 730 202
rect 393 130 527 146
rect 393 96 414 130
rect 448 112 527 130
rect 568 130 634 156
rect 448 96 470 112
rect 123 17 204 86
rect 393 80 470 96
rect 568 96 584 130
rect 618 96 634 130
rect 568 17 634 96
rect 675 152 696 186
rect 675 118 730 152
rect 675 84 696 118
rect 675 68 730 84
rect 766 186 832 202
rect 766 152 782 186
rect 816 152 832 186
rect 766 118 832 152
rect 766 84 782 118
rect 816 84 832 118
rect 766 17 832 84
rect 866 186 932 202
rect 866 152 882 186
rect 916 152 932 186
rect 866 118 932 152
rect 978 169 1012 426
rect 1046 376 1112 392
rect 1046 342 1062 376
rect 1096 342 1112 376
rect 1046 308 1112 342
rect 1046 274 1062 308
rect 1096 274 1112 308
rect 1046 258 1112 274
rect 978 153 1044 169
rect 978 119 994 153
rect 1028 119 1044 153
rect 866 84 882 118
rect 916 85 932 118
rect 1078 85 1112 258
rect 1146 160 1180 459
rect 1214 467 1248 581
rect 1282 535 1397 649
rect 1282 501 1322 535
rect 1356 501 1397 535
rect 1431 581 1633 615
rect 1431 467 1465 581
rect 1214 433 1465 467
rect 1499 520 1565 547
rect 1499 486 1515 520
rect 1549 486 1565 520
rect 1499 459 1565 486
rect 1214 312 1261 433
rect 1499 399 1533 459
rect 1599 444 1633 581
rect 1667 531 1733 649
rect 1667 497 1683 531
rect 1717 497 1733 531
rect 1667 478 1733 497
rect 1785 580 1851 596
rect 1785 546 1801 580
rect 1835 546 1851 580
rect 1785 476 1851 546
rect 1885 562 1935 649
rect 1885 528 1901 562
rect 1885 494 1935 528
rect 1975 581 2221 615
rect 1975 580 2025 581
rect 1975 546 1991 580
rect 1599 410 1713 444
rect 1785 442 1801 476
rect 1835 460 1851 476
rect 1975 470 2025 546
rect 2155 580 2221 581
rect 2155 546 2171 580
rect 2205 546 2221 580
rect 1975 460 1991 470
rect 1835 442 1991 460
rect 1785 436 1991 442
rect 1785 426 2025 436
rect 1975 420 2025 426
rect 2065 509 2115 540
rect 2065 475 2081 509
rect 2155 510 2221 546
rect 2155 476 2171 510
rect 2205 476 2221 510
rect 2273 577 2548 611
rect 2273 527 2324 577
rect 2482 567 2548 577
rect 2273 493 2289 527
rect 2323 493 2324 527
rect 2273 477 2324 493
rect 2364 514 2444 543
rect 2364 480 2380 514
rect 2414 480 2444 514
rect 2482 533 2498 567
rect 2532 533 2548 567
rect 2482 504 2548 533
rect 2588 567 2622 649
rect 2588 504 2622 533
rect 2662 567 2728 596
rect 2662 533 2678 567
rect 2712 533 2728 567
rect 2065 442 2115 475
rect 2364 462 2444 480
rect 2662 462 2728 533
rect 2774 556 2863 582
rect 2774 522 2790 556
rect 2824 522 2863 556
rect 2774 496 2863 522
rect 2364 446 2795 462
rect 2364 442 2745 446
rect 2065 428 2745 442
rect 1327 390 1533 399
rect 1327 356 1343 390
rect 1377 356 1533 390
rect 1327 347 1533 356
rect 1567 360 1645 376
rect 1567 350 1595 360
rect 1629 326 1645 360
rect 1601 316 1645 326
rect 1214 278 1220 312
rect 1254 278 1261 312
rect 1214 244 1261 278
rect 1214 210 1220 244
rect 1254 210 1261 244
rect 1214 194 1261 210
rect 1295 292 1533 313
rect 1567 310 1645 316
rect 1295 279 1487 292
rect 1295 160 1329 279
rect 1471 258 1487 279
rect 1521 276 1533 292
rect 1679 303 1713 410
rect 2065 408 2478 428
rect 1747 376 1813 392
rect 1747 342 1763 376
rect 1797 374 1813 376
rect 1797 342 2410 374
rect 1747 340 2410 342
rect 1747 337 1813 340
rect 2076 303 2278 306
rect 1679 290 2278 303
rect 1521 258 1610 276
rect 1679 269 2092 290
rect 1363 237 1429 245
rect 1471 242 1610 258
rect 1363 203 1379 237
rect 1413 208 1429 237
rect 1576 235 1610 242
rect 2076 256 2092 269
rect 2126 256 2160 290
rect 2194 256 2228 290
rect 2262 256 2278 290
rect 2076 240 2278 256
rect 1576 230 1772 235
rect 1413 203 1542 208
rect 1363 174 1542 203
rect 1576 196 1722 230
rect 1756 196 1772 230
rect 1576 180 1772 196
rect 1806 201 2042 235
rect 2344 230 2410 340
rect 1806 190 1856 201
rect 1146 144 1329 160
rect 1146 110 1180 144
rect 1214 110 1329 144
rect 1146 94 1329 110
rect 1363 124 1430 140
rect 916 84 1112 85
rect 866 51 1112 84
rect 1397 90 1430 124
rect 1363 17 1430 90
rect 1476 133 1542 174
rect 1840 156 1856 190
rect 1992 190 2042 201
rect 1476 99 1492 133
rect 1526 99 1542 133
rect 1476 70 1542 99
rect 1640 120 1706 136
rect 1640 86 1656 120
rect 1690 86 1706 120
rect 1640 17 1706 86
rect 1806 120 1856 156
rect 1840 86 1856 120
rect 1806 70 1856 86
rect 1890 135 1956 167
rect 1890 101 1906 135
rect 1940 101 1956 135
rect 1890 17 1956 101
rect 2026 156 2042 190
rect 1992 120 2042 156
rect 2026 86 2042 120
rect 2076 179 2310 206
rect 2344 196 2360 230
rect 2394 196 2410 230
rect 2344 180 2410 196
rect 2076 145 2092 179
rect 2126 172 2310 179
rect 2126 145 2142 172
rect 2076 119 2142 145
rect 2276 146 2310 172
rect 2444 146 2478 408
rect 2729 412 2745 428
rect 2779 412 2795 446
rect 2513 376 2579 392
rect 2513 342 2529 376
rect 2563 342 2579 376
rect 2513 308 2579 342
rect 2513 274 2529 308
rect 2563 274 2579 308
rect 2513 226 2579 274
rect 2617 378 2687 394
rect 2617 350 2637 378
rect 2617 316 2623 350
rect 2671 344 2687 378
rect 2657 316 2687 344
rect 2617 310 2687 316
rect 2617 276 2637 310
rect 2671 276 2687 310
rect 2617 260 2687 276
rect 2729 378 2795 412
rect 2729 344 2745 378
rect 2779 344 2795 378
rect 2729 310 2795 344
rect 2729 276 2745 310
rect 2779 276 2795 310
rect 2729 260 2795 276
rect 2829 226 2863 496
rect 2897 580 2931 649
rect 2897 497 2931 546
rect 2897 414 2931 463
rect 2897 364 2931 380
rect 2970 580 3021 596
rect 2970 546 2987 580
rect 2970 497 3021 546
rect 2970 463 2987 497
rect 2970 414 3021 463
rect 2970 380 2987 414
rect 2513 192 2863 226
rect 2970 282 3021 380
rect 3061 580 3127 649
rect 3061 546 3077 580
rect 3111 546 3127 580
rect 3283 580 3333 649
rect 3061 497 3127 546
rect 3061 463 3077 497
rect 3111 463 3127 497
rect 3061 414 3127 463
rect 3061 380 3077 414
rect 3111 380 3127 414
rect 3061 364 3127 380
rect 3173 556 3239 572
rect 3173 522 3189 556
rect 3223 522 3239 556
rect 3173 485 3239 522
rect 3173 451 3189 485
rect 3223 451 3239 485
rect 3173 414 3239 451
rect 3173 380 3189 414
rect 3223 380 3239 414
rect 3173 326 3239 380
rect 3283 546 3299 580
rect 3283 497 3333 546
rect 3283 463 3299 497
rect 3283 414 3333 463
rect 3283 380 3299 414
rect 3283 364 3333 380
rect 3373 580 3445 596
rect 3373 546 3389 580
rect 3423 546 3445 580
rect 3373 497 3445 546
rect 3373 463 3389 497
rect 3423 463 3445 497
rect 3373 414 3445 463
rect 3373 380 3389 414
rect 3423 380 3445 414
rect 3373 364 3445 380
rect 3479 580 3529 649
rect 3513 546 3529 580
rect 3479 497 3529 546
rect 3513 463 3529 497
rect 3479 414 3529 463
rect 3513 380 3529 414
rect 3479 364 3529 380
rect 3173 310 3377 326
rect 2970 210 3047 282
rect 3173 276 3327 310
rect 3361 276 3377 310
rect 3173 260 3377 276
rect 2176 121 2242 138
rect 1992 85 2042 86
rect 2176 87 2192 121
rect 2226 87 2242 121
rect 2176 85 2242 87
rect 1992 51 2242 85
rect 2276 130 2478 146
rect 2276 96 2304 130
rect 2338 96 2426 130
rect 2460 96 2478 130
rect 2276 80 2478 96
rect 2652 131 2718 158
rect 2652 97 2668 131
rect 2702 97 2718 131
rect 2652 17 2718 97
rect 2754 133 2820 192
rect 2970 176 2986 210
rect 3020 176 3047 210
rect 2754 99 2770 133
rect 2804 99 2820 133
rect 2754 70 2820 99
rect 2870 142 2936 158
rect 2870 108 2886 142
rect 2920 108 2936 142
rect 2870 17 2936 108
rect 2970 120 3047 176
rect 2970 86 2986 120
rect 3020 86 3047 120
rect 2970 70 3047 86
rect 3081 210 3131 226
rect 3115 176 3131 210
rect 3081 120 3131 176
rect 3115 86 3131 120
rect 3173 210 3244 260
rect 3411 226 3445 364
rect 3173 176 3194 210
rect 3228 176 3244 210
rect 3173 140 3244 176
rect 3173 106 3194 140
rect 3228 106 3244 140
rect 3173 90 3244 106
rect 3291 210 3341 226
rect 3291 176 3307 210
rect 3291 120 3341 176
rect 3081 17 3131 86
rect 3291 86 3307 120
rect 3291 17 3341 86
rect 3377 210 3445 226
rect 3377 176 3393 210
rect 3427 176 3445 210
rect 3377 120 3445 176
rect 3377 86 3393 120
rect 3427 86 3445 120
rect 3377 70 3445 86
rect 3479 210 3529 226
rect 3513 176 3529 210
rect 3479 120 3529 176
rect 3513 86 3529 120
rect 3479 17 3529 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 1567 326 1595 350
rect 1595 326 1601 350
rect 1567 316 1601 326
rect 2623 344 2637 350
rect 2637 344 2657 350
rect 2623 316 2657 344
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
<< metal1 >>
rect 0 683 3552 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3552 683
rect 0 617 3552 649
rect 1555 350 1613 356
rect 1555 316 1567 350
rect 1601 347 1613 350
rect 2611 350 2669 356
rect 2611 347 2623 350
rect 1601 319 2623 347
rect 1601 316 1613 319
rect 1555 310 1613 316
rect 2611 316 2623 319
rect 2657 316 2669 350
rect 2611 310 2669 316
rect 0 17 3552 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
rect 0 -49 3552 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdfsbp_2
flabel comment s 1764 481 1764 481 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 1382 323 1382 323 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 1126 276 1126 276 0 FreeSans 200 0 0 0 no_jumper_check
flabel pwell s 0 0 3552 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 3552 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 2623 316 2657 350 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel metal1 s 0 617 3552 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 3552 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 3007 94 3041 128 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3007 168 3041 202 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3007 242 3041 276 0 FreeSans 340 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 3391 94 3425 128 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3391 168 3425 202 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3552 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 3602356
string GDS_START 3577448
<< end >>
