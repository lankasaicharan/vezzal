magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 19 49 627 157
rect 0 0 672 49
<< scnmos >>
rect 98 47 128 131
rect 200 47 230 131
rect 290 47 320 131
rect 404 47 434 131
rect 518 47 548 131
<< scpmoshvt >>
rect 146 479 176 607
rect 232 479 262 607
rect 318 479 348 607
rect 404 479 434 607
rect 490 479 520 607
<< ndiff >>
rect 45 106 98 131
rect 45 72 53 106
rect 87 72 98 106
rect 45 47 98 72
rect 128 106 200 131
rect 128 72 143 106
rect 177 72 200 106
rect 128 47 200 72
rect 230 47 290 131
rect 320 47 404 131
rect 434 47 518 131
rect 548 106 601 131
rect 548 72 559 106
rect 593 72 601 106
rect 548 47 601 72
<< pdiff >>
rect 93 595 146 607
rect 93 561 101 595
rect 135 561 146 595
rect 93 525 146 561
rect 93 491 101 525
rect 135 491 146 525
rect 93 479 146 491
rect 176 595 232 607
rect 176 561 187 595
rect 221 561 232 595
rect 176 525 232 561
rect 176 491 187 525
rect 221 491 232 525
rect 176 479 232 491
rect 262 595 318 607
rect 262 561 273 595
rect 307 561 318 595
rect 262 525 318 561
rect 262 491 273 525
rect 307 491 318 525
rect 262 479 318 491
rect 348 595 404 607
rect 348 561 359 595
rect 393 561 404 595
rect 348 525 404 561
rect 348 491 359 525
rect 393 491 404 525
rect 348 479 404 491
rect 434 595 490 607
rect 434 561 445 595
rect 479 561 490 595
rect 434 525 490 561
rect 434 491 445 525
rect 479 491 490 525
rect 434 479 490 491
rect 520 595 573 607
rect 520 561 531 595
rect 565 561 573 595
rect 520 525 573 561
rect 520 491 531 525
rect 565 491 573 525
rect 520 479 573 491
<< ndiffc >>
rect 53 72 87 106
rect 143 72 177 106
rect 559 72 593 106
<< pdiffc >>
rect 101 561 135 595
rect 101 491 135 525
rect 187 561 221 595
rect 187 491 221 525
rect 273 561 307 595
rect 273 491 307 525
rect 359 561 393 595
rect 359 491 393 525
rect 445 561 479 595
rect 445 491 479 525
rect 531 561 565 595
rect 531 491 565 525
<< poly >>
rect 146 607 176 633
rect 232 607 262 633
rect 318 607 348 633
rect 404 607 434 633
rect 490 607 520 633
rect 146 377 176 479
rect 232 377 262 479
rect 98 347 176 377
rect 218 347 262 377
rect 98 299 128 347
rect 218 299 248 347
rect 318 299 348 479
rect 404 299 434 479
rect 490 377 520 479
rect 490 347 548 377
rect 518 317 548 347
rect 518 301 584 317
rect 34 283 128 299
rect 34 249 50 283
rect 84 249 128 283
rect 34 215 128 249
rect 34 181 50 215
rect 84 181 128 215
rect 34 165 128 181
rect 176 283 248 299
rect 176 249 198 283
rect 232 249 248 283
rect 176 215 248 249
rect 176 181 198 215
rect 232 181 248 215
rect 176 165 248 181
rect 290 283 356 299
rect 290 249 306 283
rect 340 249 356 283
rect 290 215 356 249
rect 290 181 306 215
rect 340 181 356 215
rect 290 165 356 181
rect 404 283 470 299
rect 404 249 420 283
rect 454 249 470 283
rect 404 215 470 249
rect 404 181 420 215
rect 454 181 470 215
rect 404 165 470 181
rect 518 267 534 301
rect 568 267 584 301
rect 518 233 584 267
rect 518 199 534 233
rect 568 199 584 233
rect 518 183 584 199
rect 98 131 128 165
rect 200 131 230 165
rect 290 131 320 165
rect 404 131 434 165
rect 518 131 548 183
rect 98 21 128 47
rect 200 21 230 47
rect 290 21 320 47
rect 404 21 434 47
rect 518 21 548 47
<< polycont >>
rect 50 249 84 283
rect 50 181 84 215
rect 198 249 232 283
rect 198 181 232 215
rect 306 249 340 283
rect 306 181 340 215
rect 420 249 454 283
rect 420 181 454 215
rect 534 267 568 301
rect 534 199 568 233
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 85 595 144 611
rect 85 561 101 595
rect 135 561 144 595
rect 85 525 144 561
rect 85 491 101 525
rect 135 491 144 525
rect 85 371 144 491
rect 178 595 230 611
rect 178 561 187 595
rect 221 561 230 595
rect 178 525 230 561
rect 178 491 187 525
rect 221 491 230 525
rect 178 441 230 491
rect 264 595 315 649
rect 264 561 273 595
rect 307 561 315 595
rect 264 525 315 561
rect 264 491 273 525
rect 307 491 315 525
rect 264 475 315 491
rect 349 595 401 611
rect 349 561 359 595
rect 393 561 401 595
rect 349 525 401 561
rect 349 491 359 525
rect 393 491 401 525
rect 349 441 401 491
rect 435 595 489 649
rect 435 561 445 595
rect 479 561 489 595
rect 435 525 489 561
rect 435 491 445 525
rect 479 491 489 525
rect 435 475 489 491
rect 523 595 581 611
rect 523 561 531 595
rect 565 561 581 595
rect 523 525 581 561
rect 523 491 531 525
rect 565 491 581 525
rect 523 441 581 491
rect 178 405 581 441
rect 85 337 164 371
rect 17 283 90 299
rect 17 249 50 283
rect 84 249 90 283
rect 17 215 90 249
rect 17 181 50 215
rect 84 181 90 215
rect 17 165 90 181
rect 124 131 164 337
rect 198 283 272 368
rect 232 249 272 283
rect 198 215 272 249
rect 232 181 272 215
rect 198 165 272 181
rect 306 283 371 368
rect 340 249 371 283
rect 306 215 371 249
rect 340 181 371 215
rect 306 165 371 181
rect 405 283 471 368
rect 405 249 420 283
rect 454 249 471 283
rect 405 215 471 249
rect 405 181 420 215
rect 454 181 471 215
rect 505 301 655 368
rect 505 267 534 301
rect 568 267 655 301
rect 505 233 655 267
rect 505 199 534 233
rect 568 199 655 233
rect 405 165 471 181
rect 49 106 90 122
rect 49 72 53 106
rect 87 72 90 106
rect 49 17 90 72
rect 124 106 483 131
rect 124 72 143 106
rect 177 72 483 106
rect 124 56 483 72
rect 543 106 609 122
rect 543 72 559 106
rect 593 72 609 106
rect 543 17 609 72
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a41oi_0
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1392164
string GDS_START 1384508
<< end >>
