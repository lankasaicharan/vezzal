magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 36 49 856 248
rect 0 0 864 49
<< scnmos >>
rect 115 94 145 222
rect 213 74 243 222
rect 299 74 329 222
rect 489 74 519 222
rect 575 74 605 222
rect 661 74 691 222
rect 747 74 777 222
<< scpmoshvt >>
rect 102 392 132 592
rect 296 368 326 592
rect 386 368 416 592
rect 476 368 506 592
rect 566 368 596 592
rect 656 368 686 592
rect 750 368 780 592
<< ndiff >>
rect 62 210 115 222
rect 62 176 70 210
rect 104 176 115 210
rect 62 140 115 176
rect 62 106 70 140
rect 104 106 115 140
rect 62 94 115 106
rect 145 188 213 222
rect 145 154 168 188
rect 202 154 213 188
rect 145 120 213 154
rect 145 94 168 120
rect 160 86 168 94
rect 202 86 213 120
rect 160 74 213 86
rect 243 210 299 222
rect 243 176 254 210
rect 288 176 299 210
rect 243 120 299 176
rect 243 86 254 120
rect 288 86 299 120
rect 243 74 299 86
rect 329 146 382 222
rect 329 112 340 146
rect 374 112 382 146
rect 329 74 382 112
rect 436 120 489 222
rect 436 86 444 120
rect 478 86 489 120
rect 436 74 489 86
rect 519 199 575 222
rect 519 165 530 199
rect 564 165 575 199
rect 519 74 575 165
rect 605 194 661 222
rect 605 160 616 194
rect 650 160 661 194
rect 605 120 661 160
rect 605 86 616 120
rect 650 86 661 120
rect 605 74 661 86
rect 691 127 747 222
rect 691 93 702 127
rect 736 93 747 127
rect 691 74 747 93
rect 777 210 830 222
rect 777 176 788 210
rect 822 176 830 210
rect 777 120 830 176
rect 777 86 788 120
rect 822 86 830 120
rect 777 74 830 86
<< pdiff >>
rect 47 580 102 592
rect 47 546 55 580
rect 89 546 102 580
rect 47 510 102 546
rect 47 476 55 510
rect 89 476 102 510
rect 47 440 102 476
rect 47 406 55 440
rect 89 406 102 440
rect 47 392 102 406
rect 132 580 187 592
rect 132 546 145 580
rect 179 546 187 580
rect 132 509 187 546
rect 132 475 145 509
rect 179 475 187 509
rect 132 438 187 475
rect 132 404 145 438
rect 179 404 187 438
rect 132 392 187 404
rect 241 580 296 592
rect 241 546 249 580
rect 283 546 296 580
rect 241 497 296 546
rect 241 463 249 497
rect 283 463 296 497
rect 241 414 296 463
rect 241 380 249 414
rect 283 380 296 414
rect 241 368 296 380
rect 326 547 386 592
rect 326 513 339 547
rect 373 513 386 547
rect 326 479 386 513
rect 326 445 339 479
rect 373 445 386 479
rect 326 410 386 445
rect 326 376 339 410
rect 373 376 386 410
rect 326 368 386 376
rect 416 580 476 592
rect 416 546 429 580
rect 463 546 476 580
rect 416 497 476 546
rect 416 463 429 497
rect 463 463 476 497
rect 416 414 476 463
rect 416 380 429 414
rect 463 380 476 414
rect 416 368 476 380
rect 506 580 566 592
rect 506 546 519 580
rect 553 546 566 580
rect 506 492 566 546
rect 506 458 519 492
rect 553 458 566 492
rect 506 368 566 458
rect 596 580 656 592
rect 596 546 609 580
rect 643 546 656 580
rect 596 497 656 546
rect 596 463 609 497
rect 643 463 656 497
rect 596 414 656 463
rect 596 380 609 414
rect 643 380 656 414
rect 596 368 656 380
rect 686 582 750 592
rect 686 548 701 582
rect 735 548 750 582
rect 686 514 750 548
rect 686 480 701 514
rect 735 480 750 514
rect 686 446 750 480
rect 686 412 701 446
rect 735 412 750 446
rect 686 368 750 412
rect 780 580 835 592
rect 780 546 793 580
rect 827 546 835 580
rect 780 497 835 546
rect 780 463 793 497
rect 827 463 835 497
rect 780 414 835 463
rect 780 380 793 414
rect 827 380 835 414
rect 780 368 835 380
<< ndiffc >>
rect 70 176 104 210
rect 70 106 104 140
rect 168 154 202 188
rect 168 86 202 120
rect 254 176 288 210
rect 254 86 288 120
rect 340 112 374 146
rect 444 86 478 120
rect 530 165 564 199
rect 616 160 650 194
rect 616 86 650 120
rect 702 93 736 127
rect 788 176 822 210
rect 788 86 822 120
<< pdiffc >>
rect 55 546 89 580
rect 55 476 89 510
rect 55 406 89 440
rect 145 546 179 580
rect 145 475 179 509
rect 145 404 179 438
rect 249 546 283 580
rect 249 463 283 497
rect 249 380 283 414
rect 339 513 373 547
rect 339 445 373 479
rect 339 376 373 410
rect 429 546 463 580
rect 429 463 463 497
rect 429 380 463 414
rect 519 546 553 580
rect 519 458 553 492
rect 609 546 643 580
rect 609 463 643 497
rect 609 380 643 414
rect 701 548 735 582
rect 701 480 735 514
rect 701 412 735 446
rect 793 546 827 580
rect 793 463 827 497
rect 793 380 827 414
<< poly >>
rect 102 592 132 618
rect 296 592 326 618
rect 386 592 416 618
rect 476 592 506 618
rect 566 592 596 618
rect 656 592 686 618
rect 750 592 780 618
rect 102 377 132 392
rect 99 356 135 377
rect 29 340 145 356
rect 296 353 326 368
rect 386 353 416 368
rect 476 353 506 368
rect 566 353 596 368
rect 656 353 686 368
rect 750 353 780 368
rect 29 306 45 340
rect 79 306 145 340
rect 293 330 419 353
rect 29 290 145 306
rect 115 222 145 290
rect 213 323 419 330
rect 473 330 509 353
rect 563 330 599 353
rect 213 314 329 323
rect 213 280 229 314
rect 263 280 329 314
rect 213 264 329 280
rect 473 314 599 330
rect 473 280 513 314
rect 547 294 599 314
rect 653 310 689 353
rect 747 310 783 353
rect 653 294 783 310
rect 547 280 605 294
rect 473 264 605 280
rect 213 222 243 264
rect 299 222 329 264
rect 489 222 519 264
rect 575 222 605 264
rect 653 260 669 294
rect 703 260 783 294
rect 653 244 783 260
rect 661 222 691 244
rect 747 222 777 244
rect 115 68 145 94
rect 213 48 243 74
rect 299 48 329 74
rect 489 48 519 74
rect 575 48 605 74
rect 661 48 691 74
rect 747 48 777 74
<< polycont >>
rect 45 306 79 340
rect 229 280 263 314
rect 513 280 547 314
rect 669 260 703 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 39 580 89 649
rect 39 546 55 580
rect 39 510 89 546
rect 39 476 55 510
rect 39 440 89 476
rect 39 406 55 440
rect 39 390 89 406
rect 129 580 195 596
rect 129 546 145 580
rect 179 546 195 580
rect 129 509 195 546
rect 129 475 145 509
rect 179 475 195 509
rect 129 438 195 475
rect 129 404 145 438
rect 179 404 195 438
rect 129 388 195 404
rect 25 340 95 356
rect 25 306 45 340
rect 79 306 95 340
rect 25 290 95 306
rect 161 330 195 388
rect 233 581 463 615
rect 233 580 283 581
rect 233 546 249 580
rect 423 580 463 581
rect 233 497 283 546
rect 233 463 249 497
rect 233 414 283 463
rect 233 380 249 414
rect 233 364 283 380
rect 323 513 339 547
rect 373 513 389 547
rect 323 479 389 513
rect 323 445 339 479
rect 373 445 389 479
rect 323 410 389 445
rect 323 376 339 410
rect 373 376 389 410
rect 161 314 279 330
rect 161 280 229 314
rect 263 280 279 314
rect 161 264 279 280
rect 323 282 389 376
rect 423 546 429 580
rect 423 497 463 546
rect 423 463 429 497
rect 423 424 463 463
rect 503 580 569 649
rect 503 546 519 580
rect 553 546 569 580
rect 503 492 569 546
rect 503 458 519 492
rect 553 458 569 492
rect 609 580 643 596
rect 609 497 643 546
rect 609 424 643 463
rect 423 414 643 424
rect 423 380 429 414
rect 463 390 609 414
rect 423 364 463 380
rect 683 582 753 649
rect 683 548 701 582
rect 735 548 753 582
rect 683 514 753 548
rect 683 480 701 514
rect 735 480 753 514
rect 683 446 753 480
rect 683 412 701 446
rect 735 412 753 446
rect 793 580 843 596
rect 827 546 843 580
rect 793 497 843 546
rect 827 463 843 497
rect 793 414 843 463
rect 609 378 643 380
rect 827 380 843 414
rect 793 378 843 380
rect 497 314 563 356
rect 609 344 843 378
rect 161 256 195 264
rect 54 222 195 256
rect 323 230 455 282
rect 497 280 513 314
rect 547 280 563 314
rect 497 264 563 280
rect 653 294 743 310
rect 653 260 669 294
rect 703 260 743 294
rect 653 244 743 260
rect 697 236 743 244
rect 54 210 104 222
rect 54 176 70 210
rect 254 210 580 230
rect 788 210 838 226
rect 54 140 104 176
rect 54 106 70 140
rect 54 90 104 106
rect 152 154 168 188
rect 202 154 218 188
rect 152 120 218 154
rect 152 86 168 120
rect 202 86 218 120
rect 152 17 218 86
rect 288 199 580 210
rect 288 196 530 199
rect 254 120 288 176
rect 514 165 530 196
rect 564 165 580 199
rect 254 70 288 86
rect 324 146 390 162
rect 514 154 580 165
rect 616 202 650 210
rect 616 194 788 202
rect 650 176 788 194
rect 822 176 838 210
rect 650 168 838 176
rect 324 112 340 146
rect 374 112 390 146
rect 616 120 650 160
rect 324 17 390 112
rect 428 86 444 120
rect 478 86 616 120
rect 428 70 650 86
rect 686 127 752 134
rect 686 93 702 127
rect 736 93 752 127
rect 686 17 752 93
rect 788 120 838 168
rect 822 86 838 120
rect 788 70 838 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a21boi_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 3558870
string GDS_START 3550878
<< end >>
