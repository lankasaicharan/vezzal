magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 331 998 704
<< pwell >>
rect 665 157 939 241
rect 41 49 939 157
rect 0 0 960 49
<< scnmos >>
rect 120 47 150 131
rect 214 47 244 131
rect 300 47 330 131
rect 555 47 585 131
rect 627 47 657 131
rect 744 47 774 215
rect 830 47 860 215
<< scpmoshvt >>
rect 120 367 150 495
rect 192 367 222 495
rect 300 367 330 495
rect 496 367 526 495
rect 582 367 612 495
rect 744 367 774 619
rect 830 367 860 619
<< ndiff >>
rect 691 187 744 215
rect 691 153 699 187
rect 733 153 744 187
rect 691 131 744 153
rect 67 106 120 131
rect 67 72 75 106
rect 109 72 120 106
rect 67 47 120 72
rect 150 93 214 131
rect 150 59 165 93
rect 199 59 214 93
rect 150 47 214 59
rect 244 106 300 131
rect 244 72 255 106
rect 289 72 300 106
rect 244 47 300 72
rect 330 106 383 131
rect 330 72 341 106
rect 375 72 383 106
rect 330 47 383 72
rect 502 106 555 131
rect 502 72 510 106
rect 544 72 555 106
rect 502 47 555 72
rect 585 47 627 131
rect 657 93 744 131
rect 657 59 685 93
rect 719 59 744 93
rect 657 47 744 59
rect 774 203 830 215
rect 774 169 785 203
rect 819 169 830 203
rect 774 101 830 169
rect 774 67 785 101
rect 819 67 830 101
rect 774 47 830 67
rect 860 203 913 215
rect 860 169 871 203
rect 905 169 913 203
rect 860 93 913 169
rect 860 59 871 93
rect 905 59 913 93
rect 860 47 913 59
<< pdiff >>
rect 691 607 744 619
rect 691 573 699 607
rect 733 573 744 607
rect 691 524 744 573
rect 691 495 699 524
rect 67 483 120 495
rect 67 449 75 483
rect 109 449 120 483
rect 67 413 120 449
rect 67 379 75 413
rect 109 379 120 413
rect 67 367 120 379
rect 150 367 192 495
rect 222 487 300 495
rect 222 453 244 487
rect 278 453 300 487
rect 222 413 300 453
rect 222 379 244 413
rect 278 379 300 413
rect 222 367 300 379
rect 330 461 496 495
rect 330 427 381 461
rect 415 427 496 461
rect 330 367 496 427
rect 526 481 582 495
rect 526 447 537 481
rect 571 447 582 481
rect 526 413 582 447
rect 526 379 537 413
rect 571 379 582 413
rect 526 367 582 379
rect 612 490 699 495
rect 733 490 744 524
rect 612 439 744 490
rect 612 405 691 439
rect 725 405 744 439
rect 612 367 744 405
rect 774 599 830 619
rect 774 565 785 599
rect 819 565 830 599
rect 774 502 830 565
rect 774 468 785 502
rect 819 468 830 502
rect 774 413 830 468
rect 774 379 785 413
rect 819 379 830 413
rect 774 367 830 379
rect 860 607 913 619
rect 860 573 871 607
rect 905 573 913 607
rect 860 509 913 573
rect 860 475 871 509
rect 905 475 913 509
rect 860 413 913 475
rect 860 379 871 413
rect 905 379 913 413
rect 860 367 913 379
<< ndiffc >>
rect 699 153 733 187
rect 75 72 109 106
rect 165 59 199 93
rect 255 72 289 106
rect 341 72 375 106
rect 510 72 544 106
rect 685 59 719 93
rect 785 169 819 203
rect 785 67 819 101
rect 871 169 905 203
rect 871 59 905 93
<< pdiffc >>
rect 699 573 733 607
rect 75 449 109 483
rect 75 379 109 413
rect 244 453 278 487
rect 244 379 278 413
rect 381 427 415 461
rect 537 447 571 481
rect 537 379 571 413
rect 699 490 733 524
rect 691 405 725 439
rect 785 565 819 599
rect 785 468 819 502
rect 785 379 819 413
rect 871 573 905 607
rect 871 475 905 509
rect 871 379 905 413
<< poly >>
rect 744 619 774 645
rect 830 619 860 645
rect 120 495 150 521
rect 192 495 222 521
rect 300 495 330 521
rect 496 495 526 521
rect 582 495 612 521
rect 120 333 150 367
rect 84 317 150 333
rect 84 283 100 317
rect 134 283 150 317
rect 84 249 150 283
rect 84 215 100 249
rect 134 215 150 249
rect 84 199 150 215
rect 192 333 222 367
rect 300 333 330 367
rect 192 317 258 333
rect 192 283 208 317
rect 242 283 258 317
rect 192 249 258 283
rect 192 215 208 249
rect 242 215 258 249
rect 192 199 258 215
rect 300 317 429 333
rect 300 283 379 317
rect 413 283 429 317
rect 300 267 429 283
rect 120 131 150 199
rect 214 131 244 199
rect 300 131 330 267
rect 496 219 526 367
rect 582 303 612 367
rect 744 303 774 367
rect 830 303 860 367
rect 582 287 657 303
rect 582 253 607 287
rect 641 253 657 287
rect 582 237 657 253
rect 699 287 860 303
rect 699 253 715 287
rect 749 253 860 287
rect 699 237 860 253
rect 408 203 526 219
rect 408 169 424 203
rect 458 183 526 203
rect 458 169 585 183
rect 408 153 585 169
rect 555 131 585 153
rect 627 131 657 237
rect 744 215 774 237
rect 830 215 860 237
rect 120 21 150 47
rect 214 21 244 47
rect 300 21 330 47
rect 555 21 585 47
rect 627 21 657 47
rect 744 21 774 47
rect 830 21 860 47
<< polycont >>
rect 100 283 134 317
rect 100 215 134 249
rect 208 283 242 317
rect 208 215 242 249
rect 379 283 413 317
rect 607 253 641 287
rect 715 253 749 287
rect 424 169 458 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 59 483 125 649
rect 59 449 75 483
rect 109 449 125 483
rect 59 413 125 449
rect 59 379 75 413
rect 109 379 125 413
rect 59 367 125 379
rect 228 487 331 503
rect 228 453 244 487
rect 278 453 331 487
rect 228 413 331 453
rect 365 461 431 649
rect 675 607 749 649
rect 675 573 699 607
rect 733 573 749 607
rect 365 427 381 461
rect 415 427 431 461
rect 365 419 431 427
rect 465 533 641 567
rect 228 379 244 413
rect 278 385 331 413
rect 465 385 499 533
rect 278 379 499 385
rect 228 367 499 379
rect 293 351 499 367
rect 533 481 571 497
rect 533 447 537 481
rect 533 413 571 447
rect 533 379 537 413
rect 84 317 168 333
rect 84 283 100 317
rect 134 283 168 317
rect 84 249 168 283
rect 84 215 100 249
rect 134 215 168 249
rect 84 199 168 215
rect 202 317 259 333
rect 202 283 208 317
rect 242 283 259 317
rect 202 249 259 283
rect 202 215 208 249
rect 242 215 259 249
rect 202 199 259 215
rect 293 233 329 351
rect 533 317 571 379
rect 607 371 641 533
rect 675 524 749 573
rect 675 490 699 524
rect 733 490 749 524
rect 675 439 749 490
rect 675 405 691 439
rect 725 405 749 439
rect 783 599 837 615
rect 783 565 785 599
rect 819 565 837 599
rect 783 502 837 565
rect 783 468 785 502
rect 819 468 837 502
rect 783 413 837 468
rect 783 379 785 413
rect 819 379 837 413
rect 607 337 749 371
rect 363 283 379 317
rect 413 283 571 317
rect 363 267 571 283
rect 293 199 379 233
rect 59 131 298 165
rect 59 106 115 131
rect 59 72 75 106
rect 109 72 115 106
rect 249 106 298 131
rect 59 56 115 72
rect 149 93 215 97
rect 149 59 165 93
rect 199 59 215 93
rect 149 17 215 59
rect 249 72 255 106
rect 289 72 298 106
rect 249 56 298 72
rect 332 106 379 199
rect 332 72 341 106
rect 375 72 379 106
rect 332 56 379 72
rect 413 203 460 219
rect 413 169 424 203
rect 458 169 460 203
rect 413 69 460 169
rect 494 106 571 267
rect 494 72 510 106
rect 544 72 571 106
rect 605 287 647 303
rect 605 253 607 287
rect 641 253 647 287
rect 605 94 647 253
rect 699 287 749 337
rect 699 253 715 287
rect 699 237 749 253
rect 783 203 837 379
rect 871 607 921 649
rect 905 573 921 607
rect 871 509 921 573
rect 905 475 921 509
rect 871 413 921 475
rect 905 379 921 413
rect 871 363 921 379
rect 681 187 749 203
rect 681 153 699 187
rect 733 153 749 187
rect 494 56 571 72
rect 681 93 749 153
rect 681 59 685 93
rect 719 59 749 93
rect 681 17 749 59
rect 783 169 785 203
rect 819 169 837 203
rect 783 101 837 169
rect 783 67 785 101
rect 819 67 837 101
rect 783 51 837 67
rect 871 203 921 219
rect 905 169 921 203
rect 871 93 921 169
rect 905 59 921 93
rect 871 17 921 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o2bb2a_2
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 799 94 833 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 799 538 833 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3658750
string GDS_START 3650114
<< end >>
