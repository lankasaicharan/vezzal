magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 48 49 764 157
rect 0 0 768 49
<< scnmos >>
rect 226 47 256 131
rect 304 47 334 131
rect 392 47 422 131
rect 490 47 520 131
rect 579 47 609 131
rect 651 47 681 131
<< scpmoshvt >>
rect 98 419 148 619
rect 196 419 246 619
rect 360 419 410 619
rect 496 419 546 619
rect 610 419 660 619
<< ndiff >>
rect 74 93 226 131
rect 74 59 86 93
rect 120 59 226 93
rect 74 47 226 59
rect 256 47 304 131
rect 334 105 392 131
rect 334 71 346 105
rect 380 71 392 105
rect 334 47 392 71
rect 422 47 490 131
rect 520 100 579 131
rect 520 66 532 100
rect 566 66 579 100
rect 520 47 579 66
rect 609 47 651 131
rect 681 111 738 131
rect 681 77 692 111
rect 726 77 738 111
rect 681 47 738 77
<< pdiff >>
rect 39 607 98 619
rect 39 573 51 607
rect 85 573 98 607
rect 39 505 98 573
rect 39 471 51 505
rect 85 471 98 505
rect 39 419 98 471
rect 148 419 196 619
rect 246 597 360 619
rect 246 563 315 597
rect 349 563 360 597
rect 246 516 360 563
rect 246 482 315 516
rect 349 482 360 516
rect 246 419 360 482
rect 410 419 496 619
rect 546 607 610 619
rect 546 573 557 607
rect 591 573 610 607
rect 546 536 610 573
rect 546 502 557 536
rect 591 502 610 536
rect 546 465 610 502
rect 546 431 557 465
rect 591 431 610 465
rect 546 419 610 431
rect 660 597 717 619
rect 660 563 671 597
rect 705 563 717 597
rect 660 465 717 563
rect 660 431 671 465
rect 705 431 717 465
rect 660 419 717 431
<< ndiffc >>
rect 86 59 120 93
rect 346 71 380 105
rect 532 66 566 100
rect 692 77 726 111
<< pdiffc >>
rect 51 573 85 607
rect 51 471 85 505
rect 315 563 349 597
rect 315 482 349 516
rect 557 573 591 607
rect 557 502 591 536
rect 557 431 591 465
rect 671 563 705 597
rect 671 431 705 465
<< poly >>
rect 98 619 148 645
rect 196 619 246 645
rect 360 619 410 645
rect 496 619 546 645
rect 610 619 660 645
rect 98 349 148 419
rect 196 359 246 419
rect 360 387 410 419
rect 360 371 448 387
rect 88 333 154 349
rect 88 299 104 333
rect 138 299 154 333
rect 88 265 154 299
rect 196 343 262 359
rect 360 351 398 371
rect 196 309 212 343
rect 246 309 262 343
rect 196 293 262 309
rect 304 337 398 351
rect 432 337 448 371
rect 304 321 448 337
rect 496 333 546 419
rect 88 231 104 265
rect 138 245 154 265
rect 138 231 256 245
rect 88 215 256 231
rect 226 131 256 215
rect 304 131 334 321
rect 496 317 562 333
rect 496 283 512 317
rect 546 283 562 317
rect 382 263 448 279
rect 382 229 398 263
rect 432 229 448 263
rect 382 213 448 229
rect 496 267 562 283
rect 392 131 422 213
rect 496 176 526 267
rect 610 231 660 419
rect 610 219 640 231
rect 490 146 526 176
rect 574 203 640 219
rect 574 169 590 203
rect 624 183 640 203
rect 624 169 681 183
rect 574 153 681 169
rect 490 131 520 146
rect 579 131 609 153
rect 651 131 681 153
rect 226 21 256 47
rect 304 21 334 47
rect 392 21 422 47
rect 490 21 520 47
rect 579 21 609 47
rect 651 21 681 47
<< polycont >>
rect 104 299 138 333
rect 212 309 246 343
rect 398 337 432 371
rect 104 231 138 265
rect 512 283 546 317
rect 398 229 432 263
rect 590 169 624 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 35 607 85 649
rect 35 573 51 607
rect 35 505 85 573
rect 35 471 51 505
rect 35 455 85 471
rect 121 597 365 613
rect 121 579 315 597
rect 121 419 263 579
rect 299 563 315 579
rect 349 563 365 597
rect 299 516 365 563
rect 299 482 315 516
rect 349 482 365 516
rect 299 466 365 482
rect 541 607 607 649
rect 541 573 557 607
rect 591 573 607 607
rect 541 536 607 573
rect 541 502 557 536
rect 591 502 607 536
rect 541 465 607 502
rect 541 431 557 465
rect 591 431 607 465
rect 18 385 155 419
rect 18 179 52 385
rect 382 371 455 430
rect 541 415 607 431
rect 655 597 742 613
rect 655 563 671 597
rect 705 563 742 597
rect 655 465 742 563
rect 655 431 671 465
rect 705 431 742 465
rect 88 333 154 349
rect 88 299 104 333
rect 138 299 154 333
rect 88 265 154 299
rect 196 343 346 359
rect 196 309 212 343
rect 246 309 346 343
rect 382 337 398 371
rect 432 337 455 371
rect 382 321 455 337
rect 655 333 742 431
rect 196 293 346 309
rect 88 231 104 265
rect 138 249 154 265
rect 312 279 346 293
rect 496 317 742 333
rect 496 283 512 317
rect 546 283 742 317
rect 312 263 448 279
rect 496 267 742 283
rect 138 231 276 249
rect 88 215 276 231
rect 18 145 206 179
rect 70 93 136 109
rect 70 59 86 93
rect 120 59 136 93
rect 70 17 136 59
rect 172 107 206 145
rect 242 177 276 215
rect 312 229 398 263
rect 432 229 448 263
rect 312 213 448 229
rect 505 203 640 219
rect 505 177 590 203
rect 242 169 590 177
rect 624 169 640 203
rect 242 143 640 169
rect 676 111 742 267
rect 172 105 396 107
rect 172 71 346 105
rect 380 71 396 105
rect 172 53 396 71
rect 516 100 582 107
rect 516 66 532 100
rect 566 66 582 100
rect 516 17 582 66
rect 676 77 692 111
rect 726 77 742 111
rect 676 53 742 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2i_lp2
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 223 538 257 572 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3875840
string GDS_START 3869518
<< end >>
