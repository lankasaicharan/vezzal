magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 66 49 718 248
rect 0 0 768 49
<< scpmos >>
rect 88 368 118 592
rect 318 368 348 592
rect 408 368 438 592
rect 504 368 534 592
rect 612 368 642 592
<< nmoslvt >>
rect 213 74 243 222
rect 321 74 351 222
rect 393 74 423 222
rect 537 74 567 222
rect 609 74 639 222
<< ndiff >>
rect 92 210 213 222
rect 92 176 100 210
rect 134 176 168 210
rect 202 176 213 210
rect 92 120 213 176
rect 92 86 100 120
rect 134 86 168 120
rect 202 86 213 120
rect 92 74 213 86
rect 243 152 321 222
rect 243 118 272 152
rect 306 118 321 152
rect 243 74 321 118
rect 351 74 393 222
rect 423 214 537 222
rect 423 180 458 214
rect 492 180 537 214
rect 423 116 537 180
rect 423 82 458 116
rect 492 82 537 116
rect 423 74 537 82
rect 567 74 609 222
rect 639 197 692 222
rect 639 163 650 197
rect 684 163 692 197
rect 639 120 692 163
rect 639 86 650 120
rect 684 86 692 120
rect 639 74 692 86
<< pdiff >>
rect 33 580 88 592
rect 33 546 41 580
rect 75 546 88 580
rect 33 497 88 546
rect 33 463 41 497
rect 75 463 88 497
rect 33 414 88 463
rect 33 380 41 414
rect 75 380 88 414
rect 33 368 88 380
rect 118 580 173 592
rect 118 546 131 580
rect 165 546 173 580
rect 118 510 173 546
rect 118 476 131 510
rect 165 476 173 510
rect 118 440 173 476
rect 118 406 131 440
rect 165 406 173 440
rect 118 368 173 406
rect 263 531 318 592
rect 263 497 271 531
rect 305 497 318 531
rect 263 424 318 497
rect 263 390 271 424
rect 305 390 318 424
rect 263 368 318 390
rect 348 584 408 592
rect 348 550 361 584
rect 395 550 408 584
rect 348 497 408 550
rect 348 463 361 497
rect 395 463 408 497
rect 348 368 408 463
rect 438 580 504 592
rect 438 546 451 580
rect 485 546 504 580
rect 438 505 504 546
rect 438 471 451 505
rect 485 471 504 505
rect 438 424 504 471
rect 438 390 451 424
rect 485 390 504 424
rect 438 368 504 390
rect 534 584 612 592
rect 534 550 553 584
rect 587 550 612 584
rect 534 497 612 550
rect 534 463 553 497
rect 587 463 612 497
rect 534 368 612 463
rect 642 580 697 592
rect 642 546 655 580
rect 689 546 697 580
rect 642 497 697 546
rect 642 463 655 497
rect 689 463 697 497
rect 642 414 697 463
rect 642 380 655 414
rect 689 380 697 414
rect 642 368 697 380
<< ndiffc >>
rect 100 176 134 210
rect 168 176 202 210
rect 100 86 134 120
rect 168 86 202 120
rect 272 118 306 152
rect 458 180 492 214
rect 458 82 492 116
rect 650 163 684 197
rect 650 86 684 120
<< pdiffc >>
rect 41 546 75 580
rect 41 463 75 497
rect 41 380 75 414
rect 131 546 165 580
rect 131 476 165 510
rect 131 406 165 440
rect 271 497 305 531
rect 271 390 305 424
rect 361 550 395 584
rect 361 463 395 497
rect 451 546 485 580
rect 451 471 485 505
rect 451 390 485 424
rect 553 550 587 584
rect 553 463 587 497
rect 655 546 689 580
rect 655 463 689 497
rect 655 380 689 414
<< poly >>
rect 88 592 118 618
rect 318 592 348 618
rect 408 592 438 618
rect 504 592 534 618
rect 612 592 642 618
rect 88 353 118 368
rect 318 353 348 368
rect 408 353 438 368
rect 504 353 534 368
rect 612 353 642 368
rect 85 336 121 353
rect 315 336 351 353
rect 405 336 441 353
rect 501 336 537 353
rect 85 332 175 336
rect 85 320 243 332
rect 85 286 125 320
rect 159 286 243 320
rect 85 270 243 286
rect 285 320 351 336
rect 285 286 301 320
rect 335 286 351 320
rect 285 270 351 286
rect 213 222 243 270
rect 321 222 351 270
rect 393 320 459 336
rect 393 286 409 320
rect 443 286 459 320
rect 393 270 459 286
rect 501 320 567 336
rect 501 286 517 320
rect 551 286 567 320
rect 501 270 567 286
rect 393 222 423 270
rect 537 222 567 270
rect 609 310 645 353
rect 609 294 675 310
rect 609 260 625 294
rect 659 260 675 294
rect 609 244 675 260
rect 609 222 639 244
rect 213 48 243 74
rect 321 48 351 74
rect 393 48 423 74
rect 537 48 567 74
rect 609 48 639 74
<< polycont >>
rect 125 286 159 320
rect 301 286 335 320
rect 409 286 443 320
rect 517 286 551 320
rect 625 260 659 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 25 580 75 596
rect 25 546 41 580
rect 25 497 75 546
rect 25 463 41 497
rect 25 414 75 463
rect 25 380 41 414
rect 115 584 411 615
rect 115 581 361 584
rect 115 580 181 581
rect 115 546 131 580
rect 165 546 181 580
rect 345 550 361 581
rect 395 550 411 584
rect 115 510 181 546
rect 115 476 131 510
rect 165 476 181 510
rect 115 440 181 476
rect 115 406 131 440
rect 165 406 181 440
rect 115 390 181 406
rect 255 531 309 547
rect 255 497 271 531
rect 305 497 309 531
rect 255 424 309 497
rect 345 497 411 550
rect 345 463 361 497
rect 395 463 411 497
rect 345 458 411 463
rect 451 580 501 596
rect 485 546 501 580
rect 451 505 501 546
rect 485 471 501 505
rect 451 424 501 471
rect 535 584 605 649
rect 535 550 553 584
rect 587 550 605 584
rect 535 497 605 550
rect 535 463 553 497
rect 587 463 605 497
rect 535 458 605 463
rect 639 580 705 596
rect 639 546 655 580
rect 689 546 705 580
rect 639 497 705 546
rect 639 463 655 497
rect 689 463 705 497
rect 639 424 705 463
rect 255 390 271 424
rect 305 390 451 424
rect 485 414 705 424
rect 485 390 655 414
rect 25 236 75 380
rect 639 380 655 390
rect 689 380 705 414
rect 639 364 705 380
rect 109 320 175 356
rect 109 286 125 320
rect 159 286 175 320
rect 109 270 175 286
rect 217 320 359 356
rect 217 286 301 320
rect 335 286 359 320
rect 217 270 359 286
rect 393 320 459 356
rect 393 286 409 320
rect 443 286 459 320
rect 393 270 459 286
rect 501 320 567 356
rect 501 286 517 320
rect 551 286 567 320
rect 501 270 567 286
rect 601 294 743 310
rect 601 260 625 294
rect 659 260 743 294
rect 601 236 743 260
rect 25 214 515 236
rect 25 210 458 214
rect 25 176 100 210
rect 134 176 168 210
rect 202 202 458 210
rect 202 176 218 202
rect 25 120 218 176
rect 432 180 458 202
rect 492 180 515 214
rect 25 86 100 120
rect 134 86 168 120
rect 202 86 218 120
rect 25 70 218 86
rect 252 152 326 165
rect 252 118 272 152
rect 306 118 326 152
rect 252 17 326 118
rect 432 116 515 180
rect 432 82 458 116
rect 492 82 515 116
rect 432 70 515 82
rect 634 197 700 202
rect 634 163 650 197
rect 684 163 700 197
rect 634 120 700 163
rect 634 86 650 120
rect 684 86 700 120
rect 634 17 700 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a221oi_1
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 2901968
string GDS_START 2894110
<< end >>
