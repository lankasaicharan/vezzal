magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2678 1852
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 14 21 1368 203
rect 29 -17 63 21
<< scnmos >>
rect 96 47 126 177
rect 190 47 220 177
rect 284 47 314 177
rect 388 47 418 177
rect 586 47 616 177
rect 670 47 700 177
rect 774 47 804 177
rect 868 47 898 177
rect 978 47 1008 177
rect 1062 47 1092 177
rect 1166 47 1196 177
rect 1260 47 1290 177
<< scpmoshvt >>
rect 98 297 134 497
rect 192 297 228 497
rect 286 297 322 497
rect 380 297 416 497
rect 578 297 614 497
rect 672 297 708 497
rect 766 297 802 497
rect 860 297 896 497
rect 970 297 1006 497
rect 1064 297 1100 497
rect 1158 297 1194 497
rect 1252 297 1288 497
<< ndiff >>
rect 40 95 96 177
rect 40 61 52 95
rect 86 61 96 95
rect 40 47 96 61
rect 126 163 190 177
rect 126 129 146 163
rect 180 129 190 163
rect 126 95 190 129
rect 126 61 146 95
rect 180 61 190 95
rect 126 47 190 61
rect 220 95 284 177
rect 220 61 240 95
rect 274 61 284 95
rect 220 47 284 61
rect 314 163 388 177
rect 314 129 334 163
rect 368 129 388 163
rect 314 95 388 129
rect 314 61 334 95
rect 368 61 388 95
rect 314 47 388 61
rect 418 95 470 177
rect 418 61 428 95
rect 462 61 470 95
rect 418 47 470 61
rect 524 95 586 177
rect 524 61 532 95
rect 566 61 586 95
rect 524 47 586 61
rect 616 163 670 177
rect 616 129 626 163
rect 660 129 670 163
rect 616 47 670 129
rect 700 95 774 177
rect 700 61 720 95
rect 754 61 774 95
rect 700 47 774 61
rect 804 163 868 177
rect 804 129 814 163
rect 848 129 868 163
rect 804 47 868 129
rect 898 163 978 177
rect 898 129 917 163
rect 951 129 978 163
rect 898 95 978 129
rect 898 61 917 95
rect 951 61 978 95
rect 898 47 978 61
rect 1008 95 1062 177
rect 1008 61 1018 95
rect 1052 61 1062 95
rect 1008 47 1062 61
rect 1092 163 1166 177
rect 1092 129 1112 163
rect 1146 129 1166 163
rect 1092 95 1166 129
rect 1092 61 1112 95
rect 1146 61 1166 95
rect 1092 47 1166 61
rect 1196 95 1260 177
rect 1196 61 1206 95
rect 1240 61 1260 95
rect 1196 47 1260 61
rect 1290 163 1342 177
rect 1290 129 1300 163
rect 1334 129 1342 163
rect 1290 95 1342 129
rect 1290 61 1300 95
rect 1334 61 1342 95
rect 1290 47 1342 61
<< pdiff >>
rect 40 483 98 497
rect 40 449 52 483
rect 86 449 98 483
rect 40 415 98 449
rect 40 381 52 415
rect 86 381 98 415
rect 40 297 98 381
rect 134 477 192 497
rect 134 443 146 477
rect 180 443 192 477
rect 134 409 192 443
rect 134 375 146 409
rect 180 375 192 409
rect 134 341 192 375
rect 134 307 146 341
rect 180 307 192 341
rect 134 297 192 307
rect 228 483 286 497
rect 228 449 240 483
rect 274 449 286 483
rect 228 415 286 449
rect 228 381 240 415
rect 274 381 286 415
rect 228 297 286 381
rect 322 477 380 497
rect 322 443 334 477
rect 368 443 380 477
rect 322 409 380 443
rect 322 375 334 409
rect 368 375 380 409
rect 322 341 380 375
rect 322 307 334 341
rect 368 307 380 341
rect 322 297 380 307
rect 416 477 578 497
rect 416 443 428 477
rect 462 443 532 477
rect 566 443 578 477
rect 416 297 578 443
rect 614 477 672 497
rect 614 443 626 477
rect 660 443 672 477
rect 614 297 672 443
rect 708 409 766 497
rect 708 375 720 409
rect 754 375 766 409
rect 708 297 766 375
rect 802 477 860 497
rect 802 443 814 477
rect 848 443 860 477
rect 802 297 860 443
rect 896 477 970 497
rect 896 443 908 477
rect 942 443 970 477
rect 896 297 970 443
rect 1006 477 1064 497
rect 1006 443 1018 477
rect 1052 443 1064 477
rect 1006 297 1064 443
rect 1100 409 1158 497
rect 1100 375 1112 409
rect 1146 375 1158 409
rect 1100 297 1158 375
rect 1194 477 1252 497
rect 1194 443 1206 477
rect 1240 443 1252 477
rect 1194 409 1252 443
rect 1194 375 1206 409
rect 1240 375 1252 409
rect 1194 297 1252 375
rect 1288 477 1347 497
rect 1288 443 1301 477
rect 1335 443 1347 477
rect 1288 409 1347 443
rect 1288 375 1301 409
rect 1335 375 1347 409
rect 1288 341 1347 375
rect 1288 307 1301 341
rect 1335 307 1347 341
rect 1288 297 1347 307
<< ndiffc >>
rect 52 61 86 95
rect 146 129 180 163
rect 146 61 180 95
rect 240 61 274 95
rect 334 129 368 163
rect 334 61 368 95
rect 428 61 462 95
rect 532 61 566 95
rect 626 129 660 163
rect 720 61 754 95
rect 814 129 848 163
rect 917 129 951 163
rect 917 61 951 95
rect 1018 61 1052 95
rect 1112 129 1146 163
rect 1112 61 1146 95
rect 1206 61 1240 95
rect 1300 129 1334 163
rect 1300 61 1334 95
<< pdiffc >>
rect 52 449 86 483
rect 52 381 86 415
rect 146 443 180 477
rect 146 375 180 409
rect 146 307 180 341
rect 240 449 274 483
rect 240 381 274 415
rect 334 443 368 477
rect 334 375 368 409
rect 334 307 368 341
rect 428 443 462 477
rect 532 443 566 477
rect 626 443 660 477
rect 720 375 754 409
rect 814 443 848 477
rect 908 443 942 477
rect 1018 443 1052 477
rect 1112 375 1146 409
rect 1206 443 1240 477
rect 1206 375 1240 409
rect 1301 443 1335 477
rect 1301 375 1335 409
rect 1301 307 1335 341
<< poly >>
rect 98 497 134 523
rect 192 497 228 523
rect 286 497 322 523
rect 380 497 416 523
rect 578 497 614 523
rect 672 497 708 523
rect 766 497 802 523
rect 860 497 896 523
rect 970 497 1006 523
rect 1064 497 1100 523
rect 1158 497 1194 523
rect 1252 497 1288 523
rect 98 282 134 297
rect 192 282 228 297
rect 286 282 322 297
rect 380 282 416 297
rect 578 282 614 297
rect 672 282 708 297
rect 766 282 802 297
rect 860 282 896 297
rect 970 282 1006 297
rect 1064 282 1100 297
rect 1158 282 1194 297
rect 1252 282 1288 297
rect 96 265 136 282
rect 190 265 230 282
rect 284 265 324 282
rect 378 265 418 282
rect 576 265 616 282
rect 670 265 710 282
rect 764 265 804 282
rect 858 265 898 282
rect 968 265 1008 282
rect 1062 265 1102 282
rect 1156 265 1196 282
rect 1250 265 1290 282
rect 96 249 418 265
rect 96 215 124 249
rect 158 215 202 249
rect 236 215 280 249
rect 314 215 358 249
rect 392 215 418 249
rect 96 199 418 215
rect 564 249 628 265
rect 564 215 574 249
rect 608 215 628 249
rect 564 199 628 215
rect 670 249 804 265
rect 670 215 720 249
rect 754 215 804 249
rect 670 199 804 215
rect 846 249 910 265
rect 846 215 856 249
rect 890 215 910 249
rect 846 199 910 215
rect 956 249 1020 265
rect 956 215 966 249
rect 1000 215 1020 249
rect 956 199 1020 215
rect 1062 249 1196 265
rect 1062 215 1112 249
rect 1146 215 1196 249
rect 1062 199 1196 215
rect 1238 249 1302 265
rect 1238 215 1248 249
rect 1282 215 1302 249
rect 1238 199 1302 215
rect 96 177 126 199
rect 190 177 220 199
rect 284 177 314 199
rect 388 177 418 199
rect 586 177 616 199
rect 670 177 700 199
rect 774 177 804 199
rect 868 177 898 199
rect 978 177 1008 199
rect 1062 177 1092 199
rect 1166 177 1196 199
rect 1260 177 1290 199
rect 96 21 126 47
rect 190 21 220 47
rect 284 21 314 47
rect 388 21 418 47
rect 586 21 616 47
rect 670 21 700 47
rect 774 21 804 47
rect 868 21 898 47
rect 978 21 1008 47
rect 1062 21 1092 47
rect 1166 21 1196 47
rect 1260 21 1290 47
<< polycont >>
rect 124 215 158 249
rect 202 215 236 249
rect 280 215 314 249
rect 358 215 392 249
rect 574 215 608 249
rect 720 215 754 249
rect 856 215 890 249
rect 966 215 1000 249
rect 1112 215 1146 249
rect 1248 215 1282 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 44 483 94 527
rect 44 449 52 483
rect 86 449 94 483
rect 44 415 94 449
rect 44 381 52 415
rect 86 381 94 415
rect 44 365 94 381
rect 138 477 188 493
rect 138 443 146 477
rect 180 443 188 477
rect 138 409 188 443
rect 138 375 146 409
rect 180 375 188 409
rect 138 341 188 375
rect 232 483 282 527
rect 232 449 240 483
rect 274 449 282 483
rect 232 415 282 449
rect 232 381 240 415
rect 274 381 282 415
rect 232 359 282 381
rect 326 477 376 493
rect 326 443 334 477
rect 368 443 376 477
rect 326 409 376 443
rect 420 477 574 527
rect 420 443 428 477
rect 462 443 532 477
rect 566 443 574 477
rect 420 425 574 443
rect 618 477 856 493
rect 618 443 626 477
rect 660 459 814 477
rect 660 443 668 459
rect 618 425 668 443
rect 806 443 814 459
rect 848 443 856 477
rect 806 425 856 443
rect 900 477 966 527
rect 900 443 908 477
rect 942 443 966 477
rect 900 425 966 443
rect 1010 477 1248 493
rect 1010 443 1018 477
rect 1052 459 1206 477
rect 1052 443 1060 459
rect 1010 425 1060 443
rect 1198 443 1206 459
rect 1240 443 1248 477
rect 326 375 334 409
rect 368 375 376 409
rect 712 409 762 425
rect 712 391 720 409
rect 138 323 146 341
rect 17 307 146 323
rect 180 323 188 341
rect 326 341 376 375
rect 326 323 334 341
rect 180 307 334 323
rect 368 307 376 341
rect 17 289 376 307
rect 420 375 720 391
rect 754 391 762 409
rect 1104 409 1154 425
rect 1104 391 1112 409
rect 754 375 1112 391
rect 1146 375 1154 409
rect 420 357 1154 375
rect 1198 409 1248 443
rect 1198 375 1206 409
rect 1240 375 1248 409
rect 1198 357 1248 375
rect 1301 477 1342 527
rect 1335 443 1342 477
rect 1301 409 1342 443
rect 1335 375 1342 409
rect 17 181 74 289
rect 420 255 486 357
rect 1301 341 1342 375
rect 108 249 486 255
rect 108 215 124 249
rect 158 215 202 249
rect 236 215 280 249
rect 314 215 358 249
rect 392 215 486 249
rect 524 289 908 323
rect 524 249 636 289
rect 524 215 574 249
rect 608 215 636 249
rect 670 249 806 255
rect 670 215 720 249
rect 754 215 806 249
rect 840 249 908 289
rect 840 215 856 249
rect 890 215 908 249
rect 942 289 1257 323
rect 1335 307 1342 341
rect 1301 291 1342 307
rect 942 249 1026 289
rect 1215 255 1257 289
rect 942 215 966 249
rect 1000 215 1026 249
rect 1070 249 1181 255
rect 1070 215 1112 249
rect 1146 215 1181 249
rect 1215 249 1363 255
rect 1215 215 1248 249
rect 1282 215 1363 249
rect 428 181 486 215
rect 17 163 384 181
rect 17 145 146 163
rect 120 129 146 145
rect 180 145 334 163
rect 180 129 196 145
rect 52 95 86 111
rect 52 17 86 61
rect 120 95 196 129
rect 308 129 334 145
rect 368 129 384 163
rect 428 163 864 181
rect 428 147 626 163
rect 523 129 626 147
rect 660 129 814 163
rect 848 129 864 163
rect 908 163 1350 181
rect 908 129 917 163
rect 951 147 1112 163
rect 951 129 974 147
rect 120 61 146 95
rect 180 61 196 95
rect 120 53 196 61
rect 240 95 274 111
rect 240 17 274 61
rect 308 95 384 129
rect 308 61 334 95
rect 368 61 384 95
rect 308 51 384 61
rect 428 95 462 111
rect 908 95 974 129
rect 1086 129 1112 147
rect 1146 145 1300 163
rect 1146 129 1162 145
rect 428 17 462 61
rect 516 61 532 95
rect 566 61 720 95
rect 754 61 917 95
rect 951 61 974 95
rect 516 51 974 61
rect 1018 95 1052 111
rect 1018 17 1052 61
rect 1086 95 1162 129
rect 1274 129 1300 145
rect 1334 129 1350 163
rect 1086 61 1112 95
rect 1146 61 1162 95
rect 1086 51 1162 61
rect 1206 95 1240 111
rect 1206 17 1240 61
rect 1274 95 1350 129
rect 1274 61 1300 95
rect 1334 61 1350 95
rect 1274 51 1350 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 737 221 771 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 533 221 567 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 1248 221 1282 255 0 FreeSans 400 180 0 0 A1
port 1 nsew signal input
flabel locali s 1070 215 1181 255 0 FreeSans 400 180 0 0 A2
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o22a_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1380 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 958290
string GDS_START 948120
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
