magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 1 49 1151 248
rect 0 0 1152 49
<< scpmos >>
rect 83 384 119 584
rect 173 384 209 584
rect 274 388 310 588
rect 358 388 394 588
rect 586 388 622 588
rect 763 368 799 592
rect 853 368 889 592
rect 943 368 979 592
rect 1033 368 1069 592
<< nmoslvt >>
rect 84 74 114 222
rect 162 74 192 222
rect 248 74 278 222
rect 334 74 364 222
rect 572 74 602 222
rect 770 74 800 222
rect 866 74 896 222
rect 952 74 982 222
rect 1038 74 1068 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 74 162 222
rect 192 120 248 222
rect 192 86 203 120
rect 237 86 248 120
rect 192 74 248 86
rect 278 188 334 222
rect 278 154 289 188
rect 323 154 334 188
rect 278 74 334 154
rect 364 132 414 222
rect 522 218 572 222
rect 515 187 572 218
rect 515 153 527 187
rect 561 153 572 187
rect 364 120 421 132
rect 515 123 572 153
rect 364 86 375 120
rect 409 86 421 120
rect 364 74 421 86
rect 522 74 572 123
rect 602 166 652 222
rect 602 137 659 166
rect 720 138 770 222
rect 602 103 613 137
rect 647 103 659 137
rect 602 74 659 103
rect 713 123 770 138
rect 713 89 725 123
rect 759 89 770 123
rect 713 74 770 89
rect 800 210 866 222
rect 800 176 816 210
rect 850 176 866 210
rect 800 74 866 176
rect 896 123 952 222
rect 896 89 907 123
rect 941 89 952 123
rect 896 74 952 89
rect 982 210 1038 222
rect 982 176 993 210
rect 1027 176 1038 210
rect 982 120 1038 176
rect 982 86 993 120
rect 1027 86 1038 120
rect 982 74 1038 86
rect 1068 210 1125 222
rect 1068 176 1079 210
rect 1113 176 1125 210
rect 1068 120 1125 176
rect 1068 86 1079 120
rect 1113 86 1125 120
rect 1068 74 1125 86
<< pdiff >>
rect 644 588 763 592
rect 224 584 274 588
rect 27 572 83 584
rect 27 538 39 572
rect 73 538 83 572
rect 27 384 83 538
rect 119 430 173 584
rect 119 396 129 430
rect 163 396 173 430
rect 119 384 173 396
rect 209 572 274 584
rect 209 538 224 572
rect 258 538 274 572
rect 209 388 274 538
rect 310 388 358 588
rect 394 434 586 588
rect 394 400 542 434
rect 576 400 586 434
rect 394 388 586 400
rect 622 580 763 588
rect 622 546 632 580
rect 666 546 719 580
rect 753 546 763 580
rect 622 388 763 546
rect 209 384 259 388
rect 713 368 763 388
rect 799 416 853 592
rect 799 382 809 416
rect 843 382 853 416
rect 799 368 853 382
rect 889 575 943 592
rect 889 541 899 575
rect 933 541 943 575
rect 889 368 943 541
rect 979 416 1033 592
rect 979 382 989 416
rect 1023 382 1033 416
rect 979 368 1033 382
rect 1069 575 1125 592
rect 1069 541 1079 575
rect 1113 541 1125 575
rect 1069 368 1125 541
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 203 86 237 120
rect 289 154 323 188
rect 527 153 561 187
rect 375 86 409 120
rect 613 103 647 137
rect 725 89 759 123
rect 816 176 850 210
rect 907 89 941 123
rect 993 176 1027 210
rect 993 86 1027 120
rect 1079 176 1113 210
rect 1079 86 1113 120
<< pdiffc >>
rect 39 538 73 572
rect 129 396 163 430
rect 224 538 258 572
rect 542 400 576 434
rect 632 546 666 580
rect 719 546 753 580
rect 809 382 843 416
rect 899 541 933 575
rect 989 382 1023 416
rect 1079 541 1113 575
<< poly >>
rect 83 584 119 610
rect 173 584 209 610
rect 274 588 310 614
rect 358 588 394 614
rect 586 588 622 614
rect 763 592 799 618
rect 853 592 889 618
rect 943 592 979 618
rect 1033 592 1069 618
rect 83 358 119 384
rect 83 326 114 358
rect 44 310 114 326
rect 173 352 209 384
rect 274 352 310 388
rect 173 336 310 352
rect 173 310 228 336
rect 44 276 60 310
rect 94 276 114 310
rect 44 260 114 276
rect 84 222 114 260
rect 162 302 228 310
rect 262 322 310 336
rect 358 356 394 388
rect 586 358 622 388
rect 358 340 424 356
rect 262 302 278 322
rect 162 280 278 302
rect 162 222 192 280
rect 248 222 278 280
rect 358 306 374 340
rect 408 306 424 340
rect 586 322 616 358
rect 358 290 424 306
rect 473 306 616 322
rect 763 310 799 368
rect 853 310 889 368
rect 943 326 979 368
rect 1033 326 1069 368
rect 943 322 1111 326
rect 358 267 388 290
rect 334 237 388 267
rect 473 272 489 306
rect 523 272 557 306
rect 591 272 616 306
rect 473 256 616 272
rect 664 294 889 310
rect 664 260 680 294
rect 714 260 748 294
rect 782 260 816 294
rect 850 274 889 294
rect 949 310 1111 322
rect 949 276 1061 310
rect 1095 276 1111 310
rect 850 260 896 274
rect 949 260 1111 276
rect 334 222 364 237
rect 572 222 602 256
rect 664 244 896 260
rect 770 222 800 244
rect 866 222 896 244
rect 952 222 982 260
rect 1038 222 1068 260
rect 84 48 114 74
rect 162 48 192 74
rect 248 48 278 74
rect 334 48 364 74
rect 572 48 602 74
rect 770 48 800 74
rect 866 48 896 74
rect 952 48 982 74
rect 1038 48 1068 74
<< polycont >>
rect 60 276 94 310
rect 228 302 262 336
rect 374 306 408 340
rect 489 272 523 306
rect 557 272 591 306
rect 680 260 714 294
rect 748 260 782 294
rect 816 260 850 294
rect 1061 276 1095 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 23 572 89 649
rect 23 538 39 572
rect 73 538 89 572
rect 203 572 280 649
rect 203 538 224 572
rect 258 538 280 572
rect 616 580 769 649
rect 616 546 632 580
rect 666 546 719 580
rect 753 546 769 580
rect 616 536 769 546
rect 883 575 949 649
rect 883 541 899 575
rect 933 541 949 575
rect 883 536 949 541
rect 1063 575 1129 649
rect 1063 541 1079 575
rect 1113 541 1129 575
rect 1063 536 1129 541
rect 25 464 424 504
rect 25 326 59 464
rect 113 396 129 430
rect 163 396 179 430
rect 25 310 110 326
rect 25 276 60 310
rect 94 276 110 310
rect 25 260 110 276
rect 144 256 178 396
rect 212 336 278 356
rect 212 302 228 336
rect 262 302 278 336
rect 212 290 278 302
rect 358 340 424 464
rect 358 306 374 340
rect 408 306 424 340
rect 358 290 424 306
rect 458 468 1111 502
rect 458 322 492 468
rect 526 400 542 434
rect 576 400 698 434
rect 526 384 698 400
rect 458 306 607 322
rect 458 272 489 306
rect 523 272 557 306
rect 591 272 607 306
rect 458 256 607 272
rect 664 310 698 384
rect 793 416 935 434
rect 793 382 809 416
rect 843 382 935 416
rect 793 364 935 382
rect 973 416 1039 434
rect 973 382 989 416
rect 1023 382 1039 416
rect 973 364 1039 382
rect 664 294 866 310
rect 664 260 680 294
rect 714 260 748 294
rect 782 260 816 294
rect 850 260 866 294
rect 144 226 492 256
rect 23 222 492 226
rect 664 244 866 260
rect 664 222 698 244
rect 23 210 178 222
rect 23 176 39 210
rect 73 192 178 210
rect 73 176 89 192
rect 527 188 698 222
rect 901 210 935 364
rect 23 120 89 176
rect 273 154 289 188
rect 323 154 493 188
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 187 86 203 120
rect 237 86 253 120
rect 187 17 253 86
rect 359 86 375 120
rect 409 86 425 120
rect 359 17 425 86
rect 459 85 493 154
rect 527 187 561 188
rect 795 176 816 210
rect 850 176 935 210
rect 977 226 1011 364
rect 1077 326 1111 468
rect 1045 310 1111 326
rect 1045 276 1061 310
rect 1095 276 1111 310
rect 1045 260 1111 276
rect 977 210 1043 226
rect 977 176 993 210
rect 1027 176 1043 210
rect 527 119 561 153
rect 597 137 663 154
rect 597 103 613 137
rect 647 103 663 137
rect 597 85 663 103
rect 459 51 663 85
rect 709 123 775 142
rect 709 89 725 123
rect 759 89 775 123
rect 709 17 775 89
rect 891 123 941 142
rect 891 89 907 123
rect 891 17 941 89
rect 977 120 1043 176
rect 977 86 993 120
rect 1027 86 1043 120
rect 977 70 1043 86
rect 1079 210 1129 226
rect 1113 176 1129 210
rect 1079 120 1129 176
rect 1113 86 1129 120
rect 1079 17 1129 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ha_2
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 SUM
port 8 nsew signal output
flabel locali s 991 94 1025 128 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
flabel locali s 991 168 1025 202 0 FreeSans 340 0 0 0 COUT
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 3754810
string GDS_START 3746058
<< end >>
