magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 29 49 817 265
rect 0 0 864 49
<< scnmos >>
rect 108 155 138 239
rect 216 71 246 239
rect 302 71 332 239
rect 404 71 434 239
rect 528 71 558 239
rect 614 71 644 239
rect 708 71 738 239
<< scpmoshvt >>
rect 108 367 138 451
rect 220 367 250 619
rect 306 367 336 619
rect 424 367 454 619
rect 510 367 540 619
rect 622 367 652 619
rect 708 367 738 619
<< ndiff >>
rect 55 215 108 239
rect 55 181 63 215
rect 97 181 108 215
rect 55 155 108 181
rect 138 158 216 239
rect 138 155 171 158
rect 163 124 171 155
rect 205 124 216 158
rect 163 71 216 124
rect 246 151 302 239
rect 246 117 257 151
rect 291 117 302 151
rect 246 71 302 117
rect 332 159 404 239
rect 332 125 357 159
rect 391 125 404 159
rect 332 71 404 125
rect 434 227 528 239
rect 434 193 464 227
rect 498 193 528 227
rect 434 71 528 193
rect 558 161 614 239
rect 558 127 569 161
rect 603 127 614 161
rect 558 71 614 127
rect 644 151 708 239
rect 644 117 659 151
rect 693 117 708 151
rect 644 71 708 117
rect 738 161 791 239
rect 738 127 749 161
rect 783 127 791 161
rect 738 71 791 127
<< pdiff >>
rect 160 607 220 619
rect 160 573 168 607
rect 202 573 220 607
rect 160 520 220 573
rect 160 486 168 520
rect 202 486 220 520
rect 160 451 220 486
rect 55 424 108 451
rect 55 390 63 424
rect 97 390 108 424
rect 55 367 108 390
rect 138 434 220 451
rect 138 400 158 434
rect 192 400 220 434
rect 138 367 220 400
rect 250 607 306 619
rect 250 573 261 607
rect 295 573 306 607
rect 250 517 306 573
rect 250 483 261 517
rect 295 483 306 517
rect 250 367 306 483
rect 336 601 424 619
rect 336 567 363 601
rect 397 567 424 601
rect 336 367 424 567
rect 454 607 510 619
rect 454 573 465 607
rect 499 573 510 607
rect 454 517 510 573
rect 454 483 465 517
rect 499 483 510 517
rect 454 367 510 483
rect 540 601 622 619
rect 540 567 564 601
rect 598 567 622 601
rect 540 367 622 567
rect 652 607 708 619
rect 652 573 663 607
rect 697 573 708 607
rect 652 517 708 573
rect 652 483 663 517
rect 697 483 708 517
rect 652 367 708 483
rect 738 601 791 619
rect 738 567 749 601
rect 783 567 791 601
rect 738 367 791 567
<< ndiffc >>
rect 63 181 97 215
rect 171 124 205 158
rect 257 117 291 151
rect 357 125 391 159
rect 464 193 498 227
rect 569 127 603 161
rect 659 117 693 151
rect 749 127 783 161
<< pdiffc >>
rect 168 573 202 607
rect 168 486 202 520
rect 63 390 97 424
rect 158 400 192 434
rect 261 573 295 607
rect 261 483 295 517
rect 363 567 397 601
rect 465 573 499 607
rect 465 483 499 517
rect 564 567 598 601
rect 663 573 697 607
rect 663 483 697 517
rect 749 567 783 601
<< poly >>
rect 220 619 250 645
rect 306 619 336 645
rect 424 619 454 645
rect 510 619 540 645
rect 622 619 652 645
rect 708 619 738 645
rect 108 451 138 477
rect 108 335 138 367
rect 220 335 250 367
rect 306 335 336 367
rect 72 319 138 335
rect 72 285 88 319
rect 122 285 138 319
rect 72 269 138 285
rect 184 319 250 335
rect 184 285 200 319
rect 234 285 250 319
rect 184 269 250 285
rect 292 319 358 335
rect 424 327 454 367
rect 510 327 540 367
rect 622 335 652 367
rect 708 335 738 367
rect 292 285 308 319
rect 342 285 358 319
rect 292 269 358 285
rect 404 311 540 327
rect 404 277 420 311
rect 454 291 540 311
rect 600 319 666 335
rect 454 277 558 291
rect 108 239 138 269
rect 216 239 246 269
rect 302 239 332 269
rect 404 261 558 277
rect 600 285 616 319
rect 650 285 666 319
rect 600 269 666 285
rect 708 319 774 335
rect 708 285 724 319
rect 758 285 774 319
rect 708 269 774 285
rect 404 239 434 261
rect 528 239 558 261
rect 614 239 644 269
rect 708 239 738 269
rect 108 129 138 155
rect 216 45 246 71
rect 302 45 332 71
rect 404 45 434 71
rect 528 45 558 71
rect 614 45 644 71
rect 708 45 738 71
<< polycont >>
rect 88 285 122 319
rect 200 285 234 319
rect 308 285 342 319
rect 420 277 454 311
rect 616 285 650 319
rect 724 285 758 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 147 607 204 649
rect 147 573 168 607
rect 202 573 204 607
rect 147 520 204 573
rect 147 486 168 520
rect 202 486 204 520
rect 18 424 113 440
rect 18 390 63 424
rect 97 390 113 424
rect 18 384 113 390
rect 147 434 204 486
rect 245 607 311 615
rect 245 573 261 607
rect 295 573 311 607
rect 245 517 311 573
rect 347 601 413 649
rect 347 567 363 601
rect 397 567 413 601
rect 347 551 413 567
rect 449 607 515 615
rect 449 573 465 607
rect 499 573 515 607
rect 449 517 515 573
rect 549 601 613 649
rect 549 567 564 601
rect 598 567 613 601
rect 549 551 613 567
rect 647 607 713 615
rect 647 573 663 607
rect 697 573 713 607
rect 647 517 713 573
rect 747 601 799 649
rect 747 567 749 601
rect 783 567 799 601
rect 747 551 799 567
rect 245 483 261 517
rect 295 483 465 517
rect 499 483 663 517
rect 697 483 847 517
rect 147 400 158 434
rect 192 400 204 434
rect 147 384 204 400
rect 238 415 758 449
rect 18 235 52 384
rect 238 350 272 415
rect 86 319 166 350
rect 86 285 88 319
rect 122 285 166 319
rect 86 269 166 285
rect 200 319 272 350
rect 234 285 272 319
rect 200 269 272 285
rect 306 347 666 381
rect 306 319 344 347
rect 306 285 308 319
rect 342 285 344 319
rect 504 319 666 347
rect 306 269 344 285
rect 378 311 470 313
rect 378 277 420 311
rect 454 277 470 311
rect 378 269 470 277
rect 504 285 616 319
rect 650 285 666 319
rect 504 269 666 285
rect 708 319 758 415
rect 708 285 724 319
rect 708 269 758 285
rect 378 235 412 269
rect 792 235 847 483
rect 18 215 412 235
rect 18 181 63 215
rect 97 201 412 215
rect 448 227 847 235
rect 97 181 113 201
rect 448 193 464 227
rect 498 201 847 227
rect 498 193 514 201
rect 448 187 514 193
rect 18 165 113 181
rect 155 158 221 167
rect 155 124 171 158
rect 205 124 221 158
rect 155 17 221 124
rect 255 151 307 167
rect 255 117 257 151
rect 291 117 307 151
rect 341 159 407 167
rect 341 125 357 159
rect 391 153 407 159
rect 553 161 619 167
rect 553 153 569 161
rect 391 127 569 153
rect 603 127 619 161
rect 391 125 619 127
rect 341 119 619 125
rect 653 151 699 167
rect 255 85 307 117
rect 653 117 659 151
rect 693 117 699 151
rect 653 85 699 117
rect 255 51 699 85
rect 733 161 799 167
rect 733 127 749 161
rect 783 127 799 161
rect 733 17 799 127
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand3b_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 799 464 833 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3730184
string GDS_START 3723048
<< end >>
