magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1682 1975
<< nwell >>
rect -38 331 422 704
<< pwell >>
rect 23 49 383 157
rect 0 0 384 49
<< scnmos >>
rect 102 47 132 131
rect 188 47 218 131
rect 274 47 304 131
<< scpmoshvt >>
rect 116 397 146 481
rect 188 397 218 481
rect 274 397 304 481
<< ndiff >>
rect 49 93 102 131
rect 49 59 57 93
rect 91 59 102 93
rect 49 47 102 59
rect 132 119 188 131
rect 132 85 143 119
rect 177 85 188 119
rect 132 47 188 85
rect 218 93 274 131
rect 218 59 229 93
rect 263 59 274 93
rect 218 47 274 59
rect 304 119 357 131
rect 304 85 315 119
rect 349 85 357 119
rect 304 47 357 85
<< pdiff >>
rect 63 443 116 481
rect 63 409 71 443
rect 105 409 116 443
rect 63 397 116 409
rect 146 397 188 481
rect 218 469 274 481
rect 218 435 229 469
rect 263 435 274 469
rect 218 397 274 435
rect 304 443 357 481
rect 304 409 315 443
rect 349 409 357 443
rect 304 397 357 409
<< ndiffc >>
rect 57 59 91 93
rect 143 85 177 119
rect 229 59 263 93
rect 315 85 349 119
<< pdiffc >>
rect 71 409 105 443
rect 229 435 263 469
rect 315 409 349 443
<< poly >>
rect 123 605 189 621
rect 123 571 139 605
rect 173 585 189 605
rect 173 571 304 585
rect 123 555 304 571
rect 116 481 146 507
rect 188 481 218 507
rect 274 481 304 555
rect 116 375 146 397
rect 57 345 146 375
rect 57 287 87 345
rect 188 297 218 397
rect 21 271 87 287
rect 21 237 37 271
rect 71 237 87 271
rect 21 203 87 237
rect 139 281 218 297
rect 139 247 155 281
rect 189 247 218 281
rect 139 231 218 247
rect 21 169 37 203
rect 71 183 87 203
rect 71 169 132 183
rect 21 153 132 169
rect 102 131 132 153
rect 188 131 218 231
rect 274 131 304 397
rect 102 21 132 47
rect 188 21 218 47
rect 274 21 304 47
<< polycont >>
rect 139 571 173 605
rect 37 237 71 271
rect 155 247 189 281
rect 37 169 71 203
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 123 571 139 605
rect 173 571 189 605
rect 123 459 189 571
rect 67 443 189 459
rect 67 409 71 443
rect 105 409 189 443
rect 225 469 267 649
rect 225 435 229 469
rect 263 435 267 469
rect 225 419 267 435
rect 311 443 353 572
rect 67 383 189 409
rect 311 409 315 443
rect 349 409 353 443
rect 67 349 275 383
rect 31 271 71 287
rect 31 237 37 271
rect 127 247 155 281
rect 189 247 205 281
rect 127 242 205 247
rect 31 203 71 237
rect 31 169 37 203
rect 241 179 275 349
rect 31 153 71 169
rect 139 145 275 179
rect 139 119 181 145
rect 53 93 95 109
rect 53 59 57 93
rect 91 59 95 93
rect 139 85 143 119
rect 177 85 181 119
rect 311 119 353 409
rect 139 69 181 85
rect 225 93 267 109
rect 53 17 95 59
rect 225 59 229 93
rect 263 59 267 93
rect 311 85 315 119
rect 349 85 353 119
rect 311 69 353 85
rect 225 17 267 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 683 384 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 384 683
rect 0 617 384 649
rect 0 17 384 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -49 384 -17
<< labels >>
flabel pwell s 0 0 384 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 384 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or2_m
flabel metal1 s 0 617 384 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 384 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 384 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6165684
string GDS_START 6160860
<< end >>
