magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 331 1478 704
rect 959 300 1171 331
<< pwell >>
rect 1163 241 1437 258
rect 31 157 321 240
rect 957 157 1437 241
rect 31 49 1437 157
rect 0 0 1440 49
<< scnmos >>
rect 110 130 140 214
rect 212 130 242 214
rect 553 47 583 131
rect 639 47 669 131
rect 711 47 741 131
rect 819 47 849 131
rect 927 47 957 131
rect 1036 47 1066 215
rect 1242 64 1272 232
rect 1328 64 1358 232
<< scpmoshvt >>
rect 126 481 156 609
rect 212 481 242 609
rect 402 481 432 609
rect 561 481 591 609
rect 633 481 663 609
rect 741 481 771 565
rect 849 481 879 565
rect 1052 336 1082 588
rect 1242 367 1272 619
rect 1328 367 1358 619
<< ndiff >>
rect 57 189 110 214
rect 57 155 65 189
rect 99 155 110 189
rect 57 130 110 155
rect 140 200 212 214
rect 140 166 151 200
rect 185 166 212 200
rect 140 130 212 166
rect 242 202 295 214
rect 242 168 253 202
rect 287 168 295 202
rect 242 130 295 168
rect 983 202 1036 215
rect 983 168 991 202
rect 1025 168 1036 202
rect 983 131 1036 168
rect 500 105 553 131
rect 500 71 508 105
rect 542 71 553 105
rect 500 47 553 71
rect 583 89 639 131
rect 583 55 594 89
rect 628 55 639 89
rect 583 47 639 55
rect 669 47 711 131
rect 741 91 819 131
rect 741 57 774 91
rect 808 57 819 91
rect 741 47 819 57
rect 849 47 927 131
rect 957 93 1036 131
rect 957 59 991 93
rect 1025 59 1036 93
rect 957 47 1036 59
rect 1066 202 1119 215
rect 1066 168 1077 202
rect 1111 168 1119 202
rect 1066 101 1119 168
rect 1066 67 1077 101
rect 1111 67 1119 101
rect 1066 47 1119 67
rect 1189 204 1242 232
rect 1189 170 1197 204
rect 1231 170 1242 204
rect 1189 110 1242 170
rect 1189 76 1197 110
rect 1231 76 1242 110
rect 1189 64 1242 76
rect 1272 220 1328 232
rect 1272 186 1283 220
rect 1317 186 1328 220
rect 1272 110 1328 186
rect 1272 76 1283 110
rect 1317 76 1328 110
rect 1272 64 1328 76
rect 1358 220 1411 232
rect 1358 186 1369 220
rect 1403 186 1411 220
rect 1358 110 1411 186
rect 1358 76 1369 110
rect 1403 76 1411 110
rect 1358 64 1411 76
<< pdiff >>
rect 73 595 126 609
rect 73 561 81 595
rect 115 561 126 595
rect 73 527 126 561
rect 73 493 81 527
rect 115 493 126 527
rect 73 481 126 493
rect 156 601 212 609
rect 156 567 167 601
rect 201 567 212 601
rect 156 533 212 567
rect 156 499 167 533
rect 201 499 212 533
rect 156 481 212 499
rect 242 597 295 609
rect 242 563 253 597
rect 287 563 295 597
rect 242 529 295 563
rect 242 495 253 529
rect 287 495 295 529
rect 242 481 295 495
rect 349 531 402 609
rect 349 497 357 531
rect 391 497 402 531
rect 349 481 402 497
rect 432 593 561 609
rect 432 559 497 593
rect 531 559 561 593
rect 432 481 561 559
rect 591 481 633 609
rect 663 593 716 609
rect 663 559 674 593
rect 708 565 716 593
rect 1189 604 1242 619
rect 995 580 1052 588
rect 995 565 1007 580
rect 708 559 741 565
rect 663 481 741 559
rect 771 481 849 565
rect 879 549 1007 565
rect 879 515 895 549
rect 929 546 1007 549
rect 1041 546 1052 580
rect 929 515 1052 546
rect 879 512 1052 515
rect 879 481 1007 512
rect 995 478 1007 481
rect 1041 478 1052 512
rect 995 444 1052 478
rect 995 410 1007 444
rect 1041 410 1052 444
rect 995 336 1052 410
rect 1082 576 1135 588
rect 1082 542 1093 576
rect 1127 542 1135 576
rect 1082 478 1135 542
rect 1082 444 1093 478
rect 1127 444 1135 478
rect 1082 382 1135 444
rect 1082 348 1093 382
rect 1127 348 1135 382
rect 1189 570 1197 604
rect 1231 570 1242 604
rect 1189 509 1242 570
rect 1189 475 1197 509
rect 1231 475 1242 509
rect 1189 413 1242 475
rect 1189 379 1197 413
rect 1231 379 1242 413
rect 1189 367 1242 379
rect 1272 599 1328 619
rect 1272 565 1283 599
rect 1317 565 1328 599
rect 1272 505 1328 565
rect 1272 471 1283 505
rect 1317 471 1328 505
rect 1272 409 1328 471
rect 1272 375 1283 409
rect 1317 375 1328 409
rect 1272 367 1328 375
rect 1358 604 1411 619
rect 1358 570 1369 604
rect 1403 570 1411 604
rect 1358 509 1411 570
rect 1358 475 1369 509
rect 1403 475 1411 509
rect 1358 413 1411 475
rect 1358 379 1369 413
rect 1403 379 1411 413
rect 1358 367 1411 379
rect 1082 336 1135 348
<< ndiffc >>
rect 65 155 99 189
rect 151 166 185 200
rect 253 168 287 202
rect 991 168 1025 202
rect 508 71 542 105
rect 594 55 628 89
rect 774 57 808 91
rect 991 59 1025 93
rect 1077 168 1111 202
rect 1077 67 1111 101
rect 1197 170 1231 204
rect 1197 76 1231 110
rect 1283 186 1317 220
rect 1283 76 1317 110
rect 1369 186 1403 220
rect 1369 76 1403 110
<< pdiffc >>
rect 81 561 115 595
rect 81 493 115 527
rect 167 567 201 601
rect 167 499 201 533
rect 253 563 287 597
rect 253 495 287 529
rect 357 497 391 531
rect 497 559 531 593
rect 674 559 708 593
rect 895 515 929 549
rect 1007 546 1041 580
rect 1007 478 1041 512
rect 1007 410 1041 444
rect 1093 542 1127 576
rect 1093 444 1127 478
rect 1093 348 1127 382
rect 1197 570 1231 604
rect 1197 475 1231 509
rect 1197 379 1231 413
rect 1283 565 1317 599
rect 1283 471 1317 505
rect 1283 375 1317 409
rect 1369 570 1403 604
rect 1369 475 1403 509
rect 1369 379 1403 413
<< poly >>
rect 126 609 156 635
rect 212 609 242 635
rect 402 609 432 635
rect 561 609 591 635
rect 633 609 663 635
rect 1242 619 1272 645
rect 1328 619 1358 645
rect 741 565 771 591
rect 849 565 879 591
rect 1052 588 1082 614
rect 126 302 156 481
rect 98 286 164 302
rect 98 252 114 286
rect 148 252 164 286
rect 98 236 164 252
rect 212 266 242 481
rect 402 298 432 481
rect 561 387 591 481
rect 519 371 591 387
rect 519 337 535 371
rect 569 337 591 371
rect 519 303 591 337
rect 402 282 468 298
rect 212 236 340 266
rect 110 214 140 236
rect 212 214 242 236
rect 110 104 140 130
rect 212 104 242 130
rect 310 105 340 236
rect 402 248 418 282
rect 452 248 468 282
rect 519 269 535 303
rect 569 269 591 303
rect 633 441 663 481
rect 741 449 771 481
rect 849 449 879 481
rect 633 425 699 441
rect 633 391 649 425
rect 683 391 699 425
rect 633 357 699 391
rect 741 433 807 449
rect 741 399 757 433
rect 791 399 807 433
rect 849 433 963 449
rect 849 419 913 433
rect 741 383 807 399
rect 897 399 913 419
rect 947 399 963 433
rect 633 323 649 357
rect 683 327 699 357
rect 897 365 963 399
rect 897 331 913 365
rect 947 331 963 365
rect 683 323 849 327
rect 633 297 849 323
rect 897 315 963 331
rect 519 255 591 269
rect 819 267 849 297
rect 519 253 669 255
rect 402 214 468 248
rect 555 225 669 253
rect 402 180 418 214
rect 452 183 468 214
rect 452 180 583 183
rect 402 153 583 180
rect 553 131 583 153
rect 639 131 669 225
rect 711 233 777 249
rect 711 199 727 233
rect 761 199 777 233
rect 711 183 777 199
rect 819 218 885 267
rect 819 184 835 218
rect 869 184 885 218
rect 711 131 741 183
rect 819 168 885 184
rect 819 131 849 168
rect 927 131 957 315
rect 1052 304 1082 336
rect 1242 320 1272 367
rect 1005 288 1082 304
rect 1005 254 1021 288
rect 1055 254 1082 288
rect 1167 314 1272 320
rect 1328 314 1358 367
rect 1167 304 1358 314
rect 1167 270 1183 304
rect 1217 284 1358 304
rect 1217 270 1272 284
rect 1167 254 1272 270
rect 1005 238 1082 254
rect 1036 215 1066 238
rect 1242 232 1272 254
rect 1328 232 1358 284
rect 310 89 376 105
rect 310 55 326 89
rect 360 55 376 89
rect 310 39 376 55
rect 553 21 583 47
rect 639 21 669 47
rect 711 21 741 47
rect 819 21 849 47
rect 927 21 957 47
rect 1036 21 1066 47
rect 1242 38 1272 64
rect 1328 38 1358 64
<< polycont >>
rect 114 252 148 286
rect 535 337 569 371
rect 418 248 452 282
rect 535 269 569 303
rect 649 391 683 425
rect 757 399 791 433
rect 913 399 947 433
rect 649 323 683 357
rect 913 331 947 365
rect 418 180 452 214
rect 727 199 761 233
rect 835 184 869 218
rect 1021 254 1055 288
rect 1183 270 1217 304
rect 326 55 360 89
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 28 595 125 611
rect 28 561 81 595
rect 115 561 125 595
rect 28 527 125 561
rect 28 493 81 527
rect 115 493 125 527
rect 28 371 125 493
rect 159 601 209 649
rect 159 567 167 601
rect 201 567 209 601
rect 159 533 209 567
rect 159 499 167 533
rect 201 499 209 533
rect 159 483 209 499
rect 243 597 461 615
rect 243 563 253 597
rect 287 581 461 597
rect 287 563 303 581
rect 243 529 303 563
rect 243 495 253 529
rect 287 495 303 529
rect 243 479 303 495
rect 341 531 391 547
rect 341 497 357 531
rect 341 441 391 497
rect 427 509 461 581
rect 495 593 547 649
rect 495 559 497 593
rect 531 559 547 593
rect 495 543 547 559
rect 658 593 861 613
rect 658 559 674 593
rect 708 559 861 593
rect 658 543 861 559
rect 427 475 793 509
rect 341 425 699 441
rect 341 407 649 425
rect 633 391 649 407
rect 683 391 699 425
rect 28 337 535 371
rect 569 337 585 371
rect 28 332 585 337
rect 28 205 62 332
rect 519 303 585 332
rect 633 357 699 391
rect 633 323 649 357
rect 683 323 699 357
rect 633 307 699 323
rect 741 433 793 475
rect 741 399 757 433
rect 791 399 793 433
rect 741 383 793 399
rect 98 286 371 298
rect 98 252 114 286
rect 148 252 371 286
rect 98 240 371 252
rect 405 282 468 298
rect 405 248 418 282
rect 452 248 468 282
rect 519 269 535 303
rect 569 269 585 303
rect 405 233 468 248
rect 741 233 785 383
rect 827 290 861 543
rect 895 580 1049 649
rect 1181 604 1240 649
rect 895 549 1007 580
rect 929 546 1007 549
rect 1041 546 1049 580
rect 929 515 1049 546
rect 895 512 1049 515
rect 895 499 1007 512
rect 1003 478 1007 499
rect 1041 478 1049 512
rect 897 433 963 449
rect 897 399 913 433
rect 947 399 963 433
rect 897 365 963 399
rect 1003 444 1049 478
rect 1003 410 1007 444
rect 1041 410 1049 444
rect 1003 392 1049 410
rect 1083 576 1141 592
rect 1083 542 1093 576
rect 1127 542 1141 576
rect 1083 478 1141 542
rect 1083 444 1093 478
rect 1127 444 1141 478
rect 897 331 913 365
rect 947 358 963 365
rect 1083 382 1141 444
rect 1083 358 1093 382
rect 947 348 1093 358
rect 1127 348 1141 382
rect 1181 570 1197 604
rect 1231 570 1240 604
rect 1181 509 1240 570
rect 1181 475 1197 509
rect 1231 475 1240 509
rect 1181 413 1240 475
rect 1181 379 1197 413
rect 1231 379 1240 413
rect 1181 363 1240 379
rect 1274 599 1327 615
rect 1274 565 1283 599
rect 1317 565 1327 599
rect 1274 505 1327 565
rect 1274 471 1283 505
rect 1317 471 1327 505
rect 1274 409 1327 471
rect 1274 375 1283 409
rect 1317 375 1327 409
rect 947 331 1141 348
rect 897 324 1141 331
rect 1107 320 1141 324
rect 1107 304 1233 320
rect 827 288 1071 290
rect 827 254 1021 288
rect 1055 254 1071 288
rect 405 214 727 233
rect 405 206 418 214
rect 28 189 99 205
rect 28 155 65 189
rect 28 139 99 155
rect 135 200 201 205
rect 135 166 151 200
rect 185 166 201 200
rect 135 162 201 166
rect 237 202 418 206
rect 237 168 253 202
rect 287 180 418 202
rect 452 199 727 214
rect 761 199 785 233
rect 921 252 1071 254
rect 1107 270 1183 304
rect 1217 270 1233 304
rect 1107 254 1233 270
rect 819 218 885 220
rect 452 180 458 199
rect 287 168 458 180
rect 237 162 458 168
rect 819 184 835 218
rect 869 184 885 218
rect 819 163 885 184
rect 135 17 169 162
rect 492 129 885 163
rect 203 89 458 128
rect 203 55 326 89
rect 360 55 458 89
rect 492 105 544 129
rect 492 71 508 105
rect 542 71 544 105
rect 921 95 955 252
rect 1107 218 1141 254
rect 1274 220 1327 375
rect 1361 604 1419 649
rect 1361 570 1369 604
rect 1403 570 1419 604
rect 1361 509 1419 570
rect 1361 475 1369 509
rect 1403 475 1419 509
rect 1361 413 1419 475
rect 1361 379 1369 413
rect 1403 379 1419 413
rect 1361 363 1419 379
rect 492 55 544 71
rect 578 89 644 95
rect 578 55 594 89
rect 628 55 644 89
rect 578 17 644 55
rect 758 91 955 95
rect 758 57 774 91
rect 808 57 955 91
rect 758 51 955 57
rect 989 202 1034 218
rect 989 168 991 202
rect 1025 168 1034 202
rect 989 93 1034 168
rect 989 59 991 93
rect 1025 59 1034 93
rect 989 17 1034 59
rect 1068 202 1141 218
rect 1068 168 1077 202
rect 1111 168 1141 202
rect 1068 101 1141 168
rect 1068 67 1077 101
rect 1111 67 1141 101
rect 1068 51 1141 67
rect 1181 204 1240 220
rect 1181 170 1197 204
rect 1231 170 1240 204
rect 1181 110 1240 170
rect 1181 76 1197 110
rect 1231 76 1240 110
rect 1181 17 1240 76
rect 1274 186 1283 220
rect 1317 186 1327 220
rect 1274 110 1327 186
rect 1274 76 1283 110
rect 1317 76 1327 110
rect 1274 60 1327 76
rect 1361 220 1419 236
rect 1361 186 1369 220
rect 1403 186 1419 220
rect 1361 110 1419 186
rect 1361 76 1369 110
rect 1403 76 1419 110
rect 1361 17 1419 76
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlxtn_2
flabel comment s 755 316 755 316 0 FreeSans 200 0 0 0 no_jumper_check
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 415 94 449 128 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1279 94 1313 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 168 1313 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 464 1313 498 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1279 538 1313 572 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 638314
string GDS_START 626158
<< end >>
