magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 331 2150 704
<< pwell >>
rect 329 195 1840 251
rect 21 176 1840 195
rect 21 49 2111 176
rect 0 0 2112 49
<< scnmos >>
rect 104 85 134 169
rect 176 85 206 169
rect 428 141 458 225
rect 547 141 577 225
rect 625 141 655 225
rect 739 141 769 225
rect 857 141 887 225
rect 975 141 1005 225
rect 1093 141 1123 225
rect 1458 141 1488 225
rect 1544 141 1574 225
rect 1656 141 1686 225
rect 1734 141 1764 225
rect 1829 66 1859 150
rect 1926 66 1956 150
rect 1998 66 2028 150
<< scpmoshvt >>
rect 84 383 134 583
rect 302 409 352 609
rect 408 409 458 609
rect 661 419 711 619
rect 767 419 817 619
rect 893 419 943 619
rect 999 419 1049 619
rect 1105 419 1155 619
rect 1458 419 1508 619
rect 1564 419 1614 619
rect 1670 419 1720 619
rect 1768 419 1818 619
rect 1872 419 1922 619
rect 1978 419 2028 619
<< ndiff >>
rect 47 144 104 169
rect 47 110 59 144
rect 93 110 104 144
rect 47 85 104 110
rect 134 85 176 169
rect 206 144 263 169
rect 206 110 217 144
rect 251 110 263 144
rect 206 85 263 110
rect 355 187 428 225
rect 355 153 367 187
rect 401 153 428 187
rect 355 141 428 153
rect 458 200 547 225
rect 458 166 469 200
rect 503 166 547 200
rect 458 141 547 166
rect 577 141 625 225
rect 655 191 739 225
rect 655 157 666 191
rect 700 157 739 191
rect 655 141 739 157
rect 769 141 857 225
rect 887 141 975 225
rect 1005 141 1093 225
rect 1123 187 1458 225
rect 1123 153 1134 187
rect 1168 153 1458 187
rect 1123 141 1458 153
rect 1488 187 1544 225
rect 1488 153 1499 187
rect 1533 153 1544 187
rect 1488 141 1544 153
rect 1574 198 1656 225
rect 1574 164 1611 198
rect 1645 164 1656 198
rect 1574 141 1656 164
rect 1686 141 1734 225
rect 1764 150 1814 225
rect 1764 141 1829 150
rect 784 114 842 141
rect 784 80 796 114
rect 830 80 842 114
rect 784 68 842 80
rect 902 114 960 141
rect 902 80 914 114
rect 948 80 960 114
rect 902 68 960 80
rect 1020 114 1078 141
rect 1020 80 1032 114
rect 1066 80 1078 114
rect 1020 68 1078 80
rect 1779 66 1829 141
rect 1859 125 1926 150
rect 1859 91 1870 125
rect 1904 91 1926 125
rect 1859 66 1926 91
rect 1956 66 1998 150
rect 2028 125 2085 150
rect 2028 91 2039 125
rect 2073 91 2085 125
rect 2028 66 2085 91
<< pdiff >>
rect 245 597 302 609
rect 27 571 84 583
rect 27 537 39 571
rect 73 537 84 571
rect 27 500 84 537
rect 27 466 39 500
rect 73 466 84 500
rect 27 429 84 466
rect 27 395 39 429
rect 73 395 84 429
rect 27 383 84 395
rect 134 571 191 583
rect 134 537 145 571
rect 179 537 191 571
rect 134 500 191 537
rect 134 466 145 500
rect 179 466 191 500
rect 134 429 191 466
rect 134 395 145 429
rect 179 395 191 429
rect 245 563 257 597
rect 291 563 302 597
rect 245 526 302 563
rect 245 492 257 526
rect 291 492 302 526
rect 245 455 302 492
rect 245 421 257 455
rect 291 421 302 455
rect 245 409 302 421
rect 352 597 408 609
rect 352 563 363 597
rect 397 563 408 597
rect 352 499 408 563
rect 352 465 363 499
rect 397 465 408 499
rect 352 409 408 465
rect 458 568 515 609
rect 458 534 469 568
rect 503 534 515 568
rect 458 409 515 534
rect 569 498 661 619
rect 569 464 581 498
rect 615 464 661 498
rect 569 419 661 464
rect 711 525 767 619
rect 711 491 722 525
rect 756 491 767 525
rect 711 419 767 491
rect 817 575 893 619
rect 817 541 828 575
rect 862 541 893 575
rect 817 419 893 541
rect 943 580 999 619
rect 943 546 954 580
rect 988 546 999 580
rect 943 419 999 546
rect 1049 575 1105 619
rect 1049 541 1060 575
rect 1094 541 1105 575
rect 1049 419 1105 541
rect 1155 607 1458 619
rect 1155 573 1166 607
rect 1200 573 1458 607
rect 1155 419 1458 573
rect 1508 575 1564 619
rect 1508 541 1519 575
rect 1553 541 1564 575
rect 1508 419 1564 541
rect 1614 575 1670 619
rect 1614 541 1625 575
rect 1659 541 1670 575
rect 1614 419 1670 541
rect 1720 419 1768 619
rect 1818 419 1872 619
rect 1922 607 1978 619
rect 1922 573 1933 607
rect 1967 573 1978 607
rect 1922 536 1978 573
rect 1922 502 1933 536
rect 1967 502 1978 536
rect 1922 465 1978 502
rect 1922 431 1933 465
rect 1967 431 1978 465
rect 1922 419 1978 431
rect 2028 597 2085 619
rect 2028 563 2039 597
rect 2073 563 2085 597
rect 2028 465 2085 563
rect 2028 431 2039 465
rect 2073 431 2085 465
rect 2028 419 2085 431
rect 134 383 191 395
<< ndiffc >>
rect 59 110 93 144
rect 217 110 251 144
rect 367 153 401 187
rect 469 166 503 200
rect 666 157 700 191
rect 1134 153 1168 187
rect 1499 153 1533 187
rect 1611 164 1645 198
rect 796 80 830 114
rect 914 80 948 114
rect 1032 80 1066 114
rect 1870 91 1904 125
rect 2039 91 2073 125
<< pdiffc >>
rect 39 537 73 571
rect 39 466 73 500
rect 39 395 73 429
rect 145 537 179 571
rect 145 466 179 500
rect 145 395 179 429
rect 257 563 291 597
rect 257 492 291 526
rect 257 421 291 455
rect 363 563 397 597
rect 363 465 397 499
rect 469 534 503 568
rect 581 464 615 498
rect 722 491 756 525
rect 828 541 862 575
rect 954 546 988 580
rect 1060 541 1094 575
rect 1166 573 1200 607
rect 1519 541 1553 575
rect 1625 541 1659 575
rect 1933 573 1967 607
rect 1933 502 1967 536
rect 1933 431 1967 465
rect 2039 563 2073 597
rect 2039 431 2073 465
<< poly >>
rect 302 609 352 635
rect 408 609 458 635
rect 661 619 711 645
rect 767 619 817 645
rect 893 619 943 645
rect 999 619 1049 645
rect 1105 619 1155 645
rect 1458 619 1508 645
rect 1564 619 1614 645
rect 1670 619 1720 645
rect 1768 619 1818 645
rect 1872 619 1922 645
rect 1978 619 2028 645
rect 84 583 134 609
rect 84 343 134 383
rect 84 327 206 343
rect 84 293 156 327
rect 190 293 206 327
rect 84 259 206 293
rect 84 225 156 259
rect 190 225 206 259
rect 84 209 206 225
rect 104 169 134 209
rect 176 169 206 209
rect 302 281 352 409
rect 408 281 458 409
rect 661 318 711 419
rect 767 384 817 419
rect 893 404 943 419
rect 999 404 1049 419
rect 767 368 845 384
rect 767 334 795 368
rect 829 334 845 368
rect 767 318 845 334
rect 893 374 1049 404
rect 1105 384 1155 419
rect 661 313 691 318
rect 302 251 458 281
rect 625 297 691 313
rect 625 263 641 297
rect 675 263 691 297
rect 767 270 797 318
rect 893 313 923 374
rect 1105 368 1416 384
rect 1105 334 1366 368
rect 1400 334 1416 368
rect 1105 326 1416 334
rect 1093 318 1416 326
rect 1458 375 1508 419
rect 887 297 1005 313
rect 887 270 903 297
rect 104 59 134 85
rect 176 59 206 85
rect 302 51 332 251
rect 428 225 458 251
rect 547 225 577 251
rect 625 247 691 263
rect 625 225 655 247
rect 739 240 797 270
rect 857 263 903 270
rect 937 263 1005 297
rect 857 240 1005 263
rect 739 225 769 240
rect 857 225 887 240
rect 975 225 1005 240
rect 1093 296 1135 318
rect 1093 225 1123 296
rect 1458 225 1488 375
rect 1564 327 1614 419
rect 1670 387 1720 419
rect 1768 387 1818 419
rect 1656 371 1722 387
rect 1656 337 1672 371
rect 1706 337 1722 371
rect 1536 311 1602 327
rect 1536 277 1552 311
rect 1586 277 1602 311
rect 1536 261 1602 277
rect 1656 321 1722 337
rect 1764 371 1830 387
rect 1764 337 1780 371
rect 1814 337 1830 371
rect 1764 321 1830 337
rect 1544 225 1574 261
rect 1656 225 1686 321
rect 1770 273 1800 321
rect 1872 273 1922 419
rect 1978 378 2028 419
rect 1734 243 1800 273
rect 1848 243 1922 273
rect 1964 362 2030 378
rect 1964 328 1980 362
rect 2014 328 2030 362
rect 1964 294 2030 328
rect 1964 260 1980 294
rect 2014 260 2030 294
rect 1964 244 2030 260
rect 1734 225 1764 243
rect 1848 195 1878 243
rect 1998 195 2028 244
rect 1829 165 1878 195
rect 1926 165 2028 195
rect 1829 150 1859 165
rect 1926 150 1956 165
rect 1998 150 2028 165
rect 428 115 458 141
rect 547 51 577 141
rect 625 115 655 141
rect 739 115 769 141
rect 857 115 887 141
rect 975 115 1005 141
rect 1093 115 1123 141
rect 1458 119 1488 141
rect 1381 103 1488 119
rect 1544 115 1574 141
rect 1656 115 1686 141
rect 1734 115 1764 141
rect 1381 69 1397 103
rect 1431 69 1488 103
rect 1381 51 1488 69
rect 1829 51 1859 66
rect 302 21 1859 51
rect 1926 40 1956 66
rect 1998 40 2028 66
<< polycont >>
rect 156 293 190 327
rect 156 225 190 259
rect 795 334 829 368
rect 641 263 675 297
rect 1366 334 1400 368
rect 903 263 937 297
rect 1672 337 1706 371
rect 1552 277 1586 311
rect 1780 337 1814 371
rect 1980 328 2014 362
rect 1980 260 2014 294
rect 1397 69 1431 103
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 23 571 89 587
rect 23 537 39 571
rect 73 537 89 571
rect 23 500 89 537
rect 23 466 39 500
rect 73 466 89 500
rect 23 429 89 466
rect 23 395 39 429
rect 73 395 89 429
rect 23 173 89 395
rect 129 571 195 649
rect 129 537 145 571
rect 179 537 195 571
rect 129 500 195 537
rect 129 466 145 500
rect 179 466 195 500
rect 129 429 195 466
rect 129 395 145 429
rect 179 395 195 429
rect 129 379 195 395
rect 241 597 307 613
rect 241 563 257 597
rect 291 563 307 597
rect 241 526 307 563
rect 241 492 257 526
rect 291 492 307 526
rect 241 455 307 492
rect 241 421 257 455
rect 291 421 307 455
rect 347 597 413 649
rect 347 563 363 597
rect 397 563 413 597
rect 347 499 413 563
rect 347 465 363 499
rect 397 465 413 499
rect 453 579 878 613
rect 453 568 519 579
rect 453 534 469 568
rect 503 534 519 568
rect 812 575 878 579
rect 453 489 519 534
rect 565 498 615 543
rect 347 449 413 465
rect 565 464 581 498
rect 565 453 615 464
rect 241 413 307 421
rect 449 419 615 453
rect 651 525 772 543
rect 651 491 722 525
rect 756 491 772 525
rect 812 541 828 575
rect 862 541 878 575
rect 812 503 878 541
rect 938 580 1004 649
rect 938 546 954 580
rect 988 546 1004 580
rect 938 503 1004 546
rect 1044 575 1110 613
rect 1044 541 1060 575
rect 1094 541 1110 575
rect 1150 607 1216 649
rect 1150 573 1166 607
rect 1200 573 1216 607
rect 1503 575 1569 613
rect 1044 537 1110 541
rect 1503 541 1519 575
rect 1553 541 1569 575
rect 1503 537 1569 541
rect 1044 503 1569 537
rect 1609 575 1675 613
rect 1609 541 1625 575
rect 1659 541 1675 575
rect 1609 537 1675 541
rect 1933 607 1983 649
rect 1967 573 1983 607
rect 1609 503 1897 537
rect 651 490 772 491
rect 449 413 483 419
rect 241 379 483 413
rect 651 383 685 490
rect 808 454 1827 467
rect 555 349 685 383
rect 721 433 1827 454
rect 721 420 842 433
rect 555 343 589 349
rect 140 327 589 343
rect 140 293 156 327
rect 190 309 589 327
rect 721 313 755 420
rect 878 384 1722 397
rect 791 371 1722 384
rect 791 368 1672 371
rect 791 334 795 368
rect 829 363 1366 368
rect 829 350 912 363
rect 829 334 845 350
rect 791 318 845 334
rect 1360 334 1366 363
rect 1400 363 1672 368
rect 1400 334 1416 363
rect 190 293 206 309
rect 140 259 206 293
rect 140 225 156 259
rect 190 225 206 259
rect 140 209 206 225
rect 281 239 519 273
rect 281 173 315 239
rect 23 144 109 173
rect 23 110 59 144
rect 93 110 109 144
rect 23 81 109 110
rect 201 144 315 173
rect 201 110 217 144
rect 251 110 315 144
rect 201 17 315 110
rect 351 187 417 203
rect 351 153 367 187
rect 401 153 417 187
rect 351 98 417 153
rect 453 200 519 239
rect 453 166 469 200
rect 503 166 519 200
rect 555 211 589 309
rect 625 297 755 313
rect 625 263 641 297
rect 675 281 755 297
rect 887 297 942 313
rect 887 281 903 297
rect 675 263 903 281
rect 937 263 942 297
rect 625 247 942 263
rect 887 236 942 247
rect 978 293 1324 327
rect 1360 310 1416 334
rect 1656 337 1672 363
rect 1706 337 1722 371
rect 1452 311 1602 327
rect 1656 321 1722 337
rect 1764 371 1827 433
rect 1764 337 1780 371
rect 1814 337 1827 371
rect 1764 321 1827 337
rect 555 200 721 211
rect 978 200 1012 293
rect 1290 274 1324 293
rect 1452 277 1552 311
rect 1586 277 1602 311
rect 1863 278 1897 503
rect 1933 536 1983 573
rect 1967 502 1983 536
rect 1933 465 1983 502
rect 1967 431 1983 465
rect 1933 415 1983 431
rect 2023 597 2094 613
rect 2023 563 2039 597
rect 2073 563 2094 597
rect 2023 465 2094 563
rect 2023 431 2039 465
rect 2073 431 2094 465
rect 2023 415 2094 431
rect 1964 362 2024 378
rect 1964 328 1980 362
rect 2014 328 2024 362
rect 1964 294 2024 328
rect 1964 278 1980 294
rect 1452 274 1602 277
rect 1290 261 1602 274
rect 555 191 1012 200
rect 555 166 666 191
rect 453 137 519 166
rect 650 157 666 166
rect 700 166 1012 191
rect 1048 223 1254 257
rect 1290 240 1486 261
rect 1638 260 1980 278
rect 2014 260 2024 294
rect 1638 244 2024 260
rect 1638 225 1672 244
rect 700 157 716 166
rect 650 137 716 157
rect 1048 130 1082 223
rect 1220 204 1254 223
rect 1220 187 1549 204
rect 780 114 846 130
rect 780 98 796 114
rect 351 80 796 98
rect 830 80 846 114
rect 351 64 846 80
rect 898 114 964 130
rect 898 80 914 114
rect 948 80 964 114
rect 898 17 964 80
rect 1016 114 1082 130
rect 1016 80 1032 114
rect 1066 80 1082 114
rect 1016 64 1082 80
rect 1118 153 1134 187
rect 1168 153 1184 187
rect 1220 170 1499 187
rect 1118 17 1184 153
rect 1483 153 1499 170
rect 1533 153 1549 187
rect 1483 137 1549 153
rect 1595 198 1672 225
rect 2060 208 2094 415
rect 1595 164 1611 198
rect 1645 164 1672 198
rect 1595 137 1672 164
rect 1273 103 1447 134
rect 1273 88 1397 103
rect 1381 69 1397 88
rect 1431 69 1447 103
rect 1381 53 1447 69
rect 1854 125 1920 154
rect 1854 91 1870 125
rect 1904 91 1920 125
rect 1854 17 1920 91
rect 2023 125 2094 208
rect 2023 91 2039 125
rect 2073 91 2094 125
rect 2023 62 2094 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 fa_lp
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 CIN
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1279 94 1313 128 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1375 94 1409 128 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 2047 94 2081 128 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 2047 168 2081 202 0 FreeSans 340 0 0 0 SUM
port 9 nsew signal output
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 COUT
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2408608
string GDS_START 2395050
<< end >>
