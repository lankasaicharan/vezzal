magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3506 1975
<< nwell >>
rect -38 331 2246 704
rect 476 305 1400 331
<< pwell >>
rect 431 185 1591 235
rect 1941 185 2207 202
rect 431 167 2207 185
rect 1 49 2207 167
rect 0 0 2208 49
<< scnmos >>
rect 82 57 112 141
rect 154 57 184 141
rect 240 57 270 141
rect 312 57 342 141
rect 513 125 543 209
rect 599 125 629 209
rect 717 79 747 163
rect 872 125 902 209
rect 1005 125 1035 209
rect 1325 125 1355 209
rect 1397 125 1427 209
rect 1485 125 1515 209
rect 1596 75 1626 159
rect 1668 75 1698 159
rect 1754 75 1784 159
rect 1826 75 1856 159
rect 2024 92 2054 176
rect 2096 92 2126 176
<< scpmoshvt >>
rect 107 409 157 609
rect 213 409 263 609
rect 585 341 635 541
rect 774 341 824 541
rect 912 371 962 571
rect 1027 341 1077 541
rect 1241 341 1291 541
rect 1379 383 1429 583
rect 1485 383 1535 583
rect 1583 383 1633 583
rect 1817 383 1867 583
rect 2074 396 2124 596
<< ndiff >>
rect 27 116 82 141
rect 27 82 37 116
rect 71 82 82 116
rect 27 57 82 82
rect 112 57 154 141
rect 184 108 240 141
rect 184 74 195 108
rect 229 74 240 108
rect 184 57 240 74
rect 270 57 312 141
rect 342 116 397 141
rect 342 82 353 116
rect 387 82 397 116
rect 342 57 397 82
rect 457 176 513 209
rect 457 142 468 176
rect 502 142 513 176
rect 457 125 513 142
rect 543 125 599 209
rect 629 163 702 209
rect 804 163 872 209
rect 629 158 717 163
rect 629 125 656 158
rect 644 124 656 125
rect 690 124 717 158
rect 644 79 717 124
rect 747 131 872 163
rect 747 97 758 131
rect 792 125 872 131
rect 902 125 1005 209
rect 1035 125 1325 209
rect 1355 125 1397 209
rect 1427 181 1485 209
rect 1427 147 1439 181
rect 1473 147 1485 181
rect 1427 125 1485 147
rect 1515 159 1565 209
rect 1515 125 1596 159
rect 792 97 804 125
rect 1252 121 1310 125
rect 747 79 804 97
rect 1252 87 1264 121
rect 1298 87 1310 121
rect 1539 121 1596 125
rect 1252 75 1310 87
rect 1539 87 1551 121
rect 1585 87 1596 121
rect 1539 75 1596 87
rect 1626 75 1668 159
rect 1698 134 1754 159
rect 1698 100 1709 134
rect 1743 100 1754 134
rect 1698 75 1754 100
rect 1784 75 1826 159
rect 1856 125 1913 159
rect 1856 91 1867 125
rect 1901 91 1913 125
rect 1967 151 2024 176
rect 1967 117 1979 151
rect 2013 117 2024 151
rect 1967 92 2024 117
rect 2054 92 2096 176
rect 2126 151 2181 176
rect 2126 117 2137 151
rect 2171 117 2181 151
rect 2126 92 2181 117
rect 1856 75 1913 91
<< pdiff >>
rect 50 597 107 609
rect 50 563 62 597
rect 96 563 107 597
rect 50 526 107 563
rect 50 492 62 526
rect 96 492 107 526
rect 50 455 107 492
rect 50 421 62 455
rect 96 421 107 455
rect 50 409 107 421
rect 157 597 213 609
rect 157 563 168 597
rect 202 563 213 597
rect 157 526 213 563
rect 157 492 168 526
rect 202 492 213 526
rect 157 455 213 492
rect 157 421 168 455
rect 202 421 213 455
rect 157 409 213 421
rect 263 597 320 609
rect 263 563 274 597
rect 308 563 320 597
rect 263 526 320 563
rect 263 492 274 526
rect 308 492 320 526
rect 263 455 320 492
rect 263 421 274 455
rect 308 421 320 455
rect 263 409 320 421
rect 2017 584 2074 596
rect 1306 571 1379 583
rect 661 541 719 542
rect 839 559 912 571
rect 839 541 851 559
rect 512 529 585 541
rect 512 495 524 529
rect 558 495 585 529
rect 512 456 585 495
rect 512 422 524 456
rect 558 422 585 456
rect 512 341 585 422
rect 635 530 774 541
rect 635 496 673 530
rect 707 496 774 530
rect 635 395 774 496
rect 635 361 673 395
rect 707 361 774 395
rect 635 341 774 361
rect 824 525 851 541
rect 885 525 912 559
rect 824 473 912 525
rect 824 439 851 473
rect 885 439 912 473
rect 824 387 912 439
rect 824 353 851 387
rect 885 371 912 387
rect 962 541 1012 571
rect 1306 541 1318 571
rect 962 371 1027 541
rect 885 353 897 371
rect 824 341 897 353
rect 977 341 1027 371
rect 1077 497 1241 541
rect 1077 463 1088 497
rect 1122 463 1241 497
rect 1077 341 1241 463
rect 1291 537 1318 541
rect 1352 537 1379 571
rect 1291 479 1379 537
rect 1291 445 1318 479
rect 1352 445 1379 479
rect 1291 387 1379 445
rect 1291 353 1318 387
rect 1352 383 1379 387
rect 1429 571 1485 583
rect 1429 537 1440 571
rect 1474 537 1485 571
rect 1429 465 1485 537
rect 1429 431 1440 465
rect 1474 431 1485 465
rect 1429 383 1485 431
rect 1535 383 1583 583
rect 1633 571 1817 583
rect 1633 537 1723 571
rect 1757 537 1817 571
rect 1633 471 1817 537
rect 1633 437 1723 471
rect 1757 437 1817 471
rect 1633 383 1817 437
rect 1867 571 1940 583
rect 1867 537 1894 571
rect 1928 537 1940 571
rect 1867 500 1940 537
rect 1867 466 1894 500
rect 1928 466 1940 500
rect 1867 429 1940 466
rect 1867 395 1894 429
rect 1928 395 1940 429
rect 2017 550 2029 584
rect 2063 550 2074 584
rect 2017 513 2074 550
rect 2017 479 2029 513
rect 2063 479 2074 513
rect 2017 442 2074 479
rect 2017 408 2029 442
rect 2063 408 2074 442
rect 2017 396 2074 408
rect 2124 584 2181 596
rect 2124 550 2135 584
rect 2169 550 2181 584
rect 2124 513 2181 550
rect 2124 479 2135 513
rect 2169 479 2181 513
rect 2124 442 2181 479
rect 2124 408 2135 442
rect 2169 408 2181 442
rect 2124 396 2181 408
rect 1867 383 1940 395
rect 1352 353 1364 383
rect 1291 341 1364 353
<< ndiffc >>
rect 37 82 71 116
rect 195 74 229 108
rect 353 82 387 116
rect 468 142 502 176
rect 656 124 690 158
rect 758 97 792 131
rect 1439 147 1473 181
rect 1264 87 1298 121
rect 1551 87 1585 121
rect 1709 100 1743 134
rect 1867 91 1901 125
rect 1979 117 2013 151
rect 2137 117 2171 151
<< pdiffc >>
rect 62 563 96 597
rect 62 492 96 526
rect 62 421 96 455
rect 168 563 202 597
rect 168 492 202 526
rect 168 421 202 455
rect 274 563 308 597
rect 274 492 308 526
rect 274 421 308 455
rect 524 495 558 529
rect 524 422 558 456
rect 673 496 707 530
rect 673 361 707 395
rect 851 525 885 559
rect 851 439 885 473
rect 851 353 885 387
rect 1088 463 1122 497
rect 1318 537 1352 571
rect 1318 445 1352 479
rect 1318 353 1352 387
rect 1440 537 1474 571
rect 1440 431 1474 465
rect 1723 537 1757 571
rect 1723 437 1757 471
rect 1894 537 1928 571
rect 1894 466 1928 500
rect 1894 395 1928 429
rect 2029 550 2063 584
rect 2029 479 2063 513
rect 2029 408 2063 442
rect 2135 550 2169 584
rect 2135 479 2169 513
rect 2135 408 2169 442
<< poly >>
rect 107 609 157 635
rect 213 609 263 635
rect 399 615 1429 645
rect 107 369 157 409
rect 82 353 157 369
rect 82 319 107 353
rect 141 319 157 353
rect 82 285 157 319
rect 213 313 263 409
rect 82 251 107 285
rect 141 265 157 285
rect 233 299 263 313
rect 233 283 299 299
rect 141 251 184 265
rect 82 235 184 251
rect 82 141 112 235
rect 154 141 184 235
rect 233 249 249 283
rect 283 249 299 283
rect 233 215 299 249
rect 233 181 249 215
rect 283 186 299 215
rect 399 186 429 615
rect 912 571 962 615
rect 1379 583 1429 615
rect 1485 583 1535 609
rect 1583 583 1633 609
rect 1817 583 1867 609
rect 2074 596 2124 622
rect 585 541 635 567
rect 774 541 824 567
rect 1027 541 1077 567
rect 1241 541 1291 567
rect 912 345 962 371
rect 1379 357 1429 383
rect 1485 357 1535 383
rect 477 284 543 300
rect 477 250 493 284
rect 527 264 543 284
rect 585 264 635 341
rect 774 315 824 341
rect 774 309 804 315
rect 677 293 804 309
rect 1027 297 1077 341
rect 1241 309 1291 341
rect 1505 309 1535 357
rect 527 250 629 264
rect 477 234 629 250
rect 677 259 693 293
rect 727 267 804 293
rect 872 281 957 297
rect 872 267 907 281
rect 727 259 907 267
rect 677 247 907 259
rect 941 247 957 281
rect 677 237 957 247
rect 513 209 543 234
rect 599 209 629 234
rect 872 231 957 237
rect 1005 281 1101 297
rect 1005 247 1051 281
rect 1085 247 1101 281
rect 1005 231 1101 247
rect 1200 293 1355 309
rect 1200 259 1216 293
rect 1250 273 1355 293
rect 1469 293 1535 309
rect 1250 259 1427 273
rect 1200 243 1427 259
rect 1469 259 1485 293
rect 1519 259 1535 293
rect 1583 351 1633 383
rect 1583 335 1769 351
rect 1583 301 1719 335
rect 1753 301 1769 335
rect 1817 315 1867 383
rect 2074 351 2124 396
rect 2017 335 2124 351
rect 1583 285 1769 301
rect 1811 299 1877 315
rect 1469 243 1535 259
rect 872 209 902 231
rect 1005 209 1035 231
rect 1325 209 1355 243
rect 1397 209 1427 243
rect 1485 209 1515 243
rect 283 181 442 186
rect 233 156 442 181
rect 240 141 270 156
rect 312 141 342 156
rect 82 31 112 57
rect 154 31 184 57
rect 240 31 270 57
rect 312 31 342 57
rect 412 51 442 156
rect 717 163 747 189
rect 513 99 543 125
rect 599 99 629 125
rect 1596 159 1626 185
rect 1668 159 1698 285
rect 1811 265 1827 299
rect 1861 265 1877 299
rect 1811 231 1877 265
rect 1811 211 1827 231
rect 1754 197 1827 211
rect 1861 197 1877 231
rect 2017 301 2033 335
rect 2067 301 2124 335
rect 2017 267 2124 301
rect 2017 233 2033 267
rect 2067 247 2124 267
rect 2067 233 2126 247
rect 2017 217 2126 233
rect 1754 181 1877 197
rect 1754 159 1784 181
rect 1826 159 1856 181
rect 2024 176 2054 217
rect 2096 176 2126 217
rect 872 99 902 125
rect 1005 99 1035 125
rect 1325 99 1355 125
rect 1397 99 1427 125
rect 1485 99 1515 125
rect 717 51 747 79
rect 1596 51 1626 75
rect 412 21 1626 51
rect 1668 49 1698 75
rect 1754 49 1784 75
rect 1826 49 1856 75
rect 2024 66 2054 92
rect 2096 66 2126 92
<< polycont >>
rect 107 319 141 353
rect 107 251 141 285
rect 249 249 283 283
rect 249 181 283 215
rect 493 250 527 284
rect 693 259 727 293
rect 907 247 941 281
rect 1051 247 1085 281
rect 1216 259 1250 293
rect 1485 259 1519 293
rect 1719 301 1753 335
rect 1827 265 1861 299
rect 1827 197 1861 231
rect 2033 301 2067 335
rect 2033 233 2067 267
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 21 597 112 613
rect 21 563 62 597
rect 96 563 112 597
rect 21 526 112 563
rect 21 492 62 526
rect 96 492 112 526
rect 21 455 112 492
rect 21 421 62 455
rect 96 421 112 455
rect 21 405 112 421
rect 152 597 218 649
rect 152 563 168 597
rect 202 563 218 597
rect 152 526 218 563
rect 152 492 168 526
rect 202 492 218 526
rect 152 455 218 492
rect 152 421 168 455
rect 202 421 218 455
rect 152 405 218 421
rect 258 597 369 613
rect 258 563 274 597
rect 308 563 369 597
rect 258 526 369 563
rect 258 492 274 526
rect 308 492 369 526
rect 258 455 369 492
rect 258 421 274 455
rect 308 421 369 455
rect 258 405 369 421
rect 508 529 574 649
rect 835 559 901 575
rect 508 495 524 529
rect 558 495 574 529
rect 508 456 574 495
rect 508 422 524 456
rect 558 422 574 456
rect 508 406 574 422
rect 657 530 723 546
rect 657 496 673 530
rect 707 496 723 530
rect 21 199 55 405
rect 335 370 369 405
rect 657 395 723 496
rect 91 353 167 369
rect 91 319 107 353
rect 141 319 167 353
rect 91 285 167 319
rect 335 336 621 370
rect 657 361 673 395
rect 707 379 723 395
rect 835 525 851 559
rect 885 525 901 559
rect 835 473 901 525
rect 835 439 851 473
rect 885 439 901 473
rect 835 387 901 439
rect 1072 497 1138 649
rect 1072 463 1088 497
rect 1122 463 1138 497
rect 1072 415 1138 463
rect 1302 571 1368 587
rect 1302 537 1318 571
rect 1352 537 1368 571
rect 1302 479 1368 537
rect 1302 445 1318 479
rect 1352 445 1368 479
rect 707 361 799 379
rect 657 345 799 361
rect 91 251 107 285
rect 141 251 167 285
rect 91 235 167 251
rect 233 283 299 299
rect 233 249 249 283
rect 283 249 299 283
rect 233 215 299 249
rect 233 199 249 215
rect 21 181 249 199
rect 283 181 299 215
rect 21 165 299 181
rect 21 116 87 165
rect 335 145 369 336
rect 587 309 621 336
rect 409 284 551 300
rect 409 250 493 284
rect 527 250 551 284
rect 409 234 551 250
rect 587 293 729 309
rect 587 259 693 293
rect 727 259 729 293
rect 587 243 729 259
rect 765 207 799 345
rect 452 176 518 198
rect 21 82 37 116
rect 71 82 87 116
rect 21 53 87 82
rect 179 108 245 129
rect 179 74 195 108
rect 229 74 245 108
rect 179 17 245 74
rect 335 116 403 145
rect 335 82 353 116
rect 387 82 403 116
rect 335 53 403 82
rect 452 142 468 176
rect 502 142 518 176
rect 452 17 518 142
rect 640 173 799 207
rect 835 353 851 387
rect 885 371 901 387
rect 1302 387 1368 445
rect 1424 571 1490 587
rect 1424 537 1440 571
rect 1474 537 1490 571
rect 1424 465 1490 537
rect 1424 431 1440 465
rect 1474 449 1490 465
rect 1707 571 1773 649
rect 1707 537 1723 571
rect 1757 537 1773 571
rect 1707 471 1773 537
rect 1474 431 1671 449
rect 1424 415 1671 431
rect 1707 437 1723 471
rect 1757 437 1773 471
rect 1707 421 1773 437
rect 1878 571 1944 587
rect 1878 537 1894 571
rect 1928 537 1944 571
rect 1878 500 1944 537
rect 1878 466 1894 500
rect 1928 466 1944 500
rect 1878 429 1944 466
rect 1302 379 1318 387
rect 885 353 1013 371
rect 835 337 1013 353
rect 640 158 706 173
rect 640 124 656 158
rect 690 124 706 158
rect 835 137 869 337
rect 640 75 706 124
rect 742 131 869 137
rect 742 97 758 131
rect 792 97 869 131
rect 742 75 869 97
rect 905 281 943 297
rect 905 247 907 281
rect 941 247 943 281
rect 905 125 943 247
rect 979 195 1013 337
rect 1049 353 1318 379
rect 1352 379 1368 387
rect 1352 353 1601 379
rect 1049 345 1601 353
rect 1049 281 1088 345
rect 1302 337 1368 345
rect 1049 247 1051 281
rect 1085 247 1088 281
rect 1049 231 1088 247
rect 1124 293 1266 309
rect 1124 259 1216 293
rect 1250 259 1266 293
rect 1469 293 1531 309
rect 1469 277 1485 293
rect 1124 243 1266 259
rect 1302 259 1485 277
rect 1519 259 1531 293
rect 1302 243 1531 259
rect 1124 195 1158 243
rect 1302 207 1336 243
rect 1567 207 1601 345
rect 979 161 1158 195
rect 1194 173 1336 207
rect 1423 181 1601 207
rect 1194 125 1228 173
rect 1423 147 1439 181
rect 1473 173 1601 181
rect 1637 233 1671 415
rect 1878 395 1894 429
rect 1928 395 1944 429
rect 1878 385 1944 395
rect 2013 584 2079 649
rect 2013 550 2029 584
rect 2063 550 2079 584
rect 2013 513 2079 550
rect 2013 479 2029 513
rect 2063 479 2079 513
rect 2013 442 2079 479
rect 2013 408 2029 442
rect 2063 408 2079 442
rect 2013 392 2079 408
rect 2119 584 2185 600
rect 2119 550 2135 584
rect 2169 550 2185 584
rect 2119 513 2185 550
rect 2119 479 2135 513
rect 2169 479 2185 513
rect 2119 442 2185 479
rect 2119 408 2135 442
rect 2169 408 2185 442
rect 1707 351 1944 385
rect 2119 356 2185 408
rect 1707 335 1769 351
rect 1707 301 1719 335
rect 1753 301 1769 335
rect 1909 335 2083 351
rect 1909 317 2033 335
rect 1707 285 1769 301
rect 1811 299 1873 315
rect 1811 265 1827 299
rect 1861 265 1873 299
rect 1811 233 1873 265
rect 1637 231 1873 233
rect 1637 199 1827 231
rect 1473 147 1489 173
rect 905 91 1228 125
rect 1264 121 1314 137
rect 1423 121 1489 147
rect 1637 137 1671 199
rect 1811 197 1827 199
rect 1861 197 1873 231
rect 1811 181 1873 197
rect 1535 121 1671 137
rect 1298 87 1314 121
rect 1264 17 1314 87
rect 1535 87 1551 121
rect 1585 87 1671 121
rect 1535 71 1671 87
rect 1709 134 1759 163
rect 1909 145 1943 317
rect 2017 301 2033 317
rect 2067 301 2083 335
rect 2017 267 2083 301
rect 2017 233 2033 267
rect 2067 233 2083 267
rect 2017 217 2083 233
rect 1743 100 1759 134
rect 1709 17 1759 100
rect 1851 125 1943 145
rect 1851 91 1867 125
rect 1901 91 1943 125
rect 1851 71 1943 91
rect 1979 151 2029 180
rect 2013 117 2029 151
rect 1979 17 2029 117
rect 2119 151 2187 356
rect 2119 117 2137 151
rect 2171 117 2187 151
rect 2119 88 2187 117
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfxtp_lp
flabel comment s 814 261 814 261 0 FreeSans 200 180 0 0 no_jumper_check
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2143 94 2177 128 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2143 168 2177 202 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2143 242 2177 276 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 2143 316 2177 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 846998
string GDS_START 832924
<< end >>
