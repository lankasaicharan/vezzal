magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 1 49 419 203
rect 0 0 576 49
<< scnmos >>
rect 80 67 110 177
rect 152 67 182 177
rect 238 67 268 177
rect 310 67 340 177
<< scpmoshvt >>
rect 80 396 130 596
rect 186 396 236 596
rect 292 396 342 596
rect 398 396 448 596
<< ndiff >>
rect 27 139 80 177
rect 27 105 35 139
rect 69 105 80 139
rect 27 67 80 105
rect 110 67 152 177
rect 182 126 238 177
rect 182 92 193 126
rect 227 92 238 126
rect 182 67 238 92
rect 268 67 310 177
rect 340 139 393 177
rect 340 105 351 139
rect 385 105 393 139
rect 340 67 393 105
<< pdiff >>
rect 27 584 80 596
rect 27 550 35 584
rect 69 550 80 584
rect 27 513 80 550
rect 27 479 35 513
rect 69 479 80 513
rect 27 442 80 479
rect 27 408 35 442
rect 69 408 80 442
rect 27 396 80 408
rect 130 584 186 596
rect 130 550 141 584
rect 175 550 186 584
rect 130 513 186 550
rect 130 479 141 513
rect 175 479 186 513
rect 130 442 186 479
rect 130 408 141 442
rect 175 408 186 442
rect 130 396 186 408
rect 236 584 292 596
rect 236 550 247 584
rect 281 550 292 584
rect 236 513 292 550
rect 236 479 247 513
rect 281 479 292 513
rect 236 442 292 479
rect 236 408 247 442
rect 281 408 292 442
rect 236 396 292 408
rect 342 584 398 596
rect 342 550 353 584
rect 387 550 398 584
rect 342 513 398 550
rect 342 479 353 513
rect 387 479 398 513
rect 342 442 398 479
rect 342 408 353 442
rect 387 408 398 442
rect 342 396 398 408
rect 448 584 501 596
rect 448 550 459 584
rect 493 550 501 584
rect 448 513 501 550
rect 448 479 459 513
rect 493 479 501 513
rect 448 442 501 479
rect 448 408 459 442
rect 493 408 501 442
rect 448 396 501 408
<< ndiffc >>
rect 35 105 69 139
rect 193 92 227 126
rect 351 105 385 139
<< pdiffc >>
rect 35 550 69 584
rect 35 479 69 513
rect 35 408 69 442
rect 141 550 175 584
rect 141 479 175 513
rect 141 408 175 442
rect 247 550 281 584
rect 247 479 281 513
rect 247 408 281 442
rect 353 550 387 584
rect 353 479 387 513
rect 353 408 387 442
rect 459 550 493 584
rect 459 479 493 513
rect 459 408 493 442
<< poly >>
rect 80 596 130 622
rect 186 596 236 622
rect 292 596 342 622
rect 398 596 448 622
rect 80 316 130 396
rect 31 313 130 316
rect 186 313 236 396
rect 292 313 342 396
rect 398 313 448 396
rect 31 300 448 313
rect 31 266 47 300
rect 81 266 448 300
rect 31 250 448 266
rect 80 247 448 250
rect 80 177 110 247
rect 152 177 182 247
rect 238 177 268 247
rect 310 177 340 247
rect 80 41 110 67
rect 152 41 182 67
rect 238 41 268 67
rect 310 41 340 67
<< polycont >>
rect 47 266 81 300
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 19 584 85 649
rect 19 550 35 584
rect 69 550 85 584
rect 19 513 85 550
rect 19 479 35 513
rect 69 479 85 513
rect 19 442 85 479
rect 19 408 35 442
rect 69 408 85 442
rect 19 392 85 408
rect 125 584 191 600
rect 125 550 141 584
rect 175 550 191 584
rect 125 513 191 550
rect 125 479 141 513
rect 175 479 191 513
rect 125 442 191 479
rect 125 408 141 442
rect 175 408 191 442
rect 20 300 91 356
rect 20 266 47 300
rect 81 266 91 300
rect 20 221 91 266
rect 125 313 191 408
rect 231 584 297 649
rect 231 550 247 584
rect 281 550 297 584
rect 231 513 297 550
rect 231 479 247 513
rect 281 479 297 513
rect 231 442 297 479
rect 231 408 247 442
rect 281 408 297 442
rect 231 392 297 408
rect 337 584 403 600
rect 337 550 353 584
rect 387 550 403 584
rect 337 513 403 550
rect 337 479 353 513
rect 387 479 403 513
rect 337 442 403 479
rect 337 408 353 442
rect 387 408 403 442
rect 337 313 403 408
rect 443 584 509 649
rect 443 550 459 584
rect 493 550 509 584
rect 443 513 509 550
rect 443 479 459 513
rect 493 479 509 513
rect 443 442 509 479
rect 443 408 459 442
rect 493 408 509 442
rect 443 392 509 408
rect 125 247 403 313
rect 125 156 191 247
rect 19 139 85 155
rect 19 105 35 139
rect 69 105 85 139
rect 19 17 85 105
rect 125 126 243 156
rect 125 92 193 126
rect 227 92 243 126
rect 125 63 243 92
rect 335 139 401 155
rect 335 105 351 139
rect 385 105 401 139
rect 335 17 401 105
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkinvlp_4
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2230934
string GDS_START 2225862
<< end >>
