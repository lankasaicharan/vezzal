magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3122 1975
<< nwell >>
rect -38 331 1862 704
<< pwell >>
rect 999 245 1813 259
rect 1 49 1813 245
rect 0 0 1824 49
<< scnmos >>
rect 80 51 110 219
rect 270 51 300 219
rect 356 51 386 219
rect 442 51 472 219
rect 528 51 558 219
rect 614 51 644 219
rect 716 51 746 219
rect 802 51 832 219
rect 888 51 918 219
rect 1082 65 1112 233
rect 1168 65 1198 233
rect 1254 65 1284 233
rect 1356 65 1386 233
rect 1442 65 1472 233
rect 1528 65 1558 233
rect 1614 65 1644 233
rect 1700 65 1730 233
<< scpmoshvt >>
rect 150 367 180 619
rect 238 367 268 619
rect 324 367 354 619
rect 426 367 456 619
rect 512 367 542 619
rect 602 367 632 619
rect 688 367 718 619
rect 774 367 804 619
rect 860 367 890 619
rect 1014 367 1044 619
rect 1100 367 1130 619
rect 1186 367 1216 619
rect 1272 367 1302 619
rect 1432 367 1462 619
rect 1518 367 1548 619
rect 1604 367 1634 619
rect 1690 367 1720 619
<< ndiff >>
rect 27 207 80 219
rect 27 173 35 207
rect 69 173 80 207
rect 27 101 80 173
rect 27 67 35 101
rect 69 67 80 101
rect 27 51 80 67
rect 110 171 163 219
rect 110 137 121 171
rect 155 137 163 171
rect 110 97 163 137
rect 110 63 121 97
rect 155 63 163 97
rect 110 51 163 63
rect 217 207 270 219
rect 217 173 225 207
rect 259 173 270 207
rect 217 97 270 173
rect 217 63 225 97
rect 259 63 270 97
rect 217 51 270 63
rect 300 169 356 219
rect 300 135 311 169
rect 345 135 356 169
rect 300 51 356 135
rect 386 179 442 219
rect 386 145 397 179
rect 431 145 442 179
rect 386 97 442 145
rect 386 63 397 97
rect 431 63 442 97
rect 386 51 442 63
rect 472 169 528 219
rect 472 135 483 169
rect 517 135 528 169
rect 472 51 528 135
rect 558 179 614 219
rect 558 145 569 179
rect 603 145 614 179
rect 558 97 614 145
rect 558 63 569 97
rect 603 63 614 97
rect 558 51 614 63
rect 644 175 716 219
rect 644 141 671 175
rect 705 141 716 175
rect 644 51 716 141
rect 746 97 802 219
rect 746 63 757 97
rect 791 63 802 97
rect 746 51 802 63
rect 832 175 888 219
rect 832 141 843 175
rect 877 141 888 175
rect 832 51 888 141
rect 918 97 971 219
rect 918 63 929 97
rect 963 63 971 97
rect 1025 107 1082 233
rect 1025 73 1037 107
rect 1071 73 1082 107
rect 1025 65 1082 73
rect 1112 195 1168 233
rect 1112 161 1123 195
rect 1157 161 1168 195
rect 1112 65 1168 161
rect 1198 181 1254 233
rect 1198 147 1209 181
rect 1243 147 1254 181
rect 1198 107 1254 147
rect 1198 73 1209 107
rect 1243 73 1254 107
rect 1198 65 1254 73
rect 1284 225 1356 233
rect 1284 191 1311 225
rect 1345 191 1356 225
rect 1284 155 1356 191
rect 1284 121 1311 155
rect 1345 121 1356 155
rect 1284 65 1356 121
rect 1386 225 1442 233
rect 1386 191 1397 225
rect 1431 191 1442 225
rect 1386 111 1442 191
rect 1386 77 1397 111
rect 1431 77 1442 111
rect 1386 65 1442 77
rect 1472 179 1528 233
rect 1472 145 1483 179
rect 1517 145 1528 179
rect 1472 107 1528 145
rect 1472 73 1483 107
rect 1517 73 1528 107
rect 1472 65 1528 73
rect 1558 221 1614 233
rect 1558 187 1569 221
rect 1603 187 1614 221
rect 1558 111 1614 187
rect 1558 77 1569 111
rect 1603 77 1614 111
rect 1558 65 1614 77
rect 1644 175 1700 233
rect 1644 141 1655 175
rect 1689 141 1700 175
rect 1644 107 1700 141
rect 1644 73 1655 107
rect 1689 73 1700 107
rect 1644 65 1700 73
rect 1730 221 1787 233
rect 1730 187 1741 221
rect 1775 187 1787 221
rect 1730 111 1787 187
rect 1730 77 1741 111
rect 1775 77 1787 111
rect 1730 65 1787 77
rect 918 51 971 63
<< pdiff >>
rect 97 599 150 619
rect 97 565 105 599
rect 139 565 150 599
rect 97 515 150 565
rect 97 481 105 515
rect 139 481 150 515
rect 97 436 150 481
rect 97 402 105 436
rect 139 402 150 436
rect 97 367 150 402
rect 180 607 238 619
rect 180 573 193 607
rect 227 573 238 607
rect 180 511 238 573
rect 180 477 193 511
rect 227 477 238 511
rect 180 413 238 477
rect 180 379 193 413
rect 227 379 238 413
rect 180 367 238 379
rect 268 599 324 619
rect 268 565 279 599
rect 313 565 324 599
rect 268 509 324 565
rect 268 475 279 509
rect 313 475 324 509
rect 268 413 324 475
rect 268 379 279 413
rect 313 379 324 413
rect 268 367 324 379
rect 354 611 426 619
rect 354 577 373 611
rect 407 577 426 611
rect 354 537 426 577
rect 354 503 373 537
rect 407 503 426 537
rect 354 459 426 503
rect 354 425 373 459
rect 407 425 426 459
rect 354 367 426 425
rect 456 599 512 619
rect 456 565 467 599
rect 501 565 512 599
rect 456 509 512 565
rect 456 475 467 509
rect 501 475 512 509
rect 456 413 512 475
rect 456 379 467 413
rect 501 379 512 413
rect 456 367 512 379
rect 542 611 602 619
rect 542 577 553 611
rect 587 577 602 611
rect 542 537 602 577
rect 542 503 553 537
rect 587 503 602 537
rect 542 457 602 503
rect 542 423 553 457
rect 587 423 602 457
rect 542 367 602 423
rect 632 599 688 619
rect 632 565 643 599
rect 677 565 688 599
rect 632 509 688 565
rect 632 475 643 509
rect 677 475 688 509
rect 632 413 688 475
rect 632 379 643 413
rect 677 379 688 413
rect 632 367 688 379
rect 718 607 774 619
rect 718 573 729 607
rect 763 573 774 607
rect 718 492 774 573
rect 718 458 729 492
rect 763 458 774 492
rect 718 367 774 458
rect 804 599 860 619
rect 804 565 815 599
rect 849 565 860 599
rect 804 514 860 565
rect 804 480 815 514
rect 849 480 860 514
rect 804 440 860 480
rect 804 406 815 440
rect 849 406 860 440
rect 804 367 860 406
rect 890 607 1014 619
rect 890 573 901 607
rect 935 573 969 607
rect 1003 573 1014 607
rect 890 492 1014 573
rect 890 458 901 492
rect 935 458 969 492
rect 1003 458 1014 492
rect 890 367 1014 458
rect 1044 599 1100 619
rect 1044 565 1055 599
rect 1089 565 1100 599
rect 1044 514 1100 565
rect 1044 480 1055 514
rect 1089 480 1100 514
rect 1044 440 1100 480
rect 1044 406 1055 440
rect 1089 406 1100 440
rect 1044 367 1100 406
rect 1130 607 1186 619
rect 1130 573 1141 607
rect 1175 573 1186 607
rect 1130 492 1186 573
rect 1130 458 1141 492
rect 1175 458 1186 492
rect 1130 367 1186 458
rect 1216 599 1272 619
rect 1216 565 1227 599
rect 1261 565 1272 599
rect 1216 512 1272 565
rect 1216 478 1227 512
rect 1261 478 1272 512
rect 1216 424 1272 478
rect 1216 390 1227 424
rect 1261 390 1272 424
rect 1216 367 1272 390
rect 1302 611 1432 619
rect 1302 577 1319 611
rect 1353 577 1387 611
rect 1421 577 1432 611
rect 1302 543 1432 577
rect 1302 509 1319 543
rect 1353 536 1432 543
rect 1353 509 1387 536
rect 1302 502 1387 509
rect 1421 502 1432 536
rect 1302 471 1432 502
rect 1302 437 1319 471
rect 1353 455 1432 471
rect 1353 437 1387 455
rect 1302 421 1387 437
rect 1421 421 1432 455
rect 1302 367 1432 421
rect 1462 599 1518 619
rect 1462 565 1473 599
rect 1507 565 1518 599
rect 1462 507 1518 565
rect 1462 473 1473 507
rect 1507 473 1518 507
rect 1462 413 1518 473
rect 1462 379 1473 413
rect 1507 379 1518 413
rect 1462 367 1518 379
rect 1548 607 1604 619
rect 1548 573 1559 607
rect 1593 573 1604 607
rect 1548 488 1604 573
rect 1548 454 1559 488
rect 1593 454 1604 488
rect 1548 367 1604 454
rect 1634 599 1690 619
rect 1634 565 1645 599
rect 1679 565 1690 599
rect 1634 512 1690 565
rect 1634 478 1645 512
rect 1679 478 1690 512
rect 1634 436 1690 478
rect 1634 402 1645 436
rect 1679 402 1690 436
rect 1634 367 1690 402
rect 1720 607 1773 619
rect 1720 573 1731 607
rect 1765 573 1773 607
rect 1720 510 1773 573
rect 1720 476 1731 510
rect 1765 476 1773 510
rect 1720 418 1773 476
rect 1720 384 1731 418
rect 1765 384 1773 418
rect 1720 367 1773 384
<< ndiffc >>
rect 35 173 69 207
rect 35 67 69 101
rect 121 137 155 171
rect 121 63 155 97
rect 225 173 259 207
rect 225 63 259 97
rect 311 135 345 169
rect 397 145 431 179
rect 397 63 431 97
rect 483 135 517 169
rect 569 145 603 179
rect 569 63 603 97
rect 671 141 705 175
rect 757 63 791 97
rect 843 141 877 175
rect 929 63 963 97
rect 1037 73 1071 107
rect 1123 161 1157 195
rect 1209 147 1243 181
rect 1209 73 1243 107
rect 1311 191 1345 225
rect 1311 121 1345 155
rect 1397 191 1431 225
rect 1397 77 1431 111
rect 1483 145 1517 179
rect 1483 73 1517 107
rect 1569 187 1603 221
rect 1569 77 1603 111
rect 1655 141 1689 175
rect 1655 73 1689 107
rect 1741 187 1775 221
rect 1741 77 1775 111
<< pdiffc >>
rect 105 565 139 599
rect 105 481 139 515
rect 105 402 139 436
rect 193 573 227 607
rect 193 477 227 511
rect 193 379 227 413
rect 279 565 313 599
rect 279 475 313 509
rect 279 379 313 413
rect 373 577 407 611
rect 373 503 407 537
rect 373 425 407 459
rect 467 565 501 599
rect 467 475 501 509
rect 467 379 501 413
rect 553 577 587 611
rect 553 503 587 537
rect 553 423 587 457
rect 643 565 677 599
rect 643 475 677 509
rect 643 379 677 413
rect 729 573 763 607
rect 729 458 763 492
rect 815 565 849 599
rect 815 480 849 514
rect 815 406 849 440
rect 901 573 935 607
rect 969 573 1003 607
rect 901 458 935 492
rect 969 458 1003 492
rect 1055 565 1089 599
rect 1055 480 1089 514
rect 1055 406 1089 440
rect 1141 573 1175 607
rect 1141 458 1175 492
rect 1227 565 1261 599
rect 1227 478 1261 512
rect 1227 390 1261 424
rect 1319 577 1353 611
rect 1387 577 1421 611
rect 1319 509 1353 543
rect 1387 502 1421 536
rect 1319 437 1353 471
rect 1387 421 1421 455
rect 1473 565 1507 599
rect 1473 473 1507 507
rect 1473 379 1507 413
rect 1559 573 1593 607
rect 1559 454 1593 488
rect 1645 565 1679 599
rect 1645 478 1679 512
rect 1645 402 1679 436
rect 1731 573 1765 607
rect 1731 476 1765 510
rect 1731 384 1765 418
<< poly >>
rect 150 619 180 645
rect 238 619 268 645
rect 324 619 354 645
rect 426 619 456 645
rect 512 619 542 645
rect 602 619 632 645
rect 688 619 718 645
rect 774 619 804 645
rect 860 619 890 645
rect 1014 619 1044 645
rect 1100 619 1130 645
rect 1186 619 1216 645
rect 1272 619 1302 645
rect 1432 619 1462 645
rect 1518 619 1548 645
rect 1604 619 1634 645
rect 1690 619 1720 645
rect 150 325 180 367
rect 238 335 268 367
rect 324 335 354 367
rect 426 335 456 367
rect 512 335 542 367
rect 602 335 632 367
rect 688 335 718 367
rect 774 335 804 367
rect 860 335 890 367
rect 1014 335 1044 367
rect 1100 335 1130 367
rect 1186 335 1216 367
rect 1272 335 1302 367
rect 1432 335 1462 367
rect 1518 335 1548 367
rect 1604 335 1634 367
rect 1690 335 1720 367
rect 21 309 180 325
rect 21 275 37 309
rect 71 275 180 309
rect 21 259 180 275
rect 222 319 560 335
rect 222 285 238 319
rect 272 285 306 319
rect 340 285 374 319
rect 408 285 442 319
rect 476 285 510 319
rect 544 285 560 319
rect 222 269 560 285
rect 602 319 940 335
rect 602 285 618 319
rect 652 285 686 319
rect 720 285 754 319
rect 788 285 822 319
rect 856 285 890 319
rect 924 285 940 319
rect 602 269 940 285
rect 1014 319 1386 335
rect 1014 285 1062 319
rect 1096 285 1130 319
rect 1164 285 1198 319
rect 1232 285 1266 319
rect 1300 285 1334 319
rect 1368 285 1386 319
rect 1432 319 1780 335
rect 1432 305 1458 319
rect 1014 269 1386 285
rect 80 219 110 259
rect 270 219 300 269
rect 356 219 386 269
rect 442 219 472 269
rect 528 219 558 269
rect 614 219 644 269
rect 716 219 746 269
rect 802 219 832 269
rect 888 219 918 269
rect 1082 233 1112 269
rect 1168 233 1198 269
rect 1254 233 1284 269
rect 1356 233 1386 269
rect 1442 285 1458 305
rect 1492 285 1526 319
rect 1560 285 1594 319
rect 1628 285 1662 319
rect 1696 285 1730 319
rect 1764 285 1780 319
rect 1442 269 1780 285
rect 1442 233 1472 269
rect 1528 233 1558 269
rect 1614 233 1644 269
rect 1700 233 1730 269
rect 80 25 110 51
rect 270 25 300 51
rect 356 25 386 51
rect 442 25 472 51
rect 528 25 558 51
rect 614 25 644 51
rect 716 25 746 51
rect 802 25 832 51
rect 888 25 918 51
rect 1082 39 1112 65
rect 1168 39 1198 65
rect 1254 39 1284 65
rect 1356 39 1386 65
rect 1442 39 1472 65
rect 1528 39 1558 65
rect 1614 39 1644 65
rect 1700 39 1730 65
<< polycont >>
rect 37 275 71 309
rect 238 285 272 319
rect 306 285 340 319
rect 374 285 408 319
rect 442 285 476 319
rect 510 285 544 319
rect 618 285 652 319
rect 686 285 720 319
rect 754 285 788 319
rect 822 285 856 319
rect 890 285 924 319
rect 1062 285 1096 319
rect 1130 285 1164 319
rect 1198 285 1232 319
rect 1266 285 1300 319
rect 1334 285 1368 319
rect 1458 285 1492 319
rect 1526 285 1560 319
rect 1594 285 1628 319
rect 1662 285 1696 319
rect 1730 285 1764 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 89 599 155 615
rect 89 565 105 599
rect 139 565 155 599
rect 89 515 155 565
rect 89 481 105 515
rect 139 481 155 515
rect 89 436 155 481
rect 89 402 105 436
rect 139 402 155 436
rect 89 386 155 402
rect 21 309 87 352
rect 21 275 37 309
rect 71 275 87 309
rect 21 273 87 275
rect 121 319 155 386
rect 189 607 235 649
rect 189 573 193 607
rect 227 573 235 607
rect 189 511 235 573
rect 189 477 193 511
rect 227 477 235 511
rect 189 413 235 477
rect 189 379 193 413
rect 227 379 235 413
rect 189 363 235 379
rect 269 599 323 615
rect 269 565 279 599
rect 313 565 323 599
rect 269 509 323 565
rect 269 475 279 509
rect 313 475 323 509
rect 269 413 323 475
rect 357 611 423 649
rect 357 577 373 611
rect 407 577 423 611
rect 357 537 423 577
rect 357 503 373 537
rect 407 503 423 537
rect 357 459 423 503
rect 357 425 373 459
rect 407 425 423 459
rect 457 599 503 615
rect 457 565 467 599
rect 501 565 503 599
rect 457 509 503 565
rect 457 475 467 509
rect 501 475 503 509
rect 269 379 279 413
rect 313 389 323 413
rect 457 413 503 475
rect 537 611 603 649
rect 537 577 553 611
rect 587 577 603 611
rect 537 537 603 577
rect 537 503 553 537
rect 587 503 603 537
rect 537 457 603 503
rect 537 423 553 457
rect 587 423 603 457
rect 637 599 679 615
rect 637 565 643 599
rect 677 565 679 599
rect 637 509 679 565
rect 637 475 643 509
rect 677 475 679 509
rect 637 424 679 475
rect 713 607 779 649
rect 713 573 729 607
rect 763 573 779 607
rect 713 492 779 573
rect 713 458 729 492
rect 763 458 779 492
rect 813 599 851 615
rect 813 565 815 599
rect 849 565 851 599
rect 813 514 851 565
rect 813 480 815 514
rect 849 480 851 514
rect 813 440 851 480
rect 885 607 1019 649
rect 885 573 901 607
rect 935 573 969 607
rect 1003 573 1019 607
rect 885 492 1019 573
rect 885 458 901 492
rect 935 458 969 492
rect 1003 458 1019 492
rect 1053 599 1091 615
rect 1053 565 1055 599
rect 1089 565 1091 599
rect 1053 514 1091 565
rect 1053 480 1055 514
rect 1089 480 1091 514
rect 813 424 815 440
rect 457 389 467 413
rect 313 379 467 389
rect 501 389 503 413
rect 637 413 815 424
rect 637 389 643 413
rect 501 379 643 389
rect 677 406 815 413
rect 849 424 851 440
rect 1053 440 1091 480
rect 1125 607 1191 649
rect 1125 573 1141 607
rect 1175 573 1191 607
rect 1125 492 1191 573
rect 1125 458 1141 492
rect 1175 458 1191 492
rect 1225 599 1285 615
rect 1225 565 1227 599
rect 1261 565 1285 599
rect 1225 512 1285 565
rect 1225 478 1227 512
rect 1261 478 1285 512
rect 1053 424 1055 440
rect 849 406 1055 424
rect 1089 424 1091 440
rect 1225 424 1285 478
rect 1089 406 1227 424
rect 677 390 1227 406
rect 1261 390 1285 424
rect 1319 611 1437 649
rect 1353 577 1387 611
rect 1421 577 1437 611
rect 1319 543 1437 577
rect 1353 536 1437 543
rect 1353 509 1387 536
rect 1319 502 1387 509
rect 1421 502 1437 536
rect 1319 471 1437 502
rect 1353 455 1437 471
rect 1353 437 1387 455
rect 1319 421 1387 437
rect 1421 421 1437 455
rect 1471 599 1507 615
rect 1471 565 1473 599
rect 1471 507 1507 565
rect 1471 473 1473 507
rect 677 379 734 390
rect 269 355 734 379
rect 976 387 1285 390
rect 1471 420 1507 473
rect 1543 607 1609 649
rect 1543 573 1559 607
rect 1593 573 1609 607
rect 1543 488 1609 573
rect 1543 454 1559 488
rect 1593 454 1609 488
rect 1643 599 1681 615
rect 1643 565 1645 599
rect 1679 565 1681 599
rect 1643 512 1681 565
rect 1643 478 1645 512
rect 1679 478 1681 512
rect 1643 436 1681 478
rect 1643 420 1645 436
rect 1471 413 1645 420
rect 1471 387 1473 413
rect 976 384 1473 387
rect 769 321 940 356
rect 602 319 940 321
rect 121 285 238 319
rect 272 285 306 319
rect 340 285 374 319
rect 408 285 442 319
rect 476 285 510 319
rect 544 285 560 319
rect 602 285 618 319
rect 652 285 686 319
rect 720 285 754 319
rect 788 285 822 319
rect 856 285 890 319
rect 924 285 940 319
rect 121 239 171 285
rect 976 251 1010 384
rect 1251 379 1473 384
rect 1507 402 1645 413
rect 1679 402 1681 436
rect 1507 386 1681 402
rect 1715 607 1781 649
rect 1715 573 1731 607
rect 1765 573 1781 607
rect 1715 510 1781 573
rect 1715 476 1731 510
rect 1765 476 1781 510
rect 1715 418 1781 476
rect 1507 379 1523 386
rect 1715 384 1731 418
rect 1765 384 1781 418
rect 1251 353 1523 379
rect 1046 319 1217 350
rect 1557 319 1804 350
rect 1046 285 1062 319
rect 1096 285 1130 319
rect 1164 285 1198 319
rect 1232 285 1266 319
rect 1300 285 1334 319
rect 1368 285 1384 319
rect 1442 285 1458 319
rect 1492 285 1526 319
rect 1560 285 1594 319
rect 1628 285 1662 319
rect 1696 285 1730 319
rect 1764 285 1804 319
rect 19 207 171 239
rect 19 173 35 207
rect 69 205 171 207
rect 209 207 268 223
rect 19 101 69 173
rect 209 173 225 207
rect 259 173 268 207
rect 19 67 35 101
rect 19 51 69 67
rect 105 137 121 171
rect 155 137 171 171
rect 105 97 171 137
rect 105 63 121 97
rect 155 63 171 97
rect 105 17 171 63
rect 209 97 268 173
rect 302 215 1010 251
rect 1106 225 1361 251
rect 1106 215 1311 225
rect 302 169 347 215
rect 302 135 311 169
rect 345 135 347 169
rect 302 119 347 135
rect 381 179 447 181
rect 381 145 397 179
rect 431 145 447 179
rect 209 63 225 97
rect 259 85 268 97
rect 381 97 447 145
rect 481 169 519 215
rect 1106 195 1159 215
rect 1106 181 1123 195
rect 481 135 483 169
rect 517 135 519 169
rect 481 119 519 135
rect 553 179 619 181
rect 553 145 569 179
rect 603 145 619 179
rect 381 85 397 97
rect 259 63 397 85
rect 431 85 447 97
rect 553 103 619 145
rect 655 175 1123 181
rect 655 141 671 175
rect 705 141 843 175
rect 877 161 1123 175
rect 1157 161 1159 195
rect 1295 191 1311 215
rect 1345 191 1361 225
rect 877 145 1159 161
rect 1193 147 1209 181
rect 1243 147 1259 181
rect 877 141 893 145
rect 655 137 893 141
rect 1193 111 1259 147
rect 1295 155 1361 191
rect 1295 121 1311 155
rect 1345 121 1361 155
rect 1395 225 1791 249
rect 1395 191 1397 225
rect 1431 221 1791 225
rect 1431 215 1569 221
rect 1431 191 1433 215
rect 1021 107 1259 111
rect 553 97 979 103
rect 553 85 569 97
rect 431 63 569 85
rect 603 63 757 97
rect 791 63 929 97
rect 963 63 979 97
rect 209 51 979 63
rect 1021 73 1037 107
rect 1071 73 1209 107
rect 1243 87 1259 107
rect 1395 111 1433 191
rect 1567 187 1569 215
rect 1603 215 1741 221
rect 1603 187 1605 215
rect 1395 87 1397 111
rect 1243 77 1397 87
rect 1431 77 1433 111
rect 1243 73 1433 77
rect 1021 51 1433 73
rect 1467 179 1533 181
rect 1467 145 1483 179
rect 1517 145 1533 179
rect 1467 107 1533 145
rect 1467 73 1483 107
rect 1517 73 1533 107
rect 1467 17 1533 73
rect 1567 111 1605 187
rect 1739 187 1741 215
rect 1775 187 1791 221
rect 1567 77 1569 111
rect 1603 77 1605 111
rect 1567 61 1605 77
rect 1639 175 1705 179
rect 1639 141 1655 175
rect 1689 141 1705 175
rect 1639 107 1705 141
rect 1639 73 1655 107
rect 1689 73 1705 107
rect 1639 17 1705 73
rect 1739 111 1791 187
rect 1739 77 1741 111
rect 1775 77 1791 111
rect 1739 61 1791 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4b_4
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 1759 316 1793 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1087 390 1121 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1183 390 1217 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 761840
string GDS_START 746138
<< end >>
