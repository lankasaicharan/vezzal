magic
tech sky130A
magscale 1 2
timestamp 1627202617
<< checkpaint >>
rect -1298 -1308 2034 1852
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 9 67 735 203
rect 30 -17 64 67
rect 285 21 735 67
<< scnmos >>
rect 87 93 117 177
rect 175 93 205 177
rect 363 47 393 177
rect 447 47 477 177
rect 543 47 573 177
rect 627 47 657 177
<< scpmoshvt >>
rect 79 410 109 494
rect 176 297 206 381
rect 363 297 393 497
rect 447 297 477 497
rect 543 297 573 497
rect 627 297 657 497
<< ndiff >>
rect 35 149 87 177
rect 35 115 43 149
rect 77 115 87 149
rect 35 93 87 115
rect 117 149 175 177
rect 117 115 131 149
rect 165 115 175 149
rect 117 93 175 115
rect 205 149 257 177
rect 205 115 215 149
rect 249 115 257 149
rect 205 93 257 115
rect 311 93 363 177
rect 311 59 319 93
rect 353 59 363 93
rect 311 47 363 59
rect 393 116 447 177
rect 393 82 403 116
rect 437 82 447 116
rect 393 47 447 82
rect 477 95 543 177
rect 477 61 493 95
rect 527 61 543 95
rect 477 47 543 61
rect 573 116 627 177
rect 573 82 583 116
rect 617 82 627 116
rect 573 47 627 82
rect 657 163 709 177
rect 657 129 667 163
rect 701 129 709 163
rect 657 95 709 129
rect 657 61 667 95
rect 701 61 709 95
rect 657 47 709 61
<< pdiff >>
rect 27 475 79 494
rect 27 441 35 475
rect 69 441 79 475
rect 27 410 79 441
rect 109 482 161 494
rect 109 448 119 482
rect 153 448 161 482
rect 109 410 161 448
rect 124 381 161 410
rect 311 425 363 497
rect 311 391 319 425
rect 353 391 363 425
rect 124 297 176 381
rect 206 353 257 381
rect 311 379 363 391
rect 206 343 258 353
rect 206 309 216 343
rect 250 309 258 343
rect 206 297 258 309
rect 313 297 363 379
rect 393 297 447 497
rect 477 297 543 497
rect 573 297 627 497
rect 657 485 709 497
rect 657 451 667 485
rect 701 451 709 485
rect 657 417 709 451
rect 657 383 667 417
rect 701 383 709 417
rect 657 297 709 383
<< ndiffc >>
rect 43 115 77 149
rect 131 115 165 149
rect 215 115 249 149
rect 319 59 353 93
rect 403 82 437 116
rect 493 61 527 95
rect 583 82 617 116
rect 667 129 701 163
rect 667 61 701 95
<< pdiffc >>
rect 35 441 69 475
rect 119 448 153 482
rect 319 391 353 425
rect 216 309 250 343
rect 667 451 701 485
rect 667 383 701 417
<< poly >>
rect 79 494 109 520
rect 363 497 393 523
rect 447 497 477 523
rect 543 497 573 523
rect 627 497 657 523
rect 79 265 109 410
rect 176 381 206 407
rect 176 265 206 297
rect 363 265 393 297
rect 447 265 477 297
rect 543 265 573 297
rect 627 265 657 297
rect 76 249 130 265
rect 76 215 86 249
rect 120 215 130 249
rect 76 199 130 215
rect 174 249 240 265
rect 174 215 190 249
rect 224 215 240 249
rect 174 199 240 215
rect 293 249 393 265
rect 293 215 303 249
rect 337 215 393 249
rect 293 199 393 215
rect 435 249 489 265
rect 435 215 445 249
rect 479 215 489 249
rect 435 199 489 215
rect 531 249 585 265
rect 531 215 541 249
rect 575 215 585 249
rect 531 199 585 215
rect 627 249 694 265
rect 627 215 643 249
rect 677 215 694 249
rect 627 199 694 215
rect 87 177 117 199
rect 175 177 205 199
rect 363 177 393 199
rect 447 177 477 199
rect 543 177 573 199
rect 627 177 657 199
rect 87 67 117 93
rect 175 67 205 93
rect 363 21 393 47
rect 447 21 477 47
rect 543 21 573 47
rect 627 21 657 47
<< polycont >>
rect 86 215 120 249
rect 190 215 224 249
rect 303 215 337 249
rect 445 215 479 249
rect 541 215 575 249
rect 643 215 677 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 475 69 491
rect 17 441 35 475
rect 103 482 169 527
rect 103 448 119 482
rect 153 448 169 482
rect 207 459 479 493
rect 651 485 717 527
rect 17 414 69 441
rect 207 414 241 459
rect 17 377 241 414
rect 294 391 319 425
rect 353 391 411 425
rect 17 165 52 377
rect 86 249 156 339
rect 199 309 216 343
rect 250 309 318 343
rect 199 305 318 309
rect 282 265 318 305
rect 120 215 156 249
rect 86 199 156 215
rect 190 249 248 265
rect 224 215 248 249
rect 190 199 248 215
rect 282 249 337 265
rect 282 215 303 249
rect 282 199 337 215
rect 282 165 318 199
rect 17 149 81 165
rect 17 115 43 149
rect 77 115 81 149
rect 17 90 81 115
rect 131 149 165 165
rect 131 17 165 115
rect 215 149 318 165
rect 249 131 318 149
rect 371 165 411 391
rect 445 249 479 459
rect 565 326 617 482
rect 651 451 667 485
rect 701 451 717 485
rect 651 417 717 451
rect 651 383 667 417
rect 701 383 717 417
rect 651 375 717 383
rect 445 199 479 215
rect 523 289 617 326
rect 523 249 589 289
rect 659 255 719 341
rect 523 215 541 249
rect 575 215 589 249
rect 523 199 589 215
rect 623 249 719 255
rect 623 215 643 249
rect 677 215 719 249
rect 623 199 719 215
rect 371 131 617 165
rect 215 90 249 115
rect 403 116 443 131
rect 303 93 369 96
rect 303 59 319 93
rect 353 59 369 93
rect 437 82 443 116
rect 577 116 617 131
rect 403 60 443 82
rect 477 95 543 97
rect 477 61 493 95
rect 527 61 543 95
rect 577 82 583 116
rect 577 62 617 82
rect 651 163 717 165
rect 651 129 667 163
rect 701 129 717 163
rect 651 95 717 129
rect 303 17 369 59
rect 477 17 543 61
rect 651 61 667 95
rect 701 61 717 95
rect 651 17 717 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 673 221 707 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 122 289 156 323 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 581 289 615 323 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 581 85 615 119 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor4bb_1
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 1726292
string GDS_START 1719932
string path 0.000 0.000 18.400 0.000 
<< end >>
