magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3138 1852
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 1 21 1825 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 173 47 203 177
rect 267 47 297 177
rect 371 47 401 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 747 47 777 177
rect 945 47 975 177
rect 1039 47 1069 177
rect 1133 47 1163 177
rect 1227 47 1257 177
rect 1311 47 1341 177
rect 1405 47 1435 177
rect 1499 47 1529 177
rect 1614 47 1644 177
rect 1717 47 1747 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 937 297 973 497
rect 1031 297 1067 497
rect 1125 297 1161 497
rect 1219 297 1255 497
rect 1313 297 1349 497
rect 1407 297 1443 497
rect 1501 297 1537 497
rect 1606 297 1642 497
rect 1709 297 1745 497
<< ndiff >>
rect 27 97 79 177
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 165 173 177
rect 109 131 129 165
rect 163 131 173 165
rect 109 47 173 131
rect 203 97 267 177
rect 203 63 223 97
rect 257 63 267 97
rect 203 47 267 63
rect 297 165 371 177
rect 297 131 317 165
rect 351 131 371 165
rect 297 47 371 131
rect 401 97 455 177
rect 401 63 411 97
rect 445 63 455 97
rect 401 47 455 63
rect 485 165 549 177
rect 485 131 505 165
rect 539 131 549 165
rect 485 47 549 131
rect 579 97 643 177
rect 579 63 599 97
rect 633 63 643 97
rect 579 47 643 63
rect 673 165 747 177
rect 673 131 693 165
rect 727 131 747 165
rect 673 47 747 131
rect 777 97 829 177
rect 777 63 787 97
rect 821 63 829 97
rect 777 47 829 63
rect 883 93 945 177
rect 883 59 891 93
rect 925 59 945 93
rect 883 47 945 59
rect 975 101 1039 177
rect 975 67 985 101
rect 1019 67 1039 101
rect 975 47 1039 67
rect 1069 93 1133 177
rect 1069 59 1079 93
rect 1113 59 1133 93
rect 1069 47 1133 59
rect 1163 101 1227 177
rect 1163 67 1173 101
rect 1207 67 1227 101
rect 1163 47 1227 67
rect 1257 102 1311 177
rect 1257 68 1267 102
rect 1301 68 1311 102
rect 1257 47 1311 68
rect 1341 101 1405 177
rect 1341 67 1361 101
rect 1395 67 1405 101
rect 1341 47 1405 67
rect 1435 93 1499 177
rect 1435 59 1455 93
rect 1489 59 1499 93
rect 1435 47 1499 59
rect 1529 152 1614 177
rect 1529 118 1549 152
rect 1583 118 1614 152
rect 1529 47 1614 118
rect 1644 93 1717 177
rect 1644 59 1663 93
rect 1697 59 1717 93
rect 1644 47 1717 59
rect 1747 101 1799 177
rect 1747 67 1757 101
rect 1791 67 1799 101
rect 1747 47 1799 67
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 297 81 451
rect 117 349 175 497
rect 117 315 129 349
rect 163 315 175 349
rect 117 297 175 315
rect 211 485 269 497
rect 211 451 223 485
rect 257 451 269 485
rect 211 297 269 451
rect 305 349 363 497
rect 305 315 317 349
rect 351 315 363 349
rect 305 297 363 315
rect 399 485 457 497
rect 399 451 411 485
rect 445 451 457 485
rect 399 297 457 451
rect 493 417 551 497
rect 493 383 505 417
rect 539 383 551 417
rect 493 297 551 383
rect 587 485 645 497
rect 587 451 599 485
rect 633 451 645 485
rect 587 297 645 451
rect 681 417 739 497
rect 681 383 693 417
rect 727 383 739 417
rect 681 297 739 383
rect 775 485 829 497
rect 775 451 787 485
rect 821 451 829 485
rect 775 297 829 451
rect 883 485 937 497
rect 883 451 891 485
rect 925 451 937 485
rect 883 297 937 451
rect 973 349 1031 497
rect 973 315 985 349
rect 1019 315 1031 349
rect 973 297 1031 315
rect 1067 485 1125 497
rect 1067 451 1079 485
rect 1113 451 1125 485
rect 1067 297 1125 451
rect 1161 349 1219 497
rect 1161 315 1173 349
rect 1207 315 1219 349
rect 1161 297 1219 315
rect 1255 485 1313 497
rect 1255 451 1267 485
rect 1301 451 1313 485
rect 1255 297 1313 451
rect 1349 477 1407 497
rect 1349 443 1361 477
rect 1395 443 1407 477
rect 1349 409 1407 443
rect 1349 375 1361 409
rect 1395 375 1407 409
rect 1349 297 1407 375
rect 1443 485 1501 497
rect 1443 451 1455 485
rect 1489 451 1501 485
rect 1443 297 1501 451
rect 1537 477 1606 497
rect 1537 443 1549 477
rect 1583 443 1606 477
rect 1537 409 1606 443
rect 1537 375 1549 409
rect 1583 375 1606 409
rect 1537 297 1606 375
rect 1642 485 1709 497
rect 1642 451 1663 485
rect 1697 451 1709 485
rect 1642 297 1709 451
rect 1745 477 1799 497
rect 1745 443 1757 477
rect 1791 443 1799 477
rect 1745 409 1799 443
rect 1745 375 1757 409
rect 1791 375 1799 409
rect 1745 297 1799 375
<< ndiffc >>
rect 35 63 69 97
rect 129 131 163 165
rect 223 63 257 97
rect 317 131 351 165
rect 411 63 445 97
rect 505 131 539 165
rect 599 63 633 97
rect 693 131 727 165
rect 787 63 821 97
rect 891 59 925 93
rect 985 67 1019 101
rect 1079 59 1113 93
rect 1173 67 1207 101
rect 1267 68 1301 102
rect 1361 67 1395 101
rect 1455 59 1489 93
rect 1549 118 1583 152
rect 1663 59 1697 93
rect 1757 67 1791 101
<< pdiffc >>
rect 35 451 69 485
rect 129 315 163 349
rect 223 451 257 485
rect 317 315 351 349
rect 411 451 445 485
rect 505 383 539 417
rect 599 451 633 485
rect 693 383 727 417
rect 787 451 821 485
rect 891 451 925 485
rect 985 315 1019 349
rect 1079 451 1113 485
rect 1173 315 1207 349
rect 1267 451 1301 485
rect 1361 443 1395 477
rect 1361 375 1395 409
rect 1455 451 1489 485
rect 1549 443 1583 477
rect 1549 375 1583 409
rect 1663 451 1697 485
rect 1757 443 1791 477
rect 1757 375 1791 409
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 937 497 973 523
rect 1031 497 1067 523
rect 1125 497 1161 523
rect 1219 497 1255 523
rect 1313 497 1349 523
rect 1407 497 1443 523
rect 1501 497 1537 523
rect 1606 497 1642 523
rect 1709 497 1745 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 937 282 973 297
rect 1031 282 1067 297
rect 1125 282 1161 297
rect 1219 282 1255 297
rect 1313 282 1349 297
rect 1407 282 1443 297
rect 1501 282 1537 297
rect 1606 282 1642 297
rect 1709 282 1745 297
rect 79 265 119 282
rect 173 265 213 282
rect 267 265 307 282
rect 361 265 401 282
rect 79 249 401 265
rect 79 215 122 249
rect 156 215 190 249
rect 224 215 401 249
rect 79 199 401 215
rect 79 177 109 199
rect 173 177 203 199
rect 267 177 297 199
rect 371 177 401 199
rect 455 265 495 282
rect 549 265 589 282
rect 643 265 683 282
rect 737 265 777 282
rect 935 265 975 282
rect 1029 265 1069 282
rect 1123 265 1163 282
rect 1217 265 1257 282
rect 455 249 777 265
rect 455 215 471 249
rect 505 215 549 249
rect 583 215 627 249
rect 661 215 705 249
rect 739 215 777 249
rect 455 199 777 215
rect 878 249 1257 265
rect 878 215 895 249
rect 929 215 963 249
rect 997 215 1041 249
rect 1075 215 1119 249
rect 1153 215 1197 249
rect 1231 215 1257 249
rect 878 199 1257 215
rect 455 177 485 199
rect 549 177 579 199
rect 643 177 673 199
rect 747 177 777 199
rect 945 177 975 199
rect 1039 177 1069 199
rect 1133 177 1163 199
rect 1227 177 1257 199
rect 1311 265 1351 282
rect 1405 265 1445 282
rect 1499 265 1539 282
rect 1604 265 1644 282
rect 1707 265 1747 282
rect 1311 249 1644 265
rect 1311 215 1502 249
rect 1536 215 1584 249
rect 1618 215 1644 249
rect 1311 199 1644 215
rect 1686 249 1750 265
rect 1686 215 1696 249
rect 1730 215 1750 249
rect 1686 199 1750 215
rect 1311 177 1341 199
rect 1405 177 1435 199
rect 1499 177 1529 199
rect 1614 177 1644 199
rect 1717 177 1747 199
rect 79 21 109 47
rect 173 21 203 47
rect 267 21 297 47
rect 371 21 401 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 747 21 777 47
rect 945 21 975 47
rect 1039 21 1069 47
rect 1133 21 1163 47
rect 1227 21 1257 47
rect 1311 21 1341 47
rect 1405 21 1435 47
rect 1499 21 1529 47
rect 1614 21 1644 47
rect 1717 21 1747 47
<< polycont >>
rect 122 215 156 249
rect 190 215 224 249
rect 471 215 505 249
rect 549 215 583 249
rect 627 215 661 249
rect 705 215 739 249
rect 895 215 929 249
rect 963 215 997 249
rect 1041 215 1075 249
rect 1119 215 1153 249
rect 1197 215 1231 249
rect 1502 215 1536 249
rect 1584 215 1618 249
rect 1696 215 1730 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 875 485 941 527
rect 19 451 35 485
rect 69 451 223 485
rect 257 451 411 485
rect 445 451 599 485
rect 633 451 787 485
rect 821 451 837 485
rect 875 451 891 485
rect 925 451 941 485
rect 1053 485 1129 527
rect 1053 451 1079 485
rect 1113 451 1129 485
rect 1241 485 1317 527
rect 1241 451 1267 485
rect 1301 451 1317 485
rect 1361 477 1395 493
rect 19 97 64 451
rect 1429 485 1505 527
rect 1429 451 1455 485
rect 1489 451 1505 485
rect 1549 477 1583 493
rect 1361 417 1395 443
rect 1647 485 1713 527
rect 1647 451 1663 485
rect 1697 451 1713 485
rect 1757 477 1809 493
rect 1549 417 1583 443
rect 479 383 505 417
rect 539 383 693 417
rect 727 409 1583 417
rect 727 383 1361 409
rect 1395 383 1549 409
rect 1361 359 1395 375
rect 1549 359 1583 375
rect 1791 443 1809 477
rect 1757 409 1809 443
rect 1791 375 1809 409
rect 1757 359 1809 375
rect 103 315 129 349
rect 163 315 317 349
rect 351 315 985 349
rect 1019 315 1173 349
rect 1207 315 1226 349
rect 1272 285 1730 319
rect 118 249 247 265
rect 118 215 122 249
rect 156 215 190 249
rect 224 215 247 249
rect 118 199 247 215
rect 471 249 810 265
rect 1272 258 1306 285
rect 505 215 549 249
rect 583 215 627 249
rect 661 215 705 249
rect 739 215 810 249
rect 849 249 1306 258
rect 1696 249 1730 285
rect 849 215 895 249
rect 929 215 963 249
rect 997 215 1041 249
rect 1075 215 1119 249
rect 1153 215 1197 249
rect 1231 215 1306 249
rect 1486 215 1502 249
rect 1536 215 1584 249
rect 471 199 810 215
rect 291 165 336 187
rect 103 131 129 165
rect 163 131 317 165
rect 351 131 370 153
rect 479 131 505 165
rect 539 131 693 165
rect 727 131 1207 165
rect 985 101 1019 131
rect 19 63 35 97
rect 69 63 223 97
rect 257 63 411 97
rect 445 63 599 97
rect 633 63 787 97
rect 821 63 837 97
rect 875 59 891 93
rect 925 59 941 93
rect 875 17 941 59
rect 1173 101 1207 131
rect 1394 181 1420 187
rect 1394 153 1583 181
rect 1360 152 1583 153
rect 1360 143 1549 152
rect 985 51 1019 67
rect 1053 59 1079 93
rect 1113 59 1129 93
rect 1053 17 1129 59
rect 1173 51 1207 67
rect 1241 102 1316 118
rect 1241 68 1267 102
rect 1301 68 1316 102
rect 1241 17 1316 68
rect 1360 101 1395 143
rect 1618 165 1662 249
rect 1696 199 1730 215
rect 1774 165 1809 359
rect 1618 131 1809 165
rect 1360 67 1361 101
rect 1360 51 1395 67
rect 1449 93 1499 109
rect 1549 102 1583 118
rect 1757 101 1809 131
rect 1449 59 1455 93
rect 1489 59 1499 93
rect 1449 17 1499 59
rect 1647 59 1663 93
rect 1697 59 1713 93
rect 1647 17 1713 59
rect 1791 67 1809 101
rect 1757 51 1809 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 336 165 370 187
rect 336 153 351 165
rect 351 153 370 165
rect 1360 153 1394 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 324 187 382 193
rect 324 153 336 187
rect 370 184 382 187
rect 1338 187 1406 193
rect 1338 184 1360 187
rect 370 156 1360 184
rect 370 153 382 156
rect 324 147 382 153
rect 1338 153 1360 156
rect 1394 153 1406 187
rect 1338 147 1406 153
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel locali s 1041 221 1075 255 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 764 221 799 255 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 S
port 3 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 A0
port 1 nsew signal input
flabel locali s 29 425 63 459 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 29 357 63 391 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 A1
port 2 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2i_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2172184
string GDS_START 2159226
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
