magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3026 1975
<< nwell >>
rect -38 331 1766 704
rect 285 319 771 331
<< pwell >>
rect 343 241 453 243
rect 343 235 769 241
rect 1 229 769 235
rect 1 49 1664 229
rect 0 0 1728 49
<< scnmos >>
rect 80 125 110 209
rect 166 125 196 209
rect 449 131 479 215
rect 574 47 604 215
rect 660 47 690 215
rect 795 119 825 203
rect 867 119 897 203
rect 953 119 983 203
rect 1047 119 1077 203
rect 1193 119 1223 203
rect 1265 119 1295 203
rect 1351 119 1381 203
rect 1445 119 1475 203
rect 1531 119 1561 203
<< scpmoshvt >>
rect 80 397 110 525
rect 166 397 196 525
rect 393 355 423 483
rect 566 355 596 607
rect 652 355 682 607
rect 787 419 817 547
rect 859 419 889 547
rect 945 419 975 547
rect 1017 419 1047 547
rect 1193 419 1223 547
rect 1265 419 1295 547
rect 1370 419 1400 547
rect 1472 419 1502 547
rect 1558 419 1588 547
<< ndiff >>
rect 369 215 427 217
rect 369 209 449 215
rect 27 184 80 209
rect 27 150 35 184
rect 69 150 80 184
rect 27 125 80 150
rect 110 184 166 209
rect 110 150 121 184
rect 155 150 166 184
rect 110 125 166 150
rect 196 174 249 209
rect 196 140 207 174
rect 241 140 249 174
rect 196 125 249 140
rect 369 175 381 209
rect 415 175 449 209
rect 369 131 449 175
rect 479 131 574 215
rect 501 69 574 131
rect 501 35 513 69
rect 547 47 574 69
rect 604 203 660 215
rect 604 169 615 203
rect 649 169 660 203
rect 604 101 660 169
rect 604 67 615 101
rect 649 67 660 101
rect 604 47 660 67
rect 690 203 743 215
rect 690 179 795 203
rect 690 145 750 179
rect 784 145 795 179
rect 690 119 795 145
rect 825 119 867 203
rect 897 163 953 203
rect 897 129 908 163
rect 942 129 953 163
rect 897 119 953 129
rect 983 119 1047 203
rect 1077 161 1193 203
rect 1077 127 1113 161
rect 1147 127 1193 161
rect 1077 119 1193 127
rect 1223 119 1265 203
rect 1295 161 1351 203
rect 1295 127 1306 161
rect 1340 127 1351 161
rect 1295 119 1351 127
rect 1381 119 1445 203
rect 1475 161 1531 203
rect 1475 127 1486 161
rect 1520 127 1531 161
rect 1475 119 1531 127
rect 1561 178 1638 203
rect 1561 144 1572 178
rect 1606 144 1638 178
rect 1561 119 1638 144
rect 690 93 743 119
rect 690 59 701 93
rect 735 59 743 93
rect 690 47 743 59
rect 547 35 559 47
rect 501 27 559 35
<< pdiff >>
rect 513 595 566 607
rect 27 513 80 525
rect 27 479 35 513
rect 69 479 80 513
rect 27 445 80 479
rect 27 411 35 445
rect 69 411 80 445
rect 27 397 80 411
rect 110 511 166 525
rect 110 477 121 511
rect 155 477 166 511
rect 110 443 166 477
rect 110 409 121 443
rect 155 409 166 443
rect 110 397 166 409
rect 196 511 249 525
rect 196 477 207 511
rect 241 477 249 511
rect 513 561 521 595
rect 555 561 566 595
rect 513 483 566 561
rect 196 443 249 477
rect 196 409 207 443
rect 241 409 249 443
rect 196 397 249 409
rect 321 451 393 483
rect 321 417 329 451
rect 363 417 393 451
rect 321 405 393 417
rect 343 355 393 405
rect 423 355 566 483
rect 596 437 652 607
rect 596 403 607 437
rect 641 403 652 437
rect 596 355 652 403
rect 682 595 735 607
rect 682 561 693 595
rect 727 561 735 595
rect 682 547 735 561
rect 682 419 787 547
rect 817 419 859 547
rect 889 533 945 547
rect 889 499 900 533
rect 934 499 945 533
rect 889 465 945 499
rect 889 431 900 465
rect 934 431 945 465
rect 889 419 945 431
rect 975 419 1017 547
rect 1047 535 1193 547
rect 1047 501 1058 535
rect 1092 508 1193 535
rect 1092 501 1148 508
rect 1047 474 1148 501
rect 1182 474 1193 508
rect 1047 467 1193 474
rect 1047 433 1058 467
rect 1092 433 1193 467
rect 1047 419 1193 433
rect 1223 419 1265 547
rect 1295 533 1370 547
rect 1295 499 1316 533
rect 1350 499 1370 533
rect 1295 465 1370 499
rect 1295 431 1316 465
rect 1350 431 1370 465
rect 1295 419 1370 431
rect 1400 419 1472 547
rect 1502 535 1558 547
rect 1502 501 1513 535
rect 1547 501 1558 535
rect 1502 467 1558 501
rect 1502 433 1513 467
rect 1547 433 1558 467
rect 1502 419 1558 433
rect 1588 533 1641 547
rect 1588 499 1599 533
rect 1633 499 1641 533
rect 1588 465 1641 499
rect 1588 431 1599 465
rect 1633 431 1641 465
rect 1588 419 1641 431
rect 682 355 735 419
<< ndiffc >>
rect 35 150 69 184
rect 121 150 155 184
rect 207 140 241 174
rect 381 175 415 209
rect 513 35 547 69
rect 615 169 649 203
rect 615 67 649 101
rect 750 145 784 179
rect 908 129 942 163
rect 1113 127 1147 161
rect 1306 127 1340 161
rect 1486 127 1520 161
rect 1572 144 1606 178
rect 701 59 735 93
<< pdiffc >>
rect 35 479 69 513
rect 35 411 69 445
rect 121 477 155 511
rect 121 409 155 443
rect 207 477 241 511
rect 521 561 555 595
rect 207 409 241 443
rect 329 417 363 451
rect 607 403 641 437
rect 693 561 727 595
rect 900 499 934 533
rect 900 431 934 465
rect 1058 501 1092 535
rect 1148 474 1182 508
rect 1058 433 1092 467
rect 1316 499 1350 533
rect 1316 431 1350 465
rect 1513 501 1547 535
rect 1513 433 1547 467
rect 1599 499 1633 533
rect 1599 431 1633 465
<< poly >>
rect 566 607 596 633
rect 652 607 682 633
rect 945 615 1588 645
rect 80 525 110 551
rect 166 547 423 577
rect 166 525 196 547
rect 393 483 423 547
rect 80 323 110 397
rect 166 371 196 397
rect 245 349 311 365
rect 787 547 817 573
rect 859 547 889 573
rect 945 547 975 615
rect 1017 547 1047 573
rect 1193 547 1223 573
rect 1265 547 1295 573
rect 1370 547 1400 615
rect 1472 547 1502 573
rect 1558 547 1588 615
rect 245 323 261 349
rect 80 315 261 323
rect 295 315 311 349
rect 80 293 311 315
rect 166 281 311 293
rect 166 247 261 281
rect 295 247 311 281
rect 393 323 423 355
rect 393 307 479 323
rect 393 273 415 307
rect 449 273 479 307
rect 566 304 596 355
rect 652 304 682 355
rect 566 303 682 304
rect 787 303 817 419
rect 859 381 889 419
rect 945 393 975 419
rect 1017 385 1047 419
rect 1193 387 1223 419
rect 859 351 897 381
rect 1017 369 1113 385
rect 1017 355 1063 369
rect 867 307 897 351
rect 1047 335 1063 355
rect 1097 335 1113 369
rect 1047 319 1113 335
rect 1157 371 1223 387
rect 1157 337 1173 371
rect 1207 337 1223 371
rect 393 257 479 273
rect 80 209 110 235
rect 166 231 311 247
rect 166 209 196 231
rect 449 215 479 257
rect 521 287 682 303
rect 521 253 537 287
rect 571 267 682 287
rect 759 287 825 303
rect 571 253 690 267
rect 521 237 690 253
rect 759 253 775 287
rect 809 253 825 287
rect 867 280 1005 307
rect 867 277 955 280
rect 759 237 825 253
rect 574 215 604 237
rect 660 215 690 237
rect 80 51 110 125
rect 166 99 196 125
rect 449 51 479 131
rect 80 21 479 51
rect 795 203 825 237
rect 939 246 955 277
rect 989 246 1005 280
rect 939 230 1005 246
rect 1047 277 1083 319
rect 1157 303 1223 337
rect 867 203 897 229
rect 953 203 983 230
rect 1047 203 1077 277
rect 1157 269 1173 303
rect 1207 269 1223 303
rect 1265 307 1295 419
rect 1370 393 1400 419
rect 1472 387 1502 419
rect 1445 371 1511 387
rect 1445 337 1461 371
rect 1495 337 1511 371
rect 1445 321 1511 337
rect 1558 385 1588 419
rect 1558 369 1624 385
rect 1558 335 1574 369
rect 1608 335 1624 369
rect 1265 280 1403 307
rect 1265 277 1353 280
rect 1157 253 1223 269
rect 1193 203 1223 253
rect 1337 246 1353 277
rect 1387 246 1403 280
rect 1337 230 1403 246
rect 1265 203 1295 229
rect 1351 203 1381 230
rect 1445 203 1475 321
rect 1558 301 1624 335
rect 1558 273 1574 301
rect 1531 267 1574 273
rect 1608 267 1624 301
rect 1531 243 1624 267
rect 1531 203 1561 243
rect 795 93 825 119
rect 867 51 897 119
rect 953 93 983 119
rect 1047 93 1077 119
rect 1193 93 1223 119
rect 1265 51 1295 119
rect 1351 93 1381 119
rect 1445 93 1475 119
rect 1531 51 1561 119
rect 574 21 604 47
rect 660 21 690 47
rect 867 21 1561 51
<< polycont >>
rect 261 315 295 349
rect 261 247 295 281
rect 415 273 449 307
rect 1063 335 1097 369
rect 1173 337 1207 371
rect 537 253 571 287
rect 775 253 809 287
rect 955 246 989 280
rect 1173 269 1207 303
rect 1461 337 1495 371
rect 1574 335 1608 369
rect 1353 246 1387 280
rect 1574 267 1608 301
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 19 563 327 597
rect 19 513 77 563
rect 19 479 35 513
rect 69 479 77 513
rect 19 445 77 479
rect 19 411 35 445
rect 69 411 77 445
rect 19 184 77 411
rect 19 150 35 184
rect 69 150 77 184
rect 19 134 77 150
rect 111 511 155 527
rect 293 521 327 563
rect 505 595 571 649
rect 505 561 521 595
rect 555 561 571 595
rect 505 557 571 561
rect 677 595 743 649
rect 677 561 693 595
rect 727 561 743 595
rect 677 557 743 561
rect 884 533 950 549
rect 884 521 900 533
rect 111 477 121 511
rect 111 443 155 477
rect 111 409 121 443
rect 111 184 155 409
rect 111 150 121 184
rect 111 99 155 150
rect 191 511 259 515
rect 191 477 207 511
rect 241 498 259 511
rect 191 464 223 477
rect 257 464 259 498
rect 293 499 900 521
rect 934 499 950 533
rect 293 487 950 499
rect 191 443 259 464
rect 869 465 950 487
rect 191 409 207 443
rect 241 409 259 443
rect 191 399 259 409
rect 313 451 379 453
rect 313 417 329 451
rect 363 417 379 451
rect 605 437 651 453
rect 191 179 225 399
rect 313 365 379 417
rect 259 349 379 365
rect 259 315 261 349
rect 295 315 379 349
rect 259 281 379 315
rect 259 247 261 281
rect 295 247 379 281
rect 413 307 465 424
rect 413 273 415 307
rect 449 273 465 307
rect 605 403 607 437
rect 641 403 651 437
rect 413 257 465 273
rect 521 287 571 303
rect 259 223 379 247
rect 521 253 537 287
rect 259 213 431 223
rect 345 209 431 213
rect 191 174 257 179
rect 191 140 207 174
rect 241 140 257 174
rect 345 175 381 209
rect 415 175 431 209
rect 345 173 431 175
rect 191 133 257 140
rect 521 139 571 253
rect 293 105 571 139
rect 605 203 651 403
rect 685 287 833 453
rect 685 253 775 287
rect 809 253 833 287
rect 685 229 833 253
rect 869 431 900 465
rect 934 431 950 465
rect 869 415 950 431
rect 1042 535 1198 649
rect 1042 501 1058 535
rect 1092 508 1198 535
rect 1092 501 1148 508
rect 1042 474 1148 501
rect 1182 474 1198 508
rect 1042 467 1198 474
rect 1042 433 1058 467
rect 1092 458 1198 467
rect 1267 533 1366 549
rect 1267 499 1316 533
rect 1350 499 1366 533
rect 1267 498 1366 499
rect 1267 464 1279 498
rect 1313 465 1366 498
rect 1313 464 1316 465
rect 1092 433 1108 458
rect 1042 415 1108 433
rect 1267 431 1316 464
rect 1350 431 1366 465
rect 605 169 615 203
rect 649 169 651 203
rect 293 99 327 105
rect 111 65 327 99
rect 605 101 651 169
rect 497 69 563 71
rect 497 35 513 69
rect 547 35 563 69
rect 605 67 615 101
rect 649 67 651 101
rect 605 51 651 67
rect 685 179 803 195
rect 685 145 750 179
rect 784 145 803 179
rect 685 93 803 145
rect 869 165 903 415
rect 937 369 1123 381
rect 937 335 1063 369
rect 1097 335 1123 369
rect 937 314 1123 335
rect 1157 371 1233 424
rect 1157 337 1173 371
rect 1207 337 1233 371
rect 1157 303 1233 337
rect 939 246 955 280
rect 989 246 1005 280
rect 1157 269 1173 303
rect 1207 269 1233 303
rect 1267 415 1366 431
rect 1497 535 1563 649
rect 1497 501 1513 535
rect 1547 501 1563 535
rect 1497 467 1563 501
rect 1497 433 1513 467
rect 1547 433 1563 467
rect 1497 417 1563 433
rect 1597 533 1694 549
rect 1597 499 1599 533
rect 1633 499 1694 533
rect 1597 465 1694 499
rect 1597 431 1599 465
rect 1633 431 1694 465
rect 1597 415 1694 431
rect 939 233 1005 246
rect 939 199 1231 233
rect 869 163 958 165
rect 869 129 908 163
rect 942 129 958 163
rect 869 113 958 129
rect 1097 161 1163 165
rect 1097 127 1113 161
rect 1147 127 1163 161
rect 685 59 701 93
rect 735 59 803 93
rect 497 17 563 35
rect 685 17 803 59
rect 1097 17 1163 127
rect 1197 87 1231 199
rect 1267 163 1303 415
rect 1337 337 1461 371
rect 1495 337 1524 371
rect 1337 314 1524 337
rect 1558 369 1624 381
rect 1558 335 1574 369
rect 1608 335 1624 369
rect 1558 301 1624 335
rect 1337 246 1353 280
rect 1387 246 1426 280
rect 1558 267 1574 301
rect 1608 267 1624 301
rect 1558 265 1624 267
rect 1337 231 1426 246
rect 1660 231 1694 415
rect 1337 197 1694 231
rect 1267 161 1356 163
rect 1267 127 1306 161
rect 1340 127 1356 161
rect 1267 121 1356 127
rect 1392 87 1426 197
rect 1570 178 1622 197
rect 1197 53 1426 87
rect 1470 161 1536 163
rect 1470 127 1486 161
rect 1520 127 1536 161
rect 1570 144 1572 178
rect 1606 144 1622 178
rect 1570 128 1622 144
rect 1470 17 1536 127
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 223 477 241 498
rect 241 477 257 498
rect 223 464 257 477
rect 1279 464 1313 498
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
<< metal1 >>
rect 0 683 1728 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1728 683
rect 0 617 1728 649
rect 211 498 269 504
rect 211 464 223 498
rect 257 495 269 498
rect 1267 498 1325 504
rect 1267 495 1279 498
rect 257 467 1279 495
rect 257 464 269 467
rect 211 458 269 464
rect 1267 464 1279 467
rect 1313 464 1325 498
rect 1267 458 1325 464
rect 0 17 1728 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1728 17
rect 0 -49 1728 -17
<< labels >>
flabel pwell s 0 0 1728 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 1728 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux4_2
flabel metal1 s 0 617 1728 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 1728 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 607 94 641 128 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 1183 390 1217 424 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1728 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1405712
string GDS_START 1392220
<< end >>
