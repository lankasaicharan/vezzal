magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 331 1190 704
<< pwell >>
rect 57 241 553 263
rect 57 49 1149 241
rect 0 0 1152 49
<< scnmos >>
rect 140 69 170 237
rect 242 69 272 237
rect 328 69 358 237
rect 430 69 460 237
rect 696 47 726 215
rect 782 47 812 215
rect 868 47 898 215
rect 954 47 984 215
rect 1040 47 1070 215
<< scpmoshvt >>
rect 140 367 170 619
rect 242 367 272 619
rect 328 367 358 619
rect 430 367 460 619
rect 516 367 546 619
rect 602 367 632 619
rect 688 367 718 619
rect 774 367 804 619
rect 1040 367 1070 619
<< ndiff >>
rect 83 225 140 237
rect 83 191 91 225
rect 125 191 140 225
rect 83 115 140 191
rect 83 81 91 115
rect 125 81 140 115
rect 83 69 140 81
rect 170 229 242 237
rect 170 195 181 229
rect 215 195 242 229
rect 170 153 242 195
rect 170 119 181 153
rect 215 119 242 153
rect 170 69 242 119
rect 272 179 328 237
rect 272 145 283 179
rect 317 145 328 179
rect 272 111 328 145
rect 272 77 283 111
rect 317 77 328 111
rect 272 69 328 77
rect 358 229 430 237
rect 358 195 385 229
rect 419 195 430 229
rect 358 153 430 195
rect 358 119 385 153
rect 419 119 430 153
rect 358 69 430 119
rect 460 225 527 237
rect 460 191 485 225
rect 519 191 527 225
rect 460 115 527 191
rect 460 81 485 115
rect 519 81 527 115
rect 460 69 527 81
rect 643 102 696 215
rect 643 68 651 102
rect 685 68 696 102
rect 643 47 696 68
rect 726 203 782 215
rect 726 169 737 203
rect 771 169 782 203
rect 726 101 782 169
rect 726 67 737 101
rect 771 67 782 101
rect 726 47 782 67
rect 812 177 868 215
rect 812 143 823 177
rect 857 143 868 177
rect 812 89 868 143
rect 812 55 823 89
rect 857 55 868 89
rect 812 47 868 55
rect 898 203 954 215
rect 898 169 909 203
rect 943 169 954 203
rect 898 101 954 169
rect 898 67 909 101
rect 943 67 954 101
rect 898 47 954 67
rect 984 207 1040 215
rect 984 173 995 207
rect 1029 173 1040 207
rect 984 93 1040 173
rect 984 59 995 93
rect 1029 59 1040 93
rect 984 47 1040 59
rect 1070 203 1123 215
rect 1070 169 1081 203
rect 1115 169 1123 203
rect 1070 101 1123 169
rect 1070 67 1081 101
rect 1115 67 1123 101
rect 1070 47 1123 67
<< pdiff >>
rect 87 599 140 619
rect 87 565 95 599
rect 129 565 140 599
rect 87 513 140 565
rect 87 479 95 513
rect 129 479 140 513
rect 87 438 140 479
rect 87 404 95 438
rect 129 404 140 438
rect 87 367 140 404
rect 170 547 242 619
rect 170 513 197 547
rect 231 513 242 547
rect 170 436 242 513
rect 170 402 197 436
rect 231 402 242 436
rect 170 367 242 402
rect 272 574 328 619
rect 272 540 283 574
rect 317 540 328 574
rect 272 502 328 540
rect 272 468 283 502
rect 317 468 328 502
rect 272 367 328 468
rect 358 547 430 619
rect 358 513 385 547
rect 419 513 430 547
rect 358 436 430 513
rect 358 402 385 436
rect 419 402 430 436
rect 358 367 430 402
rect 460 599 516 619
rect 460 565 471 599
rect 505 565 516 599
rect 460 504 516 565
rect 460 470 471 504
rect 505 470 516 504
rect 460 413 516 470
rect 460 379 471 413
rect 505 379 516 413
rect 460 367 516 379
rect 546 607 602 619
rect 546 573 557 607
rect 591 573 602 607
rect 546 530 602 573
rect 546 496 557 530
rect 591 496 602 530
rect 546 453 602 496
rect 546 419 557 453
rect 591 419 602 453
rect 546 367 602 419
rect 632 599 688 619
rect 632 565 643 599
rect 677 565 688 599
rect 632 504 688 565
rect 632 470 643 504
rect 677 470 688 504
rect 632 413 688 470
rect 632 379 643 413
rect 677 379 688 413
rect 632 367 688 379
rect 718 607 774 619
rect 718 573 729 607
rect 763 573 774 607
rect 718 530 774 573
rect 718 496 729 530
rect 763 496 774 530
rect 718 453 774 496
rect 718 419 729 453
rect 763 419 774 453
rect 718 367 774 419
rect 804 599 857 619
rect 804 565 815 599
rect 849 565 857 599
rect 804 504 857 565
rect 804 470 815 504
rect 849 470 857 504
rect 987 607 1040 619
rect 987 573 995 607
rect 1029 573 1040 607
rect 987 504 1040 573
rect 804 413 857 470
rect 804 379 815 413
rect 849 379 857 413
rect 804 367 857 379
rect 987 470 995 504
rect 1029 470 1040 504
rect 987 413 1040 470
rect 987 379 995 413
rect 1029 379 1040 413
rect 987 367 1040 379
rect 1070 599 1123 619
rect 1070 565 1081 599
rect 1115 565 1123 599
rect 1070 504 1123 565
rect 1070 470 1081 504
rect 1115 470 1123 504
rect 1070 413 1123 470
rect 1070 379 1081 413
rect 1115 379 1123 413
rect 1070 367 1123 379
<< ndiffc >>
rect 91 191 125 225
rect 91 81 125 115
rect 181 195 215 229
rect 181 119 215 153
rect 283 145 317 179
rect 283 77 317 111
rect 385 195 419 229
rect 385 119 419 153
rect 485 191 519 225
rect 485 81 519 115
rect 651 68 685 102
rect 737 169 771 203
rect 737 67 771 101
rect 823 143 857 177
rect 823 55 857 89
rect 909 169 943 203
rect 909 67 943 101
rect 995 173 1029 207
rect 995 59 1029 93
rect 1081 169 1115 203
rect 1081 67 1115 101
<< pdiffc >>
rect 95 565 129 599
rect 95 479 129 513
rect 95 404 129 438
rect 197 513 231 547
rect 197 402 231 436
rect 283 540 317 574
rect 283 468 317 502
rect 385 513 419 547
rect 385 402 419 436
rect 471 565 505 599
rect 471 470 505 504
rect 471 379 505 413
rect 557 573 591 607
rect 557 496 591 530
rect 557 419 591 453
rect 643 565 677 599
rect 643 470 677 504
rect 643 379 677 413
rect 729 573 763 607
rect 729 496 763 530
rect 729 419 763 453
rect 815 565 849 599
rect 815 470 849 504
rect 995 573 1029 607
rect 815 379 849 413
rect 995 470 1029 504
rect 995 379 1029 413
rect 1081 565 1115 599
rect 1081 470 1115 504
rect 1081 379 1115 413
<< poly >>
rect 140 619 170 645
rect 242 619 272 645
rect 328 619 358 645
rect 430 619 460 645
rect 516 619 546 645
rect 602 619 632 645
rect 688 619 718 645
rect 774 619 804 645
rect 1040 619 1070 645
rect 889 467 955 483
rect 889 433 905 467
rect 939 433 955 467
rect 889 399 955 433
rect 140 335 170 367
rect 242 335 272 367
rect 328 335 358 367
rect 430 335 460 367
rect 140 319 460 335
rect 140 285 156 319
rect 190 285 226 319
rect 260 285 303 319
rect 337 285 460 319
rect 516 345 546 367
rect 602 345 632 367
rect 688 345 718 367
rect 774 345 804 367
rect 889 365 905 399
rect 939 365 955 399
rect 889 345 955 365
rect 1040 345 1070 367
rect 516 315 1070 345
rect 140 269 460 285
rect 140 259 272 269
rect 140 237 170 259
rect 242 237 272 259
rect 328 237 358 269
rect 430 237 460 269
rect 555 251 984 267
rect 555 217 571 251
rect 605 237 984 251
rect 605 217 621 237
rect 555 201 621 217
rect 696 215 726 237
rect 782 215 812 237
rect 868 215 898 237
rect 954 215 984 237
rect 1040 215 1070 315
rect 140 43 170 69
rect 242 43 272 69
rect 328 43 358 69
rect 430 43 460 69
rect 696 21 726 47
rect 782 21 812 47
rect 868 21 898 47
rect 954 21 984 47
rect 1040 21 1070 47
<< polycont >>
rect 905 433 939 467
rect 156 285 190 319
rect 226 285 260 319
rect 303 285 337 319
rect 905 365 939 399
rect 571 217 605 251
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 79 599 507 615
rect 79 565 95 599
rect 129 581 471 599
rect 129 565 133 581
rect 79 513 133 565
rect 281 574 335 581
rect 79 479 95 513
rect 129 479 133 513
rect 79 438 133 479
rect 79 404 95 438
rect 129 404 133 438
rect 79 384 133 404
rect 181 513 197 547
rect 231 513 247 547
rect 181 436 247 513
rect 281 540 283 574
rect 317 540 335 574
rect 469 565 471 581
rect 505 565 507 599
rect 281 502 335 540
rect 281 468 283 502
rect 317 468 335 502
rect 281 452 335 468
rect 369 513 385 547
rect 419 513 435 547
rect 181 402 197 436
rect 231 418 247 436
rect 369 436 435 513
rect 369 418 385 436
rect 231 402 385 418
rect 419 402 435 436
rect 181 384 435 402
rect 31 319 353 350
rect 31 285 156 319
rect 190 285 226 319
rect 260 285 303 319
rect 337 285 353 319
rect 389 300 435 384
rect 469 504 507 565
rect 469 470 471 504
rect 505 470 507 504
rect 469 413 507 470
rect 541 607 607 649
rect 541 573 557 607
rect 591 573 607 607
rect 541 530 607 573
rect 541 496 557 530
rect 591 496 607 530
rect 541 453 607 496
rect 541 419 557 453
rect 591 419 607 453
rect 641 599 679 615
rect 641 565 643 599
rect 677 565 679 599
rect 641 504 679 565
rect 641 470 643 504
rect 677 470 679 504
rect 469 379 471 413
rect 505 385 507 413
rect 641 413 679 470
rect 713 607 779 649
rect 713 573 729 607
rect 763 573 779 607
rect 713 530 779 573
rect 713 496 729 530
rect 763 496 779 530
rect 713 453 779 496
rect 713 419 729 453
rect 763 419 779 453
rect 813 599 860 615
rect 813 565 815 599
rect 849 565 860 599
rect 979 607 1036 649
rect 979 573 995 607
rect 1029 573 1036 607
rect 813 504 860 565
rect 813 470 815 504
rect 849 470 860 504
rect 641 385 643 413
rect 505 379 643 385
rect 677 385 679 413
rect 813 413 860 470
rect 813 385 815 413
rect 677 379 815 385
rect 849 379 860 413
rect 469 351 860 379
rect 894 467 945 572
rect 894 433 905 467
rect 939 433 945 467
rect 894 399 945 433
rect 894 365 905 399
rect 939 365 945 399
rect 894 349 945 365
rect 979 504 1036 573
rect 979 470 995 504
rect 1029 470 1036 504
rect 979 413 1036 470
rect 979 379 995 413
rect 1029 379 1036 413
rect 979 363 1036 379
rect 1070 599 1131 615
rect 1070 565 1081 599
rect 1115 565 1131 599
rect 1070 504 1131 565
rect 1070 470 1081 504
rect 1115 470 1131 504
rect 1070 413 1131 470
rect 1070 379 1081 413
rect 1115 379 1131 413
rect 1070 315 1131 379
rect 389 249 449 300
rect 555 279 1131 315
rect 75 225 129 241
rect 75 191 91 225
rect 125 191 129 225
rect 75 115 129 191
rect 165 229 449 249
rect 165 195 181 229
rect 215 215 385 229
rect 215 195 231 215
rect 165 153 231 195
rect 369 195 385 215
rect 419 195 449 229
rect 165 119 181 153
rect 215 119 231 153
rect 267 145 283 179
rect 317 145 333 179
rect 75 81 91 115
rect 125 85 129 115
rect 267 111 333 145
rect 369 153 449 195
rect 369 119 385 153
rect 419 119 449 153
rect 483 225 521 253
rect 483 191 485 225
rect 519 191 521 225
rect 555 251 621 279
rect 555 217 571 251
rect 605 217 621 251
rect 555 213 621 217
rect 483 179 521 191
rect 721 211 945 245
rect 721 203 773 211
rect 721 179 737 203
rect 483 169 737 179
rect 771 169 773 203
rect 907 203 945 211
rect 483 145 773 169
rect 267 85 283 111
rect 125 81 283 85
rect 75 77 283 81
rect 317 85 333 111
rect 483 115 535 145
rect 483 85 485 115
rect 317 81 485 85
rect 519 81 535 115
rect 317 77 535 81
rect 75 51 535 77
rect 635 102 701 111
rect 635 68 651 102
rect 685 68 701 102
rect 635 17 701 68
rect 735 101 773 145
rect 735 67 737 101
rect 771 67 773 101
rect 735 51 773 67
rect 807 143 823 177
rect 857 143 873 177
rect 807 89 873 143
rect 807 55 823 89
rect 857 55 873 89
rect 807 17 873 55
rect 907 169 909 203
rect 943 169 945 203
rect 907 101 945 169
rect 907 67 909 101
rect 943 67 945 101
rect 907 51 945 67
rect 979 207 1045 223
rect 979 173 995 207
rect 1029 173 1045 207
rect 979 93 1045 173
rect 979 59 995 93
rect 1029 59 1045 93
rect 979 17 1045 59
rect 1079 203 1131 279
rect 1079 169 1081 203
rect 1115 169 1131 203
rect 1079 101 1131 169
rect 1079 67 1081 101
rect 1115 67 1131 101
rect 1079 51 1131 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 einvn_4
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 895 464 929 498 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 895 538 929 572 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4223164
string GDS_START 4213354
<< end >>
