magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2738 1975
<< nwell >>
rect -38 331 1478 704
<< pwell >>
rect 1 183 419 201
rect 1 49 1159 183
rect 0 0 1440 49
<< scnmos >>
rect 80 47 110 175
rect 152 47 182 175
rect 238 47 268 175
rect 310 47 340 175
rect 504 47 534 157
rect 576 47 606 157
rect 662 47 692 157
rect 734 47 764 157
rect 820 47 850 157
rect 892 47 922 157
rect 978 47 1008 157
rect 1050 47 1080 157
<< scpmoshvt >>
rect 80 417 130 617
rect 186 417 236 617
rect 292 417 342 617
rect 398 417 448 617
rect 504 417 554 617
rect 610 417 660 617
rect 716 417 766 617
rect 822 417 872 617
rect 928 417 978 617
rect 1034 417 1084 617
rect 1140 417 1190 617
rect 1246 417 1296 617
<< ndiff >>
rect 27 162 80 175
rect 27 128 35 162
rect 69 128 80 162
rect 27 94 80 128
rect 27 60 35 94
rect 69 60 80 94
rect 27 47 80 60
rect 110 47 152 175
rect 182 162 238 175
rect 182 128 193 162
rect 227 128 238 162
rect 182 94 238 128
rect 182 60 193 94
rect 227 60 238 94
rect 182 47 238 60
rect 268 47 310 175
rect 340 162 393 175
rect 340 128 351 162
rect 385 157 393 162
rect 385 128 504 157
rect 340 119 504 128
rect 340 94 459 119
rect 340 60 351 94
rect 385 85 459 94
rect 493 85 504 119
rect 385 60 504 85
rect 340 47 504 60
rect 534 47 576 157
rect 606 119 662 157
rect 606 85 617 119
rect 651 85 662 119
rect 606 47 662 85
rect 692 47 734 157
rect 764 105 820 157
rect 764 71 775 105
rect 809 71 820 105
rect 764 47 820 71
rect 850 47 892 157
rect 922 119 978 157
rect 922 85 933 119
rect 967 85 978 119
rect 922 47 978 85
rect 1008 47 1050 157
rect 1080 119 1133 157
rect 1080 85 1091 119
rect 1125 85 1133 119
rect 1080 47 1133 85
<< pdiff >>
rect 27 599 80 617
rect 27 565 35 599
rect 69 565 80 599
rect 27 531 80 565
rect 27 497 35 531
rect 69 497 80 531
rect 27 463 80 497
rect 27 429 35 463
rect 69 429 80 463
rect 27 417 80 429
rect 130 599 186 617
rect 130 565 141 599
rect 175 565 186 599
rect 130 531 186 565
rect 130 497 141 531
rect 175 497 186 531
rect 130 463 186 497
rect 130 429 141 463
rect 175 429 186 463
rect 130 417 186 429
rect 236 599 292 617
rect 236 565 247 599
rect 281 565 292 599
rect 236 531 292 565
rect 236 497 247 531
rect 281 497 292 531
rect 236 463 292 497
rect 236 429 247 463
rect 281 429 292 463
rect 236 417 292 429
rect 342 599 398 617
rect 342 565 353 599
rect 387 565 398 599
rect 342 531 398 565
rect 342 497 353 531
rect 387 497 398 531
rect 342 463 398 497
rect 342 429 353 463
rect 387 429 398 463
rect 342 417 398 429
rect 448 599 504 617
rect 448 565 459 599
rect 493 565 504 599
rect 448 531 504 565
rect 448 497 459 531
rect 493 497 504 531
rect 448 463 504 497
rect 448 429 459 463
rect 493 429 504 463
rect 448 417 504 429
rect 554 599 610 617
rect 554 565 565 599
rect 599 565 610 599
rect 554 531 610 565
rect 554 497 565 531
rect 599 497 610 531
rect 554 463 610 497
rect 554 429 565 463
rect 599 429 610 463
rect 554 417 610 429
rect 660 599 716 617
rect 660 565 671 599
rect 705 565 716 599
rect 660 531 716 565
rect 660 497 671 531
rect 705 497 716 531
rect 660 463 716 497
rect 660 429 671 463
rect 705 429 716 463
rect 660 417 716 429
rect 766 599 822 617
rect 766 565 777 599
rect 811 565 822 599
rect 766 531 822 565
rect 766 497 777 531
rect 811 497 822 531
rect 766 463 822 497
rect 766 429 777 463
rect 811 429 822 463
rect 766 417 822 429
rect 872 599 928 617
rect 872 565 883 599
rect 917 565 928 599
rect 872 531 928 565
rect 872 497 883 531
rect 917 497 928 531
rect 872 463 928 497
rect 872 429 883 463
rect 917 429 928 463
rect 872 417 928 429
rect 978 599 1034 617
rect 978 565 989 599
rect 1023 565 1034 599
rect 978 531 1034 565
rect 978 497 989 531
rect 1023 497 1034 531
rect 978 463 1034 497
rect 978 429 989 463
rect 1023 429 1034 463
rect 978 417 1034 429
rect 1084 599 1140 617
rect 1084 565 1095 599
rect 1129 565 1140 599
rect 1084 531 1140 565
rect 1084 497 1095 531
rect 1129 497 1140 531
rect 1084 463 1140 497
rect 1084 429 1095 463
rect 1129 429 1140 463
rect 1084 417 1140 429
rect 1190 599 1246 617
rect 1190 565 1201 599
rect 1235 565 1246 599
rect 1190 531 1246 565
rect 1190 497 1201 531
rect 1235 497 1246 531
rect 1190 463 1246 497
rect 1190 429 1201 463
rect 1235 429 1246 463
rect 1190 417 1246 429
rect 1296 599 1349 617
rect 1296 565 1307 599
rect 1341 565 1349 599
rect 1296 531 1349 565
rect 1296 497 1307 531
rect 1341 497 1349 531
rect 1296 463 1349 497
rect 1296 429 1307 463
rect 1341 429 1349 463
rect 1296 417 1349 429
<< ndiffc >>
rect 35 128 69 162
rect 35 60 69 94
rect 193 128 227 162
rect 193 60 227 94
rect 351 128 385 162
rect 351 60 385 94
rect 459 85 493 119
rect 617 85 651 119
rect 775 71 809 105
rect 933 85 967 119
rect 1091 85 1125 119
<< pdiffc >>
rect 35 565 69 599
rect 35 497 69 531
rect 35 429 69 463
rect 141 565 175 599
rect 141 497 175 531
rect 141 429 175 463
rect 247 565 281 599
rect 247 497 281 531
rect 247 429 281 463
rect 353 565 387 599
rect 353 497 387 531
rect 353 429 387 463
rect 459 565 493 599
rect 459 497 493 531
rect 459 429 493 463
rect 565 565 599 599
rect 565 497 599 531
rect 565 429 599 463
rect 671 565 705 599
rect 671 497 705 531
rect 671 429 705 463
rect 777 565 811 599
rect 777 497 811 531
rect 777 429 811 463
rect 883 565 917 599
rect 883 497 917 531
rect 883 429 917 463
rect 989 565 1023 599
rect 989 497 1023 531
rect 989 429 1023 463
rect 1095 565 1129 599
rect 1095 497 1129 531
rect 1095 429 1129 463
rect 1201 565 1235 599
rect 1201 497 1235 531
rect 1201 429 1235 463
rect 1307 565 1341 599
rect 1307 497 1341 531
rect 1307 429 1341 463
<< poly >>
rect 80 617 130 645
rect 186 617 236 645
rect 292 617 342 645
rect 398 617 448 645
rect 504 617 554 645
rect 610 617 660 645
rect 716 617 766 645
rect 822 617 872 645
rect 928 617 978 645
rect 1034 617 1084 645
rect 1140 617 1190 645
rect 1246 617 1296 645
rect 80 313 130 417
rect 186 313 236 417
rect 292 313 342 417
rect 398 313 448 417
rect 80 297 448 313
rect 80 263 96 297
rect 130 263 448 297
rect 80 247 448 263
rect 504 309 554 417
rect 610 309 660 417
rect 716 309 766 417
rect 822 309 872 417
rect 928 309 978 417
rect 1034 309 1084 417
rect 1140 309 1190 417
rect 1246 309 1296 417
rect 504 291 1296 309
rect 504 257 520 291
rect 554 257 588 291
rect 622 257 656 291
rect 690 257 724 291
rect 758 257 1296 291
rect 80 175 110 247
rect 152 175 182 247
rect 238 175 268 247
rect 310 175 340 247
rect 504 241 1296 257
rect 504 157 534 241
rect 576 157 606 241
rect 662 157 692 241
rect 734 157 764 241
rect 820 157 850 241
rect 892 157 922 241
rect 978 157 1008 241
rect 1050 157 1080 241
rect 80 21 110 47
rect 152 21 182 47
rect 238 21 268 47
rect 310 21 340 47
rect 504 21 534 47
rect 576 21 606 47
rect 662 21 692 47
rect 734 21 764 47
rect 820 21 850 47
rect 892 21 922 47
rect 978 21 1008 47
rect 1050 21 1080 47
<< polycont >>
rect 96 263 130 297
rect 520 257 554 291
rect 588 257 622 291
rect 656 257 690 291
rect 724 257 758 291
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 19 599 85 649
rect 19 565 35 599
rect 69 565 85 599
rect 19 531 85 565
rect 19 497 35 531
rect 69 497 85 531
rect 19 463 85 497
rect 19 429 35 463
rect 69 429 85 463
rect 19 413 85 429
rect 125 599 191 615
rect 125 565 141 599
rect 175 565 191 599
rect 125 531 191 565
rect 125 497 141 531
rect 175 497 191 531
rect 125 463 191 497
rect 125 429 141 463
rect 175 429 191 463
rect 125 388 191 429
rect 231 599 297 649
rect 231 565 247 599
rect 281 565 297 599
rect 231 531 297 565
rect 231 497 247 531
rect 281 497 297 531
rect 231 463 297 497
rect 231 429 247 463
rect 281 429 297 463
rect 231 422 297 429
rect 332 599 399 615
rect 332 565 353 599
rect 387 565 399 599
rect 332 531 399 565
rect 332 497 353 531
rect 387 497 399 531
rect 332 463 399 497
rect 332 429 353 463
rect 387 429 399 463
rect 332 388 399 429
rect 443 599 509 649
rect 443 565 459 599
rect 493 565 509 599
rect 443 531 509 565
rect 443 497 459 531
rect 493 497 509 531
rect 443 463 509 497
rect 443 429 459 463
rect 493 429 509 463
rect 443 417 509 429
rect 549 599 615 615
rect 549 565 565 599
rect 599 565 615 599
rect 549 531 615 565
rect 549 497 565 531
rect 599 497 615 531
rect 549 463 615 497
rect 549 429 565 463
rect 599 429 615 463
rect 25 313 85 376
rect 125 354 399 388
rect 25 297 143 313
rect 25 263 96 297
rect 130 263 143 297
rect 25 228 143 263
rect 191 307 399 354
rect 549 377 615 429
rect 655 599 721 649
rect 655 565 671 599
rect 705 565 721 599
rect 655 531 721 565
rect 655 497 671 531
rect 705 497 721 531
rect 655 463 721 497
rect 655 429 671 463
rect 705 429 721 463
rect 655 417 721 429
rect 761 599 827 615
rect 761 565 777 599
rect 811 565 827 599
rect 761 531 827 565
rect 761 497 777 531
rect 811 497 827 531
rect 761 463 827 497
rect 761 429 777 463
rect 811 429 827 463
rect 761 377 827 429
rect 867 599 933 649
rect 867 565 883 599
rect 917 565 933 599
rect 867 531 933 565
rect 867 497 883 531
rect 917 497 933 531
rect 867 463 933 497
rect 867 429 883 463
rect 917 429 933 463
rect 867 417 933 429
rect 973 599 1039 615
rect 973 565 989 599
rect 1023 565 1039 599
rect 973 531 1039 565
rect 973 497 989 531
rect 1023 497 1039 531
rect 973 463 1039 497
rect 973 429 989 463
rect 1023 429 1039 463
rect 549 375 827 377
rect 973 375 1039 429
rect 1079 599 1145 649
rect 1079 565 1095 599
rect 1129 565 1145 599
rect 1079 531 1145 565
rect 1079 497 1095 531
rect 1129 497 1145 531
rect 1079 463 1145 497
rect 1079 429 1095 463
rect 1129 429 1145 463
rect 1079 417 1145 429
rect 1185 599 1251 615
rect 1185 565 1201 599
rect 1235 565 1251 599
rect 1185 531 1251 565
rect 1185 497 1201 531
rect 1235 497 1251 531
rect 1185 463 1251 497
rect 1185 429 1201 463
rect 1235 429 1251 463
rect 549 358 1039 375
rect 1185 358 1251 429
rect 1291 599 1357 649
rect 1291 565 1307 599
rect 1341 565 1357 599
rect 1291 531 1357 565
rect 1291 497 1307 531
rect 1341 497 1357 531
rect 1291 463 1357 497
rect 1291 429 1307 463
rect 1341 429 1357 463
rect 1291 417 1357 429
rect 549 341 1347 358
rect 191 291 774 307
rect 191 257 520 291
rect 554 257 588 291
rect 622 257 656 291
rect 690 257 724 291
rect 758 257 774 291
rect 191 241 774 257
rect 191 197 246 241
rect 820 234 1347 341
rect 820 207 992 234
rect 25 162 85 178
rect 25 128 35 162
rect 69 128 85 162
rect 25 94 85 128
rect 25 60 35 94
rect 69 60 85 94
rect 25 17 85 60
rect 177 162 246 197
rect 177 128 193 162
rect 227 128 246 162
rect 177 94 246 128
rect 177 60 193 94
rect 227 60 246 94
rect 177 51 246 60
rect 335 162 510 175
rect 335 128 351 162
rect 385 128 510 162
rect 335 119 510 128
rect 335 94 459 119
rect 335 60 351 94
rect 385 85 459 94
rect 493 85 510 119
rect 385 60 510 85
rect 601 155 992 207
rect 601 119 667 155
rect 601 85 617 119
rect 651 85 667 119
rect 601 69 667 85
rect 759 105 825 121
rect 759 71 775 105
rect 809 71 825 105
rect 335 17 510 60
rect 759 17 825 71
rect 917 119 992 155
rect 917 85 933 119
rect 967 85 992 119
rect 917 69 992 85
rect 1075 119 1141 135
rect 1075 85 1091 119
rect 1125 85 1141 119
rect 1075 17 1141 85
rect 1175 53 1347 234
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 683 1440 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 0 617 1440 649
rect 0 17 1440 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -49 1440 -17
<< labels >>
flabel pwell s 0 0 1440 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1440 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkbuflp_8
flabel metal1 s 0 617 1440 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1440 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 1183 168 1217 202 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1183 94 1217 128 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1279 94 1313 128 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 1279 168 1313 202 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1440 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5388288
string GDS_START 5377980
<< end >>
