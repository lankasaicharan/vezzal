magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 332 710 704
<< pwell >>
rect 1 49 666 248
rect 0 0 672 49
<< scpmos >>
rect 86 368 116 592
rect 186 368 216 592
rect 354 368 384 592
rect 444 368 474 592
rect 556 368 586 592
<< nmoslvt >>
rect 84 74 114 222
rect 247 74 277 222
rect 325 74 355 222
rect 439 74 469 222
rect 553 74 583 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 120 247 222
rect 114 86 125 120
rect 159 86 202 120
rect 236 86 247 120
rect 114 74 247 86
rect 277 74 325 222
rect 355 74 439 222
rect 469 74 553 222
rect 583 210 640 222
rect 583 176 594 210
rect 628 176 640 210
rect 583 120 640 176
rect 583 86 594 120
rect 628 86 640 120
rect 583 74 640 86
<< pdiff >>
rect 27 580 86 592
rect 27 546 39 580
rect 73 546 86 580
rect 27 505 86 546
rect 27 471 39 505
rect 73 471 86 505
rect 27 424 86 471
rect 27 390 39 424
rect 73 390 86 424
rect 27 368 86 390
rect 116 580 186 592
rect 116 546 139 580
rect 173 546 186 580
rect 116 492 186 546
rect 116 458 139 492
rect 173 458 186 492
rect 116 368 186 458
rect 216 578 354 592
rect 216 544 239 578
rect 273 561 354 578
rect 273 544 307 561
rect 216 527 307 544
rect 341 527 354 561
rect 216 368 354 527
rect 384 441 444 592
rect 384 407 397 441
rect 431 407 444 441
rect 384 368 444 407
rect 474 542 556 592
rect 474 508 498 542
rect 532 508 556 542
rect 474 368 556 508
rect 586 580 645 592
rect 586 546 599 580
rect 633 546 645 580
rect 586 501 645 546
rect 586 467 599 501
rect 633 467 645 501
rect 586 424 645 467
rect 586 390 599 424
rect 633 390 645 424
rect 586 368 645 390
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 86 159 120
rect 202 86 236 120
rect 594 176 628 210
rect 594 86 628 120
<< pdiffc >>
rect 39 546 73 580
rect 39 471 73 505
rect 39 390 73 424
rect 139 546 173 580
rect 139 458 173 492
rect 239 544 273 578
rect 307 527 341 561
rect 397 407 431 441
rect 498 508 532 542
rect 599 546 633 580
rect 599 467 633 501
rect 599 390 633 424
<< poly >>
rect 86 592 116 618
rect 186 592 216 618
rect 354 592 384 618
rect 444 592 474 618
rect 556 592 586 618
rect 86 353 116 368
rect 186 353 216 368
rect 354 353 384 368
rect 444 353 474 368
rect 556 353 586 368
rect 83 326 119 353
rect 21 310 119 326
rect 21 276 37 310
rect 71 276 119 310
rect 21 260 119 276
rect 183 336 219 353
rect 351 336 387 353
rect 441 336 477 353
rect 183 320 277 336
rect 183 286 217 320
rect 251 286 277 320
rect 183 270 277 286
rect 84 222 114 260
rect 247 222 277 270
rect 325 320 391 336
rect 325 286 341 320
rect 375 286 391 320
rect 325 270 391 286
rect 439 320 505 336
rect 439 286 455 320
rect 489 286 505 320
rect 439 270 505 286
rect 553 326 589 353
rect 553 310 651 326
rect 553 276 601 310
rect 635 276 651 310
rect 325 222 355 270
rect 439 222 469 270
rect 553 260 651 276
rect 553 222 583 260
rect 84 48 114 74
rect 247 48 277 74
rect 325 48 355 74
rect 439 48 469 74
rect 553 48 583 74
<< polycont >>
rect 37 276 71 310
rect 217 286 251 320
rect 341 286 375 320
rect 455 286 489 320
rect 601 276 635 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 23 580 89 596
rect 23 546 39 580
rect 73 546 89 580
rect 23 505 89 546
rect 23 471 39 505
rect 73 471 89 505
rect 23 424 89 471
rect 123 580 189 596
rect 123 546 139 580
rect 173 546 189 580
rect 123 492 189 546
rect 223 578 357 649
rect 223 544 239 578
rect 273 561 357 578
rect 273 544 307 561
rect 223 527 307 544
rect 341 527 357 561
rect 223 526 357 527
rect 289 492 357 526
rect 481 542 549 649
rect 481 508 498 542
rect 532 508 549 542
rect 481 492 549 508
rect 583 580 649 596
rect 583 546 599 580
rect 633 546 649 580
rect 583 501 649 546
rect 123 458 139 492
rect 173 458 255 492
rect 583 467 599 501
rect 633 467 649 501
rect 583 458 649 467
rect 221 441 649 458
rect 23 390 39 424
rect 73 390 167 424
rect 221 407 397 441
rect 431 424 649 441
rect 431 407 599 424
rect 221 390 599 407
rect 633 390 649 424
rect 21 310 87 356
rect 21 276 37 310
rect 71 276 87 310
rect 21 260 87 276
rect 121 226 167 390
rect 201 320 267 356
rect 201 286 217 320
rect 251 286 267 320
rect 201 270 267 286
rect 313 320 391 356
rect 313 286 341 320
rect 375 286 391 320
rect 313 270 391 286
rect 439 320 551 356
rect 439 286 455 320
rect 489 286 551 320
rect 439 270 551 286
rect 585 310 651 356
rect 585 276 601 310
rect 635 276 651 310
rect 585 260 651 276
rect 23 210 644 226
rect 23 176 39 210
rect 73 192 594 210
rect 73 176 89 192
rect 23 120 89 176
rect 578 176 594 192
rect 628 176 644 210
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 120 252 136
rect 123 86 125 120
rect 159 86 202 120
rect 236 86 252 120
rect 123 17 252 86
rect 578 120 644 176
rect 578 86 594 120
rect 628 86 644 120
rect 578 70 644 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a41oi_1
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 1270900
string GDS_START 1264914
<< end >>
