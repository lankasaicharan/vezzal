magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2834 1975
<< nwell >>
rect -38 331 1574 704
rect 799 325 1007 331
<< pwell >>
rect 506 179 994 243
rect 38 162 994 179
rect 1347 162 1535 241
rect 38 49 1535 162
rect 0 0 1536 49
<< scnmos >>
rect 124 69 154 153
rect 210 69 240 153
rect 304 69 334 153
rect 593 133 623 217
rect 691 133 721 217
rect 763 133 793 217
rect 881 49 911 217
rect 1078 52 1108 136
rect 1164 52 1194 136
rect 1236 52 1266 136
rect 1426 47 1456 215
<< scpmoshvt >>
rect 80 468 110 596
rect 152 468 182 596
rect 402 409 432 537
rect 620 463 650 547
rect 706 463 736 547
rect 778 463 808 547
rect 888 361 918 613
rect 1083 367 1113 495
rect 1201 367 1231 495
rect 1287 367 1317 495
rect 1389 367 1419 619
<< ndiff >>
rect 64 118 124 153
rect 64 84 74 118
rect 108 84 124 118
rect 64 69 124 84
rect 154 128 210 153
rect 154 94 165 128
rect 199 94 210 128
rect 154 69 210 94
rect 240 118 304 153
rect 240 84 255 118
rect 289 84 304 118
rect 240 69 304 84
rect 334 128 387 153
rect 532 192 593 217
rect 532 158 544 192
rect 578 158 593 192
rect 532 133 593 158
rect 623 192 691 217
rect 623 158 646 192
rect 680 158 691 192
rect 623 133 691 158
rect 721 133 763 217
rect 793 133 881 217
rect 334 94 345 128
rect 379 94 387 128
rect 334 69 387 94
rect 808 69 881 133
rect 808 35 820 69
rect 854 49 881 69
rect 911 207 968 217
rect 911 173 922 207
rect 956 173 968 207
rect 911 49 968 173
rect 1373 163 1426 215
rect 1025 111 1078 136
rect 1025 77 1033 111
rect 1067 77 1078 111
rect 1025 52 1078 77
rect 1108 111 1164 136
rect 1108 77 1119 111
rect 1153 77 1164 111
rect 1108 52 1164 77
rect 1194 52 1236 136
rect 1266 111 1319 136
rect 1266 77 1277 111
rect 1311 77 1319 111
rect 1266 52 1319 77
rect 1373 129 1381 163
rect 1415 129 1426 163
rect 1373 93 1426 129
rect 1373 59 1381 93
rect 1415 59 1426 93
rect 854 35 866 49
rect 808 27 866 35
rect 1373 47 1426 59
rect 1456 203 1509 215
rect 1456 169 1467 203
rect 1501 169 1509 203
rect 1456 101 1509 169
rect 1456 67 1467 101
rect 1501 67 1509 101
rect 1456 47 1509 67
<< pdiff >>
rect 27 574 80 596
rect 27 540 35 574
rect 69 540 80 574
rect 27 468 80 540
rect 110 468 152 596
rect 182 582 235 596
rect 182 548 193 582
rect 227 548 235 582
rect 182 514 235 548
rect 182 480 193 514
rect 227 480 235 514
rect 182 468 235 480
rect 835 601 888 613
rect 835 567 843 601
rect 877 567 888 601
rect 835 547 888 567
rect 299 504 402 537
rect 299 470 309 504
rect 343 470 402 504
rect 299 409 402 470
rect 432 523 489 537
rect 432 489 445 523
rect 479 489 489 523
rect 432 455 489 489
rect 567 522 620 547
rect 567 488 575 522
rect 609 488 620 522
rect 567 463 620 488
rect 650 522 706 547
rect 650 488 661 522
rect 695 488 706 522
rect 650 463 706 488
rect 736 463 778 547
rect 808 516 888 547
rect 808 482 843 516
rect 877 482 888 516
rect 808 463 888 482
rect 432 421 445 455
rect 479 421 489 455
rect 432 409 489 421
rect 835 431 888 463
rect 835 397 843 431
rect 877 397 888 431
rect 835 361 888 397
rect 918 599 971 613
rect 918 565 929 599
rect 963 565 971 599
rect 918 502 971 565
rect 1336 599 1389 619
rect 1336 565 1344 599
rect 1378 565 1389 599
rect 1128 547 1186 557
rect 918 468 929 502
rect 963 468 971 502
rect 1128 513 1140 547
rect 1174 513 1186 547
rect 1128 495 1186 513
rect 1336 495 1389 565
rect 918 407 971 468
rect 918 373 929 407
rect 963 373 971 407
rect 918 361 971 373
rect 1026 411 1083 495
rect 1026 377 1038 411
rect 1072 377 1083 411
rect 1026 367 1083 377
rect 1113 367 1201 495
rect 1231 484 1287 495
rect 1231 450 1242 484
rect 1276 450 1287 484
rect 1231 416 1287 450
rect 1231 382 1242 416
rect 1276 382 1287 416
rect 1231 367 1287 382
rect 1317 484 1389 495
rect 1317 450 1344 484
rect 1378 450 1389 484
rect 1317 367 1389 450
rect 1419 599 1472 619
rect 1419 565 1430 599
rect 1464 565 1472 599
rect 1419 503 1472 565
rect 1419 469 1430 503
rect 1464 469 1472 503
rect 1419 420 1472 469
rect 1419 386 1430 420
rect 1464 386 1472 420
rect 1419 367 1472 386
<< ndiffc >>
rect 74 84 108 118
rect 165 94 199 128
rect 255 84 289 118
rect 544 158 578 192
rect 646 158 680 192
rect 345 94 379 128
rect 820 35 854 69
rect 922 173 956 207
rect 1033 77 1067 111
rect 1119 77 1153 111
rect 1277 77 1311 111
rect 1381 129 1415 163
rect 1381 59 1415 93
rect 1467 169 1501 203
rect 1467 67 1501 101
<< pdiffc >>
rect 35 540 69 574
rect 193 548 227 582
rect 193 480 227 514
rect 843 567 877 601
rect 309 470 343 504
rect 445 489 479 523
rect 575 488 609 522
rect 661 488 695 522
rect 843 482 877 516
rect 445 421 479 455
rect 843 397 877 431
rect 929 565 963 599
rect 1344 565 1378 599
rect 929 468 963 502
rect 1140 513 1174 547
rect 929 373 963 407
rect 1038 377 1072 411
rect 1242 450 1276 484
rect 1242 382 1276 416
rect 1344 450 1378 484
rect 1430 565 1464 599
rect 1430 469 1464 503
rect 1430 386 1464 420
<< poly >>
rect 80 596 110 622
rect 152 596 182 622
rect 254 615 736 645
rect 80 309 110 468
rect 21 293 110 309
rect 21 259 37 293
rect 71 259 110 293
rect 152 309 182 468
rect 254 387 284 615
rect 402 537 432 563
rect 620 547 650 573
rect 706 547 736 615
rect 888 613 918 639
rect 1389 619 1419 645
rect 778 547 808 573
rect 620 425 650 463
rect 706 437 736 463
rect 402 387 432 409
rect 254 357 432 387
rect 510 395 650 425
rect 778 395 808 463
rect 510 377 540 395
rect 152 293 262 309
rect 152 279 212 293
rect 21 225 110 259
rect 21 191 37 225
rect 71 205 110 225
rect 196 259 212 279
rect 246 259 262 293
rect 402 269 432 357
rect 474 361 540 377
rect 474 327 490 361
rect 524 347 540 361
rect 737 379 808 395
rect 524 327 695 347
rect 737 345 753 379
rect 787 345 808 379
rect 1083 495 1113 521
rect 1201 495 1231 521
rect 1287 495 1317 521
rect 737 329 808 345
rect 474 317 695 327
rect 474 311 540 317
rect 665 281 695 317
rect 196 225 262 259
rect 71 191 154 205
rect 21 175 154 191
rect 196 191 212 225
rect 246 191 262 225
rect 196 175 262 191
rect 304 253 623 269
rect 304 239 431 253
rect 124 153 154 175
rect 210 153 240 175
rect 304 153 334 239
rect 402 219 431 239
rect 465 239 623 253
rect 665 251 721 281
rect 465 219 481 239
rect 402 185 481 219
rect 593 217 623 239
rect 691 217 721 251
rect 763 217 793 329
rect 888 305 918 361
rect 850 289 918 305
rect 1083 292 1113 367
rect 1201 292 1231 367
rect 1287 335 1317 367
rect 850 255 866 289
rect 900 255 918 289
rect 850 239 918 255
rect 1078 276 1231 292
rect 1078 242 1144 276
rect 1178 262 1231 276
rect 1273 319 1339 335
rect 1273 285 1289 319
rect 1323 285 1339 319
rect 1389 303 1419 367
rect 1273 269 1339 285
rect 1381 287 1456 303
rect 1178 242 1194 262
rect 881 217 911 239
rect 402 151 431 185
rect 465 151 481 185
rect 402 135 481 151
rect 593 107 623 133
rect 691 107 721 133
rect 763 107 793 133
rect 124 43 154 69
rect 210 43 240 69
rect 304 43 334 69
rect 1078 208 1194 242
rect 1078 174 1144 208
rect 1178 174 1194 208
rect 1273 188 1303 269
rect 1381 253 1397 287
rect 1431 253 1456 287
rect 1381 237 1456 253
rect 1426 215 1456 237
rect 1078 158 1194 174
rect 1078 136 1108 158
rect 1164 136 1194 158
rect 1236 158 1303 188
rect 1236 136 1266 158
rect 881 23 911 49
rect 1078 26 1108 52
rect 1164 26 1194 52
rect 1236 26 1266 52
rect 1426 21 1456 47
<< polycont >>
rect 37 259 71 293
rect 37 191 71 225
rect 212 259 246 293
rect 490 327 524 361
rect 753 345 787 379
rect 212 191 246 225
rect 431 219 465 253
rect 866 255 900 289
rect 1144 242 1178 276
rect 1289 285 1323 319
rect 431 151 465 185
rect 1144 174 1178 208
rect 1397 253 1431 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 19 574 85 649
rect 19 540 35 574
rect 69 540 85 574
rect 19 532 85 540
rect 142 582 243 598
rect 142 548 193 582
rect 227 548 243 582
rect 142 514 243 548
rect 17 293 93 498
rect 17 259 37 293
rect 71 259 93 293
rect 17 225 93 259
rect 17 191 37 225
rect 71 191 93 225
rect 17 168 93 191
rect 142 480 193 514
rect 227 480 243 514
rect 142 420 243 480
rect 291 504 343 649
rect 291 470 309 504
rect 291 454 343 470
rect 377 575 617 609
rect 377 420 411 575
rect 142 386 411 420
rect 445 523 495 539
rect 479 489 495 523
rect 445 455 495 489
rect 479 421 495 455
rect 142 134 176 386
rect 445 377 495 421
rect 560 522 617 575
rect 827 601 893 649
rect 827 567 843 601
rect 877 567 893 601
rect 560 488 575 522
rect 609 488 617 522
rect 445 361 526 377
rect 445 352 490 361
rect 212 293 273 352
rect 246 259 273 293
rect 212 225 273 259
rect 246 191 273 225
rect 212 168 273 191
rect 329 327 490 352
rect 524 327 526 361
rect 329 311 526 327
rect 58 118 108 134
rect 58 84 74 118
rect 58 17 108 84
rect 142 128 215 134
rect 142 94 165 128
rect 199 94 215 128
rect 142 78 215 94
rect 249 118 295 134
rect 249 84 255 118
rect 289 84 295 118
rect 249 17 295 84
rect 329 128 395 311
rect 560 300 617 488
rect 651 522 699 538
rect 651 488 661 522
rect 695 488 699 522
rect 329 94 345 128
rect 379 94 395 128
rect 329 78 395 94
rect 429 253 481 269
rect 429 219 431 253
rect 465 219 481 253
rect 429 185 481 219
rect 560 208 594 300
rect 651 295 699 488
rect 827 516 893 567
rect 827 482 843 516
rect 877 482 893 516
rect 827 431 893 482
rect 827 397 843 431
rect 877 397 893 431
rect 927 599 986 615
rect 927 565 929 599
rect 963 565 986 599
rect 927 502 986 565
rect 1124 547 1190 649
rect 1124 513 1140 547
rect 1174 513 1190 547
rect 1328 599 1394 649
rect 1328 565 1344 599
rect 1378 565 1394 599
rect 927 468 929 502
rect 963 479 986 502
rect 1226 484 1292 488
rect 963 468 1158 479
rect 927 445 1158 468
rect 927 407 986 445
rect 737 379 793 395
rect 737 345 753 379
rect 787 363 793 379
rect 927 373 929 407
rect 963 373 986 407
rect 927 363 986 373
rect 787 345 986 363
rect 737 329 986 345
rect 651 289 916 295
rect 651 266 866 289
rect 429 151 431 185
rect 465 151 481 185
rect 429 108 481 151
rect 528 192 594 208
rect 528 158 544 192
rect 578 158 594 192
rect 528 142 594 158
rect 628 255 866 266
rect 900 255 916 289
rect 628 192 699 255
rect 952 221 986 329
rect 628 158 646 192
rect 680 158 699 192
rect 906 207 986 221
rect 906 173 922 207
rect 956 173 986 207
rect 1022 377 1038 411
rect 1072 377 1088 411
rect 1022 359 1088 377
rect 628 142 699 158
rect 1022 139 1071 359
rect 1124 346 1158 445
rect 1226 450 1242 484
rect 1276 450 1292 484
rect 1328 484 1394 565
rect 1328 450 1344 484
rect 1378 450 1394 484
rect 1430 599 1519 615
rect 1464 565 1519 599
rect 1430 503 1519 565
rect 1464 469 1519 503
rect 1226 416 1292 450
rect 1430 420 1519 469
rect 1226 382 1242 416
rect 1276 382 1394 416
rect 1124 319 1326 346
rect 1124 312 1289 319
rect 1273 285 1289 312
rect 1323 285 1326 319
rect 1128 276 1239 278
rect 1128 242 1144 276
rect 1178 242 1239 276
rect 1273 269 1326 285
rect 1360 303 1394 382
rect 1464 386 1519 420
rect 1430 370 1519 386
rect 1360 287 1431 303
rect 1128 208 1239 242
rect 1360 253 1397 287
rect 1360 237 1431 253
rect 1360 231 1394 237
rect 1128 174 1144 208
rect 1178 174 1239 208
rect 1128 161 1239 174
rect 1273 197 1394 231
rect 1465 203 1519 370
rect 736 111 1071 139
rect 736 108 1033 111
rect 429 105 1033 108
rect 429 74 770 105
rect 1017 77 1033 105
rect 1067 77 1071 111
rect 804 69 870 71
rect 804 35 820 69
rect 854 35 870 69
rect 1017 61 1071 77
rect 1115 111 1157 127
rect 1115 77 1119 111
rect 1153 77 1157 111
rect 804 17 870 35
rect 1115 17 1157 77
rect 1273 111 1327 197
rect 1465 169 1467 203
rect 1501 169 1519 203
rect 1273 77 1277 111
rect 1311 77 1327 111
rect 1273 61 1327 77
rect 1365 129 1381 163
rect 1415 129 1431 163
rect 1365 93 1431 129
rect 1365 59 1381 93
rect 1415 59 1431 93
rect 1365 17 1431 59
rect 1465 101 1519 169
rect 1465 67 1467 101
rect 1501 67 1519 101
rect 1465 51 1519 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
<< metal1 >>
rect 0 683 1536 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1536 683
rect 0 617 1536 649
rect 0 17 1536 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1536 17
rect 0 -49 1536 -17
<< labels >>
flabel pwell s 0 0 1536 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1536 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdlclkp_1
flabel metal1 s 0 617 1536 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1536 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 1183 168 1217 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 SCE
port 3 nsew signal input
flabel locali s 1471 94 1505 128 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1471 168 1505 202 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1471 390 1505 424 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1471 464 1505 498 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1471 538 1505 572 0 FreeSans 340 0 0 0 GCLK
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1536 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1561250
string GDS_START 1548562
<< end >>
