magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2494 1852
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1137 203
rect 30 -17 64 21
<< scnmos >>
rect 89 47 119 177
rect 183 47 213 177
rect 277 47 307 177
rect 361 47 391 177
rect 455 47 485 177
rect 549 47 579 177
rect 643 47 673 177
rect 737 47 767 177
rect 831 47 861 177
rect 925 47 955 177
rect 1029 47 1059 177
<< scpmoshvt >>
rect 81 297 117 497
rect 175 297 211 497
rect 269 297 305 497
rect 363 297 399 497
rect 457 297 493 497
rect 551 297 587 497
rect 645 297 681 497
rect 739 297 775 497
rect 833 297 869 497
rect 927 297 963 497
rect 1021 297 1057 497
<< ndiff >>
rect 27 129 89 177
rect 27 95 35 129
rect 69 95 89 129
rect 27 47 89 95
rect 119 97 183 177
rect 119 63 129 97
rect 163 63 183 97
rect 119 47 183 63
rect 213 129 277 177
rect 213 95 223 129
rect 257 95 277 129
rect 213 47 277 95
rect 307 97 361 177
rect 307 63 317 97
rect 351 63 361 97
rect 307 47 361 63
rect 391 129 455 177
rect 391 95 411 129
rect 445 95 455 129
rect 391 47 455 95
rect 485 97 549 177
rect 485 63 505 97
rect 539 63 549 97
rect 485 47 549 63
rect 579 129 643 177
rect 579 95 599 129
rect 633 95 643 129
rect 579 47 643 95
rect 673 97 737 177
rect 673 63 693 97
rect 727 63 737 97
rect 673 47 737 63
rect 767 129 831 177
rect 767 95 787 129
rect 821 95 831 129
rect 767 47 831 95
rect 861 97 925 177
rect 861 63 881 97
rect 915 63 925 97
rect 861 47 925 63
rect 955 129 1029 177
rect 955 95 975 129
rect 1009 95 1029 129
rect 955 47 1029 95
rect 1059 161 1111 177
rect 1059 127 1069 161
rect 1103 127 1111 161
rect 1059 93 1111 127
rect 1059 59 1069 93
rect 1103 59 1111 93
rect 1059 47 1111 59
<< pdiff >>
rect 27 479 81 497
rect 27 445 35 479
rect 69 445 81 479
rect 27 411 81 445
rect 27 377 35 411
rect 69 377 81 411
rect 27 343 81 377
rect 27 309 35 343
rect 69 309 81 343
rect 27 297 81 309
rect 117 485 175 497
rect 117 451 129 485
rect 163 451 175 485
rect 117 417 175 451
rect 117 383 129 417
rect 163 383 175 417
rect 117 297 175 383
rect 211 479 269 497
rect 211 445 223 479
rect 257 445 269 479
rect 211 411 269 445
rect 211 377 223 411
rect 257 377 269 411
rect 211 343 269 377
rect 211 309 223 343
rect 257 309 269 343
rect 211 297 269 309
rect 305 485 363 497
rect 305 451 317 485
rect 351 451 363 485
rect 305 417 363 451
rect 305 383 317 417
rect 351 383 363 417
rect 305 297 363 383
rect 399 463 457 497
rect 399 429 411 463
rect 445 429 457 463
rect 399 368 457 429
rect 399 334 411 368
rect 445 334 457 368
rect 399 297 457 334
rect 493 485 551 497
rect 493 451 505 485
rect 539 451 551 485
rect 493 417 551 451
rect 493 383 505 417
rect 539 383 551 417
rect 493 297 551 383
rect 587 463 645 497
rect 587 429 599 463
rect 633 429 645 463
rect 587 368 645 429
rect 587 334 599 368
rect 633 334 645 368
rect 587 297 645 334
rect 681 485 739 497
rect 681 451 693 485
rect 727 451 739 485
rect 681 417 739 451
rect 681 383 693 417
rect 727 383 739 417
rect 681 297 739 383
rect 775 463 833 497
rect 775 429 787 463
rect 821 429 833 463
rect 775 368 833 429
rect 775 334 787 368
rect 821 334 833 368
rect 775 297 833 334
rect 869 485 927 497
rect 869 451 881 485
rect 915 451 927 485
rect 869 417 927 451
rect 869 383 881 417
rect 915 383 927 417
rect 869 297 927 383
rect 963 463 1021 497
rect 963 429 975 463
rect 1009 429 1021 463
rect 963 368 1021 429
rect 963 334 975 368
rect 1009 334 1021 368
rect 963 297 1021 334
rect 1057 485 1111 497
rect 1057 451 1069 485
rect 1103 451 1111 485
rect 1057 417 1111 451
rect 1057 383 1069 417
rect 1103 383 1111 417
rect 1057 349 1111 383
rect 1057 315 1069 349
rect 1103 315 1111 349
rect 1057 297 1111 315
<< ndiffc >>
rect 35 95 69 129
rect 129 63 163 97
rect 223 95 257 129
rect 317 63 351 97
rect 411 95 445 129
rect 505 63 539 97
rect 599 95 633 129
rect 693 63 727 97
rect 787 95 821 129
rect 881 63 915 97
rect 975 95 1009 129
rect 1069 127 1103 161
rect 1069 59 1103 93
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 129 451 163 485
rect 129 383 163 417
rect 223 445 257 479
rect 223 377 257 411
rect 223 309 257 343
rect 317 451 351 485
rect 317 383 351 417
rect 411 429 445 463
rect 411 334 445 368
rect 505 451 539 485
rect 505 383 539 417
rect 599 429 633 463
rect 599 334 633 368
rect 693 451 727 485
rect 693 383 727 417
rect 787 429 821 463
rect 787 334 821 368
rect 881 451 915 485
rect 881 383 915 417
rect 975 429 1009 463
rect 975 334 1009 368
rect 1069 451 1103 485
rect 1069 383 1103 417
rect 1069 315 1103 349
<< poly >>
rect 81 497 117 523
rect 175 497 211 523
rect 269 497 305 523
rect 363 497 399 523
rect 457 497 493 523
rect 551 497 587 523
rect 645 497 681 523
rect 739 497 775 523
rect 833 497 869 523
rect 927 497 963 523
rect 1021 497 1057 523
rect 81 282 117 297
rect 175 282 211 297
rect 269 282 305 297
rect 363 282 399 297
rect 457 282 493 297
rect 551 282 587 297
rect 645 282 681 297
rect 739 282 775 297
rect 833 282 869 297
rect 927 282 963 297
rect 1021 282 1057 297
rect 79 261 119 282
rect 28 259 119 261
rect 173 259 213 282
rect 267 259 307 282
rect 28 249 307 259
rect 28 215 44 249
rect 78 215 122 249
rect 156 215 190 249
rect 224 215 307 249
rect 28 205 307 215
rect 28 203 119 205
rect 89 177 119 203
rect 183 177 213 205
rect 277 177 307 205
rect 361 259 401 282
rect 455 259 495 282
rect 549 259 589 282
rect 643 259 683 282
rect 737 259 777 282
rect 831 259 871 282
rect 925 259 965 282
rect 1019 259 1059 282
rect 361 249 1059 259
rect 361 215 381 249
rect 415 215 459 249
rect 493 215 537 249
rect 571 215 615 249
rect 649 215 693 249
rect 727 215 761 249
rect 795 215 839 249
rect 873 215 1059 249
rect 361 205 1059 215
rect 361 177 391 205
rect 455 177 485 205
rect 549 177 579 205
rect 643 177 673 205
rect 737 177 767 205
rect 831 177 861 205
rect 925 177 955 205
rect 1029 177 1059 205
rect 89 21 119 47
rect 183 21 213 47
rect 277 21 307 47
rect 361 21 391 47
rect 455 21 485 47
rect 549 21 579 47
rect 643 21 673 47
rect 737 21 767 47
rect 831 21 861 47
rect 925 21 955 47
rect 1029 21 1059 47
<< polycont >>
rect 44 215 78 249
rect 122 215 156 249
rect 190 215 224 249
rect 381 215 415 249
rect 459 215 493 249
rect 537 215 571 249
rect 615 215 649 249
rect 693 215 727 249
rect 761 215 795 249
rect 839 215 873 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 19 479 85 493
rect 19 445 35 479
rect 69 445 85 479
rect 19 411 85 445
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 129 485 163 527
rect 129 417 163 451
rect 129 367 163 383
rect 197 479 273 493
rect 197 445 223 479
rect 257 445 273 479
rect 197 411 273 445
rect 197 377 223 411
rect 257 377 273 411
rect 19 309 35 343
rect 69 323 85 343
rect 197 343 273 377
rect 317 485 351 527
rect 317 417 351 451
rect 317 367 351 383
rect 411 463 445 493
rect 411 368 445 429
rect 197 323 223 343
rect 69 309 223 323
rect 257 323 273 343
rect 479 485 555 527
rect 479 451 505 485
rect 539 451 555 485
rect 479 417 555 451
rect 479 383 505 417
rect 539 383 555 417
rect 479 367 555 383
rect 599 463 633 493
rect 599 368 633 429
rect 411 323 445 334
rect 667 485 743 527
rect 667 451 693 485
rect 727 451 743 485
rect 667 417 743 451
rect 667 383 693 417
rect 727 383 743 417
rect 667 367 743 383
rect 787 463 821 493
rect 787 368 821 429
rect 599 323 633 334
rect 855 485 931 527
rect 855 451 881 485
rect 915 451 931 485
rect 855 417 931 451
rect 855 383 881 417
rect 915 383 931 417
rect 855 367 931 383
rect 975 463 1009 493
rect 975 368 1009 429
rect 787 323 821 334
rect 975 323 1009 334
rect 257 309 349 323
rect 19 289 349 309
rect 411 289 1009 323
rect 1043 485 1119 527
rect 1043 451 1069 485
rect 1103 451 1119 485
rect 1043 417 1119 451
rect 1043 383 1069 417
rect 1103 383 1119 417
rect 1043 349 1119 383
rect 1043 315 1069 349
rect 1103 315 1119 349
rect 1043 297 1119 315
rect 28 249 268 255
rect 28 215 44 249
rect 78 215 122 249
rect 156 215 190 249
rect 224 215 268 249
rect 314 249 349 289
rect 314 215 381 249
rect 415 215 459 249
rect 493 215 537 249
rect 571 215 615 249
rect 649 215 693 249
rect 727 215 761 249
rect 795 215 839 249
rect 873 215 899 249
rect 314 181 349 215
rect 938 181 1009 289
rect 35 147 349 181
rect 411 147 1009 181
rect 35 129 69 147
rect 223 129 257 147
rect 35 51 69 95
rect 103 97 179 113
rect 103 63 129 97
rect 163 63 179 97
rect 103 17 179 63
rect 411 129 445 147
rect 223 52 257 95
rect 291 97 367 113
rect 291 63 317 97
rect 351 63 367 97
rect 291 17 367 63
rect 599 129 633 147
rect 411 51 445 95
rect 479 97 555 113
rect 479 63 505 97
rect 539 63 555 97
rect 479 17 555 63
rect 787 129 821 147
rect 599 51 633 95
rect 667 97 743 113
rect 667 63 693 97
rect 727 63 743 97
rect 667 17 743 63
rect 975 129 1009 147
rect 787 51 821 95
rect 855 97 931 113
rect 855 63 881 97
rect 915 63 931 97
rect 855 17 931 63
rect 975 51 1009 95
rect 1043 161 1119 177
rect 1043 127 1069 161
rect 1103 127 1119 161
rect 1043 93 1119 127
rect 1043 59 1069 93
rect 1103 59 1119 93
rect 1043 17 1119 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 28 215 268 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 949 153 983 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 949 221 983 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 120 221 154 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel locali s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional
flabel locali s 949 289 983 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 buf_8
rlabel metal1 s 0 -48 1196 48 1 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 496 1196 592 1 VPWR
port 5 nsew power bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1196 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1957900
string GDS_START 1948556
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
