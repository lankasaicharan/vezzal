magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 552 241 862 249
rect 1 49 862 241
rect 0 0 864 49
<< scnmos >>
rect 96 47 126 215
rect 184 47 214 215
rect 284 47 314 215
rect 384 47 414 215
rect 635 139 665 223
rect 749 139 779 223
<< scpmoshvt >>
rect 96 367 126 619
rect 182 367 212 619
rect 268 367 298 619
rect 354 367 384 619
rect 599 427 629 555
rect 742 491 772 619
<< ndiff >>
rect 27 125 96 215
rect 27 91 39 125
rect 73 91 96 125
rect 27 47 96 91
rect 126 178 184 215
rect 126 144 139 178
rect 173 144 184 178
rect 126 47 184 144
rect 214 203 284 215
rect 214 169 239 203
rect 273 169 284 203
rect 214 101 284 169
rect 214 67 239 101
rect 273 67 284 101
rect 214 47 284 67
rect 314 117 384 215
rect 314 83 325 117
rect 359 83 384 117
rect 314 47 384 83
rect 414 203 471 215
rect 414 169 425 203
rect 459 169 471 203
rect 414 101 471 169
rect 414 67 425 101
rect 459 67 471 101
rect 414 47 471 67
rect 578 206 635 223
rect 578 172 590 206
rect 624 172 635 206
rect 578 139 635 172
rect 665 198 749 223
rect 665 164 690 198
rect 724 164 749 198
rect 665 139 749 164
rect 779 198 836 223
rect 779 164 790 198
rect 824 164 836 198
rect 779 139 836 164
<< pdiff >>
rect 39 607 96 619
rect 39 573 51 607
rect 85 573 96 607
rect 39 534 96 573
rect 39 500 51 534
rect 85 500 96 534
rect 39 461 96 500
rect 39 427 51 461
rect 85 427 96 461
rect 39 367 96 427
rect 126 531 182 619
rect 126 497 137 531
rect 171 497 182 531
rect 126 413 182 497
rect 126 379 137 413
rect 171 379 182 413
rect 126 367 182 379
rect 212 599 268 619
rect 212 565 223 599
rect 257 565 268 599
rect 212 506 268 565
rect 212 472 223 506
rect 257 472 268 506
rect 212 413 268 472
rect 212 379 223 413
rect 257 379 268 413
rect 212 367 268 379
rect 298 607 354 619
rect 298 573 309 607
rect 343 573 354 607
rect 298 481 354 573
rect 298 447 309 481
rect 343 447 354 481
rect 298 367 354 447
rect 384 599 441 619
rect 384 565 395 599
rect 429 565 441 599
rect 671 607 742 619
rect 384 506 441 565
rect 671 573 683 607
rect 717 573 742 607
rect 671 555 742 573
rect 384 472 395 506
rect 429 472 441 506
rect 384 413 441 472
rect 519 473 599 555
rect 519 439 531 473
rect 565 439 599 473
rect 519 427 599 439
rect 629 491 742 555
rect 772 568 829 619
rect 772 534 783 568
rect 817 534 829 568
rect 772 491 829 534
rect 629 427 679 491
rect 384 379 395 413
rect 429 379 441 413
rect 384 367 441 379
<< ndiffc >>
rect 39 91 73 125
rect 139 144 173 178
rect 239 169 273 203
rect 239 67 273 101
rect 325 83 359 117
rect 425 169 459 203
rect 425 67 459 101
rect 590 172 624 206
rect 690 164 724 198
rect 790 164 824 198
<< pdiffc >>
rect 51 573 85 607
rect 51 500 85 534
rect 51 427 85 461
rect 137 497 171 531
rect 137 379 171 413
rect 223 565 257 599
rect 223 472 257 506
rect 223 379 257 413
rect 309 573 343 607
rect 309 447 343 481
rect 395 565 429 599
rect 683 573 717 607
rect 395 472 429 506
rect 531 439 565 473
rect 783 534 817 568
rect 395 379 429 413
<< poly >>
rect 96 619 126 645
rect 182 619 212 645
rect 268 619 298 645
rect 354 619 384 645
rect 742 619 772 645
rect 599 555 629 581
rect 599 395 629 427
rect 742 395 772 491
rect 599 379 665 395
rect 96 325 126 367
rect 182 325 212 367
rect 268 345 298 367
rect 354 345 384 367
rect 599 345 615 379
rect 649 345 665 379
rect 96 309 214 325
rect 268 315 665 345
rect 96 275 164 309
rect 198 275 214 309
rect 96 259 214 275
rect 599 311 665 315
rect 599 277 615 311
rect 649 277 665 311
rect 96 215 126 259
rect 184 215 214 259
rect 284 237 551 267
rect 599 261 665 277
rect 713 379 779 395
rect 713 345 729 379
rect 763 345 779 379
rect 713 311 779 345
rect 713 277 729 311
rect 763 277 779 311
rect 713 261 779 277
rect 284 215 314 237
rect 384 215 414 237
rect 521 117 551 237
rect 635 223 665 261
rect 749 223 779 261
rect 521 101 587 117
rect 635 113 665 139
rect 749 113 779 139
rect 521 67 537 101
rect 571 67 587 101
rect 521 51 587 67
rect 96 21 126 47
rect 184 21 214 47
rect 284 21 314 47
rect 384 21 414 47
<< polycont >>
rect 615 345 649 379
rect 164 275 198 309
rect 615 277 649 311
rect 729 345 763 379
rect 729 277 763 311
rect 537 67 571 101
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 35 607 273 615
rect 35 573 51 607
rect 85 599 273 607
rect 85 581 223 599
rect 85 573 101 581
rect 35 534 101 573
rect 207 565 223 581
rect 257 565 273 599
rect 35 500 51 534
rect 85 500 101 534
rect 35 461 101 500
rect 35 427 51 461
rect 85 427 101 461
rect 137 531 171 547
rect 137 413 171 497
rect 25 379 137 393
rect 25 359 171 379
rect 207 506 273 565
rect 207 472 223 506
rect 257 472 273 506
rect 207 413 273 472
rect 309 607 343 649
rect 309 481 343 573
rect 309 431 343 447
rect 379 599 429 615
rect 379 565 395 599
rect 379 506 429 565
rect 667 607 733 649
rect 667 573 683 607
rect 717 573 733 607
rect 667 557 733 573
rect 767 568 847 615
rect 379 472 395 506
rect 207 379 223 413
rect 257 397 273 413
rect 379 413 429 472
rect 379 397 395 413
rect 257 379 395 397
rect 207 363 429 379
rect 463 523 633 557
rect 767 534 783 568
rect 817 534 847 568
rect 767 523 847 534
rect 25 225 71 359
rect 463 325 497 523
rect 599 489 847 523
rect 148 309 497 325
rect 148 275 164 309
rect 198 275 497 309
rect 148 259 497 275
rect 531 473 565 489
rect 767 487 847 489
rect 531 227 565 439
rect 599 379 665 430
rect 599 345 615 379
rect 649 345 665 379
rect 599 311 665 345
rect 599 277 615 311
rect 649 277 665 311
rect 599 261 665 277
rect 701 379 779 430
rect 701 345 729 379
rect 763 345 779 379
rect 701 311 779 345
rect 701 277 729 311
rect 763 277 779 311
rect 701 261 779 277
rect 813 227 847 487
rect 25 191 189 225
rect 123 178 189 191
rect 23 125 89 157
rect 23 91 39 125
rect 73 91 89 125
rect 123 144 139 178
rect 173 144 189 178
rect 123 119 189 144
rect 223 203 475 225
rect 223 169 239 203
rect 273 191 425 203
rect 273 169 289 191
rect 23 85 89 91
rect 223 101 289 169
rect 409 169 425 191
rect 459 169 475 203
rect 223 85 239 101
rect 23 67 239 85
rect 273 67 289 101
rect 23 51 289 67
rect 325 117 375 157
rect 359 83 375 117
rect 325 17 375 83
rect 409 101 475 169
rect 531 206 640 227
rect 531 172 590 206
rect 624 172 640 206
rect 531 117 640 172
rect 409 67 425 101
rect 459 67 475 101
rect 409 51 475 67
rect 521 101 640 117
rect 521 67 537 101
rect 571 67 640 101
rect 521 51 640 67
rect 674 198 740 227
rect 674 164 690 198
rect 724 164 740 198
rect 674 17 740 164
rect 774 198 847 227
rect 774 164 790 198
rect 824 164 847 198
rect 774 135 847 164
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 ebufn_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 TE_B
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3331970
string GDS_START 3324732
<< end >>
