magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 332 2054 704
<< pwell >>
rect 1 49 2015 248
rect 0 0 2016 49
<< scpmos >>
rect 83 368 119 592
rect 193 368 229 592
rect 395 368 431 592
rect 485 368 521 592
rect 575 368 611 592
rect 665 368 701 592
rect 755 368 791 592
rect 865 368 901 592
rect 955 368 991 592
rect 1045 368 1081 592
rect 1247 368 1283 592
rect 1337 368 1373 592
rect 1427 368 1463 592
rect 1517 368 1553 592
rect 1607 368 1643 592
rect 1707 368 1743 592
rect 1797 368 1833 592
rect 1897 368 1933 592
<< nmoslvt >>
rect 84 74 114 222
rect 170 74 200 222
rect 256 74 286 222
rect 356 74 386 222
rect 456 74 486 222
rect 602 74 632 222
rect 693 74 723 222
rect 779 74 809 222
rect 865 74 895 222
rect 965 74 995 222
rect 1051 74 1081 222
rect 1151 74 1181 222
rect 1237 74 1267 222
rect 1337 74 1367 222
rect 1423 74 1453 222
rect 1516 74 1546 222
rect 1613 74 1643 222
rect 1716 74 1746 222
rect 1802 74 1832 222
rect 1902 74 1932 222
<< ndiff >>
rect 27 202 84 222
rect 27 168 39 202
rect 73 168 84 202
rect 27 120 84 168
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 177 170 222
rect 114 143 125 177
rect 159 143 170 177
rect 114 74 170 143
rect 200 127 256 222
rect 200 93 211 127
rect 245 93 256 127
rect 200 74 256 93
rect 286 189 356 222
rect 286 155 311 189
rect 345 155 356 189
rect 286 74 356 155
rect 386 202 456 222
rect 386 168 411 202
rect 445 168 456 202
rect 386 120 456 168
rect 386 86 411 120
rect 445 86 456 120
rect 386 74 456 86
rect 486 120 602 222
rect 486 86 529 120
rect 563 86 602 120
rect 486 74 602 86
rect 632 202 693 222
rect 632 168 648 202
rect 682 168 693 202
rect 632 120 693 168
rect 632 86 648 120
rect 682 86 693 120
rect 632 74 693 86
rect 723 210 779 222
rect 723 176 734 210
rect 768 176 779 210
rect 723 120 779 176
rect 723 86 734 120
rect 768 86 779 120
rect 723 74 779 86
rect 809 202 865 222
rect 809 168 820 202
rect 854 168 865 202
rect 809 120 865 168
rect 809 86 820 120
rect 854 86 865 120
rect 809 74 865 86
rect 895 127 965 222
rect 895 93 920 127
rect 954 93 965 127
rect 895 74 965 93
rect 995 202 1051 222
rect 995 168 1006 202
rect 1040 168 1051 202
rect 995 120 1051 168
rect 995 86 1006 120
rect 1040 86 1051 120
rect 995 74 1051 86
rect 1081 127 1151 222
rect 1081 93 1106 127
rect 1140 93 1151 127
rect 1081 74 1151 93
rect 1181 202 1237 222
rect 1181 168 1192 202
rect 1226 168 1237 202
rect 1181 120 1237 168
rect 1181 86 1192 120
rect 1226 86 1237 120
rect 1181 74 1237 86
rect 1267 127 1337 222
rect 1267 93 1292 127
rect 1326 93 1337 127
rect 1267 74 1337 93
rect 1367 202 1423 222
rect 1367 168 1378 202
rect 1412 168 1423 202
rect 1367 120 1423 168
rect 1367 86 1378 120
rect 1412 86 1423 120
rect 1367 74 1423 86
rect 1453 127 1516 222
rect 1453 93 1464 127
rect 1498 93 1516 127
rect 1453 74 1516 93
rect 1546 202 1613 222
rect 1546 168 1557 202
rect 1591 168 1613 202
rect 1546 120 1613 168
rect 1546 86 1557 120
rect 1591 86 1613 120
rect 1546 74 1613 86
rect 1643 127 1716 222
rect 1643 93 1657 127
rect 1691 93 1716 127
rect 1643 74 1716 93
rect 1746 202 1802 222
rect 1746 168 1757 202
rect 1791 168 1802 202
rect 1746 120 1802 168
rect 1746 86 1757 120
rect 1791 86 1802 120
rect 1746 74 1802 86
rect 1832 127 1902 222
rect 1832 93 1857 127
rect 1891 93 1902 127
rect 1832 74 1902 93
rect 1932 202 1989 222
rect 1932 168 1943 202
rect 1977 168 1989 202
rect 1932 120 1989 168
rect 1932 86 1943 120
rect 1977 86 1989 120
rect 1932 74 1989 86
<< pdiff >>
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 497 83 546
rect 27 463 39 497
rect 73 463 83 497
rect 27 414 83 463
rect 27 380 39 414
rect 73 380 83 414
rect 27 368 83 380
rect 119 580 193 592
rect 119 546 139 580
rect 173 546 193 580
rect 119 497 193 546
rect 119 463 139 497
rect 173 463 193 497
rect 119 414 193 463
rect 119 380 139 414
rect 173 380 193 414
rect 119 368 193 380
rect 229 580 285 592
rect 229 546 239 580
rect 273 546 285 580
rect 229 462 285 546
rect 229 428 239 462
rect 273 428 285 462
rect 229 368 285 428
rect 339 584 395 592
rect 339 550 351 584
rect 385 550 395 584
rect 339 462 395 550
rect 339 428 351 462
rect 385 428 395 462
rect 339 368 395 428
rect 431 531 485 592
rect 431 497 441 531
rect 475 497 485 531
rect 431 410 485 497
rect 431 376 441 410
rect 475 376 485 410
rect 431 368 485 376
rect 521 584 575 592
rect 521 550 531 584
rect 565 550 575 584
rect 521 514 575 550
rect 521 480 531 514
rect 565 480 575 514
rect 521 368 575 480
rect 611 531 665 592
rect 611 497 621 531
rect 655 497 665 531
rect 611 410 665 497
rect 611 376 621 410
rect 655 376 665 410
rect 611 368 665 376
rect 701 584 755 592
rect 701 550 711 584
rect 745 550 755 584
rect 701 497 755 550
rect 701 463 711 497
rect 745 463 755 497
rect 701 410 755 463
rect 701 376 711 410
rect 745 376 755 410
rect 701 368 755 376
rect 791 531 865 592
rect 791 497 811 531
rect 845 497 865 531
rect 791 426 865 497
rect 791 392 811 426
rect 845 392 865 426
rect 791 368 865 392
rect 901 584 955 592
rect 901 550 911 584
rect 945 550 955 584
rect 901 446 955 550
rect 901 412 911 446
rect 945 412 955 446
rect 901 368 955 412
rect 991 531 1045 592
rect 991 497 1001 531
rect 1035 497 1045 531
rect 991 410 1045 497
rect 991 376 1001 410
rect 1035 376 1045 410
rect 991 368 1045 376
rect 1081 584 1137 592
rect 1081 550 1091 584
rect 1125 550 1137 584
rect 1081 446 1137 550
rect 1081 412 1091 446
rect 1125 412 1137 446
rect 1081 368 1137 412
rect 1191 584 1247 592
rect 1191 550 1203 584
rect 1237 550 1247 584
rect 1191 446 1247 550
rect 1191 412 1203 446
rect 1237 412 1247 446
rect 1191 368 1247 412
rect 1283 528 1337 592
rect 1283 494 1293 528
rect 1327 494 1337 528
rect 1283 410 1337 494
rect 1283 376 1293 410
rect 1327 376 1337 410
rect 1283 368 1337 376
rect 1373 584 1427 592
rect 1373 550 1383 584
rect 1417 550 1427 584
rect 1373 446 1427 550
rect 1373 412 1383 446
rect 1417 412 1427 446
rect 1373 368 1427 412
rect 1463 531 1517 592
rect 1463 497 1473 531
rect 1507 497 1517 531
rect 1463 426 1517 497
rect 1463 392 1473 426
rect 1507 392 1517 426
rect 1463 368 1517 392
rect 1553 584 1607 592
rect 1553 550 1563 584
rect 1597 550 1607 584
rect 1553 497 1607 550
rect 1553 463 1563 497
rect 1597 463 1607 497
rect 1553 410 1607 463
rect 1553 376 1563 410
rect 1597 376 1607 410
rect 1553 368 1607 376
rect 1643 579 1707 592
rect 1643 545 1653 579
rect 1687 545 1707 579
rect 1643 462 1707 545
rect 1643 428 1653 462
rect 1687 428 1707 462
rect 1643 368 1707 428
rect 1743 584 1797 592
rect 1743 550 1753 584
rect 1787 550 1797 584
rect 1743 497 1797 550
rect 1743 463 1753 497
rect 1787 463 1797 497
rect 1743 410 1797 463
rect 1743 376 1753 410
rect 1787 376 1797 410
rect 1743 368 1797 376
rect 1833 579 1897 592
rect 1833 545 1853 579
rect 1887 545 1897 579
rect 1833 462 1897 545
rect 1833 428 1853 462
rect 1887 428 1897 462
rect 1833 368 1897 428
rect 1933 584 1989 592
rect 1933 550 1943 584
rect 1977 550 1989 584
rect 1933 497 1989 550
rect 1933 463 1943 497
rect 1977 463 1989 497
rect 1933 410 1989 463
rect 1933 376 1943 410
rect 1977 376 1989 410
rect 1933 368 1989 376
<< ndiffc >>
rect 39 168 73 202
rect 39 86 73 120
rect 125 143 159 177
rect 211 93 245 127
rect 311 155 345 189
rect 411 168 445 202
rect 411 86 445 120
rect 529 86 563 120
rect 648 168 682 202
rect 648 86 682 120
rect 734 176 768 210
rect 734 86 768 120
rect 820 168 854 202
rect 820 86 854 120
rect 920 93 954 127
rect 1006 168 1040 202
rect 1006 86 1040 120
rect 1106 93 1140 127
rect 1192 168 1226 202
rect 1192 86 1226 120
rect 1292 93 1326 127
rect 1378 168 1412 202
rect 1378 86 1412 120
rect 1464 93 1498 127
rect 1557 168 1591 202
rect 1557 86 1591 120
rect 1657 93 1691 127
rect 1757 168 1791 202
rect 1757 86 1791 120
rect 1857 93 1891 127
rect 1943 168 1977 202
rect 1943 86 1977 120
<< pdiffc >>
rect 39 546 73 580
rect 39 463 73 497
rect 39 380 73 414
rect 139 546 173 580
rect 139 463 173 497
rect 139 380 173 414
rect 239 546 273 580
rect 239 428 273 462
rect 351 550 385 584
rect 351 428 385 462
rect 441 497 475 531
rect 441 376 475 410
rect 531 550 565 584
rect 531 480 565 514
rect 621 497 655 531
rect 621 376 655 410
rect 711 550 745 584
rect 711 463 745 497
rect 711 376 745 410
rect 811 497 845 531
rect 811 392 845 426
rect 911 550 945 584
rect 911 412 945 446
rect 1001 497 1035 531
rect 1001 376 1035 410
rect 1091 550 1125 584
rect 1091 412 1125 446
rect 1203 550 1237 584
rect 1203 412 1237 446
rect 1293 494 1327 528
rect 1293 376 1327 410
rect 1383 550 1417 584
rect 1383 412 1417 446
rect 1473 497 1507 531
rect 1473 392 1507 426
rect 1563 550 1597 584
rect 1563 463 1597 497
rect 1563 376 1597 410
rect 1653 545 1687 579
rect 1653 428 1687 462
rect 1753 550 1787 584
rect 1753 463 1787 497
rect 1753 376 1787 410
rect 1853 545 1887 579
rect 1853 428 1887 462
rect 1943 550 1977 584
rect 1943 463 1977 497
rect 1943 376 1977 410
<< poly >>
rect 83 592 119 618
rect 193 592 229 618
rect 395 592 431 618
rect 485 592 521 618
rect 575 592 611 618
rect 665 592 701 618
rect 755 592 791 618
rect 865 592 901 618
rect 955 592 991 618
rect 1045 592 1081 618
rect 1247 592 1283 618
rect 1337 592 1373 618
rect 1427 592 1463 618
rect 1517 592 1553 618
rect 1607 592 1643 618
rect 1707 592 1743 618
rect 1797 592 1833 618
rect 1897 592 1933 618
rect 83 310 119 368
rect 193 310 229 368
rect 395 345 431 368
rect 485 345 521 368
rect 575 345 611 368
rect 665 345 701 368
rect 395 315 701 345
rect 755 345 791 368
rect 865 345 901 368
rect 955 345 991 368
rect 1045 345 1081 368
rect 755 315 1081 345
rect 27 294 229 310
rect 27 260 43 294
rect 77 260 111 294
rect 145 260 179 294
rect 213 267 229 294
rect 430 294 701 315
rect 213 260 386 267
rect 27 237 386 260
rect 430 260 446 294
rect 480 260 514 294
rect 548 260 582 294
rect 616 267 701 294
rect 865 310 1081 315
rect 1247 310 1283 368
rect 1337 310 1373 368
rect 1427 310 1463 368
rect 1517 310 1553 368
rect 1607 310 1643 368
rect 1707 310 1743 368
rect 1797 310 1833 368
rect 1897 310 1933 368
rect 865 294 1149 310
rect 616 260 809 267
rect 430 237 809 260
rect 84 222 114 237
rect 170 222 200 237
rect 256 222 286 237
rect 356 222 386 237
rect 456 222 486 237
rect 602 222 632 237
rect 693 222 723 237
rect 779 222 809 237
rect 865 260 895 294
rect 929 260 963 294
rect 997 260 1031 294
rect 1065 260 1099 294
rect 1133 277 1149 294
rect 1237 294 1553 310
rect 1133 260 1181 277
rect 865 244 1181 260
rect 865 222 895 244
rect 965 222 995 244
rect 1051 222 1081 244
rect 1151 222 1181 244
rect 1237 260 1289 294
rect 1323 260 1357 294
rect 1391 260 1425 294
rect 1459 260 1493 294
rect 1527 260 1553 294
rect 1237 244 1553 260
rect 1613 294 1933 310
rect 1613 260 1673 294
rect 1707 260 1741 294
rect 1775 260 1809 294
rect 1843 260 1877 294
rect 1911 260 1933 294
rect 1613 244 1933 260
rect 1237 222 1267 244
rect 1337 222 1367 244
rect 1423 222 1453 244
rect 1516 222 1546 244
rect 1613 222 1643 244
rect 1716 222 1746 244
rect 1802 222 1832 244
rect 1902 222 1932 244
rect 84 48 114 74
rect 170 48 200 74
rect 256 48 286 74
rect 356 48 386 74
rect 456 48 486 74
rect 602 48 632 74
rect 693 48 723 74
rect 779 48 809 74
rect 865 48 895 74
rect 965 48 995 74
rect 1051 48 1081 74
rect 1151 48 1181 74
rect 1237 48 1267 74
rect 1337 48 1367 74
rect 1423 48 1453 74
rect 1516 48 1546 74
rect 1613 48 1643 74
rect 1716 48 1746 74
rect 1802 48 1832 74
rect 1902 48 1932 74
<< polycont >>
rect 43 260 77 294
rect 111 260 145 294
rect 179 260 213 294
rect 446 260 480 294
rect 514 260 548 294
rect 582 260 616 294
rect 895 260 929 294
rect 963 260 997 294
rect 1031 260 1065 294
rect 1099 260 1133 294
rect 1289 260 1323 294
rect 1357 260 1391 294
rect 1425 260 1459 294
rect 1493 260 1527 294
rect 1673 260 1707 294
rect 1741 260 1775 294
rect 1809 260 1843 294
rect 1877 260 1911 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 23 580 89 649
rect 23 546 39 580
rect 73 546 89 580
rect 23 497 89 546
rect 23 463 39 497
rect 73 463 89 497
rect 23 414 89 463
rect 23 380 39 414
rect 73 380 89 414
rect 23 364 89 380
rect 123 580 189 596
rect 123 546 139 580
rect 173 546 189 580
rect 123 497 189 546
rect 123 463 139 497
rect 173 463 189 497
rect 123 414 189 463
rect 123 380 139 414
rect 173 380 189 414
rect 223 580 289 649
rect 223 546 239 580
rect 273 546 289 580
rect 223 462 289 546
rect 223 428 239 462
rect 273 428 289 462
rect 223 412 289 428
rect 335 584 1141 615
rect 335 550 351 584
rect 385 581 531 584
rect 385 550 396 581
rect 335 462 396 550
rect 520 550 531 581
rect 565 581 711 584
rect 565 550 576 581
rect 335 428 351 462
rect 385 428 396 462
rect 335 412 396 428
rect 430 531 486 547
rect 430 497 441 531
rect 475 497 486 531
rect 430 430 486 497
rect 520 514 576 550
rect 700 550 711 581
rect 745 581 911 584
rect 745 550 761 581
rect 520 480 531 514
rect 565 480 576 514
rect 520 464 576 480
rect 610 531 666 547
rect 610 497 621 531
rect 655 497 666 531
rect 610 430 666 497
rect 123 378 189 380
rect 430 410 666 430
rect 430 378 441 410
rect 123 376 441 378
rect 475 376 621 410
rect 655 376 666 410
rect 123 344 666 376
rect 700 497 761 550
rect 895 550 911 581
rect 945 581 1091 584
rect 945 550 961 581
rect 700 463 711 497
rect 745 463 761 497
rect 700 410 761 463
rect 700 376 711 410
rect 745 376 761 410
rect 700 360 761 376
rect 795 531 861 547
rect 795 497 811 531
rect 845 497 861 531
rect 795 426 861 497
rect 795 392 811 426
rect 845 392 861 426
rect 895 446 961 550
rect 1075 550 1091 581
rect 1125 550 1141 584
rect 895 412 911 446
rect 945 412 961 446
rect 995 531 1041 547
rect 995 497 1001 531
rect 1035 497 1041 531
rect 795 378 861 392
rect 995 410 1041 497
rect 1075 446 1141 550
rect 1075 412 1091 446
rect 1125 412 1141 446
rect 1187 584 1603 615
rect 1187 550 1203 584
rect 1237 578 1383 584
rect 1237 550 1253 578
rect 1187 446 1253 550
rect 1367 550 1383 578
rect 1417 581 1563 584
rect 1417 550 1433 581
rect 1187 412 1203 446
rect 1237 412 1253 446
rect 1287 528 1333 544
rect 1287 494 1293 528
rect 1327 494 1333 528
rect 995 378 1001 410
rect 795 376 1001 378
rect 1035 378 1041 410
rect 1287 410 1333 494
rect 1367 446 1433 550
rect 1547 550 1563 581
rect 1597 550 1603 584
rect 1367 412 1383 446
rect 1417 412 1433 446
rect 1467 531 1513 547
rect 1467 497 1473 531
rect 1507 497 1513 531
rect 1467 426 1513 497
rect 1287 378 1293 410
rect 1035 376 1293 378
rect 1327 378 1333 410
rect 1467 392 1473 426
rect 1507 392 1513 426
rect 1467 378 1513 392
rect 1327 376 1513 378
rect 795 344 1513 376
rect 1547 497 1603 550
rect 1547 463 1563 497
rect 1597 463 1603 497
rect 1547 410 1603 463
rect 1637 579 1703 649
rect 1637 545 1653 579
rect 1687 545 1703 579
rect 1637 462 1703 545
rect 1637 428 1653 462
rect 1687 428 1703 462
rect 1637 412 1703 428
rect 1737 584 1803 600
rect 1737 550 1753 584
rect 1787 550 1803 584
rect 1737 497 1803 550
rect 1737 463 1753 497
rect 1787 463 1803 497
rect 1547 376 1563 410
rect 1597 378 1603 410
rect 1737 410 1803 463
rect 1837 579 1903 649
rect 1837 545 1853 579
rect 1887 545 1903 579
rect 1837 462 1903 545
rect 1837 428 1853 462
rect 1887 428 1903 462
rect 1837 412 1903 428
rect 1937 584 1993 600
rect 1937 550 1943 584
rect 1977 550 1993 584
rect 1937 497 1993 550
rect 1937 463 1943 497
rect 1977 463 1993 497
rect 1737 378 1753 410
rect 1597 376 1753 378
rect 1787 378 1803 410
rect 1937 410 1993 463
rect 1937 378 1943 410
rect 1787 376 1943 378
rect 1977 376 1993 410
rect 1547 344 1993 376
rect 25 294 229 310
rect 25 260 43 294
rect 77 260 111 294
rect 145 260 179 294
rect 213 260 229 294
rect 25 236 229 260
rect 295 202 361 344
rect 409 294 632 310
rect 879 294 1223 310
rect 409 260 446 294
rect 480 260 514 294
rect 548 260 582 294
rect 616 260 632 294
rect 409 236 632 260
rect 666 260 838 294
rect 666 202 700 260
rect 23 168 39 202
rect 73 168 89 202
rect 23 120 89 168
rect 23 86 39 120
rect 73 86 89 120
rect 125 189 361 202
rect 125 177 311 189
rect 159 168 311 177
rect 125 119 159 143
rect 295 155 311 168
rect 345 155 361 189
rect 195 127 261 134
rect 23 85 89 86
rect 195 93 211 127
rect 245 93 261 127
rect 295 119 361 155
rect 395 168 411 202
rect 445 168 648 202
rect 682 168 700 202
rect 395 120 461 168
rect 632 120 700 168
rect 195 85 261 93
rect 395 86 411 120
rect 445 86 461 120
rect 395 85 461 86
rect 23 51 461 85
rect 495 86 529 120
rect 563 86 598 120
rect 495 17 598 86
rect 632 86 648 120
rect 682 86 700 120
rect 632 70 700 86
rect 734 210 768 226
rect 734 120 768 176
rect 734 17 768 86
rect 804 202 838 260
rect 879 260 895 294
rect 929 260 963 294
rect 997 260 1031 294
rect 1065 260 1099 294
rect 1133 260 1223 294
rect 879 236 1223 260
rect 1273 294 1607 310
rect 1273 260 1289 294
rect 1323 260 1357 294
rect 1391 260 1425 294
rect 1459 260 1493 294
rect 1527 260 1607 294
rect 1273 236 1607 260
rect 1657 294 1991 310
rect 1657 260 1673 294
rect 1707 260 1741 294
rect 1775 260 1809 294
rect 1843 260 1877 294
rect 1911 260 1991 294
rect 1657 236 1991 260
rect 804 168 820 202
rect 854 168 1006 202
rect 1040 168 1192 202
rect 1226 168 1378 202
rect 1412 168 1557 202
rect 1591 168 1757 202
rect 1791 168 1943 202
rect 1977 168 1993 202
rect 804 120 870 168
rect 804 86 820 120
rect 854 86 870 120
rect 804 70 870 86
rect 904 127 970 134
rect 904 93 920 127
rect 954 93 970 127
rect 904 17 970 93
rect 1006 120 1056 168
rect 1040 86 1056 120
rect 1006 70 1056 86
rect 1090 127 1156 134
rect 1090 93 1106 127
rect 1140 93 1156 127
rect 1090 17 1156 93
rect 1192 120 1242 168
rect 1226 86 1242 120
rect 1192 70 1242 86
rect 1276 127 1342 134
rect 1276 93 1292 127
rect 1326 93 1342 127
rect 1276 17 1342 93
rect 1378 120 1412 168
rect 1378 70 1412 86
rect 1448 127 1514 134
rect 1448 93 1464 127
rect 1498 93 1514 127
rect 1448 17 1514 93
rect 1557 120 1607 168
rect 1591 86 1607 120
rect 1557 70 1607 86
rect 1641 127 1707 134
rect 1641 93 1657 127
rect 1691 93 1707 127
rect 1641 17 1707 93
rect 1741 120 1807 168
rect 1741 86 1757 120
rect 1791 86 1807 120
rect 1741 70 1807 86
rect 1841 127 1907 134
rect 1841 93 1857 127
rect 1891 93 1907 127
rect 1841 17 1907 93
rect 1943 120 1993 168
rect 1977 86 1993 120
rect 1943 70 1993 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o41ai_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A4
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B1
port 5 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 3553104
string GDS_START 3536950
<< end >>
