magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 4 49 657 241
rect 0 0 672 49
<< scnmos >>
rect 83 47 113 215
rect 169 47 199 215
rect 351 47 381 215
rect 437 47 467 215
rect 543 47 573 215
<< scpmoshvt >>
rect 83 367 113 619
rect 161 367 191 619
rect 351 367 381 619
rect 438 367 468 619
rect 548 367 578 619
<< ndiff >>
rect 30 192 83 215
rect 30 158 38 192
rect 72 158 83 192
rect 30 93 83 158
rect 30 59 38 93
rect 72 59 83 93
rect 30 47 83 59
rect 113 187 169 215
rect 113 153 124 187
rect 158 153 169 187
rect 113 101 169 153
rect 113 67 124 101
rect 158 67 169 101
rect 113 47 169 67
rect 199 127 351 215
rect 199 93 210 127
rect 244 93 306 127
rect 340 93 351 127
rect 199 47 351 93
rect 381 190 437 215
rect 381 156 392 190
rect 426 156 437 190
rect 381 101 437 156
rect 381 67 392 101
rect 426 67 437 101
rect 381 47 437 67
rect 467 47 543 215
rect 573 192 631 215
rect 573 158 589 192
rect 623 158 631 192
rect 573 93 631 158
rect 573 59 589 93
rect 623 59 631 93
rect 573 47 631 59
<< pdiff >>
rect 30 607 83 619
rect 30 573 38 607
rect 72 573 83 607
rect 30 510 83 573
rect 30 476 38 510
rect 72 476 83 510
rect 30 418 83 476
rect 30 384 38 418
rect 72 384 83 418
rect 30 367 83 384
rect 113 367 161 619
rect 191 607 244 619
rect 191 573 202 607
rect 236 573 244 607
rect 191 510 244 573
rect 191 476 202 510
rect 236 476 244 510
rect 191 413 244 476
rect 191 379 202 413
rect 236 379 244 413
rect 191 367 244 379
rect 298 599 351 619
rect 298 565 306 599
rect 340 565 351 599
rect 298 522 351 565
rect 298 488 306 522
rect 340 488 351 522
rect 298 441 351 488
rect 298 407 306 441
rect 340 407 351 441
rect 298 367 351 407
rect 381 599 438 619
rect 381 565 393 599
rect 427 565 438 599
rect 381 527 438 565
rect 381 493 393 527
rect 427 493 438 527
rect 381 367 438 493
rect 468 583 548 619
rect 468 549 492 583
rect 526 549 548 583
rect 468 367 548 549
rect 578 599 631 619
rect 578 565 589 599
rect 623 565 631 599
rect 578 517 631 565
rect 578 483 589 517
rect 623 483 631 517
rect 578 436 631 483
rect 578 402 589 436
rect 623 402 631 436
rect 578 367 631 402
<< ndiffc >>
rect 38 158 72 192
rect 38 59 72 93
rect 124 153 158 187
rect 124 67 158 101
rect 210 93 244 127
rect 306 93 340 127
rect 392 156 426 190
rect 392 67 426 101
rect 589 158 623 192
rect 589 59 623 93
<< pdiffc >>
rect 38 573 72 607
rect 38 476 72 510
rect 38 384 72 418
rect 202 573 236 607
rect 202 476 236 510
rect 202 379 236 413
rect 306 565 340 599
rect 306 488 340 522
rect 306 407 340 441
rect 393 565 427 599
rect 393 493 427 527
rect 492 549 526 583
rect 589 565 623 599
rect 589 483 623 517
rect 589 402 623 436
<< poly >>
rect 83 619 113 645
rect 161 619 191 645
rect 351 619 381 645
rect 438 619 468 645
rect 548 619 578 645
rect 83 308 113 367
rect 47 292 113 308
rect 47 258 63 292
rect 97 258 113 292
rect 47 237 113 258
rect 161 345 191 367
rect 161 303 229 345
rect 351 303 381 367
rect 438 308 468 367
rect 548 308 578 367
rect 161 287 265 303
rect 161 253 215 287
rect 249 253 265 287
rect 161 237 265 253
rect 313 287 381 303
rect 313 253 329 287
rect 363 253 381 287
rect 313 237 381 253
rect 429 292 495 308
rect 429 258 445 292
rect 479 258 495 292
rect 429 242 495 258
rect 543 292 635 308
rect 543 258 585 292
rect 619 258 635 292
rect 543 242 635 258
rect 83 215 113 237
rect 169 215 199 237
rect 351 215 381 237
rect 437 215 467 242
rect 543 215 573 242
rect 83 21 113 47
rect 169 21 199 47
rect 351 21 381 47
rect 437 21 467 47
rect 543 21 573 47
<< polycont >>
rect 63 258 97 292
rect 215 253 249 287
rect 329 253 363 287
rect 445 258 479 292
rect 585 258 619 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 22 607 88 649
rect 22 573 38 607
rect 72 573 88 607
rect 22 510 88 573
rect 22 476 38 510
rect 72 476 88 510
rect 22 418 88 476
rect 22 384 38 418
rect 72 384 88 418
rect 186 607 252 615
rect 186 573 202 607
rect 236 573 252 607
rect 186 510 252 573
rect 186 476 202 510
rect 236 476 252 510
rect 186 413 252 476
rect 186 384 202 413
rect 195 379 202 384
rect 236 379 252 413
rect 290 599 355 615
rect 290 565 306 599
rect 340 565 355 599
rect 290 522 355 565
rect 290 488 306 522
rect 340 488 355 522
rect 290 441 355 488
rect 389 599 442 615
rect 389 565 393 599
rect 427 565 442 599
rect 389 527 442 565
rect 476 583 542 649
rect 476 549 492 583
rect 526 549 542 583
rect 476 543 542 549
rect 576 599 639 615
rect 576 565 589 599
rect 623 565 639 599
rect 389 493 393 527
rect 427 509 442 527
rect 576 517 639 565
rect 576 509 589 517
rect 427 493 589 509
rect 389 483 589 493
rect 623 483 639 517
rect 389 475 639 483
rect 290 407 306 441
rect 340 407 549 441
rect 195 373 252 379
rect 17 292 161 350
rect 195 339 347 373
rect 311 303 347 339
rect 17 258 63 292
rect 97 258 161 292
rect 17 242 161 258
rect 195 287 277 303
rect 195 253 215 287
rect 249 253 277 287
rect 195 237 277 253
rect 311 287 379 303
rect 311 253 329 287
rect 363 253 379 287
rect 311 240 379 253
rect 413 292 481 350
rect 413 258 445 292
rect 479 258 481 292
rect 413 240 481 258
rect 22 192 88 208
rect 311 203 347 240
rect 515 206 549 407
rect 583 436 639 475
rect 583 402 589 436
rect 623 402 639 436
rect 583 386 639 402
rect 583 292 655 352
rect 583 258 585 292
rect 619 258 655 292
rect 583 242 655 258
rect 22 158 38 192
rect 72 158 88 192
rect 22 93 88 158
rect 22 59 38 93
rect 72 59 88 93
rect 22 17 88 59
rect 122 187 347 203
rect 122 153 124 187
rect 158 169 347 187
rect 390 190 549 206
rect 158 153 160 169
rect 122 101 160 153
rect 390 156 392 190
rect 426 172 549 190
rect 585 192 639 208
rect 426 156 430 172
rect 122 67 124 101
rect 158 67 160 101
rect 122 51 160 67
rect 194 127 356 135
rect 194 93 210 127
rect 244 93 306 127
rect 340 93 356 127
rect 194 17 356 93
rect 390 101 430 156
rect 390 67 392 101
rect 426 67 430 101
rect 390 51 430 67
rect 585 158 589 192
rect 623 158 639 192
rect 585 93 639 158
rect 585 59 589 93
rect 623 59 639 93
rect 585 17 639 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2bb2oi_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2_N
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3054260
string GDS_START 3047152
<< end >>
