magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 6 49 830 241
rect 0 0 864 49
<< scnmos >>
rect 85 47 115 215
rect 171 47 201 215
rect 325 47 355 215
rect 432 47 462 215
rect 541 47 571 215
rect 649 47 679 215
rect 721 47 751 215
<< scpmoshvt >>
rect 92 367 122 619
rect 178 367 208 619
rect 325 367 355 619
rect 397 367 427 619
rect 505 367 535 619
rect 636 367 666 619
rect 722 367 752 619
<< ndiff >>
rect 32 203 85 215
rect 32 169 40 203
rect 74 169 85 203
rect 32 93 85 169
rect 32 59 40 93
rect 74 59 85 93
rect 32 47 85 59
rect 115 207 171 215
rect 115 173 126 207
rect 160 173 171 207
rect 115 101 171 173
rect 115 67 126 101
rect 160 67 171 101
rect 115 47 171 67
rect 201 167 325 215
rect 201 133 212 167
rect 246 133 280 167
rect 314 133 325 167
rect 201 89 325 133
rect 201 55 212 89
rect 246 55 280 89
rect 314 55 325 89
rect 201 47 325 55
rect 355 167 432 215
rect 355 133 380 167
rect 414 133 432 167
rect 355 91 432 133
rect 355 57 380 91
rect 414 57 432 91
rect 355 47 432 57
rect 462 91 541 215
rect 462 57 485 91
rect 519 57 541 91
rect 462 47 541 57
rect 571 167 649 215
rect 571 133 593 167
rect 627 133 649 167
rect 571 91 649 133
rect 571 57 593 91
rect 627 57 649 91
rect 571 47 649 57
rect 679 47 721 215
rect 751 203 804 215
rect 751 169 762 203
rect 796 169 804 203
rect 751 101 804 169
rect 751 67 762 101
rect 796 67 804 101
rect 751 47 804 67
<< pdiff >>
rect 39 607 92 619
rect 39 573 47 607
rect 81 573 92 607
rect 39 512 92 573
rect 39 478 47 512
rect 81 478 92 512
rect 39 413 92 478
rect 39 379 47 413
rect 81 379 92 413
rect 39 367 92 379
rect 122 599 178 619
rect 122 565 133 599
rect 167 565 178 599
rect 122 504 178 565
rect 122 470 133 504
rect 167 470 178 504
rect 122 413 178 470
rect 122 379 133 413
rect 167 379 178 413
rect 122 367 178 379
rect 208 607 325 619
rect 208 573 247 607
rect 281 573 325 607
rect 208 512 325 573
rect 208 478 247 512
rect 281 478 325 512
rect 208 421 325 478
rect 208 387 247 421
rect 281 387 325 421
rect 208 367 325 387
rect 355 367 397 619
rect 427 367 505 619
rect 535 599 636 619
rect 535 565 583 599
rect 617 565 636 599
rect 535 514 636 565
rect 535 480 583 514
rect 617 480 636 514
rect 535 434 636 480
rect 535 400 583 434
rect 617 400 636 434
rect 535 367 636 400
rect 666 607 722 619
rect 666 573 677 607
rect 711 573 722 607
rect 666 492 722 573
rect 666 458 677 492
rect 711 458 722 492
rect 666 367 722 458
rect 752 599 805 619
rect 752 565 763 599
rect 797 565 805 599
rect 752 514 805 565
rect 752 480 763 514
rect 797 480 805 514
rect 752 436 805 480
rect 752 402 763 436
rect 797 402 805 436
rect 752 367 805 402
<< ndiffc >>
rect 40 169 74 203
rect 40 59 74 93
rect 126 173 160 207
rect 126 67 160 101
rect 212 133 246 167
rect 280 133 314 167
rect 212 55 246 89
rect 280 55 314 89
rect 380 133 414 167
rect 380 57 414 91
rect 485 57 519 91
rect 593 133 627 167
rect 593 57 627 91
rect 762 169 796 203
rect 762 67 796 101
<< pdiffc >>
rect 47 573 81 607
rect 47 478 81 512
rect 47 379 81 413
rect 133 565 167 599
rect 133 470 167 504
rect 133 379 167 413
rect 247 573 281 607
rect 247 478 281 512
rect 247 387 281 421
rect 583 565 617 599
rect 583 480 617 514
rect 583 400 617 434
rect 677 573 711 607
rect 677 458 711 492
rect 763 565 797 599
rect 763 480 797 514
rect 763 402 797 436
<< poly >>
rect 92 619 122 645
rect 178 619 208 645
rect 325 619 355 645
rect 397 619 427 645
rect 505 619 535 645
rect 636 619 666 645
rect 722 619 752 645
rect 92 303 122 367
rect 178 303 208 367
rect 325 335 355 367
rect 289 319 355 335
rect 85 287 247 303
rect 85 253 197 287
rect 231 253 247 287
rect 289 285 305 319
rect 339 285 355 319
rect 289 269 355 285
rect 85 237 247 253
rect 85 215 115 237
rect 171 215 201 237
rect 325 215 355 269
rect 397 335 427 367
rect 505 335 535 367
rect 636 335 666 367
rect 397 319 463 335
rect 397 285 413 319
rect 447 285 463 319
rect 397 269 463 285
rect 505 319 571 335
rect 505 285 521 319
rect 555 285 571 319
rect 505 269 571 285
rect 613 319 679 335
rect 613 285 629 319
rect 663 285 679 319
rect 722 325 752 367
rect 722 309 835 325
rect 722 289 785 309
rect 613 269 679 285
rect 397 264 462 269
rect 432 215 462 264
rect 541 215 571 269
rect 649 215 679 269
rect 721 275 785 289
rect 819 275 835 309
rect 721 259 835 275
rect 721 215 751 259
rect 85 21 115 47
rect 171 21 201 47
rect 325 21 355 47
rect 432 21 462 47
rect 541 21 571 47
rect 649 21 679 47
rect 721 21 751 47
<< polycont >>
rect 197 253 231 287
rect 305 285 339 319
rect 413 285 447 319
rect 521 285 555 319
rect 629 285 663 319
rect 785 275 819 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 31 607 85 649
rect 31 573 47 607
rect 81 573 85 607
rect 31 512 85 573
rect 31 478 47 512
rect 81 478 85 512
rect 31 413 85 478
rect 31 379 47 413
rect 81 379 85 413
rect 31 363 85 379
rect 119 599 183 615
rect 119 565 133 599
rect 167 565 183 599
rect 119 504 183 565
rect 119 470 133 504
rect 167 470 183 504
rect 119 413 183 470
rect 119 379 133 413
rect 167 379 183 413
rect 119 339 183 379
rect 231 607 285 649
rect 231 573 247 607
rect 281 573 285 607
rect 579 599 627 615
rect 231 512 285 573
rect 231 478 247 512
rect 281 478 285 512
rect 231 421 285 478
rect 231 387 247 421
rect 281 387 285 421
rect 231 371 285 387
rect 24 203 85 219
rect 24 169 40 203
rect 74 169 85 203
rect 24 93 85 169
rect 24 59 40 93
rect 74 59 85 93
rect 24 17 85 59
rect 119 207 162 339
rect 319 337 366 592
rect 289 319 366 337
rect 119 173 126 207
rect 160 173 162 207
rect 196 287 247 303
rect 196 253 197 287
rect 231 253 247 287
rect 289 285 305 319
rect 339 285 366 319
rect 289 269 366 285
rect 400 319 461 592
rect 400 285 413 319
rect 447 285 461 319
rect 400 269 461 285
rect 495 347 545 592
rect 579 565 583 599
rect 617 565 627 599
rect 579 514 627 565
rect 579 480 583 514
rect 617 480 627 514
rect 579 434 627 480
rect 661 607 727 649
rect 661 573 677 607
rect 711 573 727 607
rect 661 492 727 573
rect 661 458 677 492
rect 711 458 727 492
rect 661 454 727 458
rect 761 599 813 615
rect 761 565 763 599
rect 797 565 813 599
rect 761 514 813 565
rect 761 480 763 514
rect 797 480 813 514
rect 579 400 583 434
rect 617 420 627 434
rect 761 436 813 480
rect 761 420 763 436
rect 617 402 763 420
rect 797 402 813 436
rect 617 400 813 402
rect 579 386 813 400
rect 579 384 735 386
rect 495 319 562 347
rect 495 285 521 319
rect 555 285 562 319
rect 495 269 562 285
rect 596 319 663 350
rect 596 285 629 319
rect 596 269 663 285
rect 196 235 247 253
rect 697 235 735 384
rect 769 309 847 352
rect 769 275 785 309
rect 819 275 847 309
rect 769 267 847 275
rect 196 233 735 235
rect 196 203 812 233
rect 196 201 762 203
rect 119 101 162 173
rect 704 169 762 201
rect 796 169 812 203
rect 119 67 126 101
rect 160 67 162 101
rect 119 51 162 67
rect 196 133 212 167
rect 246 133 280 167
rect 314 133 330 167
rect 196 89 330 133
rect 196 55 212 89
rect 246 55 280 89
rect 314 55 330 89
rect 196 17 330 55
rect 364 133 380 167
rect 414 133 593 167
rect 627 133 643 167
rect 364 91 430 133
rect 364 57 380 91
rect 414 57 430 91
rect 364 51 430 57
rect 469 91 535 99
rect 469 57 485 91
rect 519 57 535 91
rect 469 17 535 57
rect 577 91 643 133
rect 577 57 593 91
rect 627 57 643 91
rect 577 51 643 57
rect 704 101 812 169
rect 704 67 762 101
rect 796 67 812 101
rect 704 51 812 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o311a_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4416076
string GDS_START 4406744
<< end >>
