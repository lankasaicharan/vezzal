magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 332 1094 704
<< pwell >>
rect 238 236 506 256
rect 1 228 506 236
rect 1 49 1050 228
rect 0 0 1056 49
<< scpmos >>
rect 83 392 119 592
rect 173 392 209 592
rect 392 368 428 592
rect 482 368 518 592
rect 606 368 642 568
rect 737 368 773 568
rect 827 368 863 568
rect 937 368 973 568
<< nmoslvt >>
rect 84 82 114 210
rect 162 82 192 210
rect 314 82 344 230
rect 400 82 430 230
rect 621 74 651 202
rect 745 74 775 202
rect 823 74 853 202
rect 937 74 967 202
<< ndiff >>
rect 264 210 314 230
rect 27 198 84 210
rect 27 164 39 198
rect 73 164 84 198
rect 27 128 84 164
rect 27 94 39 128
rect 73 94 84 128
rect 27 82 84 94
rect 114 82 162 210
rect 192 131 314 210
rect 192 97 203 131
rect 237 97 314 131
rect 192 82 314 97
rect 344 218 400 230
rect 344 184 355 218
rect 389 184 400 218
rect 344 82 400 184
rect 430 94 480 230
rect 571 180 621 202
rect 557 144 621 180
rect 557 110 569 144
rect 603 110 621 144
rect 430 82 503 94
rect 445 48 457 82
rect 491 48 503 82
rect 557 74 621 110
rect 651 190 745 202
rect 651 156 684 190
rect 718 156 745 190
rect 651 74 745 156
rect 775 74 823 202
rect 853 144 937 202
rect 853 110 868 144
rect 902 110 937 144
rect 853 74 937 110
rect 967 190 1024 202
rect 967 156 978 190
rect 1012 156 1024 190
rect 967 120 1024 156
rect 967 86 978 120
rect 1012 86 1024 120
rect 967 74 1024 86
rect 445 36 503 48
<< pdiff >>
rect 319 592 377 604
rect 533 592 591 604
rect 27 580 83 592
rect 27 546 39 580
rect 73 546 83 580
rect 27 510 83 546
rect 27 476 39 510
rect 73 476 83 510
rect 27 440 83 476
rect 27 406 39 440
rect 73 406 83 440
rect 27 392 83 406
rect 119 580 173 592
rect 119 546 129 580
rect 163 546 173 580
rect 119 508 173 546
rect 119 474 129 508
rect 163 474 173 508
rect 119 392 173 474
rect 209 440 265 592
rect 319 558 331 592
rect 365 558 392 592
rect 319 546 392 558
rect 209 406 219 440
rect 253 406 265 440
rect 209 392 265 406
rect 342 368 392 546
rect 428 419 482 592
rect 428 385 438 419
rect 472 385 482 419
rect 428 368 482 385
rect 518 558 545 592
rect 579 568 591 592
rect 657 592 722 604
rect 657 568 672 592
rect 579 558 606 568
rect 518 368 606 558
rect 642 558 672 568
rect 706 568 722 592
rect 706 558 737 568
rect 642 368 737 558
rect 773 531 827 568
rect 773 497 783 531
rect 817 497 827 531
rect 773 440 827 497
rect 773 406 783 440
rect 817 406 827 440
rect 773 368 827 406
rect 863 560 937 568
rect 863 526 883 560
rect 917 526 937 560
rect 863 492 937 526
rect 863 458 883 492
rect 917 458 937 492
rect 863 424 937 458
rect 863 390 883 424
rect 917 390 937 424
rect 863 368 937 390
rect 973 556 1029 568
rect 973 522 983 556
rect 1017 522 1029 556
rect 973 440 1029 522
rect 973 406 983 440
rect 1017 406 1029 440
rect 973 368 1029 406
<< ndiffc >>
rect 39 164 73 198
rect 39 94 73 128
rect 203 97 237 131
rect 355 184 389 218
rect 569 110 603 144
rect 457 48 491 82
rect 684 156 718 190
rect 868 110 902 144
rect 978 156 1012 190
rect 978 86 1012 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 129 546 163 580
rect 129 474 163 508
rect 331 558 365 592
rect 219 406 253 440
rect 438 385 472 419
rect 545 558 579 592
rect 672 558 706 592
rect 783 497 817 531
rect 783 406 817 440
rect 883 526 917 560
rect 883 458 917 492
rect 883 390 917 424
rect 983 522 1017 556
rect 983 406 1017 440
<< poly >>
rect 83 592 119 618
rect 173 592 209 618
rect 392 592 428 618
rect 482 592 518 618
rect 83 366 119 392
rect 83 326 114 366
rect 21 310 114 326
rect 173 318 209 392
rect 606 568 642 594
rect 737 568 773 594
rect 827 568 863 594
rect 937 568 973 594
rect 392 318 428 368
rect 482 318 518 368
rect 606 336 642 368
rect 737 336 773 368
rect 827 336 863 368
rect 937 336 973 368
rect 585 320 651 336
rect 21 276 37 310
rect 71 276 114 310
rect 21 260 114 276
rect 84 210 114 260
rect 162 302 228 318
rect 162 268 178 302
rect 212 268 228 302
rect 392 302 512 318
rect 392 282 462 302
rect 162 252 228 268
rect 314 268 462 282
rect 496 268 512 302
rect 585 286 601 320
rect 635 286 651 320
rect 585 270 651 286
rect 693 320 775 336
rect 693 286 709 320
rect 743 286 775 320
rect 693 270 775 286
rect 314 252 512 268
rect 162 210 192 252
rect 314 230 344 252
rect 400 230 430 252
rect 621 202 651 270
rect 745 202 775 270
rect 823 320 889 336
rect 823 286 839 320
rect 873 286 889 320
rect 823 270 889 286
rect 937 320 1003 336
rect 937 286 953 320
rect 987 286 1003 320
rect 937 270 1003 286
rect 823 202 853 270
rect 937 202 967 270
rect 84 56 114 82
rect 162 56 192 82
rect 314 56 344 82
rect 400 56 430 82
rect 621 48 651 74
rect 745 48 775 74
rect 823 48 853 74
rect 937 48 967 74
<< polycont >>
rect 37 276 71 310
rect 178 268 212 302
rect 462 268 496 302
rect 601 286 635 320
rect 709 286 743 320
rect 839 286 873 320
rect 953 286 987 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 580 73 596
rect 23 546 39 580
rect 23 510 73 546
rect 23 476 39 510
rect 23 440 73 476
rect 113 580 179 596
rect 113 546 129 580
rect 163 546 179 580
rect 113 508 179 546
rect 315 592 381 649
rect 315 558 331 592
rect 365 558 381 592
rect 315 542 381 558
rect 529 592 595 649
rect 529 558 545 592
rect 579 558 595 592
rect 529 542 595 558
rect 653 592 933 615
rect 653 558 672 592
rect 706 581 933 592
rect 706 558 726 581
rect 653 542 726 558
rect 867 560 933 581
rect 767 531 833 547
rect 767 508 783 531
rect 113 474 129 508
rect 163 497 783 508
rect 817 497 833 531
rect 163 474 833 497
rect 767 440 833 474
rect 23 406 39 440
rect 73 406 219 440
rect 253 406 305 440
rect 23 390 305 406
rect 21 310 87 356
rect 21 276 37 310
rect 71 276 87 310
rect 21 260 87 276
rect 121 302 228 356
rect 121 268 178 302
rect 212 268 228 302
rect 121 252 228 268
rect 271 218 305 390
rect 23 198 305 218
rect 23 164 39 198
rect 73 184 305 198
rect 339 419 488 440
rect 339 385 438 419
rect 472 385 488 419
rect 339 364 488 385
rect 339 218 405 364
rect 585 320 651 430
rect 767 406 783 440
rect 817 406 833 440
rect 767 390 833 406
rect 867 526 883 560
rect 917 526 933 560
rect 867 492 933 526
rect 867 458 883 492
rect 917 458 933 492
rect 867 424 933 458
rect 867 390 883 424
rect 917 390 933 424
rect 967 556 1033 649
rect 967 522 983 556
rect 1017 522 1033 556
rect 967 440 1033 522
rect 967 406 983 440
rect 1017 406 1033 440
rect 967 390 1033 406
rect 339 184 355 218
rect 389 184 405 218
rect 446 302 512 318
rect 446 268 462 302
rect 496 268 512 302
rect 585 286 601 320
rect 635 286 651 320
rect 585 270 651 286
rect 693 320 759 356
rect 693 286 709 320
rect 743 286 759 320
rect 693 270 759 286
rect 793 320 889 356
rect 793 286 839 320
rect 873 286 889 320
rect 793 270 889 286
rect 937 320 1031 356
rect 937 286 953 320
rect 987 286 1031 320
rect 937 270 1031 286
rect 446 236 512 268
rect 446 202 750 236
rect 23 128 73 164
rect 271 150 305 184
rect 446 150 480 202
rect 653 190 750 202
rect 23 94 39 128
rect 23 78 73 94
rect 187 131 237 150
rect 187 97 203 131
rect 271 116 480 150
rect 553 144 619 168
rect 187 17 237 97
rect 553 110 569 144
rect 603 110 619 144
rect 653 156 684 190
rect 718 156 750 190
rect 653 140 750 156
rect 784 202 1028 236
rect 553 104 619 110
rect 784 104 818 202
rect 962 190 1028 202
rect 441 48 457 82
rect 491 48 507 82
rect 553 70 818 104
rect 852 144 918 168
rect 852 110 868 144
rect 902 110 918 144
rect 441 17 507 48
rect 852 17 918 110
rect 962 156 978 190
rect 1012 156 1028 190
rect 962 120 1028 156
rect 962 86 978 120
rect 1012 86 1028 120
rect 962 70 1028 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a222o_2
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 C2
port 6 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 8576
string GDS_START 130
<< end >>
