magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 41 49 1055 241
rect 0 0 1056 49
<< scnmos >>
rect 124 47 154 215
rect 202 47 232 215
rect 288 47 318 215
rect 366 47 396 215
rect 452 47 482 215
rect 530 47 560 215
rect 661 47 691 215
rect 747 47 777 215
rect 840 47 870 215
rect 934 47 964 215
<< scpmoshvt >>
rect 124 367 154 619
rect 202 367 232 619
rect 288 367 318 619
rect 366 367 396 619
rect 452 367 482 619
rect 530 367 560 619
rect 644 367 674 619
rect 730 367 760 619
rect 848 367 878 619
rect 934 367 964 619
<< ndiff >>
rect 67 184 124 215
rect 67 150 79 184
rect 113 150 124 184
rect 67 103 124 150
rect 67 69 79 103
rect 113 69 124 103
rect 67 47 124 69
rect 154 47 202 215
rect 232 103 288 215
rect 232 69 243 103
rect 277 69 288 103
rect 232 47 288 69
rect 318 47 366 215
rect 396 184 452 215
rect 396 150 407 184
rect 441 150 452 184
rect 396 93 452 150
rect 396 59 407 93
rect 441 59 452 93
rect 396 47 452 59
rect 482 47 530 215
rect 560 103 661 215
rect 560 69 571 103
rect 605 69 661 103
rect 560 47 661 69
rect 691 203 747 215
rect 691 169 702 203
rect 736 169 747 203
rect 691 103 747 169
rect 691 69 702 103
rect 736 69 747 103
rect 691 47 747 69
rect 777 113 840 215
rect 777 79 788 113
rect 822 79 840 113
rect 777 47 840 79
rect 870 203 934 215
rect 870 169 881 203
rect 915 169 934 203
rect 870 103 934 169
rect 870 69 881 103
rect 915 69 934 103
rect 870 47 934 69
rect 964 113 1029 215
rect 964 79 983 113
rect 1017 79 1029 113
rect 964 47 1029 79
<< pdiff >>
rect 65 597 124 619
rect 65 563 77 597
rect 111 563 124 597
rect 65 503 124 563
rect 65 469 77 503
rect 111 469 124 503
rect 65 409 124 469
rect 65 375 77 409
rect 111 375 124 409
rect 65 367 124 375
rect 154 367 202 619
rect 232 584 288 619
rect 232 550 243 584
rect 277 550 288 584
rect 232 367 288 550
rect 318 367 366 619
rect 396 409 452 619
rect 396 375 407 409
rect 441 375 452 409
rect 396 367 452 375
rect 482 367 530 619
rect 560 603 644 619
rect 560 569 583 603
rect 617 569 644 603
rect 560 506 644 569
rect 560 472 583 506
rect 617 472 644 506
rect 560 409 644 472
rect 560 375 583 409
rect 617 375 644 409
rect 560 367 644 375
rect 674 597 730 619
rect 674 563 685 597
rect 719 563 730 597
rect 674 503 730 563
rect 674 469 685 503
rect 719 469 730 503
rect 674 409 730 469
rect 674 375 685 409
rect 719 375 730 409
rect 674 367 730 375
rect 760 603 848 619
rect 760 569 787 603
rect 821 569 848 603
rect 760 477 848 569
rect 760 443 787 477
rect 821 443 848 477
rect 760 367 848 443
rect 878 597 934 619
rect 878 563 889 597
rect 923 563 934 597
rect 878 503 934 563
rect 878 469 889 503
rect 923 469 934 503
rect 878 409 934 469
rect 878 375 889 409
rect 923 375 934 409
rect 878 367 934 375
rect 964 603 1021 619
rect 964 569 975 603
rect 1009 569 1021 603
rect 964 477 1021 569
rect 964 443 975 477
rect 1009 443 1021 477
rect 964 367 1021 443
<< ndiffc >>
rect 79 150 113 184
rect 79 69 113 103
rect 243 69 277 103
rect 407 150 441 184
rect 407 59 441 93
rect 571 69 605 103
rect 702 169 736 203
rect 702 69 736 103
rect 788 79 822 113
rect 881 169 915 203
rect 881 69 915 103
rect 983 79 1017 113
<< pdiffc >>
rect 77 563 111 597
rect 77 469 111 503
rect 77 375 111 409
rect 243 550 277 584
rect 407 375 441 409
rect 583 569 617 603
rect 583 472 617 506
rect 583 375 617 409
rect 685 563 719 597
rect 685 469 719 503
rect 685 375 719 409
rect 787 569 821 603
rect 787 443 821 477
rect 889 563 923 597
rect 889 469 923 503
rect 889 375 923 409
rect 975 569 1009 603
rect 975 443 1009 477
<< poly >>
rect 124 619 154 645
rect 202 619 232 645
rect 288 619 318 645
rect 366 619 396 645
rect 452 619 482 645
rect 530 619 560 645
rect 644 619 674 645
rect 730 619 760 645
rect 848 619 878 645
rect 934 619 964 645
rect 124 303 154 367
rect 88 287 154 303
rect 88 253 104 287
rect 138 253 154 287
rect 88 237 154 253
rect 124 215 154 237
rect 202 303 232 367
rect 288 303 318 367
rect 202 287 318 303
rect 202 253 233 287
rect 267 253 318 287
rect 202 237 318 253
rect 202 215 232 237
rect 288 215 318 237
rect 366 303 396 367
rect 452 303 482 367
rect 366 287 482 303
rect 366 253 411 287
rect 445 253 482 287
rect 366 237 482 253
rect 366 215 396 237
rect 452 215 482 237
rect 530 321 560 367
rect 644 321 674 367
rect 730 321 760 367
rect 848 321 878 367
rect 934 321 964 367
rect 530 305 596 321
rect 530 271 546 305
rect 580 271 596 305
rect 530 255 596 271
rect 644 305 964 321
rect 644 271 680 305
rect 714 271 748 305
rect 782 271 816 305
rect 850 271 884 305
rect 918 271 964 305
rect 644 255 964 271
rect 530 215 560 255
rect 661 215 691 255
rect 747 215 777 255
rect 840 215 870 255
rect 934 215 964 255
rect 124 21 154 47
rect 202 21 232 47
rect 288 21 318 47
rect 366 21 396 47
rect 452 21 482 47
rect 530 21 560 47
rect 661 21 691 47
rect 747 21 777 47
rect 840 21 870 47
rect 934 21 964 47
<< polycont >>
rect 104 253 138 287
rect 233 253 267 287
rect 411 253 445 287
rect 546 271 580 305
rect 680 271 714 305
rect 748 271 782 305
rect 816 271 850 305
rect 884 271 918 305
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 18 597 111 613
rect 18 563 77 597
rect 18 503 111 563
rect 227 584 293 649
rect 227 550 243 584
rect 277 550 293 584
rect 227 515 293 550
rect 567 603 633 649
rect 567 569 583 603
rect 617 569 633 603
rect 18 469 77 503
rect 567 506 633 569
rect 18 409 111 469
rect 18 375 77 409
rect 18 359 111 375
rect 147 445 531 479
rect 18 200 52 359
rect 147 303 181 445
rect 325 375 407 409
rect 441 375 457 409
rect 325 359 457 375
rect 88 287 181 303
rect 88 253 104 287
rect 138 253 181 287
rect 88 236 181 253
rect 217 287 283 356
rect 217 253 233 287
rect 267 253 283 287
rect 217 236 283 253
rect 325 200 359 359
rect 497 321 531 445
rect 567 472 583 506
rect 617 472 633 506
rect 567 409 633 472
rect 567 375 583 409
rect 617 375 633 409
rect 567 359 633 375
rect 669 597 735 613
rect 669 563 685 597
rect 719 563 735 597
rect 669 503 735 563
rect 669 469 685 503
rect 719 469 735 503
rect 669 409 735 469
rect 771 603 837 649
rect 771 569 787 603
rect 821 569 837 603
rect 771 477 837 569
rect 771 443 787 477
rect 821 443 837 477
rect 771 427 837 443
rect 873 597 939 613
rect 873 563 889 597
rect 923 563 939 597
rect 873 503 939 563
rect 873 469 889 503
rect 923 469 939 503
rect 669 375 685 409
rect 719 391 735 409
rect 873 409 939 469
rect 975 603 1025 649
rect 1009 569 1025 603
rect 975 477 1025 569
rect 1009 443 1025 477
rect 975 427 1025 443
rect 873 391 889 409
rect 719 375 889 391
rect 923 391 939 409
rect 923 375 1031 391
rect 669 357 1031 375
rect 497 305 596 321
rect 395 287 461 303
rect 395 253 411 287
rect 445 253 461 287
rect 497 271 546 305
rect 580 271 596 305
rect 497 255 596 271
rect 632 305 934 321
rect 632 271 680 305
rect 714 271 748 305
rect 782 271 816 305
rect 850 271 884 305
rect 918 271 934 305
rect 632 255 934 271
rect 395 236 461 253
rect 632 200 666 255
rect 985 219 1031 357
rect 18 184 666 200
rect 18 166 79 184
rect 63 150 79 166
rect 113 166 407 184
rect 113 150 129 166
rect 63 103 129 150
rect 391 150 407 166
rect 441 166 666 184
rect 702 203 1031 219
rect 736 185 881 203
rect 441 150 457 166
rect 63 69 79 103
rect 113 69 129 103
rect 63 53 129 69
rect 227 103 293 130
rect 227 69 243 103
rect 277 69 293 103
rect 227 17 293 69
rect 391 93 457 150
rect 391 59 407 93
rect 441 59 457 93
rect 555 103 621 130
rect 555 69 571 103
rect 605 69 621 103
rect 555 17 621 69
rect 702 103 736 169
rect 865 169 881 185
rect 915 185 1031 203
rect 915 169 931 185
rect 702 53 736 69
rect 772 113 822 149
rect 772 79 788 113
rect 772 17 822 79
rect 865 103 931 169
rect 865 69 881 103
rect 915 69 931 103
rect 865 53 931 69
rect 967 113 1033 149
rect 967 79 983 113
rect 1017 79 1033 113
rect 967 17 1033 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 maj3_4
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6759390
string GDS_START 6751678
<< end >>
