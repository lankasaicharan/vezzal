magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 887 235 1341 241
rect 359 180 1341 235
rect 22 49 1341 180
rect 0 0 1344 49
<< scnmos >>
rect 105 70 135 154
rect 191 70 221 154
rect 438 125 468 209
rect 524 125 554 209
rect 596 125 626 209
rect 696 125 726 209
rect 776 125 806 209
rect 966 47 996 215
rect 1038 47 1068 215
rect 1146 47 1176 215
rect 1232 47 1262 215
<< scpmoshvt >>
rect 84 464 114 592
rect 221 464 251 592
rect 444 473 474 601
rect 552 473 582 601
rect 624 473 654 601
rect 733 473 763 557
rect 805 473 835 557
rect 966 367 996 619
rect 1052 367 1082 619
rect 1146 367 1176 619
rect 1232 367 1262 619
<< ndiff >>
rect 48 129 105 154
rect 48 95 56 129
rect 90 95 105 129
rect 48 70 105 95
rect 135 118 191 154
rect 135 84 146 118
rect 180 84 191 118
rect 135 70 191 84
rect 221 118 274 154
rect 221 84 232 118
rect 266 84 274 118
rect 221 70 274 84
rect 385 184 438 209
rect 385 150 393 184
rect 427 150 438 184
rect 385 125 438 150
rect 468 184 524 209
rect 468 150 479 184
rect 513 150 524 184
rect 468 125 524 150
rect 554 125 596 209
rect 626 184 696 209
rect 626 150 651 184
rect 685 150 696 184
rect 626 125 696 150
rect 726 125 776 209
rect 806 184 859 209
rect 806 150 817 184
rect 851 150 859 184
rect 806 125 859 150
rect 913 203 966 215
rect 913 169 921 203
rect 955 169 966 203
rect 913 101 966 169
rect 913 67 921 101
rect 955 67 966 101
rect 913 47 966 67
rect 996 47 1038 215
rect 1068 93 1146 215
rect 1068 59 1087 93
rect 1121 59 1146 93
rect 1068 47 1146 59
rect 1176 203 1232 215
rect 1176 169 1187 203
rect 1221 169 1232 203
rect 1176 101 1232 169
rect 1176 67 1187 101
rect 1221 67 1232 101
rect 1176 47 1232 67
rect 1262 203 1315 215
rect 1262 169 1273 203
rect 1307 169 1315 203
rect 1262 93 1315 169
rect 1262 59 1273 93
rect 1307 59 1315 93
rect 1262 47 1315 59
<< pdiff >>
rect 913 607 966 619
rect 31 578 84 592
rect 31 544 39 578
rect 73 544 84 578
rect 31 510 84 544
rect 31 476 39 510
rect 73 476 84 510
rect 31 464 84 476
rect 114 578 221 592
rect 114 544 125 578
rect 159 544 221 578
rect 114 510 221 544
rect 114 476 125 510
rect 159 476 221 510
rect 114 464 221 476
rect 251 510 307 592
rect 251 476 265 510
rect 299 476 307 510
rect 251 464 307 476
rect 372 473 444 601
rect 474 593 552 601
rect 474 559 496 593
rect 530 559 552 593
rect 474 473 552 559
rect 582 473 624 601
rect 654 587 711 601
rect 654 553 669 587
rect 703 557 711 587
rect 913 573 921 607
rect 955 573 966 607
rect 913 557 966 573
rect 703 553 733 557
rect 654 519 733 553
rect 654 485 669 519
rect 703 485 733 519
rect 654 473 733 485
rect 763 473 805 557
rect 835 532 966 557
rect 835 498 846 532
rect 880 531 966 532
rect 880 498 921 531
rect 835 497 921 498
rect 955 497 966 531
rect 835 473 966 497
rect 372 447 422 473
rect 372 413 380 447
rect 414 413 422 447
rect 372 397 422 413
rect 913 446 966 473
rect 913 412 921 446
rect 955 412 966 446
rect 913 367 966 412
rect 996 599 1052 619
rect 996 565 1007 599
rect 1041 565 1052 599
rect 996 507 1052 565
rect 996 473 1007 507
rect 1041 473 1052 507
rect 996 413 1052 473
rect 996 379 1007 413
rect 1041 379 1052 413
rect 996 367 1052 379
rect 1082 573 1146 619
rect 1082 539 1097 573
rect 1131 539 1146 573
rect 1082 367 1146 539
rect 1176 413 1232 619
rect 1176 379 1187 413
rect 1221 379 1232 413
rect 1176 367 1232 379
rect 1262 573 1315 619
rect 1262 539 1273 573
rect 1307 539 1315 573
rect 1262 367 1315 539
<< ndiffc >>
rect 56 95 90 129
rect 146 84 180 118
rect 232 84 266 118
rect 393 150 427 184
rect 479 150 513 184
rect 651 150 685 184
rect 817 150 851 184
rect 921 169 955 203
rect 921 67 955 101
rect 1087 59 1121 93
rect 1187 169 1221 203
rect 1187 67 1221 101
rect 1273 169 1307 203
rect 1273 59 1307 93
<< pdiffc >>
rect 39 544 73 578
rect 39 476 73 510
rect 125 544 159 578
rect 125 476 159 510
rect 265 476 299 510
rect 496 559 530 593
rect 669 553 703 587
rect 921 573 955 607
rect 669 485 703 519
rect 846 498 880 532
rect 921 497 955 531
rect 380 413 414 447
rect 921 412 955 446
rect 1007 565 1041 599
rect 1007 473 1041 507
rect 1007 379 1041 413
rect 1097 539 1131 573
rect 1187 379 1221 413
rect 1273 539 1307 573
<< poly >>
rect 84 592 114 618
rect 221 592 251 618
rect 444 601 474 627
rect 552 601 582 627
rect 624 601 654 627
rect 966 619 996 645
rect 1052 619 1082 645
rect 1146 619 1176 645
rect 1232 619 1262 645
rect 733 557 763 583
rect 805 557 835 583
rect 84 310 114 464
rect 221 310 251 464
rect 444 365 474 473
rect 552 437 582 473
rect 77 294 143 310
rect 77 260 93 294
rect 127 260 143 294
rect 77 226 143 260
rect 77 192 93 226
rect 127 192 143 226
rect 77 176 143 192
rect 185 294 251 310
rect 185 260 201 294
rect 235 260 251 294
rect 185 226 251 260
rect 299 349 474 365
rect 299 315 315 349
rect 349 335 474 349
rect 516 421 582 437
rect 516 387 532 421
rect 566 387 582 421
rect 516 353 582 387
rect 624 441 654 473
rect 624 425 690 441
rect 624 391 640 425
rect 674 391 690 425
rect 624 375 690 391
rect 349 315 365 335
rect 299 281 365 315
rect 516 319 532 353
rect 566 319 582 353
rect 733 333 763 473
rect 516 303 582 319
rect 630 313 763 333
rect 624 303 763 313
rect 805 438 835 473
rect 805 422 871 438
rect 805 388 821 422
rect 855 388 871 422
rect 805 372 871 388
rect 299 247 315 281
rect 349 261 365 281
rect 349 247 468 261
rect 299 231 468 247
rect 185 192 201 226
rect 235 192 251 226
rect 185 176 251 192
rect 105 154 135 176
rect 191 154 221 176
rect 105 44 135 70
rect 191 44 221 70
rect 335 51 365 231
rect 438 209 468 231
rect 524 209 554 303
rect 624 283 660 303
rect 624 261 654 283
rect 805 261 835 372
rect 966 324 996 367
rect 596 231 654 261
rect 596 209 626 231
rect 696 209 726 235
rect 776 231 835 261
rect 882 308 996 324
rect 882 274 898 308
rect 932 274 996 308
rect 1052 303 1082 367
rect 1146 325 1176 367
rect 1232 325 1262 367
rect 1146 309 1323 325
rect 882 258 996 274
rect 776 209 806 231
rect 966 215 996 258
rect 1038 287 1104 303
rect 1038 253 1054 287
rect 1088 253 1104 287
rect 1038 237 1104 253
rect 1146 275 1273 309
rect 1307 275 1323 309
rect 1146 259 1323 275
rect 1038 215 1068 237
rect 1146 215 1176 259
rect 1232 215 1262 259
rect 438 99 468 125
rect 524 99 554 125
rect 596 51 626 125
rect 696 103 726 125
rect 335 21 626 51
rect 668 87 734 103
rect 776 99 806 125
rect 668 53 684 87
rect 718 53 734 87
rect 668 37 734 53
rect 966 21 996 47
rect 1038 21 1068 47
rect 1146 21 1176 47
rect 1232 21 1262 47
<< polycont >>
rect 93 260 127 294
rect 93 192 127 226
rect 201 260 235 294
rect 315 315 349 349
rect 532 387 566 421
rect 640 391 674 425
rect 532 319 566 353
rect 821 388 855 422
rect 315 247 349 281
rect 201 192 235 226
rect 898 274 932 308
rect 1054 253 1088 287
rect 1273 275 1307 309
rect 684 53 718 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 23 578 82 594
rect 23 544 39 578
rect 73 544 82 578
rect 23 510 82 544
rect 23 476 39 510
rect 73 476 82 510
rect 23 426 82 476
rect 116 578 161 649
rect 116 544 125 578
rect 159 544 161 578
rect 116 510 161 544
rect 116 476 125 510
rect 159 476 161 510
rect 116 460 161 476
rect 195 562 397 596
rect 195 426 229 562
rect 265 510 327 526
rect 299 476 327 510
rect 363 519 397 562
rect 480 593 546 649
rect 830 607 971 649
rect 480 559 496 593
rect 530 559 546 593
rect 480 553 546 559
rect 653 587 744 603
rect 653 553 669 587
rect 703 553 744 587
rect 653 519 744 553
rect 363 485 582 519
rect 265 460 327 476
rect 23 392 229 426
rect 23 134 57 392
rect 293 365 327 460
rect 364 447 430 451
rect 364 413 380 447
rect 414 413 430 447
rect 364 399 430 413
rect 93 294 167 358
rect 127 260 167 294
rect 93 226 167 260
rect 127 192 167 226
rect 93 168 167 192
rect 201 294 259 358
rect 235 260 259 294
rect 201 226 259 260
rect 235 192 259 226
rect 201 168 259 192
rect 293 349 351 365
rect 293 315 315 349
rect 349 315 351 349
rect 293 281 351 315
rect 293 247 315 281
rect 349 247 351 281
rect 293 231 351 247
rect 385 259 430 399
rect 516 421 582 485
rect 653 485 669 519
rect 703 485 744 519
rect 653 475 744 485
rect 830 573 921 607
rect 955 573 971 607
rect 830 532 971 573
rect 830 498 846 532
rect 880 531 971 532
rect 880 498 921 531
rect 830 497 921 498
rect 955 497 971 531
rect 830 482 971 497
rect 516 387 532 421
rect 566 387 582 421
rect 516 353 582 387
rect 516 319 532 353
rect 566 319 582 353
rect 516 303 582 319
rect 624 425 676 441
rect 624 391 640 425
rect 674 391 676 425
rect 624 259 676 391
rect 293 134 327 231
rect 385 225 676 259
rect 710 310 744 475
rect 905 446 971 482
rect 805 422 871 438
rect 805 388 821 422
rect 855 388 871 422
rect 905 412 921 446
rect 955 412 971 446
rect 1005 599 1047 615
rect 1005 565 1007 599
rect 1041 565 1047 599
rect 1005 507 1047 565
rect 1081 573 1147 649
rect 1081 539 1097 573
rect 1131 539 1147 573
rect 1081 531 1147 539
rect 1257 573 1323 649
rect 1257 539 1273 573
rect 1307 539 1323 573
rect 1257 531 1323 539
rect 1005 473 1007 507
rect 1041 497 1047 507
rect 1041 473 1323 497
rect 1005 463 1323 473
rect 1005 413 1108 463
rect 805 378 871 388
rect 1005 379 1007 413
rect 1041 379 1108 413
rect 1005 378 1108 379
rect 805 344 1108 378
rect 1181 413 1223 429
rect 1181 379 1187 413
rect 1221 379 1223 413
rect 710 308 950 310
rect 710 274 898 308
rect 932 274 950 308
rect 710 273 950 274
rect 385 199 429 225
rect 377 184 429 199
rect 377 150 393 184
rect 427 150 429 184
rect 377 134 429 150
rect 463 184 529 191
rect 463 150 479 184
rect 513 150 529 184
rect 23 129 106 134
rect 23 95 56 129
rect 90 95 106 129
rect 23 79 106 95
rect 140 118 188 134
rect 140 84 146 118
rect 180 84 188 118
rect 140 17 188 84
rect 222 118 327 134
rect 222 84 232 118
rect 266 84 327 118
rect 222 68 327 84
rect 463 17 529 150
rect 563 100 597 225
rect 710 191 744 273
rect 984 239 1018 344
rect 905 205 1018 239
rect 1052 287 1104 303
rect 1052 253 1054 287
rect 1088 253 1104 287
rect 905 203 955 205
rect 635 184 744 191
rect 635 150 651 184
rect 685 150 744 184
rect 635 134 744 150
rect 801 184 867 200
rect 801 150 817 184
rect 851 150 867 184
rect 563 87 734 100
rect 563 53 684 87
rect 718 53 734 87
rect 563 51 734 53
rect 801 17 867 150
rect 905 169 921 203
rect 1052 171 1104 253
rect 905 101 955 169
rect 905 67 921 101
rect 989 137 1104 171
rect 1181 203 1223 379
rect 1269 309 1323 463
rect 1269 275 1273 309
rect 1307 275 1323 309
rect 1269 259 1323 275
rect 1181 169 1187 203
rect 1221 169 1223 203
rect 989 75 1037 137
rect 1071 93 1137 103
rect 905 51 955 67
rect 1071 59 1087 93
rect 1121 59 1137 93
rect 1071 17 1137 59
rect 1181 101 1223 169
rect 1181 67 1187 101
rect 1221 67 1223 101
rect 1181 51 1223 67
rect 1257 203 1323 219
rect 1257 169 1273 203
rect 1307 169 1323 203
rect 1257 93 1323 169
rect 1257 59 1273 93
rect 1307 59 1323 93
rect 1257 17 1323 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrtn_2
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 991 94 1025 128 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1183 94 1217 128 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1183 168 1217 202 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1183 390 1217 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2701304
string GDS_START 2690128
<< end >>
