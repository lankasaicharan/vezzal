magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 1 49 1949 241
rect 0 0 2016 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 252 47 282 215
rect 338 47 368 215
rect 424 47 454 215
rect 510 47 540 215
rect 596 47 626 215
rect 682 47 712 215
rect 872 47 902 215
rect 958 47 988 215
rect 1044 47 1074 215
rect 1130 47 1160 215
rect 1218 47 1248 215
rect 1304 47 1334 215
rect 1390 47 1420 215
rect 1496 47 1526 215
rect 1582 47 1612 215
rect 1668 47 1698 215
rect 1754 47 1784 215
rect 1840 47 1870 215
<< scpmoshvt >>
rect 94 367 124 619
rect 180 367 210 619
rect 266 367 296 619
rect 352 367 382 619
rect 438 367 468 619
rect 524 367 554 619
rect 610 367 640 619
rect 696 367 726 619
rect 804 367 834 619
rect 890 367 920 619
rect 976 367 1006 619
rect 1062 367 1092 619
rect 1252 367 1282 619
rect 1338 367 1368 619
rect 1424 367 1454 619
rect 1510 367 1540 619
rect 1596 367 1626 619
rect 1682 367 1712 619
rect 1768 367 1798 619
rect 1854 367 1884 619
<< ndiff >>
rect 27 192 80 215
rect 27 158 35 192
rect 69 158 80 192
rect 27 101 80 158
rect 27 67 35 101
rect 69 67 80 101
rect 27 47 80 67
rect 110 132 166 215
rect 110 98 121 132
rect 155 98 166 132
rect 110 47 166 98
rect 196 192 252 215
rect 196 158 207 192
rect 241 158 252 192
rect 196 101 252 158
rect 196 67 207 101
rect 241 67 252 101
rect 196 47 252 67
rect 282 132 338 215
rect 282 98 293 132
rect 327 98 338 132
rect 282 47 338 98
rect 368 192 424 215
rect 368 158 379 192
rect 413 158 424 192
rect 368 101 424 158
rect 368 67 379 101
rect 413 67 424 101
rect 368 47 424 67
rect 454 124 510 215
rect 454 90 465 124
rect 499 90 510 124
rect 454 47 510 90
rect 540 183 596 215
rect 540 149 551 183
rect 585 149 596 183
rect 540 47 596 149
rect 626 124 682 215
rect 626 90 637 124
rect 671 90 682 124
rect 626 47 682 90
rect 712 183 765 215
rect 712 149 723 183
rect 757 149 765 183
rect 712 47 765 149
rect 819 181 872 215
rect 819 147 827 181
rect 861 147 872 181
rect 819 47 872 147
rect 902 124 958 215
rect 902 90 913 124
rect 947 90 958 124
rect 902 47 958 90
rect 988 181 1044 215
rect 988 147 999 181
rect 1033 147 1044 181
rect 988 47 1044 147
rect 1074 124 1130 215
rect 1074 90 1085 124
rect 1119 90 1130 124
rect 1074 47 1130 90
rect 1160 192 1218 215
rect 1160 158 1171 192
rect 1205 158 1218 192
rect 1160 101 1218 158
rect 1160 67 1171 101
rect 1205 67 1218 101
rect 1160 47 1218 67
rect 1248 132 1304 215
rect 1248 98 1259 132
rect 1293 98 1304 132
rect 1248 47 1304 98
rect 1334 192 1390 215
rect 1334 158 1345 192
rect 1379 158 1390 192
rect 1334 101 1390 158
rect 1334 67 1345 101
rect 1379 67 1390 101
rect 1334 47 1390 67
rect 1420 132 1496 215
rect 1420 98 1440 132
rect 1474 98 1496 132
rect 1420 47 1496 98
rect 1526 192 1582 215
rect 1526 158 1537 192
rect 1571 158 1582 192
rect 1526 101 1582 158
rect 1526 67 1537 101
rect 1571 67 1582 101
rect 1526 47 1582 67
rect 1612 132 1668 215
rect 1612 98 1623 132
rect 1657 98 1668 132
rect 1612 47 1668 98
rect 1698 192 1754 215
rect 1698 158 1709 192
rect 1743 158 1754 192
rect 1698 101 1754 158
rect 1698 67 1709 101
rect 1743 67 1754 101
rect 1698 47 1754 67
rect 1784 132 1840 215
rect 1784 98 1795 132
rect 1829 98 1840 132
rect 1784 47 1840 98
rect 1870 192 1923 215
rect 1870 158 1881 192
rect 1915 158 1923 192
rect 1870 101 1923 158
rect 1870 67 1881 101
rect 1915 67 1923 101
rect 1870 47 1923 67
<< pdiff >>
rect 41 607 94 619
rect 41 573 49 607
rect 83 573 94 607
rect 41 510 94 573
rect 41 476 49 510
rect 83 476 94 510
rect 41 413 94 476
rect 41 379 49 413
rect 83 379 94 413
rect 41 367 94 379
rect 124 599 180 619
rect 124 565 135 599
rect 169 565 180 599
rect 124 508 180 565
rect 124 474 135 508
rect 169 474 180 508
rect 124 413 180 474
rect 124 379 135 413
rect 169 379 180 413
rect 124 367 180 379
rect 210 607 266 619
rect 210 573 221 607
rect 255 573 266 607
rect 210 515 266 573
rect 210 481 221 515
rect 255 481 266 515
rect 210 423 266 481
rect 210 389 221 423
rect 255 389 266 423
rect 210 367 266 389
rect 296 599 352 619
rect 296 565 307 599
rect 341 565 352 599
rect 296 508 352 565
rect 296 474 307 508
rect 341 474 352 508
rect 296 413 352 474
rect 296 379 307 413
rect 341 379 352 413
rect 296 367 352 379
rect 382 607 438 619
rect 382 573 393 607
rect 427 573 438 607
rect 382 515 438 573
rect 382 481 393 515
rect 427 481 438 515
rect 382 423 438 481
rect 382 389 393 423
rect 427 389 438 423
rect 382 367 438 389
rect 468 599 524 619
rect 468 565 479 599
rect 513 565 524 599
rect 468 508 524 565
rect 468 474 479 508
rect 513 474 524 508
rect 468 413 524 474
rect 468 379 479 413
rect 513 379 524 413
rect 468 367 524 379
rect 554 607 610 619
rect 554 573 565 607
rect 599 573 610 607
rect 554 515 610 573
rect 554 481 565 515
rect 599 481 610 515
rect 554 423 610 481
rect 554 389 565 423
rect 599 389 610 423
rect 554 367 610 389
rect 640 599 696 619
rect 640 565 651 599
rect 685 565 696 599
rect 640 508 696 565
rect 640 474 651 508
rect 685 474 696 508
rect 640 413 696 474
rect 640 379 651 413
rect 685 379 696 413
rect 640 367 696 379
rect 726 607 804 619
rect 726 573 748 607
rect 782 573 804 607
rect 726 495 804 573
rect 726 461 748 495
rect 782 461 804 495
rect 726 367 804 461
rect 834 599 890 619
rect 834 565 845 599
rect 879 565 890 599
rect 834 520 890 565
rect 834 486 845 520
rect 879 486 890 520
rect 834 423 890 486
rect 834 389 845 423
rect 879 389 890 423
rect 834 367 890 389
rect 920 607 976 619
rect 920 573 931 607
rect 965 573 976 607
rect 920 495 976 573
rect 920 461 931 495
rect 965 461 976 495
rect 920 367 976 461
rect 1006 599 1062 619
rect 1006 565 1017 599
rect 1051 565 1062 599
rect 1006 520 1062 565
rect 1006 486 1017 520
rect 1051 486 1062 520
rect 1006 423 1062 486
rect 1006 389 1017 423
rect 1051 389 1062 423
rect 1006 367 1062 389
rect 1092 607 1145 619
rect 1092 573 1103 607
rect 1137 573 1145 607
rect 1092 495 1145 573
rect 1092 461 1103 495
rect 1137 461 1145 495
rect 1092 367 1145 461
rect 1199 607 1252 619
rect 1199 573 1207 607
rect 1241 573 1252 607
rect 1199 495 1252 573
rect 1199 461 1207 495
rect 1241 461 1252 495
rect 1199 367 1252 461
rect 1282 531 1338 619
rect 1282 497 1293 531
rect 1327 497 1338 531
rect 1282 423 1338 497
rect 1282 389 1293 423
rect 1327 389 1338 423
rect 1282 367 1338 389
rect 1368 607 1424 619
rect 1368 573 1379 607
rect 1413 573 1424 607
rect 1368 495 1424 573
rect 1368 461 1379 495
rect 1413 461 1424 495
rect 1368 367 1424 461
rect 1454 531 1510 619
rect 1454 497 1465 531
rect 1499 497 1510 531
rect 1454 439 1510 497
rect 1454 405 1465 439
rect 1499 405 1510 439
rect 1454 367 1510 405
rect 1540 607 1596 619
rect 1540 573 1551 607
rect 1585 573 1596 607
rect 1540 513 1596 573
rect 1540 479 1551 513
rect 1585 479 1596 513
rect 1540 423 1596 479
rect 1540 389 1551 423
rect 1585 389 1596 423
rect 1540 367 1596 389
rect 1626 531 1682 619
rect 1626 497 1637 531
rect 1671 497 1682 531
rect 1626 413 1682 497
rect 1626 379 1637 413
rect 1671 379 1682 413
rect 1626 367 1682 379
rect 1712 607 1768 619
rect 1712 573 1723 607
rect 1757 573 1768 607
rect 1712 513 1768 573
rect 1712 479 1723 513
rect 1757 479 1768 513
rect 1712 423 1768 479
rect 1712 389 1723 423
rect 1757 389 1768 423
rect 1712 367 1768 389
rect 1798 531 1854 619
rect 1798 497 1809 531
rect 1843 497 1854 531
rect 1798 413 1854 497
rect 1798 379 1809 413
rect 1843 379 1854 413
rect 1798 367 1854 379
rect 1884 599 1937 619
rect 1884 565 1895 599
rect 1929 565 1937 599
rect 1884 505 1937 565
rect 1884 471 1895 505
rect 1929 471 1937 505
rect 1884 413 1937 471
rect 1884 379 1895 413
rect 1929 379 1937 413
rect 1884 367 1937 379
<< ndiffc >>
rect 35 158 69 192
rect 35 67 69 101
rect 121 98 155 132
rect 207 158 241 192
rect 207 67 241 101
rect 293 98 327 132
rect 379 158 413 192
rect 379 67 413 101
rect 465 90 499 124
rect 551 149 585 183
rect 637 90 671 124
rect 723 149 757 183
rect 827 147 861 181
rect 913 90 947 124
rect 999 147 1033 181
rect 1085 90 1119 124
rect 1171 158 1205 192
rect 1171 67 1205 101
rect 1259 98 1293 132
rect 1345 158 1379 192
rect 1345 67 1379 101
rect 1440 98 1474 132
rect 1537 158 1571 192
rect 1537 67 1571 101
rect 1623 98 1657 132
rect 1709 158 1743 192
rect 1709 67 1743 101
rect 1795 98 1829 132
rect 1881 158 1915 192
rect 1881 67 1915 101
<< pdiffc >>
rect 49 573 83 607
rect 49 476 83 510
rect 49 379 83 413
rect 135 565 169 599
rect 135 474 169 508
rect 135 379 169 413
rect 221 573 255 607
rect 221 481 255 515
rect 221 389 255 423
rect 307 565 341 599
rect 307 474 341 508
rect 307 379 341 413
rect 393 573 427 607
rect 393 481 427 515
rect 393 389 427 423
rect 479 565 513 599
rect 479 474 513 508
rect 479 379 513 413
rect 565 573 599 607
rect 565 481 599 515
rect 565 389 599 423
rect 651 565 685 599
rect 651 474 685 508
rect 651 379 685 413
rect 748 573 782 607
rect 748 461 782 495
rect 845 565 879 599
rect 845 486 879 520
rect 845 389 879 423
rect 931 573 965 607
rect 931 461 965 495
rect 1017 565 1051 599
rect 1017 486 1051 520
rect 1017 389 1051 423
rect 1103 573 1137 607
rect 1103 461 1137 495
rect 1207 573 1241 607
rect 1207 461 1241 495
rect 1293 497 1327 531
rect 1293 389 1327 423
rect 1379 573 1413 607
rect 1379 461 1413 495
rect 1465 497 1499 531
rect 1465 405 1499 439
rect 1551 573 1585 607
rect 1551 479 1585 513
rect 1551 389 1585 423
rect 1637 497 1671 531
rect 1637 379 1671 413
rect 1723 573 1757 607
rect 1723 479 1757 513
rect 1723 389 1757 423
rect 1809 497 1843 531
rect 1809 379 1843 413
rect 1895 565 1929 599
rect 1895 471 1929 505
rect 1895 379 1929 413
<< poly >>
rect 94 619 124 645
rect 180 619 210 645
rect 266 619 296 645
rect 352 619 382 645
rect 438 619 468 645
rect 524 619 554 645
rect 610 619 640 645
rect 696 619 726 645
rect 804 619 834 645
rect 890 619 920 645
rect 976 619 1006 645
rect 1062 619 1092 645
rect 1252 619 1282 645
rect 1338 619 1368 645
rect 1424 619 1454 645
rect 1510 619 1540 645
rect 1596 619 1626 645
rect 1682 619 1712 645
rect 1768 619 1798 645
rect 1854 619 1884 645
rect 94 303 124 367
rect 180 303 210 367
rect 266 303 296 367
rect 352 303 382 367
rect 438 303 468 367
rect 524 303 554 367
rect 610 303 640 367
rect 696 303 726 367
rect 804 333 834 367
rect 890 333 920 367
rect 976 333 1006 367
rect 1062 333 1092 367
rect 804 303 1092 333
rect 1252 303 1282 367
rect 1338 303 1368 367
rect 1424 303 1454 367
rect 1510 303 1540 367
rect 1596 303 1626 367
rect 1682 303 1712 367
rect 1768 303 1798 367
rect 1854 303 1884 367
rect 30 287 382 303
rect 30 253 46 287
rect 80 253 114 287
rect 148 253 182 287
rect 216 253 250 287
rect 284 253 318 287
rect 352 273 382 287
rect 424 287 762 303
rect 352 253 368 273
rect 30 237 368 253
rect 80 215 110 237
rect 166 215 196 237
rect 252 215 282 237
rect 338 215 368 237
rect 424 253 440 287
rect 474 253 508 287
rect 542 253 576 287
rect 610 253 644 287
rect 678 253 712 287
rect 746 253 762 287
rect 424 237 762 253
rect 869 287 1139 303
rect 869 253 885 287
rect 919 253 953 287
rect 987 253 1021 287
rect 1055 253 1089 287
rect 1123 267 1139 287
rect 1202 287 1540 303
rect 1123 253 1160 267
rect 869 237 1160 253
rect 1202 253 1218 287
rect 1252 253 1286 287
rect 1320 253 1354 287
rect 1388 253 1422 287
rect 1456 253 1490 287
rect 1524 253 1540 287
rect 1202 237 1540 253
rect 1582 287 1988 303
rect 1582 253 1598 287
rect 1632 253 1666 287
rect 1700 253 1734 287
rect 1768 253 1802 287
rect 1836 253 1870 287
rect 1904 253 1938 287
rect 1972 253 1988 287
rect 1582 237 1988 253
rect 424 215 454 237
rect 510 215 540 237
rect 596 215 626 237
rect 682 215 712 237
rect 872 215 902 237
rect 958 215 988 237
rect 1044 215 1074 237
rect 1130 215 1160 237
rect 1218 215 1248 237
rect 1304 215 1334 237
rect 1390 215 1420 237
rect 1496 215 1526 237
rect 1582 215 1612 237
rect 1668 215 1698 237
rect 1754 215 1784 237
rect 1840 215 1870 237
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 424 21 454 47
rect 510 21 540 47
rect 596 21 626 47
rect 682 21 712 47
rect 872 21 902 47
rect 958 21 988 47
rect 1044 21 1074 47
rect 1130 21 1160 47
rect 1218 21 1248 47
rect 1304 21 1334 47
rect 1390 21 1420 47
rect 1496 21 1526 47
rect 1582 21 1612 47
rect 1668 21 1698 47
rect 1754 21 1784 47
rect 1840 21 1870 47
<< polycont >>
rect 46 253 80 287
rect 114 253 148 287
rect 182 253 216 287
rect 250 253 284 287
rect 318 253 352 287
rect 440 253 474 287
rect 508 253 542 287
rect 576 253 610 287
rect 644 253 678 287
rect 712 253 746 287
rect 885 253 919 287
rect 953 253 987 287
rect 1021 253 1055 287
rect 1089 253 1123 287
rect 1218 253 1252 287
rect 1286 253 1320 287
rect 1354 253 1388 287
rect 1422 253 1456 287
rect 1490 253 1524 287
rect 1598 253 1632 287
rect 1666 253 1700 287
rect 1734 253 1768 287
rect 1802 253 1836 287
rect 1870 253 1904 287
rect 1938 253 1972 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 33 607 99 649
rect 33 573 49 607
rect 83 573 99 607
rect 33 510 99 573
rect 33 476 49 510
rect 83 476 99 510
rect 33 413 99 476
rect 33 379 49 413
rect 83 379 99 413
rect 33 363 99 379
rect 133 599 171 615
rect 133 565 135 599
rect 169 565 171 599
rect 133 508 171 565
rect 133 474 135 508
rect 169 474 171 508
rect 133 413 171 474
rect 133 379 135 413
rect 169 379 171 413
rect 205 607 271 649
rect 205 573 221 607
rect 255 573 271 607
rect 205 515 271 573
rect 205 481 221 515
rect 255 481 271 515
rect 205 423 271 481
rect 205 389 221 423
rect 255 389 271 423
rect 305 599 343 615
rect 305 565 307 599
rect 341 565 343 599
rect 305 508 343 565
rect 305 474 307 508
rect 341 474 343 508
rect 305 413 343 474
rect 133 355 171 379
rect 305 379 307 413
rect 341 379 343 413
rect 377 607 443 649
rect 377 573 393 607
rect 427 573 443 607
rect 377 515 443 573
rect 377 481 393 515
rect 427 481 443 515
rect 377 423 443 481
rect 377 389 393 423
rect 427 389 443 423
rect 477 599 515 615
rect 477 565 479 599
rect 513 565 515 599
rect 477 508 515 565
rect 477 474 479 508
rect 513 474 515 508
rect 477 413 515 474
rect 305 355 343 379
rect 477 379 479 413
rect 513 379 515 413
rect 549 607 615 649
rect 549 573 565 607
rect 599 573 615 607
rect 549 515 615 573
rect 549 481 565 515
rect 599 481 615 515
rect 549 423 615 481
rect 549 389 565 423
rect 599 389 615 423
rect 649 599 698 615
rect 649 565 651 599
rect 685 565 698 599
rect 649 508 698 565
rect 649 474 651 508
rect 685 474 698 508
rect 649 423 698 474
rect 732 607 798 649
rect 732 573 748 607
rect 782 573 798 607
rect 732 495 798 573
rect 732 461 748 495
rect 782 461 798 495
rect 732 457 798 461
rect 832 599 881 615
rect 832 565 845 599
rect 879 565 881 599
rect 832 520 881 565
rect 832 486 845 520
rect 879 486 881 520
rect 832 423 881 486
rect 915 607 981 649
rect 915 573 931 607
rect 965 573 981 607
rect 915 495 981 573
rect 915 461 931 495
rect 965 461 981 495
rect 915 457 981 461
rect 1015 599 1053 615
rect 1015 565 1017 599
rect 1051 565 1053 599
rect 1015 520 1053 565
rect 1015 486 1017 520
rect 1051 486 1053 520
rect 1015 423 1053 486
rect 1087 607 1153 649
rect 1087 573 1103 607
rect 1137 573 1153 607
rect 1087 495 1153 573
rect 1087 461 1103 495
rect 1137 461 1153 495
rect 1087 457 1153 461
rect 1191 607 1945 615
rect 1191 573 1207 607
rect 1241 581 1379 607
rect 1241 573 1257 581
rect 1191 495 1257 573
rect 1363 573 1379 581
rect 1413 581 1551 607
rect 1413 573 1429 581
rect 1191 461 1207 495
rect 1241 461 1257 495
rect 1191 457 1257 461
rect 1291 531 1329 547
rect 1291 497 1293 531
rect 1327 497 1329 531
rect 1291 423 1329 497
rect 1363 495 1429 573
rect 1535 573 1551 581
rect 1585 581 1723 607
rect 1585 573 1601 581
rect 1363 461 1379 495
rect 1413 461 1429 495
rect 1363 457 1429 461
rect 1463 531 1501 547
rect 1463 497 1465 531
rect 1499 497 1501 531
rect 1463 439 1501 497
rect 1463 423 1465 439
rect 649 413 845 423
rect 477 355 515 379
rect 649 379 651 413
rect 685 389 845 413
rect 879 389 1017 423
rect 1051 389 1293 423
rect 1327 405 1465 423
rect 1499 405 1501 439
rect 1327 389 1501 405
rect 1535 513 1601 573
rect 1707 573 1723 581
rect 1757 599 1945 607
rect 1757 581 1895 599
rect 1757 573 1773 581
rect 1535 479 1551 513
rect 1585 479 1601 513
rect 1535 423 1601 479
rect 1535 389 1551 423
rect 1585 389 1601 423
rect 1635 531 1673 547
rect 1635 497 1637 531
rect 1671 497 1673 531
rect 1635 413 1673 497
rect 685 379 701 389
rect 649 355 701 379
rect 1635 379 1637 413
rect 1671 379 1673 413
rect 1707 513 1773 573
rect 1887 565 1895 581
rect 1929 565 1945 599
rect 1707 479 1723 513
rect 1757 479 1773 513
rect 1707 423 1773 479
rect 1707 389 1723 423
rect 1757 389 1773 423
rect 1807 531 1853 547
rect 1807 497 1809 531
rect 1843 497 1853 531
rect 1807 413 1853 497
rect 1635 355 1673 379
rect 1807 379 1809 413
rect 1843 379 1853 413
rect 1807 355 1853 379
rect 1887 505 1945 565
rect 1887 471 1895 505
rect 1929 471 1945 505
rect 1887 413 1945 471
rect 1887 379 1895 413
rect 1929 379 1945 413
rect 1887 363 1945 379
rect 133 321 701 355
rect 799 321 1853 355
rect 17 253 46 287
rect 80 253 114 287
rect 148 253 182 287
rect 216 253 250 287
rect 284 253 318 287
rect 352 253 368 287
rect 17 242 368 253
rect 402 253 440 287
rect 474 253 508 287
rect 542 253 576 287
rect 610 253 644 287
rect 678 253 712 287
rect 746 253 762 287
rect 402 242 762 253
rect 799 208 835 321
rect 869 253 885 287
rect 919 253 953 287
rect 987 253 1021 287
rect 1055 253 1089 287
rect 1123 253 1139 287
rect 869 242 1139 253
rect 1173 253 1218 287
rect 1252 253 1286 287
rect 1320 253 1354 287
rect 1388 253 1422 287
rect 1456 253 1490 287
rect 1524 253 1540 287
rect 1173 242 1540 253
rect 1582 253 1598 287
rect 1632 253 1666 287
rect 1700 253 1734 287
rect 1768 253 1802 287
rect 1836 253 1870 287
rect 1904 253 1938 287
rect 1972 253 1999 287
rect 1582 242 1999 253
rect 19 192 765 208
rect 19 158 35 192
rect 69 174 207 192
rect 69 158 71 174
rect 19 101 71 158
rect 205 158 207 174
rect 241 174 379 192
rect 241 158 243 174
rect 19 67 35 101
rect 69 67 71 101
rect 19 51 71 67
rect 105 132 171 140
rect 105 98 121 132
rect 155 98 171 132
rect 105 17 171 98
rect 205 101 243 158
rect 377 158 379 174
rect 413 183 765 192
rect 413 174 551 183
rect 413 158 423 174
rect 205 67 207 101
rect 241 67 243 101
rect 205 51 243 67
rect 277 132 343 140
rect 277 98 293 132
rect 327 98 343 132
rect 277 17 343 98
rect 377 101 423 158
rect 542 149 551 174
rect 585 174 723 183
rect 585 149 593 174
rect 377 67 379 101
rect 413 67 423 101
rect 377 51 423 67
rect 457 124 508 140
rect 542 133 593 149
rect 714 149 723 174
rect 757 149 765 183
rect 457 90 465 124
rect 499 90 508 124
rect 457 89 508 90
rect 627 124 680 140
rect 714 133 765 149
rect 799 192 1931 208
rect 799 181 1171 192
rect 799 147 827 181
rect 861 174 999 181
rect 861 147 871 174
rect 799 131 871 147
rect 990 147 999 174
rect 1033 174 1171 181
rect 1033 147 1042 174
rect 627 90 637 124
rect 671 97 680 124
rect 905 124 956 140
rect 990 131 1042 147
rect 1161 158 1171 174
rect 1205 174 1345 192
rect 1205 158 1209 174
rect 905 97 913 124
rect 671 90 913 97
rect 947 97 956 124
rect 1076 124 1127 140
rect 1076 97 1085 124
rect 947 90 1085 97
rect 1119 90 1127 124
rect 627 89 1127 90
rect 457 51 1127 89
rect 1161 101 1209 158
rect 1343 158 1345 174
rect 1379 174 1537 192
rect 1379 158 1390 174
rect 1161 67 1171 101
rect 1205 67 1209 101
rect 1161 51 1209 67
rect 1243 132 1309 140
rect 1243 98 1259 132
rect 1293 98 1309 132
rect 1243 17 1309 98
rect 1343 101 1390 158
rect 1524 158 1537 174
rect 1571 174 1709 192
rect 1571 158 1573 174
rect 1343 67 1345 101
rect 1379 67 1390 101
rect 1343 51 1390 67
rect 1424 132 1490 140
rect 1424 98 1440 132
rect 1474 98 1490 132
rect 1424 17 1490 98
rect 1524 101 1573 158
rect 1707 158 1709 174
rect 1743 174 1881 192
rect 1743 158 1745 174
rect 1524 67 1537 101
rect 1571 67 1573 101
rect 1524 51 1573 67
rect 1607 132 1673 140
rect 1607 98 1623 132
rect 1657 98 1673 132
rect 1607 17 1673 98
rect 1707 101 1745 158
rect 1879 158 1881 174
rect 1915 158 1931 192
rect 1707 67 1709 101
rect 1743 67 1745 101
rect 1707 51 1745 67
rect 1779 132 1845 140
rect 1779 98 1795 132
rect 1829 98 1845 132
rect 1779 17 1845 98
rect 1879 101 1931 158
rect 1879 67 1881 101
rect 1915 67 1931 101
rect 1879 51 1931 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a311oi_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3261568
string GDS_START 3244138
<< end >>
