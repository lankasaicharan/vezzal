magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3506 1975
<< nwell >>
rect -38 331 2246 704
<< pwell >>
rect 383 49 1861 180
rect 0 0 2208 49
<< scnmos >>
rect 462 70 492 154
rect 548 70 578 154
rect 634 70 664 154
rect 720 70 750 154
rect 806 70 836 154
rect 892 70 922 154
rect 978 70 1008 154
rect 1064 70 1094 154
rect 1150 70 1180 154
rect 1236 70 1266 154
rect 1322 70 1352 154
rect 1408 70 1438 154
rect 1494 70 1524 154
rect 1580 70 1610 154
rect 1666 70 1696 154
rect 1752 70 1782 154
<< scpmoshvt >>
rect 118 367 148 619
rect 204 367 234 619
rect 290 367 320 619
rect 376 367 406 619
rect 462 367 492 619
rect 548 367 578 619
rect 634 367 664 619
rect 720 367 750 619
rect 806 367 836 619
rect 892 367 922 619
rect 978 367 1008 619
rect 1064 367 1094 619
rect 1150 367 1180 619
rect 1236 367 1266 619
rect 1322 367 1352 619
rect 1408 367 1438 619
rect 1494 367 1524 619
rect 1580 367 1610 619
rect 1666 367 1696 619
rect 1752 367 1782 619
rect 1838 367 1868 619
rect 1924 367 1954 619
rect 2010 367 2040 619
rect 2096 367 2126 619
<< ndiff >>
rect 409 129 462 154
rect 409 95 417 129
rect 451 95 462 129
rect 409 70 462 95
rect 492 129 548 154
rect 492 95 503 129
rect 537 95 548 129
rect 492 70 548 95
rect 578 129 634 154
rect 578 95 589 129
rect 623 95 634 129
rect 578 70 634 95
rect 664 129 720 154
rect 664 95 675 129
rect 709 95 720 129
rect 664 70 720 95
rect 750 129 806 154
rect 750 95 761 129
rect 795 95 806 129
rect 750 70 806 95
rect 836 129 892 154
rect 836 95 847 129
rect 881 95 892 129
rect 836 70 892 95
rect 922 129 978 154
rect 922 95 933 129
rect 967 95 978 129
rect 922 70 978 95
rect 1008 129 1064 154
rect 1008 95 1019 129
rect 1053 95 1064 129
rect 1008 70 1064 95
rect 1094 129 1150 154
rect 1094 95 1105 129
rect 1139 95 1150 129
rect 1094 70 1150 95
rect 1180 129 1236 154
rect 1180 95 1191 129
rect 1225 95 1236 129
rect 1180 70 1236 95
rect 1266 129 1322 154
rect 1266 95 1277 129
rect 1311 95 1322 129
rect 1266 70 1322 95
rect 1352 129 1408 154
rect 1352 95 1363 129
rect 1397 95 1408 129
rect 1352 70 1408 95
rect 1438 129 1494 154
rect 1438 95 1449 129
rect 1483 95 1494 129
rect 1438 70 1494 95
rect 1524 129 1580 154
rect 1524 95 1535 129
rect 1569 95 1580 129
rect 1524 70 1580 95
rect 1610 129 1666 154
rect 1610 95 1621 129
rect 1655 95 1666 129
rect 1610 70 1666 95
rect 1696 129 1752 154
rect 1696 95 1707 129
rect 1741 95 1752 129
rect 1696 70 1752 95
rect 1782 129 1835 154
rect 1782 95 1793 129
rect 1827 95 1835 129
rect 1782 70 1835 95
<< pdiff >>
rect 61 595 118 619
rect 61 561 73 595
rect 107 561 118 595
rect 61 511 118 561
rect 61 477 73 511
rect 107 477 118 511
rect 61 425 118 477
rect 61 391 73 425
rect 107 391 118 425
rect 61 367 118 391
rect 148 595 204 619
rect 148 561 159 595
rect 193 561 204 595
rect 148 511 204 561
rect 148 477 159 511
rect 193 477 204 511
rect 148 425 204 477
rect 148 391 159 425
rect 193 391 204 425
rect 148 367 204 391
rect 234 595 290 619
rect 234 561 245 595
rect 279 561 290 595
rect 234 511 290 561
rect 234 477 245 511
rect 279 477 290 511
rect 234 425 290 477
rect 234 391 245 425
rect 279 391 290 425
rect 234 367 290 391
rect 320 595 376 619
rect 320 561 331 595
rect 365 561 376 595
rect 320 511 376 561
rect 320 477 331 511
rect 365 477 376 511
rect 320 425 376 477
rect 320 391 331 425
rect 365 391 376 425
rect 320 367 376 391
rect 406 595 462 619
rect 406 561 417 595
rect 451 561 462 595
rect 406 511 462 561
rect 406 477 417 511
rect 451 477 462 511
rect 406 425 462 477
rect 406 391 417 425
rect 451 391 462 425
rect 406 367 462 391
rect 492 595 548 619
rect 492 561 503 595
rect 537 561 548 595
rect 492 511 548 561
rect 492 477 503 511
rect 537 477 548 511
rect 492 425 548 477
rect 492 391 503 425
rect 537 391 548 425
rect 492 367 548 391
rect 578 595 634 619
rect 578 561 589 595
rect 623 561 634 595
rect 578 511 634 561
rect 578 477 589 511
rect 623 477 634 511
rect 578 425 634 477
rect 578 391 589 425
rect 623 391 634 425
rect 578 367 634 391
rect 664 595 720 619
rect 664 561 675 595
rect 709 561 720 595
rect 664 511 720 561
rect 664 477 675 511
rect 709 477 720 511
rect 664 425 720 477
rect 664 391 675 425
rect 709 391 720 425
rect 664 367 720 391
rect 750 595 806 619
rect 750 561 761 595
rect 795 561 806 595
rect 750 511 806 561
rect 750 477 761 511
rect 795 477 806 511
rect 750 425 806 477
rect 750 391 761 425
rect 795 391 806 425
rect 750 367 806 391
rect 836 595 892 619
rect 836 561 847 595
rect 881 561 892 595
rect 836 511 892 561
rect 836 477 847 511
rect 881 477 892 511
rect 836 425 892 477
rect 836 391 847 425
rect 881 391 892 425
rect 836 367 892 391
rect 922 595 978 619
rect 922 561 933 595
rect 967 561 978 595
rect 922 511 978 561
rect 922 477 933 511
rect 967 477 978 511
rect 922 425 978 477
rect 922 391 933 425
rect 967 391 978 425
rect 922 367 978 391
rect 1008 595 1064 619
rect 1008 561 1019 595
rect 1053 561 1064 595
rect 1008 511 1064 561
rect 1008 477 1019 511
rect 1053 477 1064 511
rect 1008 425 1064 477
rect 1008 391 1019 425
rect 1053 391 1064 425
rect 1008 367 1064 391
rect 1094 595 1150 619
rect 1094 561 1105 595
rect 1139 561 1150 595
rect 1094 511 1150 561
rect 1094 477 1105 511
rect 1139 477 1150 511
rect 1094 425 1150 477
rect 1094 391 1105 425
rect 1139 391 1150 425
rect 1094 367 1150 391
rect 1180 595 1236 619
rect 1180 561 1191 595
rect 1225 561 1236 595
rect 1180 511 1236 561
rect 1180 477 1191 511
rect 1225 477 1236 511
rect 1180 425 1236 477
rect 1180 391 1191 425
rect 1225 391 1236 425
rect 1180 367 1236 391
rect 1266 595 1322 619
rect 1266 561 1277 595
rect 1311 561 1322 595
rect 1266 511 1322 561
rect 1266 477 1277 511
rect 1311 477 1322 511
rect 1266 425 1322 477
rect 1266 391 1277 425
rect 1311 391 1322 425
rect 1266 367 1322 391
rect 1352 595 1408 619
rect 1352 561 1363 595
rect 1397 561 1408 595
rect 1352 511 1408 561
rect 1352 477 1363 511
rect 1397 477 1408 511
rect 1352 425 1408 477
rect 1352 391 1363 425
rect 1397 391 1408 425
rect 1352 367 1408 391
rect 1438 595 1494 619
rect 1438 561 1449 595
rect 1483 561 1494 595
rect 1438 511 1494 561
rect 1438 477 1449 511
rect 1483 477 1494 511
rect 1438 425 1494 477
rect 1438 391 1449 425
rect 1483 391 1494 425
rect 1438 367 1494 391
rect 1524 595 1580 619
rect 1524 561 1535 595
rect 1569 561 1580 595
rect 1524 511 1580 561
rect 1524 477 1535 511
rect 1569 477 1580 511
rect 1524 425 1580 477
rect 1524 391 1535 425
rect 1569 391 1580 425
rect 1524 367 1580 391
rect 1610 595 1666 619
rect 1610 561 1621 595
rect 1655 561 1666 595
rect 1610 511 1666 561
rect 1610 477 1621 511
rect 1655 477 1666 511
rect 1610 425 1666 477
rect 1610 391 1621 425
rect 1655 391 1666 425
rect 1610 367 1666 391
rect 1696 595 1752 619
rect 1696 561 1707 595
rect 1741 561 1752 595
rect 1696 511 1752 561
rect 1696 477 1707 511
rect 1741 477 1752 511
rect 1696 425 1752 477
rect 1696 391 1707 425
rect 1741 391 1752 425
rect 1696 367 1752 391
rect 1782 595 1838 619
rect 1782 561 1793 595
rect 1827 561 1838 595
rect 1782 511 1838 561
rect 1782 477 1793 511
rect 1827 477 1838 511
rect 1782 425 1838 477
rect 1782 391 1793 425
rect 1827 391 1838 425
rect 1782 367 1838 391
rect 1868 595 1924 619
rect 1868 561 1879 595
rect 1913 561 1924 595
rect 1868 511 1924 561
rect 1868 477 1879 511
rect 1913 477 1924 511
rect 1868 425 1924 477
rect 1868 391 1879 425
rect 1913 391 1924 425
rect 1868 367 1924 391
rect 1954 595 2010 619
rect 1954 561 1965 595
rect 1999 561 2010 595
rect 1954 511 2010 561
rect 1954 477 1965 511
rect 1999 477 2010 511
rect 1954 425 2010 477
rect 1954 391 1965 425
rect 1999 391 2010 425
rect 1954 367 2010 391
rect 2040 595 2096 619
rect 2040 561 2051 595
rect 2085 561 2096 595
rect 2040 511 2096 561
rect 2040 477 2051 511
rect 2085 477 2096 511
rect 2040 425 2096 477
rect 2040 391 2051 425
rect 2085 391 2096 425
rect 2040 367 2096 391
rect 2126 595 2179 619
rect 2126 561 2137 595
rect 2171 561 2179 595
rect 2126 511 2179 561
rect 2126 477 2137 511
rect 2171 477 2179 511
rect 2126 425 2179 477
rect 2126 391 2137 425
rect 2171 391 2179 425
rect 2126 367 2179 391
<< ndiffc >>
rect 417 95 451 129
rect 503 95 537 129
rect 589 95 623 129
rect 675 95 709 129
rect 761 95 795 129
rect 847 95 881 129
rect 933 95 967 129
rect 1019 95 1053 129
rect 1105 95 1139 129
rect 1191 95 1225 129
rect 1277 95 1311 129
rect 1363 95 1397 129
rect 1449 95 1483 129
rect 1535 95 1569 129
rect 1621 95 1655 129
rect 1707 95 1741 129
rect 1793 95 1827 129
<< pdiffc >>
rect 73 561 107 595
rect 73 477 107 511
rect 73 391 107 425
rect 159 561 193 595
rect 159 477 193 511
rect 159 391 193 425
rect 245 561 279 595
rect 245 477 279 511
rect 245 391 279 425
rect 331 561 365 595
rect 331 477 365 511
rect 331 391 365 425
rect 417 561 451 595
rect 417 477 451 511
rect 417 391 451 425
rect 503 561 537 595
rect 503 477 537 511
rect 503 391 537 425
rect 589 561 623 595
rect 589 477 623 511
rect 589 391 623 425
rect 675 561 709 595
rect 675 477 709 511
rect 675 391 709 425
rect 761 561 795 595
rect 761 477 795 511
rect 761 391 795 425
rect 847 561 881 595
rect 847 477 881 511
rect 847 391 881 425
rect 933 561 967 595
rect 933 477 967 511
rect 933 391 967 425
rect 1019 561 1053 595
rect 1019 477 1053 511
rect 1019 391 1053 425
rect 1105 561 1139 595
rect 1105 477 1139 511
rect 1105 391 1139 425
rect 1191 561 1225 595
rect 1191 477 1225 511
rect 1191 391 1225 425
rect 1277 561 1311 595
rect 1277 477 1311 511
rect 1277 391 1311 425
rect 1363 561 1397 595
rect 1363 477 1397 511
rect 1363 391 1397 425
rect 1449 561 1483 595
rect 1449 477 1483 511
rect 1449 391 1483 425
rect 1535 561 1569 595
rect 1535 477 1569 511
rect 1535 391 1569 425
rect 1621 561 1655 595
rect 1621 477 1655 511
rect 1621 391 1655 425
rect 1707 561 1741 595
rect 1707 477 1741 511
rect 1707 391 1741 425
rect 1793 561 1827 595
rect 1793 477 1827 511
rect 1793 391 1827 425
rect 1879 561 1913 595
rect 1879 477 1913 511
rect 1879 391 1913 425
rect 1965 561 1999 595
rect 1965 477 1999 511
rect 1965 391 1999 425
rect 2051 561 2085 595
rect 2051 477 2085 511
rect 2051 391 2085 425
rect 2137 561 2171 595
rect 2137 477 2171 511
rect 2137 391 2171 425
<< poly >>
rect 118 619 148 645
rect 204 619 234 645
rect 290 619 320 645
rect 376 619 406 645
rect 462 619 492 645
rect 548 619 578 645
rect 634 619 664 645
rect 720 619 750 645
rect 806 619 836 645
rect 892 619 922 645
rect 978 619 1008 645
rect 1064 619 1094 645
rect 1150 619 1180 645
rect 1236 619 1266 645
rect 1322 619 1352 645
rect 1408 619 1438 645
rect 1494 619 1524 645
rect 1580 619 1610 645
rect 1666 619 1696 645
rect 1752 619 1782 645
rect 1838 619 1868 645
rect 1924 619 1954 645
rect 2010 619 2040 645
rect 2096 619 2126 645
rect 118 325 148 367
rect 204 325 234 367
rect 290 325 320 367
rect 376 325 406 367
rect 462 325 492 367
rect 548 325 578 367
rect 634 325 664 367
rect 720 325 750 367
rect 806 325 836 367
rect 892 325 922 367
rect 978 325 1008 367
rect 1064 325 1094 367
rect 1150 325 1180 367
rect 1236 325 1266 367
rect 1322 325 1352 367
rect 1408 325 1438 367
rect 1494 325 1524 367
rect 1580 325 1610 367
rect 1666 325 1696 367
rect 1752 325 1782 367
rect 1838 325 1868 367
rect 1924 325 1954 367
rect 2010 325 2040 367
rect 2096 325 2126 367
rect 118 309 2126 325
rect 118 275 155 309
rect 189 275 223 309
rect 257 275 291 309
rect 325 275 359 309
rect 393 275 427 309
rect 461 275 590 309
rect 624 275 761 309
rect 795 275 934 309
rect 968 275 1105 309
rect 1139 275 1278 309
rect 1312 275 1450 309
rect 1484 275 1622 309
rect 1656 275 1787 309
rect 1821 275 1855 309
rect 1889 275 1923 309
rect 1957 275 1991 309
rect 2025 275 2059 309
rect 2093 275 2126 309
rect 118 259 2126 275
rect 462 154 492 259
rect 548 154 578 259
rect 634 154 664 259
rect 720 154 750 259
rect 806 154 836 259
rect 892 154 922 259
rect 978 154 1008 259
rect 1064 154 1094 259
rect 1150 154 1180 259
rect 1236 154 1266 259
rect 1322 154 1352 259
rect 1408 154 1438 259
rect 1494 154 1524 259
rect 1580 154 1610 259
rect 1666 154 1696 259
rect 1752 154 1782 259
rect 462 44 492 70
rect 548 44 578 70
rect 634 44 664 70
rect 720 44 750 70
rect 806 44 836 70
rect 892 44 922 70
rect 978 44 1008 70
rect 1064 44 1094 70
rect 1150 44 1180 70
rect 1236 44 1266 70
rect 1322 44 1352 70
rect 1408 44 1438 70
rect 1494 44 1524 70
rect 1580 44 1610 70
rect 1666 44 1696 70
rect 1752 44 1782 70
<< polycont >>
rect 155 275 189 309
rect 223 275 257 309
rect 291 275 325 309
rect 359 275 393 309
rect 427 275 461 309
rect 590 275 624 309
rect 761 275 795 309
rect 934 275 968 309
rect 1105 275 1139 309
rect 1278 275 1312 309
rect 1450 275 1484 309
rect 1622 275 1656 309
rect 1787 275 1821 309
rect 1855 275 1889 309
rect 1923 275 1957 309
rect 1991 275 2025 309
rect 2059 275 2093 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 64 595 116 649
rect 64 561 73 595
rect 107 561 116 595
rect 64 511 116 561
rect 64 477 73 511
rect 107 477 116 511
rect 64 425 116 477
rect 64 391 73 425
rect 107 391 116 425
rect 64 367 116 391
rect 151 595 202 611
rect 151 561 159 595
rect 193 561 202 595
rect 151 511 202 561
rect 151 477 159 511
rect 193 477 202 511
rect 151 425 202 477
rect 151 390 159 425
rect 193 390 202 425
rect 151 367 202 390
rect 236 595 288 649
rect 236 561 245 595
rect 279 561 288 595
rect 236 511 288 561
rect 236 477 245 511
rect 279 477 288 511
rect 236 425 288 477
rect 236 391 245 425
rect 279 391 288 425
rect 236 367 288 391
rect 323 595 374 611
rect 323 561 331 595
rect 365 561 374 595
rect 323 511 374 561
rect 323 477 331 511
rect 365 477 374 511
rect 323 425 374 477
rect 323 390 331 425
rect 365 390 374 425
rect 323 367 374 390
rect 408 595 460 649
rect 408 561 417 595
rect 451 561 460 595
rect 408 511 460 561
rect 408 477 417 511
rect 451 477 460 511
rect 408 425 460 477
rect 408 391 417 425
rect 451 391 460 425
rect 408 367 460 391
rect 495 595 546 611
rect 495 561 503 595
rect 537 561 546 595
rect 495 511 546 561
rect 495 477 503 511
rect 537 477 546 511
rect 495 425 546 477
rect 495 390 503 425
rect 537 390 546 425
rect 118 309 461 325
rect 118 242 155 309
rect 189 275 223 309
rect 257 276 291 309
rect 325 276 359 309
rect 393 276 427 309
rect 261 275 291 276
rect 333 275 359 276
rect 405 275 427 276
rect 189 242 227 275
rect 261 242 299 275
rect 333 242 371 275
rect 405 242 461 275
rect 118 232 461 242
rect 407 129 461 145
rect 407 95 417 129
rect 451 95 461 129
rect 407 17 461 95
rect 495 129 546 390
rect 580 595 632 649
rect 580 561 589 595
rect 623 561 632 595
rect 580 511 632 561
rect 580 477 589 511
rect 623 477 632 511
rect 580 425 632 477
rect 580 391 589 425
rect 623 391 632 425
rect 580 367 632 391
rect 667 595 718 611
rect 667 561 675 595
rect 709 561 718 595
rect 667 511 718 561
rect 667 477 675 511
rect 709 477 718 511
rect 667 425 718 477
rect 667 390 675 425
rect 709 390 718 425
rect 580 309 633 325
rect 580 242 590 309
rect 624 242 633 309
rect 580 232 633 242
rect 495 95 503 129
rect 537 95 546 129
rect 495 79 546 95
rect 580 129 633 145
rect 580 95 589 129
rect 623 95 633 129
rect 580 17 633 95
rect 667 129 718 390
rect 752 595 804 649
rect 752 561 761 595
rect 795 561 804 595
rect 752 511 804 561
rect 752 477 761 511
rect 795 477 804 511
rect 752 425 804 477
rect 752 391 761 425
rect 795 391 804 425
rect 752 367 804 391
rect 839 595 890 611
rect 839 561 847 595
rect 881 561 890 595
rect 839 511 890 561
rect 839 477 847 511
rect 881 477 890 511
rect 839 425 890 477
rect 839 390 847 425
rect 881 390 890 425
rect 752 309 805 325
rect 752 242 761 309
rect 795 242 805 309
rect 752 232 805 242
rect 667 95 675 129
rect 709 95 718 129
rect 667 79 718 95
rect 752 129 805 145
rect 752 95 761 129
rect 795 95 805 129
rect 752 17 805 95
rect 839 129 890 390
rect 924 595 976 649
rect 924 561 933 595
rect 967 561 976 595
rect 924 511 976 561
rect 924 477 933 511
rect 967 477 976 511
rect 924 425 976 477
rect 924 391 933 425
rect 967 391 976 425
rect 924 367 976 391
rect 1010 595 1062 611
rect 1010 561 1019 595
rect 1053 561 1062 595
rect 1010 511 1062 561
rect 1010 477 1019 511
rect 1053 477 1062 511
rect 1010 425 1062 477
rect 1010 390 1019 425
rect 1053 390 1062 425
rect 1010 377 1062 390
rect 924 309 977 325
rect 924 242 934 309
rect 968 242 977 309
rect 924 232 977 242
rect 839 95 847 129
rect 881 95 890 129
rect 839 79 890 95
rect 924 129 977 145
rect 924 95 933 129
rect 967 95 977 129
rect 924 17 977 95
rect 1011 129 1062 377
rect 1096 595 1148 649
rect 1096 561 1105 595
rect 1139 561 1148 595
rect 1096 511 1148 561
rect 1096 477 1105 511
rect 1139 477 1148 511
rect 1096 425 1148 477
rect 1096 391 1105 425
rect 1139 391 1148 425
rect 1096 367 1148 391
rect 1183 595 1234 611
rect 1183 561 1191 595
rect 1225 561 1234 595
rect 1183 511 1234 561
rect 1183 477 1191 511
rect 1225 477 1234 511
rect 1183 425 1234 477
rect 1183 390 1191 425
rect 1225 390 1234 425
rect 1096 309 1149 325
rect 1096 242 1105 309
rect 1139 242 1149 309
rect 1096 232 1149 242
rect 1011 95 1019 129
rect 1053 95 1062 129
rect 1011 79 1062 95
rect 1096 129 1149 145
rect 1096 95 1105 129
rect 1139 95 1149 129
rect 1096 17 1149 95
rect 1183 129 1234 390
rect 1268 595 1320 649
rect 1268 561 1277 595
rect 1311 561 1320 595
rect 1268 511 1320 561
rect 1268 477 1277 511
rect 1311 477 1320 511
rect 1268 425 1320 477
rect 1268 391 1277 425
rect 1311 391 1320 425
rect 1268 367 1320 391
rect 1355 595 1406 611
rect 1355 561 1363 595
rect 1397 561 1406 595
rect 1355 511 1406 561
rect 1355 477 1363 511
rect 1397 477 1406 511
rect 1355 425 1406 477
rect 1355 390 1363 425
rect 1397 390 1406 425
rect 1268 309 1321 325
rect 1268 242 1278 309
rect 1312 242 1321 309
rect 1268 232 1321 242
rect 1183 95 1191 129
rect 1225 95 1234 129
rect 1183 79 1234 95
rect 1268 129 1321 145
rect 1268 95 1277 129
rect 1311 95 1321 129
rect 1268 17 1321 95
rect 1355 129 1406 390
rect 1440 595 1492 649
rect 1440 561 1449 595
rect 1483 561 1492 595
rect 1440 511 1492 561
rect 1440 477 1449 511
rect 1483 477 1492 511
rect 1440 425 1492 477
rect 1440 391 1449 425
rect 1483 391 1492 425
rect 1440 367 1492 391
rect 1527 595 1578 611
rect 1527 561 1535 595
rect 1569 561 1578 595
rect 1527 511 1578 561
rect 1527 477 1535 511
rect 1569 477 1578 511
rect 1527 425 1578 477
rect 1527 390 1535 425
rect 1569 390 1578 425
rect 1440 309 1493 325
rect 1440 242 1450 309
rect 1484 242 1493 309
rect 1440 232 1493 242
rect 1355 95 1363 129
rect 1397 95 1406 129
rect 1355 79 1406 95
rect 1440 129 1493 145
rect 1440 95 1449 129
rect 1483 95 1493 129
rect 1440 17 1493 95
rect 1527 129 1578 390
rect 1612 595 1664 649
rect 1612 561 1621 595
rect 1655 561 1664 595
rect 1612 511 1664 561
rect 1612 477 1621 511
rect 1655 477 1664 511
rect 1612 425 1664 477
rect 1612 391 1621 425
rect 1655 391 1664 425
rect 1612 367 1664 391
rect 1699 595 1750 611
rect 1699 561 1707 595
rect 1741 561 1750 595
rect 1699 511 1750 561
rect 1699 477 1707 511
rect 1741 477 1750 511
rect 1699 425 1750 477
rect 1699 390 1707 425
rect 1741 390 1750 425
rect 1612 309 1665 325
rect 1612 242 1622 309
rect 1656 242 1665 309
rect 1612 232 1665 242
rect 1527 95 1535 129
rect 1569 95 1578 129
rect 1527 79 1578 95
rect 1612 129 1665 145
rect 1612 95 1621 129
rect 1655 95 1665 129
rect 1612 17 1665 95
rect 1699 129 1750 390
rect 1784 595 1836 649
rect 1784 561 1793 595
rect 1827 561 1836 595
rect 1784 511 1836 561
rect 1784 477 1793 511
rect 1827 477 1836 511
rect 1784 425 1836 477
rect 1784 391 1793 425
rect 1827 391 1836 425
rect 1784 367 1836 391
rect 1871 595 1922 611
rect 1871 561 1879 595
rect 1913 561 1922 595
rect 1871 511 1922 561
rect 1871 477 1879 511
rect 1913 477 1922 511
rect 1871 425 1922 477
rect 1871 390 1879 425
rect 1913 390 1922 425
rect 1871 367 1922 390
rect 1956 595 2008 649
rect 1956 561 1965 595
rect 1999 561 2008 595
rect 1956 511 2008 561
rect 1956 477 1965 511
rect 1999 477 2008 511
rect 1956 425 2008 477
rect 1956 391 1965 425
rect 1999 391 2008 425
rect 1956 367 2008 391
rect 2042 595 2094 611
rect 2042 561 2051 595
rect 2085 561 2094 595
rect 2042 511 2094 561
rect 2042 477 2051 511
rect 2085 477 2094 511
rect 2042 425 2094 477
rect 2042 390 2051 425
rect 2085 390 2094 425
rect 2042 367 2094 390
rect 2128 595 2179 649
rect 2128 561 2137 595
rect 2171 561 2179 595
rect 2128 511 2179 561
rect 2128 477 2137 511
rect 2171 477 2179 511
rect 2128 425 2179 477
rect 2128 391 2137 425
rect 2171 391 2179 425
rect 2128 367 2179 391
rect 1784 309 2109 325
rect 1784 275 1787 309
rect 1821 276 1855 309
rect 1889 276 1923 309
rect 1957 276 1991 309
rect 1821 275 1843 276
rect 1889 275 1915 276
rect 1957 275 1987 276
rect 2025 275 2059 309
rect 1784 242 1843 275
rect 1877 242 1915 275
rect 1949 242 1987 275
rect 2021 242 2059 275
rect 2093 242 2109 309
rect 1784 232 2109 242
rect 1699 95 1707 129
rect 1741 95 1750 129
rect 1699 79 1750 95
rect 1784 129 1837 145
rect 1784 95 1793 129
rect 1827 95 1837 129
rect 1784 17 1837 95
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 159 391 193 424
rect 159 390 193 391
rect 331 391 365 424
rect 331 390 365 391
rect 503 391 537 424
rect 503 390 537 391
rect 155 275 189 276
rect 227 275 257 276
rect 257 275 261 276
rect 299 275 325 276
rect 325 275 333 276
rect 371 275 393 276
rect 393 275 405 276
rect 155 242 189 275
rect 227 242 261 275
rect 299 242 333 275
rect 371 242 405 275
rect 675 391 709 424
rect 675 390 709 391
rect 590 275 624 276
rect 590 242 624 275
rect 847 391 881 424
rect 847 390 881 391
rect 761 275 795 276
rect 761 242 795 275
rect 1019 391 1053 424
rect 1019 390 1053 391
rect 934 275 968 276
rect 934 242 968 275
rect 1191 391 1225 424
rect 1191 390 1225 391
rect 1105 275 1139 276
rect 1105 242 1139 275
rect 1363 391 1397 424
rect 1363 390 1397 391
rect 1278 275 1312 276
rect 1278 242 1312 275
rect 1535 391 1569 424
rect 1535 390 1569 391
rect 1450 275 1484 276
rect 1450 242 1484 275
rect 1707 391 1741 424
rect 1707 390 1741 391
rect 1622 275 1656 276
rect 1622 242 1656 275
rect 1879 391 1913 424
rect 1879 390 1913 391
rect 2051 391 2085 424
rect 2051 390 2085 391
rect 1843 275 1855 276
rect 1855 275 1877 276
rect 1915 275 1923 276
rect 1923 275 1949 276
rect 1987 275 1991 276
rect 1991 275 2021 276
rect 2059 275 2093 276
rect 1843 242 1877 275
rect 1915 242 1949 275
rect 1987 242 2021 275
rect 2059 242 2093 275
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 147 424 2097 430
rect 147 390 159 424
rect 193 390 331 424
rect 365 390 503 424
rect 537 390 675 424
rect 709 390 847 424
rect 881 390 1019 424
rect 1053 390 1191 424
rect 1225 390 1363 424
rect 1397 390 1535 424
rect 1569 390 1707 424
rect 1741 390 1879 424
rect 1913 390 2051 424
rect 2085 390 2097 424
rect 147 384 2097 390
rect 143 276 2105 282
rect 143 242 155 276
rect 189 242 227 276
rect 261 242 299 276
rect 333 242 371 276
rect 405 242 590 276
rect 624 242 761 276
rect 795 242 934 276
rect 968 242 1105 276
rect 1139 242 1278 276
rect 1312 242 1450 276
rect 1484 242 1622 276
rect 1656 242 1843 276
rect 1877 242 1915 276
rect 1949 242 1987 276
rect 2021 242 2059 276
rect 2093 242 2105 276
rect 143 236 2105 242
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 clkinv_16
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 143 236 2105 282 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel metal1 s 147 384 2097 430 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4681606
string GDS_START 4664778
<< end >>
