magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2354 1975
<< nwell >>
rect -38 331 1094 704
<< pwell >>
rect 1 49 1047 241
rect 0 0 1056 49
<< scnmos >>
rect 84 47 114 215
rect 170 47 200 215
rect 256 47 286 215
rect 342 47 372 215
rect 428 47 458 215
rect 514 47 544 215
rect 600 47 630 215
rect 686 47 716 215
rect 856 47 886 215
rect 934 47 964 215
<< scpmoshvt >>
rect 84 367 114 619
rect 170 367 200 619
rect 256 367 286 619
rect 342 367 372 619
rect 442 367 472 619
rect 542 367 572 619
rect 642 367 672 619
rect 742 367 772 619
rect 856 367 886 619
rect 934 367 964 619
<< ndiff >>
rect 27 119 84 215
rect 27 85 39 119
rect 73 85 84 119
rect 27 47 84 85
rect 114 123 170 215
rect 114 89 125 123
rect 159 89 170 123
rect 114 47 170 89
rect 200 93 256 215
rect 200 59 211 93
rect 245 59 256 93
rect 200 47 256 59
rect 286 123 342 215
rect 286 89 297 123
rect 331 89 342 123
rect 286 47 342 89
rect 372 186 428 215
rect 372 152 383 186
rect 417 152 428 186
rect 372 47 428 152
rect 458 123 514 215
rect 458 89 469 123
rect 503 89 514 123
rect 458 47 514 89
rect 544 186 600 215
rect 544 152 555 186
rect 589 152 600 186
rect 544 47 600 152
rect 630 203 686 215
rect 630 169 641 203
rect 675 169 686 203
rect 630 101 686 169
rect 630 67 641 101
rect 675 67 686 101
rect 630 47 686 67
rect 716 105 856 215
rect 716 71 741 105
rect 775 71 856 105
rect 716 47 856 71
rect 886 47 934 215
rect 964 203 1021 215
rect 964 169 975 203
rect 1009 169 1021 203
rect 964 101 1021 169
rect 964 67 975 101
rect 1009 67 1021 101
rect 964 47 1021 67
<< pdiff >>
rect 27 607 84 619
rect 27 573 39 607
rect 73 573 84 607
rect 27 481 84 573
rect 27 447 39 481
rect 73 447 84 481
rect 27 367 84 447
rect 114 599 170 619
rect 114 565 125 599
rect 159 565 170 599
rect 114 481 170 565
rect 114 447 125 481
rect 159 447 170 481
rect 114 367 170 447
rect 200 578 256 619
rect 200 544 211 578
rect 245 544 256 578
rect 200 367 256 544
rect 286 599 342 619
rect 286 565 297 599
rect 331 565 342 599
rect 286 481 342 565
rect 286 447 297 481
rect 331 447 342 481
rect 286 367 342 447
rect 372 531 442 619
rect 372 497 397 531
rect 431 497 442 531
rect 372 413 442 497
rect 372 379 397 413
rect 431 379 442 413
rect 372 367 442 379
rect 472 599 542 619
rect 472 565 497 599
rect 531 565 542 599
rect 472 481 542 565
rect 472 447 497 481
rect 531 447 542 481
rect 472 367 542 447
rect 572 531 642 619
rect 572 497 597 531
rect 631 497 642 531
rect 572 413 642 497
rect 572 379 597 413
rect 631 379 642 413
rect 572 367 642 379
rect 672 599 742 619
rect 672 565 697 599
rect 731 565 742 599
rect 672 506 742 565
rect 672 472 697 506
rect 731 472 742 506
rect 672 413 742 472
rect 672 379 697 413
rect 731 379 742 413
rect 672 367 742 379
rect 772 607 856 619
rect 772 573 797 607
rect 831 573 856 607
rect 772 510 856 573
rect 772 476 797 510
rect 831 476 856 510
rect 772 413 856 476
rect 772 379 797 413
rect 831 379 856 413
rect 772 367 856 379
rect 886 367 934 619
rect 964 599 1021 619
rect 964 565 975 599
rect 1009 565 1021 599
rect 964 506 1021 565
rect 964 472 975 506
rect 1009 472 1021 506
rect 964 413 1021 472
rect 964 379 975 413
rect 1009 379 1021 413
rect 964 367 1021 379
<< ndiffc >>
rect 39 85 73 119
rect 125 89 159 123
rect 211 59 245 93
rect 297 89 331 123
rect 383 152 417 186
rect 469 89 503 123
rect 555 152 589 186
rect 641 169 675 203
rect 641 67 675 101
rect 741 71 775 105
rect 975 169 1009 203
rect 975 67 1009 101
<< pdiffc >>
rect 39 573 73 607
rect 39 447 73 481
rect 125 565 159 599
rect 125 447 159 481
rect 211 544 245 578
rect 297 565 331 599
rect 297 447 331 481
rect 397 497 431 531
rect 397 379 431 413
rect 497 565 531 599
rect 497 447 531 481
rect 597 497 631 531
rect 597 379 631 413
rect 697 565 731 599
rect 697 472 731 506
rect 697 379 731 413
rect 797 573 831 607
rect 797 476 831 510
rect 797 379 831 413
rect 975 565 1009 599
rect 975 472 1009 506
rect 975 379 1009 413
<< poly >>
rect 84 619 114 645
rect 170 619 200 645
rect 256 619 286 645
rect 342 619 372 645
rect 442 619 472 645
rect 542 619 572 645
rect 642 619 672 645
rect 742 619 772 645
rect 856 619 886 645
rect 934 619 964 645
rect 84 329 114 367
rect 170 329 200 367
rect 256 329 286 367
rect 342 329 372 367
rect 442 329 472 367
rect 542 329 572 367
rect 642 329 672 367
rect 742 329 772 367
rect 84 313 772 329
rect 84 279 165 313
rect 199 279 233 313
rect 267 279 301 313
rect 335 279 369 313
rect 403 279 437 313
rect 471 279 505 313
rect 539 279 573 313
rect 607 279 641 313
rect 675 279 709 313
rect 743 279 772 313
rect 856 303 886 367
rect 84 263 772 279
rect 820 287 886 303
rect 84 215 114 263
rect 170 215 200 263
rect 256 215 286 263
rect 342 215 372 263
rect 428 215 458 263
rect 514 215 544 263
rect 600 215 630 263
rect 686 215 716 263
rect 820 253 836 287
rect 870 267 886 287
rect 934 267 964 367
rect 870 253 964 267
rect 820 237 964 253
rect 856 215 886 237
rect 934 215 964 237
rect 84 21 114 47
rect 170 21 200 47
rect 256 21 286 47
rect 342 21 372 47
rect 428 21 458 47
rect 514 21 544 47
rect 600 21 630 47
rect 686 21 716 47
rect 856 21 886 47
rect 934 21 964 47
<< polycont >>
rect 165 279 199 313
rect 233 279 267 313
rect 301 279 335 313
rect 369 279 403 313
rect 437 279 471 313
rect 505 279 539 313
rect 573 279 607 313
rect 641 279 675 313
rect 709 279 743 313
rect 836 253 870 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 23 607 73 649
rect 23 573 39 607
rect 23 481 73 573
rect 23 447 39 481
rect 23 431 73 447
rect 109 599 175 615
rect 109 565 125 599
rect 159 565 175 599
rect 109 481 175 565
rect 211 578 245 649
rect 211 499 245 544
rect 281 599 747 615
rect 281 565 297 599
rect 331 581 497 599
rect 331 565 347 581
rect 109 447 125 481
rect 159 465 175 481
rect 281 481 347 565
rect 481 565 497 581
rect 531 581 697 599
rect 531 565 547 581
rect 281 465 297 481
rect 159 447 297 465
rect 331 447 347 481
rect 109 431 347 447
rect 381 531 447 547
rect 381 497 397 531
rect 431 497 447 531
rect 381 413 447 497
rect 481 481 547 565
rect 681 565 697 581
rect 731 565 747 599
rect 481 447 497 481
rect 531 447 547 481
rect 481 431 547 447
rect 581 531 647 547
rect 581 497 597 531
rect 631 497 647 531
rect 381 397 397 413
rect 37 379 397 397
rect 431 397 447 413
rect 581 413 647 497
rect 581 397 597 413
rect 431 379 597 397
rect 631 379 647 413
rect 37 363 647 379
rect 681 506 747 565
rect 681 472 697 506
rect 731 472 747 506
rect 681 413 747 472
rect 681 379 697 413
rect 731 379 747 413
rect 681 363 747 379
rect 781 607 847 649
rect 781 573 797 607
rect 831 573 847 607
rect 781 510 847 573
rect 781 476 797 510
rect 831 476 847 510
rect 781 413 847 476
rect 781 379 797 413
rect 831 379 847 413
rect 781 363 847 379
rect 959 599 1025 615
rect 959 565 975 599
rect 1009 565 1025 599
rect 959 506 1025 565
rect 959 472 975 506
rect 1009 472 1025 506
rect 959 413 1025 472
rect 959 379 975 413
rect 1009 379 1025 413
rect 37 356 71 363
rect 25 229 71 356
rect 149 313 759 329
rect 149 279 165 313
rect 199 279 233 313
rect 267 279 301 313
rect 335 279 369 313
rect 403 279 437 313
rect 471 279 505 313
rect 539 279 573 313
rect 607 279 641 313
rect 675 279 709 313
rect 743 279 759 313
rect 149 263 759 279
rect 25 195 589 229
rect 367 186 417 195
rect 23 119 73 161
rect 23 85 39 119
rect 23 17 73 85
rect 109 127 331 161
rect 109 123 159 127
rect 109 89 125 123
rect 297 123 331 127
rect 109 51 159 89
rect 195 59 211 93
rect 245 59 261 93
rect 195 17 261 59
rect 367 152 383 186
rect 555 186 589 195
rect 367 119 417 152
rect 453 123 519 161
rect 297 85 331 89
rect 453 89 469 123
rect 503 89 519 123
rect 555 119 589 152
rect 625 203 691 219
rect 625 169 641 203
rect 675 169 691 203
rect 453 85 519 89
rect 625 101 691 169
rect 725 202 759 263
rect 793 287 886 303
rect 793 253 836 287
rect 870 253 886 287
rect 793 236 886 253
rect 959 203 1025 379
rect 959 202 975 203
rect 725 169 975 202
rect 1009 169 1025 203
rect 725 168 1025 169
rect 625 85 641 101
rect 297 67 641 85
rect 675 67 691 101
rect 297 51 691 67
rect 725 105 791 134
rect 725 71 741 105
rect 775 71 791 105
rect 725 17 791 71
rect 959 101 1025 168
rect 959 67 975 101
rect 1009 67 1025 101
rect 959 51 1025 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 683 1056 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1056 683
rect 0 617 1056 649
rect 0 17 1056 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -49 1056 -17
<< labels >>
flabel pwell s 0 0 1056 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1056 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 buflp_4
flabel metal1 s 0 617 1056 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1056 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1056 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6981404
string GDS_START 6973716
<< end >>
