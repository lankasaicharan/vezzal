magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3230 1852
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 49 21 1929 203
rect 49 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 147 47 177 177
rect 241 47 271 177
rect 401 47 431 177
rect 495 47 525 177
rect 589 47 619 177
rect 683 47 713 177
rect 777 47 807 177
rect 871 47 901 177
rect 965 47 995 177
rect 1069 47 1099 177
rect 1153 47 1183 177
rect 1247 47 1277 177
rect 1341 47 1371 177
rect 1435 47 1465 177
rect 1529 47 1559 177
rect 1623 47 1653 177
rect 1717 47 1747 177
rect 1821 47 1851 177
<< scpmoshvt >>
rect 81 297 117 497
rect 185 297 221 497
rect 403 297 439 497
rect 497 297 533 497
rect 591 297 627 497
rect 685 297 721 497
rect 779 297 815 497
rect 873 297 909 497
rect 967 297 1003 497
rect 1061 297 1097 497
rect 1155 297 1191 497
rect 1249 297 1285 497
rect 1343 297 1379 497
rect 1437 297 1473 497
rect 1531 297 1567 497
rect 1625 297 1661 497
rect 1719 297 1755 497
rect 1813 297 1849 497
<< ndiff >>
rect 75 163 147 177
rect 75 129 97 163
rect 131 129 147 163
rect 75 95 147 129
rect 75 61 97 95
rect 131 61 147 95
rect 75 47 147 61
rect 177 163 241 177
rect 177 129 191 163
rect 225 129 241 163
rect 177 95 241 129
rect 177 61 191 95
rect 225 61 241 95
rect 177 47 241 61
rect 271 163 401 177
rect 271 61 289 163
rect 391 61 401 163
rect 271 47 401 61
rect 431 163 495 177
rect 431 129 451 163
rect 485 129 495 163
rect 431 95 495 129
rect 431 61 451 95
rect 485 61 495 95
rect 431 47 495 61
rect 525 95 589 177
rect 525 61 545 95
rect 579 61 589 95
rect 525 47 589 61
rect 619 163 683 177
rect 619 129 639 163
rect 673 129 683 163
rect 619 95 683 129
rect 619 61 639 95
rect 673 61 683 95
rect 619 47 683 61
rect 713 95 777 177
rect 713 61 733 95
rect 767 61 777 95
rect 713 47 777 61
rect 807 163 871 177
rect 807 129 827 163
rect 861 129 871 163
rect 807 95 871 129
rect 807 61 827 95
rect 861 61 871 95
rect 807 47 871 61
rect 901 95 965 177
rect 901 61 921 95
rect 955 61 965 95
rect 901 47 965 61
rect 995 163 1069 177
rect 995 129 1015 163
rect 1049 129 1069 163
rect 995 95 1069 129
rect 995 61 1015 95
rect 1049 61 1069 95
rect 995 47 1069 61
rect 1099 95 1153 177
rect 1099 61 1109 95
rect 1143 61 1153 95
rect 1099 47 1153 61
rect 1183 163 1247 177
rect 1183 129 1203 163
rect 1237 129 1247 163
rect 1183 95 1247 129
rect 1183 61 1203 95
rect 1237 61 1247 95
rect 1183 47 1247 61
rect 1277 95 1341 177
rect 1277 61 1297 95
rect 1331 61 1341 95
rect 1277 47 1341 61
rect 1371 163 1435 177
rect 1371 129 1391 163
rect 1425 129 1435 163
rect 1371 95 1435 129
rect 1371 61 1391 95
rect 1425 61 1435 95
rect 1371 47 1435 61
rect 1465 95 1529 177
rect 1465 61 1485 95
rect 1519 61 1529 95
rect 1465 47 1529 61
rect 1559 163 1623 177
rect 1559 129 1579 163
rect 1613 129 1623 163
rect 1559 95 1623 129
rect 1559 61 1579 95
rect 1613 61 1623 95
rect 1559 47 1623 61
rect 1653 95 1717 177
rect 1653 61 1673 95
rect 1707 61 1717 95
rect 1653 47 1717 61
rect 1747 163 1821 177
rect 1747 129 1767 163
rect 1801 129 1821 163
rect 1747 95 1821 129
rect 1747 61 1767 95
rect 1801 61 1821 95
rect 1747 47 1821 61
rect 1851 95 1903 177
rect 1851 61 1861 95
rect 1895 61 1903 95
rect 1851 47 1903 61
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 415 81 451
rect 27 381 35 415
rect 69 381 81 415
rect 27 345 81 381
rect 27 311 35 345
rect 69 311 81 345
rect 27 297 81 311
rect 117 477 185 497
rect 117 443 129 477
rect 163 443 185 477
rect 117 409 185 443
rect 117 375 129 409
rect 163 375 185 409
rect 117 341 185 375
rect 117 307 129 341
rect 163 307 185 341
rect 117 297 185 307
rect 221 485 287 497
rect 221 451 233 485
rect 267 451 287 485
rect 221 415 287 451
rect 221 381 233 415
rect 267 381 287 415
rect 221 345 287 381
rect 221 311 233 345
rect 267 311 287 345
rect 221 297 287 311
rect 345 477 403 497
rect 345 443 357 477
rect 391 443 403 477
rect 345 409 403 443
rect 345 375 357 409
rect 391 375 403 409
rect 345 341 403 375
rect 345 307 357 341
rect 391 307 403 341
rect 345 297 403 307
rect 439 485 497 497
rect 439 451 451 485
rect 485 451 497 485
rect 439 417 497 451
rect 439 383 451 417
rect 485 383 497 417
rect 439 297 497 383
rect 533 477 591 497
rect 533 443 545 477
rect 579 443 591 477
rect 533 409 591 443
rect 533 375 545 409
rect 579 375 591 409
rect 533 341 591 375
rect 533 307 545 341
rect 579 307 591 341
rect 533 297 591 307
rect 627 485 685 497
rect 627 451 639 485
rect 673 451 685 485
rect 627 417 685 451
rect 627 383 639 417
rect 673 383 685 417
rect 627 297 685 383
rect 721 477 779 497
rect 721 443 733 477
rect 767 443 779 477
rect 721 409 779 443
rect 721 375 733 409
rect 767 375 779 409
rect 721 341 779 375
rect 721 307 733 341
rect 767 307 779 341
rect 721 297 779 307
rect 815 485 873 497
rect 815 451 827 485
rect 861 451 873 485
rect 815 417 873 451
rect 815 383 827 417
rect 861 383 873 417
rect 815 297 873 383
rect 909 477 967 497
rect 909 443 921 477
rect 955 443 967 477
rect 909 409 967 443
rect 909 375 921 409
rect 955 375 967 409
rect 909 341 967 375
rect 909 307 921 341
rect 955 307 967 341
rect 909 297 967 307
rect 1003 485 1061 497
rect 1003 451 1015 485
rect 1049 451 1061 485
rect 1003 417 1061 451
rect 1003 383 1015 417
rect 1049 383 1061 417
rect 1003 297 1061 383
rect 1097 477 1155 497
rect 1097 443 1109 477
rect 1143 443 1155 477
rect 1097 409 1155 443
rect 1097 375 1109 409
rect 1143 375 1155 409
rect 1097 341 1155 375
rect 1097 307 1109 341
rect 1143 307 1155 341
rect 1097 297 1155 307
rect 1191 409 1249 497
rect 1191 375 1203 409
rect 1237 375 1249 409
rect 1191 341 1249 375
rect 1191 307 1203 341
rect 1237 307 1249 341
rect 1191 297 1249 307
rect 1285 477 1343 497
rect 1285 443 1297 477
rect 1331 443 1343 477
rect 1285 409 1343 443
rect 1285 375 1297 409
rect 1331 375 1343 409
rect 1285 297 1343 375
rect 1379 409 1437 497
rect 1379 375 1391 409
rect 1425 375 1437 409
rect 1379 341 1437 375
rect 1379 307 1391 341
rect 1425 307 1437 341
rect 1379 297 1437 307
rect 1473 477 1531 497
rect 1473 443 1485 477
rect 1519 443 1531 477
rect 1473 409 1531 443
rect 1473 375 1485 409
rect 1519 375 1531 409
rect 1473 297 1531 375
rect 1567 409 1625 497
rect 1567 375 1579 409
rect 1613 375 1625 409
rect 1567 341 1625 375
rect 1567 307 1579 341
rect 1613 307 1625 341
rect 1567 297 1625 307
rect 1661 477 1719 497
rect 1661 443 1673 477
rect 1707 443 1719 477
rect 1661 409 1719 443
rect 1661 375 1673 409
rect 1707 375 1719 409
rect 1661 297 1719 375
rect 1755 409 1813 497
rect 1755 375 1767 409
rect 1801 375 1813 409
rect 1755 341 1813 375
rect 1755 307 1767 341
rect 1801 307 1813 341
rect 1755 297 1813 307
rect 1849 477 1905 497
rect 1849 443 1861 477
rect 1895 443 1905 477
rect 1849 409 1905 443
rect 1849 375 1861 409
rect 1895 375 1905 409
rect 1849 297 1905 375
<< ndiffc >>
rect 97 129 131 163
rect 97 61 131 95
rect 191 129 225 163
rect 191 61 225 95
rect 289 61 391 163
rect 451 129 485 163
rect 451 61 485 95
rect 545 61 579 95
rect 639 129 673 163
rect 639 61 673 95
rect 733 61 767 95
rect 827 129 861 163
rect 827 61 861 95
rect 921 61 955 95
rect 1015 129 1049 163
rect 1015 61 1049 95
rect 1109 61 1143 95
rect 1203 129 1237 163
rect 1203 61 1237 95
rect 1297 61 1331 95
rect 1391 129 1425 163
rect 1391 61 1425 95
rect 1485 61 1519 95
rect 1579 129 1613 163
rect 1579 61 1613 95
rect 1673 61 1707 95
rect 1767 129 1801 163
rect 1767 61 1801 95
rect 1861 61 1895 95
<< pdiffc >>
rect 35 451 69 485
rect 35 381 69 415
rect 35 311 69 345
rect 129 443 163 477
rect 129 375 163 409
rect 129 307 163 341
rect 233 451 267 485
rect 233 381 267 415
rect 233 311 267 345
rect 357 443 391 477
rect 357 375 391 409
rect 357 307 391 341
rect 451 451 485 485
rect 451 383 485 417
rect 545 443 579 477
rect 545 375 579 409
rect 545 307 579 341
rect 639 451 673 485
rect 639 383 673 417
rect 733 443 767 477
rect 733 375 767 409
rect 733 307 767 341
rect 827 451 861 485
rect 827 383 861 417
rect 921 443 955 477
rect 921 375 955 409
rect 921 307 955 341
rect 1015 451 1049 485
rect 1015 383 1049 417
rect 1109 443 1143 477
rect 1109 375 1143 409
rect 1109 307 1143 341
rect 1203 375 1237 409
rect 1203 307 1237 341
rect 1297 443 1331 477
rect 1297 375 1331 409
rect 1391 375 1425 409
rect 1391 307 1425 341
rect 1485 443 1519 477
rect 1485 375 1519 409
rect 1579 375 1613 409
rect 1579 307 1613 341
rect 1673 443 1707 477
rect 1673 375 1707 409
rect 1767 375 1801 409
rect 1767 307 1801 341
rect 1861 443 1895 477
rect 1861 375 1895 409
<< poly >>
rect 81 497 117 523
rect 185 497 221 523
rect 403 497 439 523
rect 497 497 533 523
rect 591 497 627 523
rect 685 497 721 523
rect 779 497 815 523
rect 873 497 909 523
rect 967 497 1003 523
rect 1061 497 1097 523
rect 1155 497 1191 523
rect 1249 497 1285 523
rect 1343 497 1379 523
rect 1437 497 1473 523
rect 1531 497 1567 523
rect 1625 497 1661 523
rect 1719 497 1755 523
rect 1813 497 1849 523
rect 81 282 117 297
rect 185 282 221 297
rect 403 282 439 297
rect 497 282 533 297
rect 591 282 627 297
rect 685 282 721 297
rect 779 282 815 297
rect 873 282 909 297
rect 967 282 1003 297
rect 1061 282 1097 297
rect 1155 282 1191 297
rect 1249 282 1285 297
rect 1343 282 1379 297
rect 1437 282 1473 297
rect 1531 282 1567 297
rect 1625 282 1661 297
rect 1719 282 1755 297
rect 1813 282 1849 297
rect 79 265 119 282
rect 183 265 223 282
rect 401 265 441 282
rect 495 265 535 282
rect 589 265 629 282
rect 683 265 723 282
rect 777 265 817 282
rect 871 265 911 282
rect 965 265 1005 282
rect 1059 265 1099 282
rect 31 249 271 265
rect 31 215 41 249
rect 75 215 271 249
rect 31 199 271 215
rect 147 177 177 199
rect 241 177 271 199
rect 401 249 1099 265
rect 401 215 421 249
rect 455 215 499 249
rect 533 215 577 249
rect 611 215 655 249
rect 689 215 733 249
rect 767 215 801 249
rect 835 215 879 249
rect 913 215 957 249
rect 991 215 1035 249
rect 1069 215 1099 249
rect 401 199 1099 215
rect 401 177 431 199
rect 495 177 525 199
rect 589 177 619 199
rect 683 177 713 199
rect 777 177 807 199
rect 871 177 901 199
rect 965 177 995 199
rect 1069 177 1099 199
rect 1153 265 1193 282
rect 1247 265 1287 282
rect 1341 265 1381 282
rect 1435 265 1475 282
rect 1529 265 1569 282
rect 1623 265 1663 282
rect 1717 265 1757 282
rect 1811 265 1851 282
rect 1153 249 1851 265
rect 1153 215 1176 249
rect 1210 215 1254 249
rect 1288 215 1332 249
rect 1366 215 1410 249
rect 1444 215 1488 249
rect 1522 215 1556 249
rect 1590 215 1634 249
rect 1668 215 1712 249
rect 1746 215 1851 249
rect 1153 199 1851 215
rect 1153 177 1183 199
rect 1247 177 1277 199
rect 1341 177 1371 199
rect 1435 177 1465 199
rect 1529 177 1559 199
rect 1623 177 1653 199
rect 1717 177 1747 199
rect 1821 177 1851 199
rect 147 21 177 47
rect 241 21 271 47
rect 401 21 431 47
rect 495 21 525 47
rect 589 21 619 47
rect 683 21 713 47
rect 777 21 807 47
rect 871 21 901 47
rect 965 21 995 47
rect 1069 21 1099 47
rect 1153 21 1183 47
rect 1247 21 1277 47
rect 1341 21 1371 47
rect 1435 21 1465 47
rect 1529 21 1559 47
rect 1623 21 1653 47
rect 1717 21 1747 47
rect 1821 21 1851 47
<< polycont >>
rect 41 215 75 249
rect 421 215 455 249
rect 499 215 533 249
rect 577 215 611 249
rect 655 215 689 249
rect 733 215 767 249
rect 801 215 835 249
rect 879 215 913 249
rect 957 215 991 249
rect 1035 215 1069 249
rect 1176 215 1210 249
rect 1254 215 1288 249
rect 1332 215 1366 249
rect 1410 215 1444 249
rect 1488 215 1522 249
rect 1556 215 1590 249
rect 1634 215 1668 249
rect 1712 215 1746 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 25 485 69 527
rect 25 451 35 485
rect 25 415 69 451
rect 25 381 35 415
rect 25 345 69 381
rect 25 311 35 345
rect 25 291 69 311
rect 103 477 189 493
rect 103 443 129 477
rect 163 443 189 477
rect 103 409 189 443
rect 103 375 129 409
rect 163 375 189 409
rect 103 341 189 375
rect 103 307 129 341
rect 163 307 189 341
rect 103 291 189 307
rect 233 485 292 527
rect 267 451 292 485
rect 233 415 292 451
rect 267 381 292 415
rect 233 345 292 381
rect 267 311 292 345
rect 233 291 292 311
rect 335 477 399 493
rect 335 443 357 477
rect 391 443 399 477
rect 335 409 399 443
rect 335 375 357 409
rect 391 375 399 409
rect 335 341 399 375
rect 443 485 493 527
rect 443 451 451 485
rect 485 451 493 485
rect 443 417 493 451
rect 443 383 451 417
rect 485 383 493 417
rect 443 367 493 383
rect 537 477 587 493
rect 537 443 545 477
rect 579 443 587 477
rect 537 409 587 443
rect 537 375 545 409
rect 579 375 587 409
rect 335 307 357 341
rect 391 333 399 341
rect 537 341 587 375
rect 631 485 681 527
rect 631 451 639 485
rect 673 451 681 485
rect 631 417 681 451
rect 631 383 639 417
rect 673 383 681 417
rect 631 367 681 383
rect 725 477 775 493
rect 725 443 733 477
rect 767 443 775 477
rect 725 409 775 443
rect 725 375 733 409
rect 767 375 775 409
rect 537 333 545 341
rect 391 307 545 333
rect 579 333 587 341
rect 725 341 775 375
rect 819 485 869 527
rect 819 451 827 485
rect 861 451 869 485
rect 819 417 869 451
rect 819 383 827 417
rect 861 383 869 417
rect 819 367 869 383
rect 913 477 963 493
rect 913 443 921 477
rect 955 443 963 477
rect 913 409 963 443
rect 913 375 921 409
rect 955 375 963 409
rect 725 333 733 341
rect 579 307 733 333
rect 767 333 775 341
rect 913 341 963 375
rect 1007 485 1057 527
rect 1007 451 1015 485
rect 1049 451 1057 485
rect 1007 417 1057 451
rect 1007 383 1015 417
rect 1049 383 1057 417
rect 1007 367 1057 383
rect 1101 477 1903 493
rect 1101 443 1109 477
rect 1143 459 1297 477
rect 1143 443 1151 459
rect 1101 409 1151 443
rect 1289 443 1297 459
rect 1331 459 1485 477
rect 1331 443 1339 459
rect 1101 375 1109 409
rect 1143 375 1151 409
rect 913 333 921 341
rect 767 307 921 333
rect 955 333 963 341
rect 1101 341 1151 375
rect 1101 333 1109 341
rect 955 307 1109 333
rect 1143 307 1151 341
rect 335 291 1151 307
rect 1195 409 1245 425
rect 1195 375 1203 409
rect 1237 375 1245 409
rect 1195 341 1245 375
rect 1289 409 1339 443
rect 1477 443 1485 459
rect 1519 459 1673 477
rect 1519 443 1527 459
rect 1289 375 1297 409
rect 1331 375 1339 409
rect 1289 357 1339 375
rect 1383 409 1433 425
rect 1383 375 1391 409
rect 1425 375 1433 409
rect 1195 307 1203 341
rect 1237 323 1245 341
rect 1383 341 1433 375
rect 1477 409 1527 443
rect 1665 443 1673 459
rect 1707 459 1861 477
rect 1707 443 1715 459
rect 1477 375 1485 409
rect 1519 375 1527 409
rect 1477 357 1527 375
rect 1571 409 1621 425
rect 1571 375 1579 409
rect 1613 375 1621 409
rect 1383 323 1391 341
rect 1237 307 1391 323
rect 1425 323 1433 341
rect 1571 341 1621 375
rect 1665 409 1715 443
rect 1853 443 1861 459
rect 1895 443 1903 477
rect 1665 375 1673 409
rect 1707 375 1715 409
rect 1665 357 1715 375
rect 1759 409 1809 425
rect 1759 375 1767 409
rect 1801 375 1809 409
rect 1571 323 1579 341
rect 1425 307 1579 323
rect 1613 323 1621 341
rect 1759 341 1809 375
rect 1853 409 1903 443
rect 1853 375 1861 409
rect 1895 375 1903 409
rect 1853 357 1903 375
rect 1759 323 1767 341
rect 1613 307 1767 323
rect 1801 323 1809 341
rect 1801 307 1913 323
rect 145 257 189 291
rect 1195 289 1913 307
rect 17 249 101 257
rect 17 215 41 249
rect 75 215 101 249
rect 17 213 101 215
rect 145 249 1104 257
rect 145 215 421 249
rect 455 215 499 249
rect 533 215 577 249
rect 611 215 655 249
rect 689 215 733 249
rect 767 215 801 249
rect 835 215 879 249
rect 913 215 957 249
rect 991 215 1035 249
rect 1069 215 1104 249
rect 1158 249 1776 255
rect 1158 215 1176 249
rect 1210 215 1254 249
rect 1288 215 1332 249
rect 1366 215 1410 249
rect 1444 215 1488 249
rect 1522 215 1556 249
rect 1590 215 1634 249
rect 1668 215 1712 249
rect 1746 215 1776 249
rect 145 213 247 215
rect 17 51 63 213
rect 97 163 141 179
rect 131 129 141 163
rect 97 95 141 129
rect 131 61 141 95
rect 97 17 141 61
rect 175 163 247 213
rect 1810 181 1913 289
rect 175 129 191 163
rect 225 129 247 163
rect 175 95 247 129
rect 175 61 191 95
rect 225 61 247 95
rect 175 51 247 61
rect 289 163 391 181
rect 289 17 391 61
rect 425 163 1913 181
rect 425 129 451 163
rect 485 145 639 163
rect 485 129 501 145
rect 425 95 501 129
rect 613 129 639 145
rect 673 145 827 163
rect 673 129 689 145
rect 425 61 451 95
rect 485 61 501 95
rect 425 51 501 61
rect 545 95 579 111
rect 545 17 579 61
rect 613 95 689 129
rect 801 129 827 145
rect 861 145 1015 163
rect 861 129 877 145
rect 613 61 639 95
rect 673 61 689 95
rect 613 51 689 61
rect 733 95 767 111
rect 733 17 767 61
rect 801 95 877 129
rect 989 129 1015 145
rect 1049 145 1203 163
rect 1049 129 1065 145
rect 801 61 827 95
rect 861 61 877 95
rect 801 51 877 61
rect 921 95 955 111
rect 921 17 955 61
rect 989 95 1065 129
rect 1177 129 1203 145
rect 1237 145 1391 163
rect 1237 129 1253 145
rect 989 61 1015 95
rect 1049 61 1065 95
rect 989 51 1065 61
rect 1109 95 1143 111
rect 1109 17 1143 61
rect 1177 95 1253 129
rect 1365 129 1391 145
rect 1425 145 1579 163
rect 1425 129 1441 145
rect 1177 61 1203 95
rect 1237 61 1253 95
rect 1177 51 1253 61
rect 1297 95 1331 111
rect 1297 17 1331 61
rect 1365 95 1441 129
rect 1553 129 1579 145
rect 1613 145 1767 163
rect 1613 129 1629 145
rect 1365 61 1391 95
rect 1425 61 1441 95
rect 1365 51 1441 61
rect 1485 95 1519 111
rect 1485 17 1519 61
rect 1553 95 1629 129
rect 1741 129 1767 145
rect 1801 145 1913 163
rect 1801 129 1817 145
rect 1553 61 1579 95
rect 1613 61 1629 95
rect 1553 51 1629 61
rect 1673 95 1707 111
rect 1673 17 1707 61
rect 1741 95 1817 129
rect 1741 61 1767 95
rect 1801 61 1817 95
rect 1741 51 1817 61
rect 1861 95 1915 111
rect 1895 61 1915 95
rect 1861 17 1915 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 23 221 57 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 1854 289 1888 323 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel locali s 1158 215 1776 255 0 FreeSans 400 0 0 0 SLEEP
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sky130_fd_sc_hdll__lpflow_isobufsrc_8
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 112940
string GDS_START 98754
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
