magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3506 1975
<< nwell >>
rect -38 331 2246 704
<< pwell >>
rect 29 157 719 229
rect 934 217 1325 235
rect 934 173 1491 217
rect 1931 201 2205 273
rect 1738 173 2205 201
rect 934 157 2205 173
rect 29 49 2205 157
rect 0 0 2208 49
<< scnmos >>
rect 112 119 142 203
rect 226 119 256 203
rect 298 119 328 203
rect 434 119 464 203
rect 506 119 536 203
rect 610 119 640 203
rect 801 47 831 131
rect 1017 125 1047 209
rect 1119 125 1149 209
rect 1197 125 1227 209
rect 1382 63 1412 191
rect 1487 63 1517 147
rect 1640 63 1670 147
rect 1712 63 1742 147
rect 1817 47 1847 175
rect 2010 79 2040 247
rect 2096 79 2126 247
<< scpmoshvt >>
rect 124 487 154 615
rect 226 487 256 615
rect 298 487 328 615
rect 384 487 414 615
rect 478 487 508 615
rect 580 487 610 615
rect 824 469 854 597
rect 1020 451 1050 535
rect 1106 451 1136 535
rect 1178 451 1208 535
rect 1348 451 1378 619
rect 1488 451 1518 619
rect 1593 493 1623 577
rect 1665 493 1695 577
rect 1820 409 1850 577
rect 2010 367 2040 619
rect 2096 367 2126 619
<< ndiff >>
rect 55 178 112 203
rect 55 144 67 178
rect 101 144 112 178
rect 55 119 112 144
rect 142 178 226 203
rect 142 144 155 178
rect 189 144 226 178
rect 142 119 226 144
rect 256 119 298 203
rect 328 178 434 203
rect 328 144 387 178
rect 421 144 434 178
rect 328 119 434 144
rect 464 119 506 203
rect 536 178 610 203
rect 536 144 555 178
rect 589 144 610 178
rect 536 119 610 144
rect 640 190 693 203
rect 640 156 651 190
rect 685 156 693 190
rect 640 119 693 156
rect 960 175 1017 209
rect 960 141 968 175
rect 1002 141 1017 175
rect 747 99 801 131
rect 747 65 755 99
rect 789 65 801 99
rect 747 47 801 65
rect 831 106 899 131
rect 960 125 1017 141
rect 1047 184 1119 209
rect 1047 150 1058 184
rect 1092 150 1119 184
rect 1047 125 1119 150
rect 1149 125 1197 209
rect 1227 191 1299 209
rect 1227 125 1382 191
rect 831 72 842 106
rect 876 72 899 106
rect 831 47 899 72
rect 1249 109 1382 125
rect 1249 75 1259 109
rect 1293 75 1382 109
rect 1249 63 1382 75
rect 1412 169 1465 191
rect 1412 135 1423 169
rect 1457 147 1465 169
rect 1957 219 2010 247
rect 1957 185 1965 219
rect 1999 185 2010 219
rect 1764 161 1817 175
rect 1764 147 1772 161
rect 1457 135 1487 147
rect 1412 63 1487 135
rect 1517 117 1640 147
rect 1517 83 1595 117
rect 1629 83 1640 117
rect 1517 63 1640 83
rect 1670 63 1712 147
rect 1742 127 1772 147
rect 1806 127 1817 161
rect 1742 93 1817 127
rect 1742 63 1772 93
rect 1764 59 1772 63
rect 1806 59 1817 93
rect 1764 47 1817 59
rect 1847 163 1900 175
rect 1847 129 1858 163
rect 1892 129 1900 163
rect 1847 95 1900 129
rect 1847 61 1858 95
rect 1892 61 1900 95
rect 1957 125 2010 185
rect 1957 91 1965 125
rect 1999 91 2010 125
rect 1957 79 2010 91
rect 2040 235 2096 247
rect 2040 201 2051 235
rect 2085 201 2096 235
rect 2040 125 2096 201
rect 2040 91 2051 125
rect 2085 91 2096 125
rect 2040 79 2096 91
rect 2126 235 2179 247
rect 2126 201 2137 235
rect 2171 201 2179 235
rect 2126 125 2179 201
rect 2126 91 2137 125
rect 2171 91 2179 125
rect 2126 79 2179 91
rect 1847 47 1900 61
<< pdiff >>
rect 67 599 124 615
rect 67 565 79 599
rect 113 565 124 599
rect 67 529 124 565
rect 67 495 79 529
rect 113 495 124 529
rect 67 487 124 495
rect 154 571 226 615
rect 154 537 172 571
rect 206 537 226 571
rect 154 487 226 537
rect 256 487 298 615
rect 328 603 384 615
rect 328 569 339 603
rect 373 569 384 603
rect 328 533 384 569
rect 328 499 339 533
rect 373 499 384 533
rect 328 487 384 499
rect 414 487 478 615
rect 508 588 580 615
rect 508 554 531 588
rect 565 554 580 588
rect 508 487 580 554
rect 610 601 663 615
rect 610 567 621 601
rect 655 567 663 601
rect 1223 611 1348 619
rect 610 533 663 567
rect 610 499 621 533
rect 655 499 663 533
rect 610 487 663 499
rect 717 578 824 597
rect 717 544 727 578
rect 761 544 824 578
rect 717 469 824 544
rect 854 515 907 597
rect 1223 577 1235 611
rect 1269 577 1348 611
rect 1223 541 1348 577
rect 1223 535 1235 541
rect 854 481 865 515
rect 899 481 907 515
rect 854 469 907 481
rect 967 497 1020 535
rect 967 463 975 497
rect 1009 463 1020 497
rect 967 451 1020 463
rect 1050 510 1106 535
rect 1050 476 1061 510
rect 1095 476 1106 510
rect 1050 451 1106 476
rect 1136 451 1178 535
rect 1208 507 1235 535
rect 1269 507 1348 541
rect 1208 451 1348 507
rect 1378 499 1488 619
rect 1378 465 1389 499
rect 1423 465 1488 499
rect 1378 451 1488 465
rect 1518 599 1571 619
rect 1957 607 2010 619
rect 1518 565 1529 599
rect 1563 577 1571 599
rect 1563 565 1593 577
rect 1518 497 1593 565
rect 1518 463 1529 497
rect 1563 493 1593 497
rect 1623 493 1665 577
rect 1695 569 1820 577
rect 1695 552 1775 569
rect 1695 518 1706 552
rect 1740 535 1775 552
rect 1809 535 1820 569
rect 1740 518 1820 535
rect 1695 499 1820 518
rect 1695 493 1775 499
rect 1563 463 1571 493
rect 1518 451 1571 463
rect 1763 465 1775 493
rect 1809 465 1820 499
rect 1763 409 1820 465
rect 1850 565 1903 577
rect 1850 531 1861 565
rect 1895 531 1903 565
rect 1850 455 1903 531
rect 1850 421 1861 455
rect 1895 421 1903 455
rect 1850 409 1903 421
rect 1957 573 1965 607
rect 1999 573 2010 607
rect 1957 515 2010 573
rect 1957 481 1965 515
rect 1999 481 2010 515
rect 1957 419 2010 481
rect 1957 385 1965 419
rect 1999 385 2010 419
rect 1957 367 2010 385
rect 2040 599 2096 619
rect 2040 565 2051 599
rect 2085 565 2096 599
rect 2040 502 2096 565
rect 2040 468 2051 502
rect 2085 468 2096 502
rect 2040 413 2096 468
rect 2040 379 2051 413
rect 2085 379 2096 413
rect 2040 367 2096 379
rect 2126 607 2179 619
rect 2126 573 2137 607
rect 2171 573 2179 607
rect 2126 510 2179 573
rect 2126 476 2137 510
rect 2171 476 2179 510
rect 2126 413 2179 476
rect 2126 379 2137 413
rect 2171 379 2179 413
rect 2126 367 2179 379
<< ndiffc >>
rect 67 144 101 178
rect 155 144 189 178
rect 387 144 421 178
rect 555 144 589 178
rect 651 156 685 190
rect 968 141 1002 175
rect 755 65 789 99
rect 1058 150 1092 184
rect 842 72 876 106
rect 1259 75 1293 109
rect 1423 135 1457 169
rect 1965 185 1999 219
rect 1595 83 1629 117
rect 1772 127 1806 161
rect 1772 59 1806 93
rect 1858 129 1892 163
rect 1858 61 1892 95
rect 1965 91 1999 125
rect 2051 201 2085 235
rect 2051 91 2085 125
rect 2137 201 2171 235
rect 2137 91 2171 125
<< pdiffc >>
rect 79 565 113 599
rect 79 495 113 529
rect 172 537 206 571
rect 339 569 373 603
rect 339 499 373 533
rect 531 554 565 588
rect 621 567 655 601
rect 621 499 655 533
rect 727 544 761 578
rect 1235 577 1269 611
rect 865 481 899 515
rect 975 463 1009 497
rect 1061 476 1095 510
rect 1235 507 1269 541
rect 1389 465 1423 499
rect 1529 565 1563 599
rect 1529 463 1563 497
rect 1706 518 1740 552
rect 1775 535 1809 569
rect 1775 465 1809 499
rect 1861 531 1895 565
rect 1861 421 1895 455
rect 1965 573 1999 607
rect 1965 481 1999 515
rect 1965 385 1999 419
rect 2051 565 2085 599
rect 2051 468 2085 502
rect 2051 379 2085 413
rect 2137 573 2171 607
rect 2137 476 2171 510
rect 2137 379 2171 413
<< poly >>
rect 124 615 154 641
rect 226 615 256 641
rect 298 615 328 641
rect 384 615 414 641
rect 478 615 508 641
rect 580 615 610 641
rect 824 597 854 623
rect 1348 619 1378 645
rect 1488 619 1518 645
rect 2010 619 2040 645
rect 2096 619 2126 645
rect 124 465 154 487
rect 226 465 256 487
rect 106 435 256 465
rect 106 376 136 435
rect 184 377 250 393
rect 76 360 142 376
rect 76 326 92 360
rect 126 326 142 360
rect 184 343 200 377
rect 234 357 250 377
rect 234 343 256 357
rect 184 327 256 343
rect 76 292 142 326
rect 76 258 92 292
rect 126 258 142 292
rect 76 242 142 258
rect 112 203 142 242
rect 226 203 256 327
rect 298 291 328 487
rect 384 455 414 487
rect 370 439 436 455
rect 370 405 386 439
rect 420 405 436 439
rect 370 389 436 405
rect 478 341 508 487
rect 580 419 610 487
rect 1020 535 1050 561
rect 1106 535 1136 561
rect 1178 535 1208 561
rect 824 447 854 469
rect 1593 577 1623 603
rect 1665 577 1695 603
rect 1820 577 1850 603
rect 795 419 854 447
rect 1020 429 1050 451
rect 580 403 701 419
rect 580 389 651 403
rect 610 369 651 389
rect 685 369 701 403
rect 470 325 536 341
rect 470 291 486 325
rect 520 291 536 325
rect 298 275 364 291
rect 470 275 536 291
rect 298 241 314 275
rect 348 241 364 275
rect 298 225 364 241
rect 298 203 328 225
rect 434 203 464 229
rect 506 203 536 275
rect 610 335 701 369
rect 610 301 651 335
rect 685 301 701 335
rect 610 285 701 301
rect 765 417 854 419
rect 765 403 831 417
rect 765 369 781 403
rect 815 369 831 403
rect 909 399 1050 429
rect 909 369 939 399
rect 765 335 831 369
rect 765 301 781 335
rect 815 301 831 335
rect 765 285 831 301
rect 610 203 640 285
rect 801 131 831 285
rect 873 353 939 369
rect 873 319 889 353
rect 923 319 939 353
rect 1106 351 1136 451
rect 1178 429 1208 451
rect 1178 399 1271 429
rect 1197 387 1271 399
rect 1197 353 1221 387
rect 1255 353 1271 387
rect 873 285 939 319
rect 873 251 889 285
rect 923 251 939 285
rect 873 235 939 251
rect 1017 335 1149 351
rect 1017 301 1099 335
rect 1133 301 1149 335
rect 1017 285 1149 301
rect 1197 319 1271 353
rect 1197 285 1221 319
rect 1255 285 1271 319
rect 1017 209 1047 285
rect 1197 269 1271 285
rect 1348 279 1378 451
rect 1488 419 1518 451
rect 1460 403 1526 419
rect 1460 369 1476 403
rect 1510 369 1526 403
rect 1460 353 1526 369
rect 1593 307 1623 493
rect 1665 447 1695 493
rect 1665 431 1742 447
rect 1665 397 1681 431
rect 1715 397 1742 431
rect 1665 381 1742 397
rect 1119 209 1149 235
rect 1197 209 1227 269
rect 1321 263 1412 279
rect 1321 229 1337 263
rect 1371 229 1412 263
rect 1321 213 1412 229
rect 112 51 142 119
rect 226 93 256 119
rect 298 93 328 119
rect 434 51 464 119
rect 506 93 536 119
rect 610 93 640 119
rect 112 21 464 51
rect 1382 191 1412 213
rect 1487 277 1623 307
rect 1487 219 1559 277
rect 1017 99 1047 125
rect 1119 103 1149 125
rect 1089 87 1155 103
rect 1197 99 1227 125
rect 1089 53 1105 87
rect 1139 53 1155 87
rect 1487 185 1509 219
rect 1543 185 1559 219
rect 1487 169 1559 185
rect 1604 219 1670 235
rect 1604 185 1620 219
rect 1654 185 1670 219
rect 1604 169 1670 185
rect 1487 147 1517 169
rect 1640 147 1670 169
rect 1712 147 1742 381
rect 1820 361 1850 409
rect 1790 345 1856 361
rect 1790 311 1806 345
rect 1840 311 1856 345
rect 2010 335 2040 367
rect 2096 335 2126 367
rect 1790 277 1856 311
rect 1790 243 1806 277
rect 1840 243 1856 277
rect 1961 319 2126 335
rect 1961 285 1977 319
rect 2011 285 2126 319
rect 1961 269 2126 285
rect 2010 247 2040 269
rect 2096 247 2126 269
rect 1790 227 1856 243
rect 1817 175 1847 227
rect 801 21 831 47
rect 1089 37 1155 53
rect 1382 37 1412 63
rect 1487 37 1517 63
rect 1640 37 1670 63
rect 1712 37 1742 63
rect 2010 53 2040 79
rect 2096 53 2126 79
rect 1817 21 1847 47
<< polycont >>
rect 92 326 126 360
rect 200 343 234 377
rect 92 258 126 292
rect 386 405 420 439
rect 651 369 685 403
rect 486 291 520 325
rect 314 241 348 275
rect 651 301 685 335
rect 781 369 815 403
rect 781 301 815 335
rect 889 319 923 353
rect 1221 353 1255 387
rect 889 251 923 285
rect 1099 301 1133 335
rect 1221 285 1255 319
rect 1476 369 1510 403
rect 1681 397 1715 431
rect 1337 229 1371 263
rect 1105 53 1139 87
rect 1509 185 1543 219
rect 1620 185 1654 219
rect 1806 311 1840 345
rect 1806 243 1840 277
rect 1977 285 2011 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 63 599 122 615
rect 63 565 79 599
rect 113 565 122 599
rect 63 529 122 565
rect 63 495 79 529
rect 113 495 122 529
rect 156 571 222 649
rect 156 537 172 571
rect 206 537 222 571
rect 156 528 222 537
rect 323 603 389 615
rect 323 569 339 603
rect 373 569 389 603
rect 323 533 389 569
rect 525 588 569 649
rect 525 554 531 588
rect 565 554 569 588
rect 525 538 569 554
rect 605 601 671 605
rect 605 567 621 601
rect 655 567 671 601
rect 63 494 122 495
rect 323 499 339 533
rect 373 529 389 533
rect 605 533 671 567
rect 373 504 491 529
rect 373 499 545 504
rect 323 498 545 499
rect 22 460 234 494
rect 323 489 511 498
rect 22 194 56 460
rect 200 455 234 460
rect 457 464 511 489
rect 200 439 423 455
rect 90 360 166 426
rect 90 326 92 360
rect 126 326 166 360
rect 200 405 386 439
rect 420 405 423 439
rect 200 389 423 405
rect 457 424 545 464
rect 605 499 621 533
rect 655 499 671 533
rect 711 578 761 649
rect 1219 611 1275 649
rect 711 544 727 578
rect 711 528 761 544
rect 795 567 1169 601
rect 605 494 671 499
rect 795 494 829 567
rect 605 460 829 494
rect 457 390 615 424
rect 200 377 250 389
rect 234 343 250 377
rect 200 327 250 343
rect 90 292 166 326
rect 90 258 92 292
rect 126 258 166 292
rect 407 325 545 355
rect 407 291 486 325
rect 520 291 545 325
rect 90 228 166 258
rect 223 275 353 291
rect 223 241 314 275
rect 348 241 353 275
rect 581 257 615 390
rect 22 178 111 194
rect 22 144 67 178
rect 101 144 111 178
rect 22 128 111 144
rect 145 178 189 194
rect 145 144 155 178
rect 145 17 189 144
rect 223 77 353 241
rect 387 223 615 257
rect 651 403 747 424
rect 685 369 747 403
rect 651 335 747 369
rect 685 301 747 335
rect 651 240 747 301
rect 781 403 829 460
rect 815 369 829 403
rect 781 335 829 369
rect 815 301 829 335
rect 387 178 427 223
rect 781 206 829 301
rect 645 190 829 206
rect 421 144 427 178
rect 387 127 427 144
rect 539 178 605 189
rect 539 144 555 178
rect 589 144 605 178
rect 539 17 605 144
rect 645 156 651 190
rect 685 172 829 190
rect 863 515 925 533
rect 863 481 865 515
rect 899 481 925 515
rect 863 353 925 481
rect 863 319 889 353
rect 923 319 925 353
rect 863 285 925 319
rect 863 251 889 285
rect 923 251 925 285
rect 863 235 925 251
rect 959 498 1027 518
rect 959 497 991 498
rect 959 463 975 497
rect 1025 464 1027 498
rect 1009 463 1027 464
rect 959 455 1027 463
rect 1061 510 1099 526
rect 1095 476 1099 510
rect 685 156 781 172
rect 645 140 781 156
rect 863 122 907 235
rect 959 191 993 455
rect 1061 421 1099 476
rect 1029 387 1099 421
rect 1135 457 1169 567
rect 1219 577 1235 611
rect 1269 577 1275 611
rect 1527 599 1597 615
rect 1219 541 1275 577
rect 1219 507 1235 541
rect 1269 507 1275 541
rect 1219 491 1275 507
rect 1309 549 1493 583
rect 1309 457 1343 549
rect 1135 423 1343 457
rect 1377 499 1425 515
rect 1377 465 1389 499
rect 1423 465 1425 499
rect 1029 249 1063 387
rect 1135 351 1169 423
rect 1377 389 1425 465
rect 1097 335 1169 351
rect 1097 301 1099 335
rect 1133 301 1169 335
rect 1097 285 1169 301
rect 1205 387 1425 389
rect 1205 353 1221 387
rect 1255 353 1425 387
rect 1459 413 1493 549
rect 1527 565 1529 599
rect 1563 565 1597 599
rect 1527 497 1597 565
rect 1527 463 1529 497
rect 1563 463 1597 497
rect 1690 569 1825 649
rect 1949 607 2011 649
rect 1690 552 1775 569
rect 1690 518 1706 552
rect 1740 535 1775 552
rect 1809 535 1825 569
rect 1740 518 1825 535
rect 1690 499 1825 518
rect 1690 465 1775 499
rect 1809 465 1825 499
rect 1859 565 1910 581
rect 1859 531 1861 565
rect 1895 531 1910 565
rect 1527 447 1597 463
rect 1459 403 1527 413
rect 1459 369 1476 403
rect 1510 369 1527 403
rect 1459 367 1527 369
rect 1205 333 1425 353
rect 1205 319 1459 333
rect 1205 285 1221 319
rect 1255 299 1459 319
rect 1255 285 1271 299
rect 1321 263 1387 265
rect 1321 249 1337 263
rect 1029 229 1337 249
rect 1371 229 1387 263
rect 1029 215 1387 229
rect 952 181 993 191
rect 1054 184 1098 215
rect 952 175 1018 181
rect 952 141 968 175
rect 1002 141 1018 175
rect 952 131 1018 141
rect 1054 150 1058 184
rect 1092 150 1098 184
rect 1054 134 1098 150
rect 1132 145 1387 179
rect 839 106 907 122
rect 739 99 805 106
rect 739 65 755 99
rect 789 65 805 99
rect 739 17 805 65
rect 839 72 842 106
rect 876 97 907 106
rect 1132 97 1193 145
rect 876 87 1193 97
rect 876 72 1105 87
rect 839 53 1105 72
rect 1139 53 1193 87
rect 1241 109 1309 111
rect 1241 75 1259 109
rect 1293 75 1309 109
rect 1241 17 1309 75
rect 1343 85 1387 145
rect 1421 169 1459 299
rect 1493 289 1527 367
rect 1563 361 1597 447
rect 1859 455 1910 531
rect 1859 431 1861 455
rect 1665 397 1681 431
rect 1715 421 1861 431
rect 1895 421 1910 455
rect 1715 397 1910 421
rect 1665 395 1910 397
rect 1563 345 1842 361
rect 1563 327 1806 345
rect 1698 311 1806 327
rect 1840 311 1842 345
rect 1493 255 1664 289
rect 1604 219 1664 255
rect 1421 135 1423 169
rect 1457 135 1459 169
rect 1421 119 1459 135
rect 1493 185 1509 219
rect 1543 185 1559 219
rect 1493 85 1559 185
rect 1604 185 1620 219
rect 1654 185 1664 219
rect 1604 169 1664 185
rect 1698 277 1842 311
rect 1698 243 1806 277
rect 1840 243 1842 277
rect 1698 227 1842 243
rect 1876 335 1910 395
rect 1949 573 1965 607
rect 1999 573 2011 607
rect 1949 515 2011 573
rect 1949 481 1965 515
rect 1999 481 2011 515
rect 1949 419 2011 481
rect 1949 385 1965 419
rect 1999 385 2011 419
rect 1949 369 2011 385
rect 2045 599 2093 615
rect 2045 565 2051 599
rect 2085 565 2093 599
rect 2045 502 2093 565
rect 2045 468 2051 502
rect 2085 468 2093 502
rect 2045 413 2093 468
rect 2045 379 2051 413
rect 2085 379 2093 413
rect 1876 319 2011 335
rect 1876 285 1977 319
rect 1876 269 2011 285
rect 1698 133 1732 227
rect 1876 179 1910 269
rect 2045 235 2093 379
rect 2127 607 2187 649
rect 2127 573 2137 607
rect 2171 573 2187 607
rect 2127 510 2187 573
rect 2127 476 2137 510
rect 2171 476 2187 510
rect 2127 413 2187 476
rect 2127 379 2137 413
rect 2171 379 2187 413
rect 2127 363 2187 379
rect 1343 51 1559 85
rect 1595 117 1732 133
rect 1629 83 1732 117
rect 1595 67 1732 83
rect 1766 161 1808 177
rect 1766 127 1772 161
rect 1806 127 1808 161
rect 1766 93 1808 127
rect 1766 59 1772 93
rect 1806 59 1808 93
rect 1766 17 1808 59
rect 1842 163 1910 179
rect 1842 129 1858 163
rect 1892 129 1910 163
rect 1842 95 1910 129
rect 1842 61 1858 95
rect 1892 61 1910 95
rect 1842 51 1910 61
rect 1949 219 2011 235
rect 1949 185 1965 219
rect 1999 185 2011 219
rect 1949 125 2011 185
rect 1949 91 1965 125
rect 1999 91 2011 125
rect 1949 17 2011 91
rect 2045 201 2051 235
rect 2085 201 2093 235
rect 2045 125 2093 201
rect 2045 91 2051 125
rect 2085 91 2093 125
rect 2045 75 2093 91
rect 2127 235 2187 251
rect 2127 201 2137 235
rect 2171 201 2187 235
rect 2127 125 2187 201
rect 2127 91 2137 125
rect 2171 91 2187 125
rect 2127 17 2187 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 511 464 545 498
rect 991 497 1025 498
rect 991 464 1009 497
rect 1009 464 1025 497
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
<< metal1 >>
rect 0 683 2208 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2208 683
rect 0 617 2208 649
rect 499 498 557 504
rect 499 464 511 498
rect 545 495 557 498
rect 979 498 1037 504
rect 979 495 991 498
rect 545 467 991 495
rect 545 464 557 467
rect 499 458 557 464
rect 979 464 991 467
rect 1025 464 1037 498
rect 979 458 1037 464
rect 0 17 2208 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2208 17
rect 0 -49 2208 -17
<< labels >>
flabel pwell s 0 0 2208 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2208 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfxtp_2
flabel metal1 s 0 617 2208 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2208 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2047 94 2081 128 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 168 2081 202 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 242 2081 276 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 390 2081 424 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 464 2081 498 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2047 538 2081 572 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2208 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4073122
string GDS_START 4054910
<< end >>
