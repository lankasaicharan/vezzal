magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4370 1975
<< nwell >>
rect -38 331 3110 704
<< pwell >>
rect 1827 235 2133 279
rect 2660 235 3040 241
rect 63 157 635 231
rect 1054 165 1184 191
rect 1491 165 3040 235
rect 1054 157 3040 165
rect 63 49 3040 157
rect 0 0 3072 49
<< scnmos >>
rect 142 121 172 205
rect 214 121 244 205
rect 300 121 330 205
rect 372 121 402 205
rect 526 121 556 205
rect 847 47 877 131
rect 933 47 963 131
rect 1207 55 1237 139
rect 1293 55 1323 139
rect 1365 55 1395 139
rect 1578 125 1608 209
rect 1650 125 1680 209
rect 1903 125 1933 253
rect 1975 125 2005 253
rect 2129 125 2159 209
rect 2214 125 2244 209
rect 2352 125 2382 209
rect 2460 125 2490 209
rect 2739 131 2769 215
rect 2841 47 2871 215
rect 2927 47 2957 215
<< scpmoshvt >>
rect 92 481 122 609
rect 178 481 208 609
rect 250 481 280 609
rect 358 481 388 609
rect 666 462 696 590
rect 875 483 905 611
rect 961 483 991 611
rect 1211 415 1241 499
rect 1297 415 1327 499
rect 1369 415 1399 499
rect 1525 415 1555 499
rect 1630 379 1660 463
rect 1751 379 1781 547
rect 1968 463 1998 547
rect 2077 379 2107 547
rect 2273 435 2303 519
rect 2359 435 2389 519
rect 2549 483 2579 567
rect 2739 367 2769 495
rect 2841 367 2871 619
rect 2927 367 2957 619
<< ndiff >>
rect 89 180 142 205
rect 89 146 97 180
rect 131 146 142 180
rect 89 121 142 146
rect 172 121 214 205
rect 244 180 300 205
rect 244 146 255 180
rect 289 146 300 180
rect 244 121 300 146
rect 330 121 372 205
rect 402 180 526 205
rect 402 146 413 180
rect 447 146 481 180
rect 515 146 526 180
rect 402 121 526 146
rect 556 180 609 205
rect 556 146 567 180
rect 601 146 609 180
rect 556 121 609 146
rect 1080 157 1158 165
rect 794 106 847 131
rect 794 72 802 106
rect 836 72 847 106
rect 794 47 847 72
rect 877 106 933 131
rect 877 72 888 106
rect 922 72 933 106
rect 877 47 933 72
rect 963 106 1016 131
rect 963 72 974 106
rect 1008 72 1016 106
rect 963 47 1016 72
rect 1080 123 1092 157
rect 1126 139 1158 157
rect 1853 209 1903 253
rect 1517 195 1578 209
rect 1517 161 1525 195
rect 1559 161 1578 195
rect 1126 123 1207 139
rect 1080 55 1207 123
rect 1237 115 1293 139
rect 1237 81 1248 115
rect 1282 81 1293 115
rect 1237 55 1293 81
rect 1323 55 1365 139
rect 1395 106 1448 139
rect 1517 125 1578 161
rect 1608 125 1650 209
rect 1680 198 1903 209
rect 1680 164 1691 198
rect 1725 164 1777 198
rect 1811 164 1858 198
rect 1892 164 1903 198
rect 1680 125 1903 164
rect 1933 125 1975 253
rect 2005 245 2107 253
rect 2005 211 2019 245
rect 2053 211 2107 245
rect 2005 209 2107 211
rect 2005 177 2129 209
rect 2005 143 2084 177
rect 2118 143 2129 177
rect 2005 125 2129 143
rect 2159 125 2214 209
rect 2244 125 2352 209
rect 2382 183 2460 209
rect 2382 149 2393 183
rect 2427 149 2460 183
rect 2382 125 2460 149
rect 2490 183 2543 209
rect 2490 149 2501 183
rect 2535 149 2543 183
rect 2490 125 2543 149
rect 2686 190 2739 215
rect 2686 156 2694 190
rect 2728 156 2739 190
rect 2686 131 2739 156
rect 2769 203 2841 215
rect 2769 169 2784 203
rect 2818 169 2841 203
rect 2769 131 2841 169
rect 1395 72 1406 106
rect 1440 72 1448 106
rect 1395 55 1448 72
rect 2788 99 2841 131
rect 2788 65 2796 99
rect 2830 65 2841 99
rect 2788 47 2841 65
rect 2871 203 2927 215
rect 2871 169 2882 203
rect 2916 169 2927 203
rect 2871 101 2927 169
rect 2871 67 2882 101
rect 2916 67 2927 101
rect 2871 47 2927 67
rect 2957 159 3014 215
rect 2957 125 2968 159
rect 3002 125 3014 159
rect 2957 89 3014 125
rect 2957 55 2968 89
rect 3002 55 3014 89
rect 2957 47 3014 55
<< pdiff >>
rect 39 597 92 609
rect 39 563 47 597
rect 81 563 92 597
rect 39 529 92 563
rect 39 495 47 529
rect 81 495 92 529
rect 39 481 92 495
rect 122 601 178 609
rect 122 567 133 601
rect 167 567 178 601
rect 122 481 178 567
rect 208 481 250 609
rect 280 601 358 609
rect 280 567 302 601
rect 336 567 358 601
rect 280 481 358 567
rect 388 527 441 609
rect 388 493 399 527
rect 433 493 441 527
rect 388 481 441 493
rect 559 578 666 590
rect 559 544 569 578
rect 603 544 666 578
rect 559 510 666 544
rect 559 476 569 510
rect 603 476 666 510
rect 559 462 666 476
rect 696 510 749 590
rect 696 476 707 510
rect 741 476 749 510
rect 696 462 749 476
rect 803 483 875 611
rect 905 603 961 611
rect 905 569 916 603
rect 950 569 961 603
rect 905 483 961 569
rect 991 591 1044 611
rect 991 557 1002 591
rect 1036 557 1044 591
rect 991 483 1044 557
rect 803 463 853 483
rect 803 429 811 463
rect 845 429 853 463
rect 803 417 853 429
rect 1888 561 1946 569
rect 1698 535 1751 547
rect 1698 501 1706 535
rect 1740 501 1751 535
rect 1104 487 1211 499
rect 1104 453 1112 487
rect 1146 453 1211 487
rect 1104 415 1211 453
rect 1241 461 1297 499
rect 1241 427 1252 461
rect 1286 427 1297 461
rect 1241 415 1297 427
rect 1327 415 1369 499
rect 1399 491 1525 499
rect 1399 457 1412 491
rect 1446 457 1525 491
rect 1399 415 1525 457
rect 1555 463 1608 499
rect 1698 465 1751 501
rect 1698 463 1706 465
rect 1555 461 1630 463
rect 1555 427 1566 461
rect 1600 427 1630 461
rect 1555 415 1630 427
rect 1580 379 1630 415
rect 1660 431 1706 463
rect 1740 431 1751 465
rect 1660 379 1751 431
rect 1781 535 1834 547
rect 1781 501 1792 535
rect 1826 501 1834 535
rect 1781 465 1834 501
rect 1781 431 1792 465
rect 1826 431 1834 465
rect 1888 527 1900 561
rect 1934 547 1946 561
rect 1934 527 1968 547
rect 1888 463 1968 527
rect 1998 463 2077 547
rect 1781 379 1834 431
rect 2020 421 2077 463
rect 2020 387 2032 421
rect 2066 387 2077 421
rect 2020 379 2077 387
rect 2107 507 2160 547
rect 2107 473 2118 507
rect 2152 473 2160 507
rect 2107 390 2160 473
rect 2107 379 2157 390
rect 2788 607 2841 619
rect 2788 573 2796 607
rect 2830 573 2841 607
rect 2496 542 2549 567
rect 2220 505 2273 519
rect 2220 471 2228 505
rect 2262 471 2273 505
rect 2220 435 2273 471
rect 2303 505 2359 519
rect 2303 471 2314 505
rect 2348 471 2359 505
rect 2303 435 2359 471
rect 2389 494 2442 519
rect 2389 460 2400 494
rect 2434 460 2442 494
rect 2496 508 2504 542
rect 2538 508 2549 542
rect 2496 483 2549 508
rect 2579 542 2632 567
rect 2579 508 2590 542
rect 2624 508 2632 542
rect 2579 483 2632 508
rect 2788 510 2841 573
rect 2788 495 2796 510
rect 2389 435 2442 460
rect 2686 481 2739 495
rect 2686 447 2694 481
rect 2728 447 2739 481
rect 2686 413 2739 447
rect 2686 379 2694 413
rect 2728 379 2739 413
rect 2686 367 2739 379
rect 2769 476 2796 495
rect 2830 476 2841 510
rect 2769 415 2841 476
rect 2769 381 2780 415
rect 2814 381 2841 415
rect 2769 367 2841 381
rect 2871 599 2927 619
rect 2871 565 2882 599
rect 2916 565 2927 599
rect 2871 509 2927 565
rect 2871 475 2882 509
rect 2916 475 2927 509
rect 2871 415 2927 475
rect 2871 381 2882 415
rect 2916 381 2927 415
rect 2871 367 2927 381
rect 2957 607 3010 619
rect 2957 573 2968 607
rect 3002 573 3010 607
rect 2957 539 3010 573
rect 2957 505 2968 539
rect 3002 505 3010 539
rect 2957 467 3010 505
rect 2957 433 2968 467
rect 3002 433 3010 467
rect 2957 367 3010 433
<< ndiffc >>
rect 97 146 131 180
rect 255 146 289 180
rect 413 146 447 180
rect 481 146 515 180
rect 567 146 601 180
rect 802 72 836 106
rect 888 72 922 106
rect 974 72 1008 106
rect 1092 123 1126 157
rect 1525 161 1559 195
rect 1248 81 1282 115
rect 1691 164 1725 198
rect 1777 164 1811 198
rect 1858 164 1892 198
rect 2019 211 2053 245
rect 2084 143 2118 177
rect 2393 149 2427 183
rect 2501 149 2535 183
rect 2694 156 2728 190
rect 2784 169 2818 203
rect 1406 72 1440 106
rect 2796 65 2830 99
rect 2882 169 2916 203
rect 2882 67 2916 101
rect 2968 125 3002 159
rect 2968 55 3002 89
<< pdiffc >>
rect 47 563 81 597
rect 47 495 81 529
rect 133 567 167 601
rect 302 567 336 601
rect 399 493 433 527
rect 569 544 603 578
rect 569 476 603 510
rect 707 476 741 510
rect 916 569 950 603
rect 1002 557 1036 591
rect 811 429 845 463
rect 1706 501 1740 535
rect 1112 453 1146 487
rect 1252 427 1286 461
rect 1412 457 1446 491
rect 1566 427 1600 461
rect 1706 431 1740 465
rect 1792 501 1826 535
rect 1792 431 1826 465
rect 1900 527 1934 561
rect 2032 387 2066 421
rect 2118 473 2152 507
rect 2796 573 2830 607
rect 2228 471 2262 505
rect 2314 471 2348 505
rect 2400 460 2434 494
rect 2504 508 2538 542
rect 2590 508 2624 542
rect 2694 447 2728 481
rect 2694 379 2728 413
rect 2796 476 2830 510
rect 2780 381 2814 415
rect 2882 565 2916 599
rect 2882 475 2916 509
rect 2882 381 2916 415
rect 2968 573 3002 607
rect 2968 505 3002 539
rect 2968 433 3002 467
<< poly >>
rect 92 609 122 635
rect 178 609 208 635
rect 250 609 280 635
rect 358 609 388 635
rect 666 590 696 616
rect 875 611 905 637
rect 961 611 991 637
rect 1059 615 2205 645
rect 2841 619 2871 645
rect 2927 619 2957 645
rect 92 361 122 481
rect 44 345 122 361
rect 44 311 60 345
rect 94 311 122 345
rect 178 335 208 481
rect 250 449 280 481
rect 358 459 388 481
rect 250 433 316 449
rect 250 399 266 433
rect 300 399 316 433
rect 358 429 402 459
rect 250 383 316 399
rect 286 381 316 383
rect 286 351 330 381
rect 44 277 122 311
rect 172 305 244 335
rect 44 243 60 277
rect 94 257 122 277
rect 94 243 172 257
rect 44 227 172 243
rect 142 205 172 227
rect 214 205 244 305
rect 300 205 330 351
rect 372 326 402 429
rect 666 440 696 462
rect 666 410 753 440
rect 592 346 658 362
rect 592 326 608 346
rect 372 312 608 326
rect 642 312 658 346
rect 372 296 658 312
rect 372 205 402 296
rect 526 205 556 231
rect 723 187 753 410
rect 875 365 905 483
rect 961 451 991 483
rect 1059 451 1089 615
rect 1211 499 1241 525
rect 1297 499 1327 615
rect 1751 547 1781 573
rect 1369 499 1399 525
rect 1525 499 1555 525
rect 961 435 1089 451
rect 961 401 977 435
rect 1011 401 1089 435
rect 1630 463 1660 489
rect 961 367 1089 401
rect 687 171 753 187
rect 687 137 703 171
rect 737 137 753 171
rect 142 95 172 121
rect 214 53 244 121
rect 300 95 330 121
rect 372 95 402 121
rect 526 53 556 121
rect 687 103 753 137
rect 847 349 913 365
rect 847 315 863 349
rect 897 315 913 349
rect 847 281 913 315
rect 847 247 863 281
rect 897 247 913 281
rect 847 231 913 247
rect 961 333 977 367
rect 1011 333 1089 367
rect 1211 341 1241 415
rect 1297 389 1327 415
rect 1369 367 1399 415
rect 1369 351 1435 367
rect 961 299 1089 333
rect 961 265 977 299
rect 1011 265 1089 299
rect 1166 325 1315 341
rect 1166 291 1182 325
rect 1216 291 1315 325
rect 1166 275 1315 291
rect 847 131 877 231
rect 961 227 1089 265
rect 1285 253 1315 275
rect 1369 317 1385 351
rect 1419 317 1435 351
rect 1369 301 1435 317
rect 961 197 1237 227
rect 1285 223 1323 253
rect 1369 227 1399 301
rect 1525 297 1555 415
rect 1968 547 1998 573
rect 2077 547 2107 573
rect 1968 419 1998 463
rect 1922 403 2005 419
rect 1630 339 1660 379
rect 1630 309 1680 339
rect 1516 281 1582 297
rect 1516 247 1532 281
rect 1566 261 1582 281
rect 1566 247 1608 261
rect 1516 231 1608 247
rect 961 183 991 197
rect 933 153 991 183
rect 933 131 963 153
rect 687 69 703 103
rect 737 69 753 103
rect 687 53 753 69
rect 214 23 753 53
rect 1207 139 1237 197
rect 1293 139 1323 223
rect 1365 211 1431 227
rect 1365 177 1381 211
rect 1415 177 1431 211
rect 1578 209 1608 231
rect 1650 209 1680 309
rect 1751 305 1781 379
rect 1922 369 1938 403
rect 1972 369 2005 403
rect 1922 353 2005 369
rect 1751 281 1933 305
rect 1751 247 1767 281
rect 1801 275 1933 281
rect 1801 247 1817 275
rect 1903 253 1933 275
rect 1975 253 2005 353
rect 2077 357 2107 379
rect 2175 375 2205 615
rect 2549 567 2579 593
rect 2273 519 2303 545
rect 2359 519 2389 545
rect 2739 495 2769 521
rect 2549 451 2579 483
rect 2500 435 2579 451
rect 2172 357 2205 375
rect 2077 345 2205 357
rect 2077 327 2202 345
rect 1751 231 1817 247
rect 1365 161 1431 177
rect 1365 139 1395 161
rect 2129 209 2159 327
rect 2273 297 2303 435
rect 2359 367 2389 435
rect 2500 401 2516 435
rect 2550 401 2579 435
rect 2500 367 2579 401
rect 2352 351 2418 367
rect 2352 317 2368 351
rect 2402 317 2418 351
rect 2500 345 2516 367
rect 2352 301 2418 317
rect 2460 333 2516 345
rect 2550 345 2579 367
rect 2739 345 2769 367
rect 2550 333 2769 345
rect 2460 315 2769 333
rect 2841 329 2871 367
rect 2244 281 2310 297
rect 2244 261 2260 281
rect 2214 247 2260 261
rect 2294 247 2310 281
rect 2214 231 2310 247
rect 2352 267 2388 301
rect 2214 209 2244 231
rect 2352 209 2382 267
rect 2460 209 2490 315
rect 2739 215 2769 315
rect 2817 313 2883 329
rect 2817 279 2833 313
rect 2867 293 2883 313
rect 2927 293 2957 367
rect 2867 279 2957 293
rect 2817 263 2957 279
rect 2841 215 2871 263
rect 2927 215 2957 263
rect 1578 99 1608 125
rect 1650 103 1680 125
rect 1650 87 1729 103
rect 1903 99 1933 125
rect 1975 99 2005 125
rect 2129 99 2159 125
rect 2214 99 2244 125
rect 2352 99 2382 125
rect 2460 99 2490 125
rect 2739 105 2769 131
rect 847 21 877 47
rect 933 21 963 47
rect 1207 29 1237 55
rect 1293 29 1323 55
rect 1365 29 1395 55
rect 1650 53 1679 87
rect 1713 53 1729 87
rect 1650 37 1729 53
rect 2841 21 2871 47
rect 2927 21 2957 47
<< polycont >>
rect 60 311 94 345
rect 266 399 300 433
rect 60 243 94 277
rect 608 312 642 346
rect 977 401 1011 435
rect 703 137 737 171
rect 863 315 897 349
rect 863 247 897 281
rect 977 333 1011 367
rect 977 265 1011 299
rect 1182 291 1216 325
rect 1385 317 1419 351
rect 1532 247 1566 281
rect 703 69 737 103
rect 1381 177 1415 211
rect 1938 369 1972 403
rect 1767 247 1801 281
rect 2516 401 2550 435
rect 2368 317 2402 351
rect 2516 333 2550 367
rect 2260 247 2294 281
rect 2833 279 2867 313
rect 1679 53 1713 87
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 31 597 83 613
rect 31 563 47 597
rect 81 563 83 597
rect 117 601 183 649
rect 117 567 133 601
rect 167 567 183 601
rect 117 563 183 567
rect 286 601 519 615
rect 286 567 302 601
rect 336 567 519 601
rect 286 563 519 567
rect 31 529 83 563
rect 31 495 47 529
rect 81 527 449 529
rect 81 495 399 527
rect 31 493 399 495
rect 433 493 449 527
rect 31 479 449 493
rect 17 433 451 445
rect 17 399 266 433
rect 300 399 451 433
rect 17 390 451 399
rect 485 424 519 563
rect 553 578 605 649
rect 900 603 966 649
rect 553 544 569 578
rect 603 544 605 578
rect 553 510 605 544
rect 553 476 569 510
rect 603 476 605 510
rect 553 460 605 476
rect 639 560 864 594
rect 900 569 916 603
rect 950 569 966 603
rect 900 567 966 569
rect 1000 591 1358 607
rect 639 424 673 560
rect 830 533 864 560
rect 1000 557 1002 591
rect 1036 557 1358 591
rect 1000 541 1358 557
rect 485 390 673 424
rect 707 510 757 526
rect 741 476 757 510
rect 830 505 966 533
rect 830 499 1148 505
rect 17 345 110 356
rect 17 311 60 345
rect 94 311 110 345
rect 17 277 110 311
rect 485 281 519 390
rect 707 356 757 476
rect 932 487 1148 499
rect 932 471 1112 487
rect 17 243 60 277
rect 94 243 110 277
rect 17 230 110 243
rect 239 230 519 281
rect 558 346 757 356
rect 558 312 608 346
rect 642 312 757 346
rect 558 310 757 312
rect 793 463 861 465
rect 793 429 811 463
rect 845 437 861 463
rect 1076 453 1112 471
rect 1146 453 1148 487
rect 1076 437 1148 453
rect 845 435 1027 437
rect 845 429 977 435
rect 793 401 977 429
rect 1011 401 1027 435
rect 793 399 1027 401
rect 81 180 147 196
rect 81 146 97 180
rect 131 146 147 180
rect 81 17 147 146
rect 239 180 305 230
rect 239 146 255 180
rect 289 146 305 180
rect 239 130 305 146
rect 397 180 524 196
rect 397 146 413 180
rect 447 146 481 180
rect 515 146 524 180
rect 397 17 524 146
rect 558 180 617 310
rect 558 146 567 180
rect 601 146 617 180
rect 558 130 617 146
rect 687 171 753 276
rect 687 137 703 171
rect 737 137 753 171
rect 687 103 753 137
rect 687 69 703 103
rect 737 69 753 103
rect 687 53 753 69
rect 793 122 827 399
rect 971 367 1027 399
rect 861 349 937 365
rect 861 315 863 349
rect 897 315 937 349
rect 861 281 937 315
rect 861 247 863 281
rect 897 247 937 281
rect 971 333 977 367
rect 1011 333 1027 367
rect 971 299 1027 333
rect 971 265 977 299
rect 1011 265 1027 299
rect 971 249 1027 265
rect 861 156 937 247
rect 1076 157 1142 437
rect 1182 341 1218 541
rect 1076 123 1092 157
rect 1126 123 1142 157
rect 793 106 846 122
rect 793 72 802 106
rect 836 72 846 106
rect 793 56 846 72
rect 880 106 931 122
rect 880 72 888 106
rect 922 72 931 106
rect 880 17 931 72
rect 965 106 1024 122
rect 1076 119 1142 123
rect 1176 325 1218 341
rect 1176 291 1182 325
rect 1216 291 1218 325
rect 1176 275 1218 291
rect 1252 461 1290 477
rect 1286 427 1290 461
rect 1252 283 1290 427
rect 1324 421 1358 541
rect 1396 491 1462 649
rect 1396 457 1412 491
rect 1446 457 1462 491
rect 1396 455 1462 457
rect 1496 513 1670 547
rect 1496 421 1530 513
rect 1324 387 1530 421
rect 1564 461 1602 477
rect 1564 427 1566 461
rect 1600 427 1602 461
rect 1564 353 1602 427
rect 1369 351 1602 353
rect 1369 317 1385 351
rect 1419 317 1602 351
rect 1636 381 1670 513
rect 1704 535 1749 649
rect 1884 561 2272 593
rect 1704 501 1706 535
rect 1740 501 1749 535
rect 1704 465 1749 501
rect 1704 431 1706 465
rect 1740 431 1749 465
rect 1704 415 1749 431
rect 1783 535 1842 551
rect 1783 501 1792 535
rect 1826 501 1842 535
rect 1884 527 1900 561
rect 1934 559 2272 561
rect 1934 527 1950 559
rect 1884 523 1950 527
rect 1783 489 1842 501
rect 2102 507 2168 523
rect 2102 489 2118 507
rect 1783 473 2118 489
rect 2152 473 2168 507
rect 1783 465 2168 473
rect 1783 431 1792 465
rect 1826 455 2168 465
rect 2212 505 2272 559
rect 2212 471 2228 505
rect 2262 471 2272 505
rect 2212 455 2272 471
rect 2306 505 2357 649
rect 2488 542 2552 649
rect 2771 607 2844 649
rect 2771 573 2796 607
rect 2830 573 2844 607
rect 2306 471 2314 505
rect 2348 471 2357 505
rect 2306 455 2357 471
rect 2391 494 2450 510
rect 2391 460 2400 494
rect 2434 460 2450 494
rect 2488 508 2504 542
rect 2538 508 2552 542
rect 2488 492 2552 508
rect 2586 542 2640 558
rect 2586 508 2590 542
rect 2624 508 2640 542
rect 1826 431 1842 455
rect 1783 415 1842 431
rect 2391 451 2450 460
rect 2391 435 2552 451
rect 2391 421 2516 435
rect 1922 403 1982 419
rect 1922 381 1938 403
rect 1636 369 1938 381
rect 1972 369 1982 403
rect 2016 387 2032 421
rect 2066 401 2516 421
rect 2550 401 2552 435
rect 2066 387 2552 401
rect 2016 383 2140 387
rect 1636 347 1982 369
rect 1252 281 1817 283
rect 965 72 974 106
rect 1008 85 1024 106
rect 1176 85 1214 275
rect 1252 247 1532 281
rect 1566 247 1767 281
rect 1801 247 1817 281
rect 1252 245 1817 247
rect 2019 245 2140 383
rect 2500 367 2552 387
rect 1252 143 1286 245
rect 2053 211 2140 245
rect 1365 177 1381 211
rect 1415 195 1559 211
rect 1415 177 1525 195
rect 1365 161 1525 177
rect 1365 145 1559 161
rect 1593 198 1908 202
rect 1593 164 1691 198
rect 1725 164 1777 198
rect 1811 164 1858 198
rect 1892 164 1908 198
rect 1593 162 1908 164
rect 2019 177 2140 211
rect 1008 72 1214 85
rect 965 51 1214 72
rect 1248 115 1286 143
rect 1282 81 1286 115
rect 1248 65 1286 81
rect 1390 106 1456 111
rect 1390 72 1406 106
rect 1440 72 1456 106
rect 1390 17 1456 72
rect 1593 17 1627 162
rect 2019 143 2084 177
rect 2118 143 2140 177
rect 2019 134 2140 143
rect 2174 351 2418 353
rect 2174 317 2368 351
rect 2402 317 2418 351
rect 2500 333 2516 367
rect 2550 333 2552 367
rect 2500 317 2552 333
rect 1663 100 1985 128
rect 2174 100 2208 317
rect 2586 283 2640 508
rect 2771 510 2844 573
rect 2244 281 2640 283
rect 2244 247 2260 281
rect 2294 247 2640 281
rect 2678 481 2737 497
rect 2678 447 2694 481
rect 2728 447 2737 481
rect 2678 413 2737 447
rect 2678 379 2694 413
rect 2728 379 2737 413
rect 2678 329 2737 379
rect 2771 476 2796 510
rect 2830 476 2844 510
rect 2771 415 2844 476
rect 2771 381 2780 415
rect 2814 381 2844 415
rect 2771 365 2844 381
rect 2878 599 2918 615
rect 2878 565 2882 599
rect 2916 565 2918 599
rect 2878 509 2918 565
rect 2878 475 2882 509
rect 2916 475 2918 509
rect 2878 415 2918 475
rect 2952 607 3018 649
rect 2952 573 2968 607
rect 3002 573 3018 607
rect 2952 539 3018 573
rect 2952 505 2968 539
rect 3002 505 3018 539
rect 2952 467 3018 505
rect 2952 433 2968 467
rect 3002 433 3018 467
rect 2878 381 2882 415
rect 2916 399 2918 415
rect 2916 381 3055 399
rect 2878 365 3055 381
rect 2678 313 2867 329
rect 2678 279 2833 313
rect 2678 263 2867 279
rect 1663 87 2208 100
rect 1663 53 1679 87
rect 1713 53 2208 87
rect 2377 183 2443 199
rect 2377 149 2393 183
rect 2427 149 2443 183
rect 2377 17 2443 149
rect 2485 183 2551 247
rect 2485 149 2501 183
rect 2535 149 2551 183
rect 2485 133 2551 149
rect 2678 190 2734 263
rect 2911 227 3055 365
rect 2678 156 2694 190
rect 2728 156 2734 190
rect 2678 140 2734 156
rect 2768 203 2834 219
rect 2768 169 2784 203
rect 2818 169 2834 203
rect 2768 99 2834 169
rect 2768 65 2796 99
rect 2830 65 2834 99
rect 2768 17 2834 65
rect 2878 203 3055 227
rect 2878 169 2882 203
rect 2916 193 3055 203
rect 2916 169 2918 193
rect 2878 101 2918 169
rect 2878 67 2882 101
rect 2916 67 2918 101
rect 2878 51 2918 67
rect 2952 125 2968 159
rect 3002 125 3018 159
rect 2952 89 3018 125
rect 2952 55 2968 89
rect 3002 55 3018 89
rect 2952 17 3018 55
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
<< metal1 >>
rect 0 683 3072 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3072 683
rect 0 617 3072 649
rect 0 17 3072 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3072 17
rect 0 -49 3072 -17
<< labels >>
flabel pwell s 0 0 3072 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 3072 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfstp_2
flabel comment s 1382 272 1382 272 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 3072 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 3072 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 895 168 929 202 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 94 737 128 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 703 168 737 202 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2911 242 2945 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 3007 242 3041 276 0 FreeSans 340 0 0 0 Q
port 10 nsew signal output
flabel locali s 1663 94 1697 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 1759 94 1793 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 1855 94 1889 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 1951 94 1985 128 0 FreeSans 340 0 0 0 SET_B
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3072 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 152778
string GDS_START 132074
<< end >>
