magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 23 157 328 180
rect 947 157 1315 267
rect 23 49 1315 157
rect 0 0 1344 49
<< scnmos >>
rect 102 70 132 154
rect 219 70 249 154
rect 471 47 501 131
rect 557 47 587 131
rect 629 47 659 131
rect 737 47 767 131
rect 809 47 839 131
rect 1026 73 1056 241
rect 1098 73 1128 241
rect 1206 73 1236 241
<< scpmoshvt >>
rect 94 464 124 592
rect 219 464 249 592
rect 424 473 454 601
rect 593 473 623 601
rect 665 473 695 601
rect 770 473 800 557
rect 848 473 878 557
rect 1026 367 1056 619
rect 1112 367 1142 619
rect 1213 367 1243 619
<< ndiff >>
rect 49 128 102 154
rect 49 94 57 128
rect 91 94 102 128
rect 49 70 102 94
rect 132 125 219 154
rect 132 91 159 125
rect 193 91 219 125
rect 132 70 219 91
rect 249 118 302 154
rect 973 217 1026 241
rect 973 183 981 217
rect 1015 183 1026 217
rect 249 84 260 118
rect 294 84 302 118
rect 249 70 302 84
rect 414 101 471 131
rect 414 67 422 101
rect 456 67 471 101
rect 414 47 471 67
rect 501 91 557 131
rect 501 57 512 91
rect 546 57 557 91
rect 501 47 557 57
rect 587 47 629 131
rect 659 101 737 131
rect 659 67 692 101
rect 726 67 737 101
rect 659 47 737 67
rect 767 47 809 131
rect 839 95 911 131
rect 839 61 869 95
rect 903 61 911 95
rect 973 119 1026 183
rect 973 85 981 119
rect 1015 85 1026 119
rect 973 73 1026 85
rect 1056 73 1098 241
rect 1128 218 1206 241
rect 1128 184 1161 218
rect 1195 184 1206 218
rect 1128 119 1206 184
rect 1128 85 1161 119
rect 1195 85 1206 119
rect 1128 73 1206 85
rect 1236 218 1289 241
rect 1236 184 1247 218
rect 1281 184 1289 218
rect 1236 119 1289 184
rect 1236 85 1247 119
rect 1281 85 1289 119
rect 1236 73 1289 85
rect 839 47 911 61
<< pdiff >>
rect 41 580 94 592
rect 41 546 49 580
rect 83 546 94 580
rect 41 510 94 546
rect 41 476 49 510
rect 83 476 94 510
rect 41 464 94 476
rect 124 580 219 592
rect 124 546 135 580
rect 169 546 219 580
rect 124 510 219 546
rect 124 476 135 510
rect 169 476 219 510
rect 124 464 219 476
rect 249 531 313 592
rect 249 497 271 531
rect 305 497 313 531
rect 249 464 313 497
rect 371 531 424 601
rect 371 497 379 531
rect 413 497 424 531
rect 371 473 424 497
rect 454 589 593 601
rect 454 555 524 589
rect 558 555 593 589
rect 454 519 593 555
rect 454 485 524 519
rect 558 485 593 519
rect 454 473 593 485
rect 623 473 665 601
rect 695 557 748 601
rect 973 578 1026 619
rect 973 557 981 578
rect 695 531 770 557
rect 695 497 706 531
rect 740 497 770 531
rect 695 473 770 497
rect 800 473 848 557
rect 878 544 981 557
rect 1015 544 1026 578
rect 878 530 1026 544
rect 878 496 889 530
rect 923 496 1026 530
rect 878 473 1026 496
rect 973 367 1026 473
rect 1056 599 1112 619
rect 1056 565 1067 599
rect 1101 565 1112 599
rect 1056 494 1112 565
rect 1056 460 1067 494
rect 1101 460 1112 494
rect 1056 367 1112 460
rect 1142 569 1213 619
rect 1142 535 1161 569
rect 1195 535 1213 569
rect 1142 367 1213 535
rect 1243 599 1296 619
rect 1243 565 1254 599
rect 1288 565 1296 599
rect 1243 503 1296 565
rect 1243 469 1254 503
rect 1288 469 1296 503
rect 1243 420 1296 469
rect 1243 386 1254 420
rect 1288 386 1296 420
rect 1243 367 1296 386
<< ndiffc >>
rect 57 94 91 128
rect 159 91 193 125
rect 981 183 1015 217
rect 260 84 294 118
rect 422 67 456 101
rect 512 57 546 91
rect 692 67 726 101
rect 869 61 903 95
rect 981 85 1015 119
rect 1161 184 1195 218
rect 1161 85 1195 119
rect 1247 184 1281 218
rect 1247 85 1281 119
<< pdiffc >>
rect 49 546 83 580
rect 49 476 83 510
rect 135 546 169 580
rect 135 476 169 510
rect 271 497 305 531
rect 379 497 413 531
rect 524 555 558 589
rect 524 485 558 519
rect 706 497 740 531
rect 981 544 1015 578
rect 889 496 923 530
rect 1067 565 1101 599
rect 1067 460 1101 494
rect 1161 535 1195 569
rect 1254 565 1288 599
rect 1254 469 1288 503
rect 1254 386 1288 420
<< poly >>
rect 94 592 124 618
rect 219 592 249 618
rect 424 601 454 627
rect 593 601 623 627
rect 665 601 695 627
rect 1026 619 1056 645
rect 1112 619 1142 645
rect 1213 619 1243 645
rect 770 557 800 583
rect 848 557 878 583
rect 94 310 124 464
rect 219 310 249 464
rect 424 432 454 473
rect 593 441 623 473
rect 293 416 454 432
rect 293 382 309 416
rect 343 382 454 416
rect 293 366 454 382
rect 94 294 177 310
rect 94 260 127 294
rect 161 260 177 294
rect 94 226 177 260
rect 94 192 127 226
rect 161 192 177 226
rect 94 176 177 192
rect 219 294 287 310
rect 219 260 237 294
rect 271 260 287 294
rect 219 226 287 260
rect 219 192 237 226
rect 271 192 287 226
rect 219 176 287 192
rect 424 219 454 366
rect 496 425 623 441
rect 496 391 512 425
rect 546 411 623 425
rect 546 391 587 411
rect 496 357 587 391
rect 496 323 512 357
rect 546 323 587 357
rect 496 307 587 323
rect 424 203 515 219
rect 102 154 132 176
rect 219 154 249 176
rect 424 169 465 203
rect 499 169 515 203
rect 424 153 515 169
rect 471 131 501 153
rect 557 131 587 307
rect 665 333 695 473
rect 770 441 800 473
rect 848 441 878 473
rect 738 425 804 441
rect 738 391 754 425
rect 788 391 804 425
rect 738 375 804 391
rect 846 425 912 441
rect 846 391 862 425
rect 896 391 912 425
rect 846 375 912 391
rect 665 303 803 333
rect 737 285 803 303
rect 629 245 695 261
rect 629 211 645 245
rect 679 211 695 245
rect 629 195 695 211
rect 737 251 753 285
rect 787 251 803 285
rect 737 235 803 251
rect 629 131 659 195
rect 737 131 767 235
rect 846 183 876 375
rect 1026 333 1056 367
rect 1112 335 1142 367
rect 933 317 1056 333
rect 933 283 949 317
rect 983 283 1056 317
rect 933 267 1056 283
rect 1026 241 1056 267
rect 1098 319 1164 335
rect 1213 334 1243 367
rect 1098 285 1114 319
rect 1148 285 1164 319
rect 1098 269 1164 285
rect 1206 318 1272 334
rect 1206 284 1222 318
rect 1256 284 1272 318
rect 1098 241 1128 269
rect 1206 268 1272 284
rect 1206 241 1236 268
rect 809 153 876 183
rect 809 131 839 153
rect 102 44 132 70
rect 219 44 249 70
rect 1026 47 1056 73
rect 1098 47 1128 73
rect 1206 47 1236 73
rect 471 21 501 47
rect 557 21 587 47
rect 629 21 659 47
rect 737 21 767 47
rect 809 21 839 47
<< polycont >>
rect 309 382 343 416
rect 127 260 161 294
rect 127 192 161 226
rect 237 260 271 294
rect 237 192 271 226
rect 512 391 546 425
rect 512 323 546 357
rect 465 169 499 203
rect 754 391 788 425
rect 862 391 896 425
rect 645 211 679 245
rect 753 251 787 285
rect 949 283 983 317
rect 1114 285 1148 319
rect 1222 284 1256 318
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 33 580 91 596
rect 33 546 49 580
rect 83 546 91 580
rect 33 510 91 546
rect 33 476 49 510
rect 83 476 91 510
rect 33 426 91 476
rect 131 580 169 649
rect 131 546 135 580
rect 131 510 169 546
rect 131 476 135 510
rect 131 460 169 476
rect 203 581 484 615
rect 203 426 237 581
rect 271 531 345 547
rect 305 497 345 531
rect 271 481 345 497
rect 33 392 237 426
rect 309 416 345 481
rect 33 128 91 392
rect 343 382 345 416
rect 125 294 173 358
rect 125 260 127 294
rect 161 260 173 294
rect 125 226 173 260
rect 125 192 127 226
rect 161 192 173 226
rect 125 168 173 192
rect 207 294 275 358
rect 207 260 237 294
rect 271 260 275 294
rect 207 226 275 260
rect 207 192 237 226
rect 271 192 275 226
rect 207 168 275 192
rect 309 134 345 382
rect 33 94 57 128
rect 33 78 91 94
rect 143 125 209 134
rect 143 91 159 125
rect 193 91 209 125
rect 143 17 209 91
rect 244 118 345 134
rect 244 84 260 118
rect 294 84 345 118
rect 244 66 345 84
rect 379 531 416 547
rect 413 497 416 531
rect 379 273 416 497
rect 450 435 484 581
rect 518 589 564 649
rect 518 555 524 589
rect 558 555 564 589
rect 518 519 564 555
rect 518 485 524 519
rect 558 485 564 519
rect 518 469 564 485
rect 598 581 810 615
rect 450 425 562 435
rect 450 391 512 425
rect 546 391 562 425
rect 450 357 562 391
rect 450 323 512 357
rect 546 323 562 357
rect 450 307 562 323
rect 598 273 632 581
rect 668 531 740 547
rect 668 497 706 531
rect 668 481 740 497
rect 668 355 702 481
rect 776 441 810 581
rect 873 578 1017 649
rect 873 544 981 578
rect 1015 544 1017 578
rect 873 530 1017 544
rect 873 496 889 530
rect 923 528 1017 530
rect 1051 599 1111 615
rect 1051 565 1067 599
rect 1101 565 1111 599
rect 923 496 983 528
rect 873 480 983 496
rect 1051 494 1111 565
rect 1145 569 1211 649
rect 1145 535 1161 569
rect 1195 535 1211 569
rect 1145 528 1211 535
rect 1252 599 1326 615
rect 1252 565 1254 599
rect 1288 565 1326 599
rect 1252 503 1326 565
rect 1017 460 1067 494
rect 1101 460 1218 494
rect 1017 441 1051 460
rect 738 425 810 441
rect 738 391 754 425
rect 788 391 810 425
rect 738 389 810 391
rect 846 425 1051 441
rect 846 391 862 425
rect 896 391 1051 425
rect 846 389 1051 391
rect 668 321 983 355
rect 907 317 983 321
rect 731 285 803 287
rect 379 245 695 273
rect 379 239 645 245
rect 379 107 415 239
rect 629 211 645 239
rect 679 211 695 245
rect 629 209 695 211
rect 731 251 753 285
rect 787 251 803 285
rect 731 235 803 251
rect 907 283 949 317
rect 907 267 983 283
rect 449 203 515 205
rect 449 169 465 203
rect 499 175 515 203
rect 731 175 765 235
rect 907 179 941 267
rect 1017 233 1051 389
rect 499 169 765 175
rect 449 141 765 169
rect 801 145 941 179
rect 975 217 1051 233
rect 975 183 981 217
rect 1015 183 1051 217
rect 801 107 835 145
rect 975 119 1051 183
rect 379 101 472 107
rect 379 67 422 101
rect 456 67 472 101
rect 379 51 472 67
rect 506 91 562 107
rect 506 57 512 91
rect 546 57 562 91
rect 676 101 835 107
rect 676 67 692 101
rect 726 67 835 101
rect 676 63 835 67
rect 869 95 919 111
rect 506 17 562 57
rect 903 61 919 95
rect 975 85 981 119
rect 1015 85 1051 119
rect 975 69 1051 85
rect 1085 319 1148 426
rect 1085 285 1114 319
rect 1085 269 1148 285
rect 1184 334 1218 460
rect 1252 469 1254 503
rect 1288 469 1326 503
rect 1252 420 1326 469
rect 1252 386 1254 420
rect 1288 386 1326 420
rect 1252 370 1326 386
rect 1184 318 1256 334
rect 1184 284 1222 318
rect 1085 69 1121 269
rect 1184 268 1256 284
rect 1290 234 1326 370
rect 1155 218 1198 234
rect 1155 184 1161 218
rect 1195 184 1198 218
rect 1155 119 1198 184
rect 1155 85 1161 119
rect 1195 85 1198 119
rect 869 17 919 61
rect 1155 17 1198 85
rect 1232 218 1326 234
rect 1232 184 1247 218
rect 1281 184 1326 218
rect 1232 119 1326 184
rect 1232 85 1247 119
rect 1281 85 1326 119
rect 1232 69 1326 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlrtp_1
flabel comment s 432 308 432 308 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 1087 94 1121 128 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1087 390 1121 424 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 464 1313 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 1279 538 1313 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1909354
string GDS_START 1897964
<< end >>
