magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1874 1975
<< nwell >>
rect -38 331 614 704
<< pwell >>
rect 1 49 477 243
rect 0 0 576 49
<< scnmos >>
rect 80 49 110 217
rect 152 49 182 217
rect 260 49 290 217
rect 368 49 398 217
<< scpmoshvt >>
rect 80 367 110 619
rect 188 367 218 619
rect 296 367 326 619
rect 368 367 398 619
<< ndiff >>
rect 27 205 80 217
rect 27 171 35 205
rect 69 171 80 205
rect 27 95 80 171
rect 27 61 35 95
rect 69 61 80 95
rect 27 49 80 61
rect 110 49 152 217
rect 182 177 260 217
rect 182 143 209 177
rect 243 143 260 177
rect 182 101 260 143
rect 182 67 209 101
rect 243 67 260 101
rect 182 49 260 67
rect 290 165 368 217
rect 290 131 320 165
rect 354 131 368 165
rect 290 91 368 131
rect 290 57 320 91
rect 354 57 368 91
rect 290 49 368 57
rect 398 205 451 217
rect 398 171 409 205
rect 443 171 451 205
rect 398 101 451 171
rect 398 67 409 101
rect 443 67 451 101
rect 398 49 451 67
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 508 80 565
rect 27 474 35 508
rect 69 474 80 508
rect 27 420 80 474
rect 27 386 35 420
rect 69 386 80 420
rect 27 367 80 386
rect 110 607 188 619
rect 110 573 132 607
rect 166 573 188 607
rect 110 496 188 573
rect 110 462 132 496
rect 166 462 188 496
rect 110 367 188 462
rect 218 607 296 619
rect 218 573 241 607
rect 275 573 296 607
rect 218 508 296 573
rect 218 474 241 508
rect 275 474 296 508
rect 218 420 296 474
rect 218 386 241 420
rect 275 386 296 420
rect 218 367 296 386
rect 326 367 368 619
rect 398 607 451 619
rect 398 573 409 607
rect 443 573 451 607
rect 398 515 451 573
rect 398 481 409 515
rect 443 481 451 515
rect 398 419 451 481
rect 398 385 409 419
rect 443 385 451 419
rect 398 367 451 385
<< ndiffc >>
rect 35 171 69 205
rect 35 61 69 95
rect 209 143 243 177
rect 209 67 243 101
rect 320 131 354 165
rect 320 57 354 91
rect 409 171 443 205
rect 409 67 443 101
<< pdiffc >>
rect 35 565 69 599
rect 35 474 69 508
rect 35 386 69 420
rect 132 573 166 607
rect 132 462 166 496
rect 241 573 275 607
rect 241 474 275 508
rect 241 386 275 420
rect 409 573 443 607
rect 409 481 443 515
rect 409 385 443 419
<< poly >>
rect 80 619 110 645
rect 188 619 218 645
rect 296 619 326 645
rect 368 619 398 645
rect 80 308 110 367
rect 27 292 110 308
rect 188 305 218 367
rect 296 335 326 367
rect 27 258 43 292
rect 77 258 110 292
rect 27 242 110 258
rect 80 217 110 242
rect 152 289 218 305
rect 152 255 168 289
rect 202 255 218 289
rect 152 239 218 255
rect 260 319 326 335
rect 260 285 276 319
rect 310 285 326 319
rect 260 269 326 285
rect 368 325 398 367
rect 368 309 460 325
rect 368 275 410 309
rect 444 275 460 309
rect 152 217 182 239
rect 260 217 290 269
rect 368 259 460 275
rect 368 217 398 259
rect 80 23 110 49
rect 152 23 182 49
rect 260 23 290 49
rect 368 23 398 49
<< polycont >>
rect 43 258 77 292
rect 168 255 202 289
rect 276 285 310 319
rect 410 275 444 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 19 599 82 615
rect 19 565 35 599
rect 69 565 82 599
rect 19 508 82 565
rect 19 474 35 508
rect 69 474 82 508
rect 19 420 82 474
rect 116 607 182 649
rect 116 573 132 607
rect 166 573 182 607
rect 116 496 182 573
rect 116 462 132 496
rect 166 462 182 496
rect 116 454 182 462
rect 225 607 291 615
rect 225 573 241 607
rect 275 573 291 607
rect 225 508 291 573
rect 225 474 241 508
rect 275 474 291 508
rect 225 420 291 474
rect 19 386 35 420
rect 69 386 241 420
rect 275 386 291 420
rect 393 607 557 615
rect 393 573 409 607
rect 443 573 557 607
rect 393 515 557 573
rect 393 481 409 515
rect 443 481 557 515
rect 393 419 557 481
rect 393 385 409 419
rect 443 385 557 419
rect 19 292 85 352
rect 19 258 43 292
rect 77 258 85 292
rect 19 242 85 258
rect 119 305 175 352
rect 253 319 360 352
rect 119 289 202 305
rect 119 255 168 289
rect 253 285 276 319
rect 310 285 360 319
rect 253 269 360 285
rect 394 309 461 350
rect 394 275 410 309
rect 444 275 461 309
rect 394 269 461 275
rect 119 239 202 255
rect 19 205 85 208
rect 19 171 35 205
rect 69 171 85 205
rect 19 95 85 171
rect 19 61 35 95
rect 69 61 85 95
rect 119 76 169 239
rect 500 235 557 385
rect 236 205 557 235
rect 236 199 409 205
rect 236 193 270 199
rect 203 177 270 193
rect 203 143 209 177
rect 243 143 270 177
rect 404 171 409 199
rect 443 177 557 205
rect 443 171 459 177
rect 203 101 270 143
rect 19 17 85 61
rect 203 67 209 101
rect 243 67 270 101
rect 203 51 270 67
rect 304 131 320 165
rect 354 131 370 165
rect 304 91 370 131
rect 304 57 320 91
rect 354 57 370 91
rect 304 17 370 57
rect 404 101 459 171
rect 404 67 409 101
rect 443 67 459 101
rect 404 51 459 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
<< metal1 >>
rect 0 683 576 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 576 683
rect 0 617 576 649
rect 0 17 576 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 576 17
rect 0 -49 576 -17
<< labels >>
flabel pwell s 0 0 576 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 576 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a211oi_1
flabel metal1 s 0 617 576 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 576 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 538 545 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 576 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 213646
string GDS_START 207526
<< end >>
