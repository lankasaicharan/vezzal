magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 1 49 812 241
rect 0 0 864 49
<< scnmos >>
rect 80 47 110 215
rect 234 47 264 215
rect 321 47 351 215
rect 511 47 541 215
rect 583 47 613 215
rect 703 47 733 215
<< scpmoshvt >>
rect 80 367 110 619
rect 234 367 264 619
rect 321 367 351 619
rect 511 367 541 619
rect 613 367 643 619
rect 703 367 733 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 94 80 169
rect 27 60 35 94
rect 69 60 80 94
rect 27 47 80 60
rect 110 200 234 215
rect 110 166 139 200
rect 173 166 234 200
rect 110 93 234 166
rect 110 59 139 93
rect 173 59 234 93
rect 110 47 234 59
rect 264 47 321 215
rect 351 185 511 215
rect 351 151 387 185
rect 421 151 466 185
rect 500 151 511 185
rect 351 101 511 151
rect 351 67 387 101
rect 421 67 466 101
rect 500 67 511 101
rect 351 47 511 67
rect 541 47 583 215
rect 613 122 703 215
rect 613 88 642 122
rect 676 88 703 122
rect 613 47 703 88
rect 733 203 786 215
rect 733 169 744 203
rect 778 169 786 203
rect 733 101 786 169
rect 733 67 744 101
rect 778 67 786 101
rect 733 47 786 67
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 509 80 565
rect 27 475 35 509
rect 69 475 80 509
rect 27 413 80 475
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 607 234 619
rect 110 573 121 607
rect 155 573 189 607
rect 223 573 234 607
rect 110 525 234 573
rect 110 491 121 525
rect 155 491 189 525
rect 223 491 234 525
rect 110 439 234 491
rect 110 405 121 439
rect 155 405 189 439
rect 223 405 234 439
rect 110 367 234 405
rect 264 599 321 619
rect 264 565 276 599
rect 310 565 321 599
rect 264 527 321 565
rect 264 493 276 527
rect 310 493 321 527
rect 264 455 321 493
rect 264 421 276 455
rect 310 421 321 455
rect 264 367 321 421
rect 351 607 404 619
rect 351 573 362 607
rect 396 573 404 607
rect 351 513 404 573
rect 351 479 362 513
rect 396 479 404 513
rect 351 367 404 479
rect 458 607 511 619
rect 458 573 466 607
rect 500 573 511 607
rect 458 513 511 573
rect 458 479 466 513
rect 500 479 511 513
rect 458 367 511 479
rect 541 542 613 619
rect 541 508 566 542
rect 600 508 613 542
rect 541 439 613 508
rect 541 405 566 439
rect 600 405 613 439
rect 541 367 613 405
rect 643 599 703 619
rect 643 565 655 599
rect 689 565 703 599
rect 643 529 703 565
rect 643 495 655 529
rect 689 495 703 529
rect 643 455 703 495
rect 643 421 655 455
rect 689 421 703 455
rect 643 367 703 421
rect 733 599 786 619
rect 733 565 744 599
rect 778 565 786 599
rect 733 504 786 565
rect 733 470 744 504
rect 778 470 786 504
rect 733 413 786 470
rect 733 379 744 413
rect 778 379 786 413
rect 733 367 786 379
<< ndiffc >>
rect 35 169 69 203
rect 35 60 69 94
rect 139 166 173 200
rect 139 59 173 93
rect 387 151 421 185
rect 466 151 500 185
rect 387 67 421 101
rect 466 67 500 101
rect 642 88 676 122
rect 744 169 778 203
rect 744 67 778 101
<< pdiffc >>
rect 35 565 69 599
rect 35 475 69 509
rect 35 379 69 413
rect 121 573 155 607
rect 189 573 223 607
rect 121 491 155 525
rect 189 491 223 525
rect 121 405 155 439
rect 189 405 223 439
rect 276 565 310 599
rect 276 493 310 527
rect 276 421 310 455
rect 362 573 396 607
rect 362 479 396 513
rect 466 573 500 607
rect 466 479 500 513
rect 566 508 600 542
rect 566 405 600 439
rect 655 565 689 599
rect 655 495 689 529
rect 655 421 689 455
rect 744 565 778 599
rect 744 470 778 504
rect 744 379 778 413
<< poly >>
rect 80 619 110 645
rect 234 619 264 645
rect 321 619 351 645
rect 511 619 541 645
rect 613 619 643 645
rect 703 619 733 645
rect 80 335 110 367
rect 80 311 153 335
rect 80 277 103 311
rect 137 277 153 311
rect 234 303 264 367
rect 80 261 153 277
rect 195 287 264 303
rect 80 215 110 261
rect 195 253 211 287
rect 245 253 264 287
rect 195 237 264 253
rect 234 215 264 237
rect 321 303 351 367
rect 511 345 541 367
rect 321 287 387 303
rect 321 253 337 287
rect 371 253 387 287
rect 321 237 387 253
rect 461 287 541 345
rect 613 303 643 367
rect 703 303 733 367
rect 461 253 477 287
rect 511 253 541 287
rect 589 287 655 303
rect 589 267 605 287
rect 461 237 541 253
rect 321 215 351 237
rect 511 215 541 237
rect 583 253 605 267
rect 639 253 655 287
rect 583 237 655 253
rect 703 287 769 303
rect 703 253 719 287
rect 753 253 769 287
rect 703 237 769 253
rect 583 215 613 237
rect 703 215 733 237
rect 80 21 110 47
rect 234 21 264 47
rect 321 21 351 47
rect 511 21 541 47
rect 583 21 613 47
rect 703 21 733 47
<< polycont >>
rect 103 277 137 311
rect 211 253 245 287
rect 337 253 371 287
rect 477 253 511 287
rect 605 253 639 287
rect 719 253 753 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 17 599 69 615
rect 17 565 35 599
rect 17 509 69 565
rect 17 475 35 509
rect 17 413 69 475
rect 17 379 35 413
rect 105 607 239 649
rect 105 573 121 607
rect 155 573 189 607
rect 223 573 239 607
rect 105 525 239 573
rect 105 491 121 525
rect 155 491 189 525
rect 223 491 239 525
rect 105 439 239 491
rect 105 405 121 439
rect 155 405 189 439
rect 223 405 239 439
rect 273 599 312 615
rect 273 565 276 599
rect 310 565 312 599
rect 273 527 312 565
rect 273 493 276 527
rect 310 493 312 527
rect 273 455 312 493
rect 346 607 412 649
rect 346 573 362 607
rect 396 573 412 607
rect 346 513 412 573
rect 346 479 362 513
rect 396 479 412 513
rect 346 473 412 479
rect 450 607 694 615
rect 450 573 466 607
rect 500 599 694 607
rect 500 581 655 599
rect 500 573 516 581
rect 450 513 516 573
rect 650 565 655 581
rect 689 565 694 599
rect 450 479 466 513
rect 500 479 516 513
rect 450 473 516 479
rect 550 542 616 547
rect 550 508 566 542
rect 600 508 616 542
rect 273 421 276 455
rect 310 439 312 455
rect 550 439 616 508
rect 310 421 566 439
rect 273 405 566 421
rect 600 405 616 439
rect 650 529 694 565
rect 650 495 655 529
rect 689 495 694 529
rect 650 455 694 495
rect 650 421 655 455
rect 689 421 694 455
rect 650 405 694 421
rect 728 599 794 615
rect 728 565 744 599
rect 778 565 794 599
rect 728 504 794 565
rect 728 470 744 504
rect 778 470 794 504
rect 728 413 794 470
rect 17 215 69 379
rect 728 379 744 413
rect 778 379 794 413
rect 728 371 794 379
rect 103 337 794 371
rect 103 311 153 337
rect 137 277 153 311
rect 103 261 153 277
rect 211 287 273 303
rect 245 253 273 287
rect 211 237 273 253
rect 17 203 85 215
rect 17 169 35 203
rect 69 169 85 203
rect 17 94 85 169
rect 17 60 35 94
rect 69 60 85 94
rect 17 51 85 60
rect 123 200 189 203
rect 123 166 139 200
rect 173 166 189 200
rect 123 93 189 166
rect 123 59 139 93
rect 173 59 189 93
rect 223 66 273 237
rect 307 287 371 303
rect 307 253 337 287
rect 307 237 371 253
rect 307 66 353 237
rect 405 203 441 337
rect 477 287 557 303
rect 511 253 557 287
rect 477 237 557 253
rect 591 287 658 303
rect 591 253 605 287
rect 639 253 658 287
rect 591 237 658 253
rect 692 253 719 287
rect 753 253 847 287
rect 692 237 847 253
rect 387 185 744 203
rect 421 151 466 185
rect 500 169 744 185
rect 778 169 794 203
rect 500 167 794 169
rect 500 151 516 167
rect 387 101 516 151
rect 421 67 466 101
rect 500 67 516 101
rect 123 17 189 59
rect 387 51 516 67
rect 626 122 692 133
rect 626 88 642 122
rect 676 88 692 122
rect 626 17 692 88
rect 740 101 794 167
rect 740 67 744 101
rect 778 67 794 101
rect 740 51 794 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a221o_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 319 94 353 128 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 94 257 128 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 168 257 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6121196
string GDS_START 6112176
<< end >>
