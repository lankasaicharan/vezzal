magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 68 49 854 241
rect 0 0 864 49
<< scnmos >>
rect 147 131 177 215
rect 303 47 333 215
rect 389 47 419 215
rect 496 47 526 215
rect 591 47 621 215
rect 745 131 775 215
<< scpmoshvt >>
rect 80 508 110 592
rect 303 367 333 619
rect 375 367 405 619
rect 483 367 513 619
rect 591 367 621 619
rect 699 367 729 451
<< ndiff >>
rect 94 191 147 215
rect 94 157 102 191
rect 136 157 147 191
rect 94 131 147 157
rect 177 179 303 215
rect 177 145 248 179
rect 282 145 303 179
rect 177 131 303 145
rect 250 93 303 131
rect 250 59 258 93
rect 292 59 303 93
rect 250 47 303 59
rect 333 203 389 215
rect 333 169 344 203
rect 378 169 389 203
rect 333 101 389 169
rect 333 67 344 101
rect 378 67 389 101
rect 333 47 389 67
rect 419 167 496 215
rect 419 133 439 167
rect 473 133 496 167
rect 419 93 496 133
rect 419 59 439 93
rect 473 59 496 93
rect 419 47 496 59
rect 526 203 591 215
rect 526 169 537 203
rect 571 169 591 203
rect 526 101 591 169
rect 526 67 537 101
rect 571 67 591 101
rect 526 47 591 67
rect 621 183 745 215
rect 621 149 632 183
rect 666 149 700 183
rect 734 149 745 183
rect 621 131 745 149
rect 775 189 828 215
rect 775 155 786 189
rect 820 155 828 189
rect 775 131 828 155
rect 621 93 674 131
rect 621 59 632 93
rect 666 59 674 93
rect 621 47 674 59
<< pdiff >>
rect 250 599 303 619
rect 27 568 80 592
rect 27 534 35 568
rect 69 534 80 568
rect 27 508 80 534
rect 110 568 163 592
rect 110 534 121 568
rect 155 534 163 568
rect 110 508 163 534
rect 250 565 258 599
rect 292 565 303 599
rect 250 505 303 565
rect 250 471 258 505
rect 292 471 303 505
rect 250 413 303 471
rect 250 379 258 413
rect 292 379 303 413
rect 250 367 303 379
rect 333 367 375 619
rect 405 367 483 619
rect 513 367 591 619
rect 621 607 674 619
rect 621 573 632 607
rect 666 573 674 607
rect 621 501 674 573
rect 621 467 632 501
rect 666 467 674 501
rect 621 451 674 467
rect 621 367 699 451
rect 729 424 782 451
rect 729 390 740 424
rect 774 390 782 424
rect 729 367 782 390
<< ndiffc >>
rect 102 157 136 191
rect 248 145 282 179
rect 258 59 292 93
rect 344 169 378 203
rect 344 67 378 101
rect 439 133 473 167
rect 439 59 473 93
rect 537 169 571 203
rect 537 67 571 101
rect 632 149 666 183
rect 700 149 734 183
rect 786 155 820 189
rect 632 59 666 93
<< pdiffc >>
rect 35 534 69 568
rect 121 534 155 568
rect 258 565 292 599
rect 258 471 292 505
rect 258 379 292 413
rect 632 573 666 607
rect 632 467 666 501
rect 740 390 774 424
<< poly >>
rect 303 619 333 645
rect 375 619 405 645
rect 483 619 513 645
rect 591 619 621 645
rect 80 592 110 618
rect 80 376 110 508
rect 80 360 177 376
rect 699 451 729 477
rect 80 326 96 360
rect 130 326 177 360
rect 303 345 333 367
rect 80 292 177 326
rect 255 303 333 345
rect 80 258 96 292
rect 130 258 177 292
rect 80 242 177 258
rect 147 215 177 242
rect 219 287 333 303
rect 219 253 235 287
rect 269 253 333 287
rect 375 335 405 367
rect 483 335 513 367
rect 375 319 441 335
rect 375 285 391 319
rect 425 285 441 319
rect 375 269 441 285
rect 483 319 549 335
rect 483 285 499 319
rect 533 285 549 319
rect 483 269 549 285
rect 591 303 621 367
rect 699 335 729 367
rect 699 319 813 335
rect 699 305 763 319
rect 591 287 657 303
rect 219 237 333 253
rect 303 215 333 237
rect 389 215 419 269
rect 496 215 526 269
rect 591 253 607 287
rect 641 253 657 287
rect 591 237 657 253
rect 745 285 763 305
rect 797 285 813 319
rect 745 269 813 285
rect 591 215 621 237
rect 745 215 775 269
rect 147 105 177 131
rect 745 105 775 131
rect 303 21 333 47
rect 389 21 419 47
rect 496 21 526 47
rect 591 21 621 47
<< polycont >>
rect 96 326 130 360
rect 96 258 130 292
rect 235 253 269 287
rect 391 285 425 319
rect 499 285 533 319
rect 607 253 641 287
rect 763 285 797 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 19 568 71 584
rect 19 534 35 568
rect 69 534 71 568
rect 19 492 71 534
rect 105 568 171 649
rect 105 534 121 568
rect 155 534 171 568
rect 105 526 171 534
rect 242 599 339 615
rect 242 565 258 599
rect 292 565 339 599
rect 242 505 339 565
rect 19 458 206 492
rect 17 360 130 424
rect 17 326 96 360
rect 17 292 130 326
rect 17 258 96 292
rect 17 241 130 258
rect 164 303 206 458
rect 242 471 258 505
rect 292 471 339 505
rect 242 413 339 471
rect 616 607 682 649
rect 616 573 632 607
rect 666 573 682 607
rect 616 501 682 573
rect 616 467 632 501
rect 666 467 682 501
rect 616 463 682 467
rect 242 379 258 413
rect 292 379 339 413
rect 242 363 339 379
rect 164 287 271 303
rect 164 253 235 287
rect 269 253 271 287
rect 164 237 271 253
rect 305 251 339 363
rect 375 424 790 429
rect 375 390 740 424
rect 774 390 790 424
rect 375 386 790 390
rect 375 319 441 386
rect 375 285 391 319
rect 425 285 441 319
rect 483 319 549 352
rect 483 285 499 319
rect 533 285 549 319
rect 605 287 643 352
rect 605 253 607 287
rect 641 253 643 287
rect 164 207 198 237
rect 305 217 571 251
rect 605 221 643 253
rect 677 251 711 386
rect 747 319 847 352
rect 747 285 763 319
rect 797 285 847 319
rect 677 217 832 251
rect 305 213 389 217
rect 86 191 198 207
rect 86 157 102 191
rect 136 157 198 191
rect 342 203 389 213
rect 86 141 198 157
rect 232 145 248 179
rect 282 145 308 179
rect 232 93 308 145
rect 232 59 258 93
rect 292 59 308 93
rect 232 17 308 59
rect 342 169 344 203
rect 378 169 389 203
rect 511 203 571 217
rect 342 101 389 169
rect 342 67 344 101
rect 378 67 389 101
rect 342 51 389 67
rect 423 167 477 183
rect 423 133 439 167
rect 473 133 477 167
rect 423 93 477 133
rect 423 59 439 93
rect 473 59 477 93
rect 423 17 477 59
rect 511 169 537 203
rect 784 189 832 217
rect 511 101 571 169
rect 511 67 537 101
rect 511 51 571 67
rect 616 149 632 183
rect 666 149 700 183
rect 734 149 750 183
rect 616 93 750 149
rect 784 155 786 189
rect 820 155 832 189
rect 784 139 832 155
rect 616 59 632 93
rect 666 59 750 93
rect 616 17 750 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4bb_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 511 94 545 128 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 511 168 545 202 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3352976
string GDS_START 3345644
<< end >>
