magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 60 49 664 157
rect 0 0 672 49
<< scnmos >>
rect 143 47 173 131
rect 221 47 251 131
rect 299 47 329 131
rect 377 47 407 131
rect 479 47 509 131
rect 551 47 581 131
<< scpmoshvt >>
rect 87 409 137 609
rect 193 409 243 609
rect 299 409 349 609
rect 405 409 455 609
rect 515 409 565 609
<< ndiff >>
rect 86 108 143 131
rect 86 74 98 108
rect 132 74 143 108
rect 86 47 143 74
rect 173 47 221 131
rect 251 47 299 131
rect 329 47 377 131
rect 407 103 479 131
rect 407 69 418 103
rect 452 69 479 103
rect 407 47 479 69
rect 509 47 551 131
rect 581 111 638 131
rect 581 77 592 111
rect 626 77 638 111
rect 581 47 638 77
<< pdiff >>
rect 30 597 87 609
rect 30 563 42 597
rect 76 563 87 597
rect 30 512 87 563
rect 30 478 42 512
rect 76 478 87 512
rect 30 409 87 478
rect 137 597 193 609
rect 137 563 148 597
rect 182 563 193 597
rect 137 526 193 563
rect 137 492 148 526
rect 182 492 193 526
rect 137 455 193 492
rect 137 421 148 455
rect 182 421 193 455
rect 137 409 193 421
rect 243 597 299 609
rect 243 563 254 597
rect 288 563 299 597
rect 243 525 299 563
rect 243 491 254 525
rect 288 491 299 525
rect 243 409 299 491
rect 349 597 405 609
rect 349 563 360 597
rect 394 563 405 597
rect 349 526 405 563
rect 349 492 360 526
rect 394 492 405 526
rect 349 455 405 492
rect 349 421 360 455
rect 394 421 405 455
rect 349 409 405 421
rect 455 597 515 609
rect 455 563 466 597
rect 500 563 515 597
rect 455 526 515 563
rect 455 492 466 526
rect 500 492 515 526
rect 455 455 515 492
rect 455 421 466 455
rect 500 421 515 455
rect 455 409 515 421
rect 565 597 622 609
rect 565 563 576 597
rect 610 563 622 597
rect 565 526 622 563
rect 565 492 576 526
rect 610 492 622 526
rect 565 455 622 492
rect 565 421 576 455
rect 610 421 622 455
rect 565 409 622 421
<< ndiffc >>
rect 98 74 132 108
rect 418 69 452 103
rect 592 77 626 111
<< pdiffc >>
rect 42 563 76 597
rect 42 478 76 512
rect 148 563 182 597
rect 148 492 182 526
rect 148 421 182 455
rect 254 563 288 597
rect 254 491 288 525
rect 360 563 394 597
rect 360 492 394 526
rect 360 421 394 455
rect 466 563 500 597
rect 466 492 500 526
rect 466 421 500 455
rect 576 563 610 597
rect 576 492 610 526
rect 576 421 610 455
<< poly >>
rect 87 609 137 635
rect 193 609 243 635
rect 299 609 349 635
rect 405 609 455 635
rect 515 609 565 635
rect 87 231 137 409
rect 193 356 243 409
rect 299 369 349 409
rect 405 369 455 409
rect 515 369 565 409
rect 185 340 251 356
rect 185 306 201 340
rect 235 306 251 340
rect 185 290 251 306
rect 107 215 173 231
rect 107 181 123 215
rect 157 181 173 215
rect 107 165 173 181
rect 143 131 173 165
rect 221 131 251 290
rect 293 353 359 369
rect 293 319 309 353
rect 343 319 359 353
rect 293 285 359 319
rect 293 251 309 285
rect 343 251 359 285
rect 293 235 359 251
rect 401 353 467 369
rect 401 319 417 353
rect 451 319 467 353
rect 401 285 467 319
rect 401 251 417 285
rect 451 251 467 285
rect 401 235 467 251
rect 515 353 581 369
rect 515 319 531 353
rect 565 319 581 353
rect 515 285 581 319
rect 515 251 531 285
rect 565 251 581 285
rect 515 235 581 251
rect 299 131 329 235
rect 401 176 431 235
rect 515 176 545 235
rect 377 146 431 176
rect 479 146 581 176
rect 377 131 407 146
rect 479 131 509 146
rect 551 131 581 146
rect 143 21 173 47
rect 221 21 251 47
rect 299 21 329 47
rect 377 21 407 47
rect 479 21 509 47
rect 551 21 581 47
<< polycont >>
rect 201 306 235 340
rect 123 181 157 215
rect 309 319 343 353
rect 309 251 343 285
rect 417 319 451 353
rect 417 251 451 285
rect 531 319 565 353
rect 531 251 565 285
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 26 597 92 649
rect 26 563 42 597
rect 76 563 92 597
rect 26 512 92 563
rect 26 478 42 512
rect 76 478 92 512
rect 26 462 92 478
rect 132 597 198 613
rect 132 563 148 597
rect 182 563 198 597
rect 132 526 198 563
rect 132 492 148 526
rect 182 492 198 526
rect 132 455 198 492
rect 238 597 304 649
rect 238 563 254 597
rect 288 563 304 597
rect 238 525 304 563
rect 238 491 254 525
rect 288 491 304 525
rect 238 475 304 491
rect 344 597 410 613
rect 344 563 360 597
rect 394 563 410 597
rect 344 526 410 563
rect 344 492 360 526
rect 394 492 410 526
rect 132 426 148 455
rect 25 421 148 426
rect 182 439 198 455
rect 344 455 410 492
rect 344 439 360 455
rect 182 421 360 439
rect 394 421 410 455
rect 25 405 410 421
rect 450 597 516 649
rect 450 563 466 597
rect 500 563 516 597
rect 450 526 516 563
rect 450 492 466 526
rect 500 492 516 526
rect 450 455 516 492
rect 450 421 466 455
rect 500 421 516 455
rect 450 405 516 421
rect 560 597 651 613
rect 560 563 576 597
rect 610 563 651 597
rect 560 526 651 563
rect 560 492 576 526
rect 610 492 651 526
rect 560 455 651 492
rect 560 421 576 455
rect 610 421 651 455
rect 560 405 651 421
rect 25 392 198 405
rect 25 129 71 392
rect 121 340 251 356
rect 121 306 201 340
rect 235 306 251 340
rect 121 290 251 306
rect 293 353 359 369
rect 293 319 309 353
rect 343 319 359 353
rect 293 285 359 319
rect 293 251 309 285
rect 343 251 359 285
rect 293 235 359 251
rect 401 353 467 369
rect 401 319 417 353
rect 451 319 467 353
rect 401 285 467 319
rect 401 251 417 285
rect 451 251 467 285
rect 401 235 467 251
rect 505 353 581 369
rect 505 319 531 353
rect 565 319 581 353
rect 505 285 581 319
rect 505 251 531 285
rect 565 251 581 285
rect 505 235 581 251
rect 107 215 173 231
rect 107 181 123 215
rect 157 199 173 215
rect 617 199 651 405
rect 157 181 651 199
rect 107 165 651 181
rect 25 108 148 129
rect 25 95 98 108
rect 82 74 98 95
rect 132 74 148 108
rect 82 53 148 74
rect 402 103 468 129
rect 402 69 418 103
rect 452 69 468 103
rect 402 17 468 69
rect 576 111 642 165
rect 576 77 592 111
rect 626 77 642 111
rect 576 53 642 77
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4b_lp
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 782824
string GDS_START 776086
<< end >>
