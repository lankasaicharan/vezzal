magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2218 1852
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 12 21 897 203
rect 24 -17 58 21
<< scnmos >>
rect 121 47 151 177
rect 215 47 245 177
rect 302 47 332 177
rect 507 47 537 177
rect 601 47 631 177
rect 685 47 715 177
rect 789 47 819 177
<< scpmoshvt >>
rect 113 297 149 497
rect 219 297 255 497
rect 304 297 340 497
rect 499 297 535 497
rect 581 297 617 497
rect 687 297 723 497
rect 781 297 817 497
<< ndiff >>
rect 38 157 121 177
rect 38 123 50 157
rect 84 123 121 157
rect 38 89 121 123
rect 38 55 50 89
rect 84 55 121 89
rect 38 47 121 55
rect 151 93 215 177
rect 151 59 161 93
rect 195 59 215 93
rect 151 47 215 59
rect 245 163 302 177
rect 245 129 255 163
rect 289 129 302 163
rect 245 47 302 129
rect 332 93 391 177
rect 332 59 349 93
rect 383 59 391 93
rect 332 47 391 59
rect 445 95 507 177
rect 445 61 453 95
rect 487 61 507 95
rect 445 47 507 61
rect 537 163 601 177
rect 537 129 547 163
rect 581 129 601 163
rect 537 95 601 129
rect 537 61 547 95
rect 581 61 601 95
rect 537 47 601 61
rect 631 163 685 177
rect 631 129 641 163
rect 675 129 685 163
rect 631 95 685 129
rect 631 61 641 95
rect 675 61 685 95
rect 631 47 685 61
rect 715 163 789 177
rect 715 129 735 163
rect 769 129 789 163
rect 715 95 789 129
rect 715 61 735 95
rect 769 61 789 95
rect 715 47 789 61
rect 819 95 871 177
rect 819 61 829 95
rect 863 61 871 95
rect 819 47 871 61
<< pdiff >>
rect 46 477 113 497
rect 46 443 66 477
rect 100 443 113 477
rect 46 409 113 443
rect 46 375 66 409
rect 100 375 113 409
rect 46 341 113 375
rect 46 307 66 341
rect 100 307 113 341
rect 46 297 113 307
rect 149 488 219 497
rect 149 454 168 488
rect 202 454 219 488
rect 149 420 219 454
rect 149 386 168 420
rect 202 386 219 420
rect 149 297 219 386
rect 255 297 304 497
rect 340 477 499 497
rect 340 443 352 477
rect 386 443 453 477
rect 487 443 499 477
rect 340 409 499 443
rect 340 375 352 409
rect 386 375 453 409
rect 487 375 499 409
rect 340 297 499 375
rect 535 297 581 497
rect 617 477 687 497
rect 617 443 629 477
rect 663 443 687 477
rect 617 409 687 443
rect 617 375 629 409
rect 663 375 687 409
rect 617 297 687 375
rect 723 477 781 497
rect 723 443 735 477
rect 769 443 781 477
rect 723 409 781 443
rect 723 375 735 409
rect 769 375 781 409
rect 723 297 781 375
rect 817 477 871 497
rect 817 443 829 477
rect 863 443 871 477
rect 817 297 871 443
<< ndiffc >>
rect 50 123 84 157
rect 50 55 84 89
rect 161 59 195 93
rect 255 129 289 163
rect 349 59 383 93
rect 453 61 487 95
rect 547 129 581 163
rect 547 61 581 95
rect 641 129 675 163
rect 641 61 675 95
rect 735 129 769 163
rect 735 61 769 95
rect 829 61 863 95
<< pdiffc >>
rect 66 443 100 477
rect 66 375 100 409
rect 66 307 100 341
rect 168 454 202 488
rect 168 386 202 420
rect 352 443 386 477
rect 453 443 487 477
rect 352 375 386 409
rect 453 375 487 409
rect 629 443 663 477
rect 629 375 663 409
rect 735 443 769 477
rect 735 375 769 409
rect 829 443 863 477
<< poly >>
rect 113 497 149 523
rect 219 497 255 523
rect 304 497 340 523
rect 499 497 535 523
rect 581 497 617 523
rect 687 497 723 523
rect 781 497 817 523
rect 113 282 149 297
rect 219 282 255 297
rect 304 282 340 297
rect 499 282 535 297
rect 581 282 617 297
rect 687 282 723 297
rect 781 282 817 297
rect 111 265 151 282
rect 217 265 257 282
rect 25 249 151 265
rect 25 215 35 249
rect 69 215 151 249
rect 25 195 151 215
rect 193 249 257 265
rect 193 215 203 249
rect 237 215 257 249
rect 193 199 257 215
rect 302 265 342 282
rect 497 265 537 282
rect 302 249 375 265
rect 302 215 321 249
rect 355 215 375 249
rect 302 199 375 215
rect 453 249 537 265
rect 453 215 463 249
rect 497 215 537 249
rect 453 199 537 215
rect 579 265 619 282
rect 685 265 725 282
rect 779 265 819 282
rect 579 249 643 265
rect 579 215 589 249
rect 623 215 643 249
rect 579 199 643 215
rect 685 249 819 265
rect 685 215 725 249
rect 759 215 819 249
rect 685 199 819 215
rect 121 177 151 195
rect 215 177 245 199
rect 302 177 332 199
rect 507 177 537 199
rect 601 177 631 199
rect 685 177 715 199
rect 789 177 819 199
rect 121 21 151 47
rect 215 21 245 47
rect 302 21 332 47
rect 507 21 537 47
rect 601 21 631 47
rect 685 21 715 47
rect 789 21 819 47
<< polycont >>
rect 35 215 69 249
rect 203 215 237 249
rect 321 215 355 249
rect 463 215 497 249
rect 589 215 623 249
rect 725 215 759 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 50 477 116 493
rect 50 443 66 477
rect 100 443 116 477
rect 50 409 116 443
rect 50 375 66 409
rect 100 375 116 409
rect 50 341 116 375
rect 160 488 202 527
rect 160 454 168 488
rect 160 420 202 454
rect 160 386 168 420
rect 340 477 491 493
rect 340 443 352 477
rect 386 443 453 477
rect 487 443 491 477
rect 340 409 491 443
rect 629 477 675 527
rect 663 443 675 477
rect 629 409 675 443
rect 160 370 202 386
rect 236 375 352 409
rect 386 375 453 409
rect 487 375 593 409
rect 50 307 66 341
rect 100 334 116 341
rect 236 334 270 375
rect 100 307 270 334
rect 50 299 270 307
rect 109 289 270 299
rect 17 249 69 265
rect 17 215 35 249
rect 17 195 69 215
rect 109 161 153 289
rect 187 249 266 255
rect 187 215 203 249
rect 237 215 266 249
rect 304 249 381 341
rect 304 215 321 249
rect 355 215 381 249
rect 447 249 523 341
rect 559 325 593 375
rect 663 375 675 409
rect 709 477 769 493
rect 709 443 735 477
rect 803 477 881 527
rect 803 443 829 477
rect 863 443 881 477
rect 709 409 769 443
rect 709 375 735 409
rect 769 375 898 409
rect 629 359 675 375
rect 559 291 743 325
rect 699 257 743 291
rect 447 215 463 249
rect 497 215 523 249
rect 567 249 665 257
rect 567 215 589 249
rect 623 215 665 249
rect 699 249 775 257
rect 699 215 725 249
rect 759 215 775 249
rect 836 181 898 375
rect 34 157 153 161
rect 34 123 50 157
rect 84 127 153 157
rect 227 163 597 181
rect 227 129 255 163
rect 289 147 547 163
rect 289 129 314 147
rect 521 129 547 147
rect 581 129 597 163
rect 84 123 100 127
rect 34 89 100 123
rect 453 95 487 111
rect 34 55 50 89
rect 84 55 100 89
rect 134 59 161 93
rect 195 59 349 93
rect 383 59 401 93
rect 34 51 100 55
rect 453 17 487 61
rect 521 95 597 129
rect 521 61 547 95
rect 581 61 597 95
rect 521 54 597 61
rect 641 163 675 181
rect 641 95 675 129
rect 641 17 675 61
rect 709 163 898 181
rect 709 129 735 163
rect 769 147 898 163
rect 769 129 785 147
rect 709 95 785 129
rect 709 61 735 95
rect 769 61 785 95
rect 709 53 785 61
rect 829 95 863 113
rect 829 17 863 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 320 292 364 326 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 447 215 523 341 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 485 238 485 238 0 FreeSans 400 0 0 0 A2
port 2 nsew
flabel locali s 851 357 885 391 0 FreeSans 400 0 0 0 X
port 10 nsew signal output
flabel locali s 218 221 252 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 24 221 58 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 567 215 665 257 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 313 221 357 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel nwell s 28 527 62 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 24 -17 58 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 24 -17 58 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional
flabel metal1 s 28 527 62 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o221a_2
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2491968
string GDS_START 2484146
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
