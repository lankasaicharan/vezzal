magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1288 -1260 1704 2245
use sky130_fd_pr__hvdfm1sd2__example_5595914180829  sky130_fd_pr__hvdfm1sd2__example_5595914180829_0
timestamp 1627201311
transform 1 0 180 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808237  sky130_fd_pr__hvdfm1sd__example_55959141808237_0
timestamp 1627201311
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808237  sky130_fd_pr__hvdfm1sd__example_55959141808237_1
timestamp 1627201311
transform 1 0 416 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 444 985 444 985 0 FreeSans 300 0 0 0 S
flabel comment s 208 985 208 985 0 FreeSans 300 0 0 0 D
flabel comment s -28 985 -28 985 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 37245772
string GDS_START 37244266
<< end >>
