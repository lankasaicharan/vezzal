magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 1 49 634 241
rect 0 0 672 49
<< scnmos >>
rect 80 47 110 215
rect 169 47 199 215
rect 267 47 297 215
rect 353 47 383 215
rect 439 47 469 215
rect 525 47 555 215
<< scpmoshvt >>
rect 80 367 110 619
rect 152 367 182 619
rect 267 367 297 619
rect 353 367 383 619
rect 439 367 469 619
rect 525 367 555 619
<< ndiff >>
rect 27 203 80 215
rect 27 169 35 203
rect 69 169 80 203
rect 27 93 80 169
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 203 169 215
rect 110 169 124 203
rect 158 169 169 203
rect 110 101 169 169
rect 110 67 124 101
rect 158 67 169 101
rect 110 47 169 67
rect 199 163 267 215
rect 199 129 216 163
rect 250 129 267 163
rect 199 89 267 129
rect 199 55 216 89
rect 250 55 267 89
rect 199 47 267 55
rect 297 203 353 215
rect 297 169 308 203
rect 342 169 353 203
rect 297 101 353 169
rect 297 67 308 101
rect 342 67 353 101
rect 297 47 353 67
rect 383 179 439 215
rect 383 145 394 179
rect 428 145 439 179
rect 383 93 439 145
rect 383 59 394 93
rect 428 59 439 93
rect 383 47 439 59
rect 469 203 525 215
rect 469 169 480 203
rect 514 169 525 203
rect 469 101 525 169
rect 469 67 480 101
rect 514 67 525 101
rect 469 47 525 67
rect 555 179 608 215
rect 555 145 566 179
rect 600 145 608 179
rect 555 93 608 145
rect 555 59 566 93
rect 600 59 608 93
rect 555 47 608 59
<< pdiff >>
rect 27 607 80 619
rect 27 573 35 607
rect 69 573 80 607
rect 27 513 80 573
rect 27 479 35 513
rect 69 479 80 513
rect 27 423 80 479
rect 27 389 35 423
rect 69 389 80 423
rect 27 367 80 389
rect 110 367 152 619
rect 182 607 267 619
rect 182 573 208 607
rect 242 573 267 607
rect 182 493 267 573
rect 182 459 208 493
rect 242 459 267 493
rect 182 367 267 459
rect 297 599 353 619
rect 297 565 308 599
rect 342 565 353 599
rect 297 509 353 565
rect 297 475 308 509
rect 342 475 353 509
rect 297 413 353 475
rect 297 379 308 413
rect 342 379 353 413
rect 297 367 353 379
rect 383 611 439 619
rect 383 577 394 611
rect 428 577 439 611
rect 383 537 439 577
rect 383 503 394 537
rect 428 503 439 537
rect 383 457 439 503
rect 383 423 394 457
rect 428 423 439 457
rect 383 367 439 423
rect 469 599 525 619
rect 469 565 480 599
rect 514 565 525 599
rect 469 509 525 565
rect 469 475 480 509
rect 514 475 525 509
rect 469 413 525 475
rect 469 379 480 413
rect 514 379 525 413
rect 469 367 525 379
rect 555 607 608 619
rect 555 573 566 607
rect 600 573 608 607
rect 555 534 608 573
rect 555 500 566 534
rect 600 500 608 534
rect 555 457 608 500
rect 555 423 566 457
rect 600 423 608 457
rect 555 367 608 423
<< ndiffc >>
rect 35 169 69 203
rect 35 59 69 93
rect 124 169 158 203
rect 124 67 158 101
rect 216 129 250 163
rect 216 55 250 89
rect 308 169 342 203
rect 308 67 342 101
rect 394 145 428 179
rect 394 59 428 93
rect 480 169 514 203
rect 480 67 514 101
rect 566 145 600 179
rect 566 59 600 93
<< pdiffc >>
rect 35 573 69 607
rect 35 479 69 513
rect 35 389 69 423
rect 208 573 242 607
rect 208 459 242 493
rect 308 565 342 599
rect 308 475 342 509
rect 308 379 342 413
rect 394 577 428 611
rect 394 503 428 537
rect 394 423 428 457
rect 480 565 514 599
rect 480 475 514 509
rect 480 379 514 413
rect 566 573 600 607
rect 566 500 600 534
rect 566 423 600 457
<< poly >>
rect 80 619 110 645
rect 152 619 182 645
rect 267 619 297 645
rect 353 619 383 645
rect 439 619 469 645
rect 525 619 555 645
rect 80 345 110 367
rect 38 315 110 345
rect 152 335 182 367
rect 152 319 218 335
rect 38 292 104 315
rect 38 258 54 292
rect 88 267 104 292
rect 152 285 168 319
rect 202 285 218 319
rect 152 269 218 285
rect 267 333 297 367
rect 353 333 383 367
rect 439 333 469 367
rect 525 333 555 367
rect 267 317 555 333
rect 267 283 283 317
rect 317 283 351 317
rect 385 283 419 317
rect 453 283 487 317
rect 521 283 555 317
rect 88 258 110 267
rect 38 237 110 258
rect 80 215 110 237
rect 169 215 199 269
rect 267 267 555 283
rect 267 215 297 267
rect 353 215 383 267
rect 439 215 469 267
rect 525 215 555 267
rect 80 21 110 47
rect 169 21 199 47
rect 267 21 297 47
rect 353 21 383 47
rect 439 21 469 47
rect 525 21 555 47
<< polycont >>
rect 54 258 88 292
rect 168 285 202 319
rect 283 283 317 317
rect 351 283 385 317
rect 419 283 453 317
rect 487 283 521 317
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 19 607 85 615
rect 19 573 35 607
rect 69 573 85 607
rect 19 513 85 573
rect 19 479 35 513
rect 69 479 85 513
rect 19 423 85 479
rect 192 607 258 649
rect 192 573 208 607
rect 242 573 258 607
rect 192 493 258 573
rect 192 459 208 493
rect 242 459 258 493
rect 192 454 258 459
rect 308 599 344 615
rect 342 565 344 599
rect 308 509 344 565
rect 342 475 344 509
rect 19 389 35 423
rect 69 420 85 423
rect 69 389 272 420
rect 19 386 272 389
rect 17 292 88 352
rect 17 258 54 292
rect 122 319 204 351
rect 122 285 168 319
rect 202 285 204 319
rect 122 269 204 285
rect 238 317 272 386
rect 308 413 344 475
rect 378 611 444 649
rect 378 577 394 611
rect 428 577 444 611
rect 378 537 444 577
rect 378 503 394 537
rect 428 503 444 537
rect 378 457 444 503
rect 378 423 394 457
rect 428 423 444 457
rect 478 599 516 615
rect 478 565 480 599
rect 514 565 516 599
rect 478 509 516 565
rect 478 475 480 509
rect 514 475 516 509
rect 342 389 344 413
rect 478 413 516 475
rect 550 607 616 649
rect 550 573 566 607
rect 600 573 616 607
rect 550 534 616 573
rect 550 500 566 534
rect 600 500 616 534
rect 550 457 616 500
rect 550 423 566 457
rect 600 423 616 457
rect 478 389 480 413
rect 342 379 480 389
rect 514 389 516 413
rect 514 379 655 389
rect 308 351 655 379
rect 238 283 283 317
rect 317 283 351 317
rect 385 283 419 317
rect 453 283 487 317
rect 521 283 537 317
rect 17 242 88 258
rect 238 235 272 283
rect 571 249 655 351
rect 19 203 85 208
rect 19 169 35 203
rect 69 169 85 203
rect 19 93 85 169
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 122 203 272 235
rect 122 169 124 203
rect 158 197 272 203
rect 306 213 655 249
rect 306 203 344 213
rect 158 169 166 197
rect 122 101 166 169
rect 306 169 308 203
rect 342 169 344 203
rect 478 203 516 213
rect 122 67 124 101
rect 158 67 166 101
rect 122 51 166 67
rect 200 129 216 163
rect 250 129 266 163
rect 200 89 266 129
rect 200 55 216 89
rect 250 55 266 89
rect 200 17 266 55
rect 306 101 344 169
rect 306 67 308 101
rect 342 67 344 101
rect 306 51 344 67
rect 378 145 394 179
rect 428 145 444 179
rect 378 93 444 145
rect 378 59 394 93
rect 428 59 444 93
rect 378 17 444 59
rect 478 169 480 203
rect 514 169 516 203
rect 478 101 516 169
rect 478 67 480 101
rect 514 67 516 101
rect 478 51 516 67
rect 550 145 566 179
rect 600 145 616 179
rect 550 93 616 145
rect 550 59 566 93
rect 600 59 616 93
rect 550 17 616 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or2_4
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 6148630
string GDS_START 6142052
<< end >>
