magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 332 806 704
<< pwell >>
rect 254 281 356 290
rect 254 248 451 281
rect 2 49 756 248
rect 0 0 768 49
<< scpmos >>
rect 186 368 216 592
rect 276 368 306 592
rect 366 368 396 592
rect 468 368 498 592
rect 558 368 588 592
rect 648 368 678 592
<< nmoslvt >>
rect 81 74 111 222
rect 345 107 375 255
rect 475 74 505 222
rect 561 74 591 222
rect 647 74 677 222
<< ndiff >>
rect 280 255 330 264
rect 280 252 345 255
rect 28 210 81 222
rect 28 176 36 210
rect 70 176 81 210
rect 28 120 81 176
rect 28 86 36 120
rect 70 86 81 120
rect 28 74 81 86
rect 111 210 164 222
rect 111 176 122 210
rect 156 176 164 210
rect 111 120 164 176
rect 111 86 122 120
rect 156 86 164 120
rect 280 218 288 252
rect 322 218 345 252
rect 280 107 345 218
rect 375 222 425 255
rect 375 116 475 222
rect 375 107 416 116
rect 111 74 164 86
rect 404 82 416 107
rect 450 82 475 116
rect 404 74 475 82
rect 505 116 561 222
rect 505 82 516 116
rect 550 82 561 116
rect 505 74 561 82
rect 591 205 647 222
rect 591 171 602 205
rect 636 171 647 205
rect 591 74 647 171
rect 677 210 730 222
rect 677 176 688 210
rect 722 176 730 210
rect 677 120 730 176
rect 677 86 688 120
rect 722 86 730 120
rect 677 74 730 86
<< pdiff >>
rect 131 580 186 592
rect 131 546 139 580
rect 173 546 186 580
rect 131 510 186 546
rect 131 476 139 510
rect 173 476 186 510
rect 131 440 186 476
rect 131 406 139 440
rect 173 406 186 440
rect 131 368 186 406
rect 216 547 276 592
rect 216 513 229 547
rect 263 513 276 547
rect 216 479 276 513
rect 216 445 229 479
rect 263 445 276 479
rect 216 411 276 445
rect 216 377 229 411
rect 263 377 276 411
rect 216 368 276 377
rect 306 580 366 592
rect 306 546 319 580
rect 353 546 366 580
rect 306 508 366 546
rect 306 474 319 508
rect 353 474 366 508
rect 306 368 366 474
rect 396 578 468 592
rect 396 544 410 578
rect 444 544 468 578
rect 396 368 468 544
rect 498 580 558 592
rect 498 546 511 580
rect 545 546 558 580
rect 498 508 558 546
rect 498 474 511 508
rect 545 474 558 508
rect 498 368 558 474
rect 588 578 648 592
rect 588 544 601 578
rect 635 544 648 578
rect 588 368 648 544
rect 678 580 733 592
rect 678 546 691 580
rect 725 546 733 580
rect 678 508 733 546
rect 678 474 691 508
rect 725 474 733 508
rect 678 368 733 474
<< ndiffc >>
rect 36 176 70 210
rect 36 86 70 120
rect 122 176 156 210
rect 122 86 156 120
rect 288 218 322 252
rect 416 82 450 116
rect 516 82 550 116
rect 602 171 636 205
rect 688 176 722 210
rect 688 86 722 120
<< pdiffc >>
rect 139 546 173 580
rect 139 476 173 510
rect 139 406 173 440
rect 229 513 263 547
rect 229 445 263 479
rect 229 377 263 411
rect 319 546 353 580
rect 319 474 353 508
rect 410 544 444 578
rect 511 546 545 580
rect 511 474 545 508
rect 601 544 635 578
rect 691 546 725 580
rect 691 474 725 508
<< poly >>
rect 186 592 216 618
rect 276 592 306 618
rect 366 592 396 618
rect 468 592 498 618
rect 558 592 588 618
rect 648 592 678 618
rect 186 353 216 368
rect 276 353 306 368
rect 366 353 396 368
rect 468 353 498 368
rect 558 353 588 368
rect 648 353 678 368
rect 21 337 309 353
rect 21 303 37 337
rect 71 323 309 337
rect 363 336 399 353
rect 465 336 501 353
rect 555 336 591 353
rect 645 336 681 353
rect 71 303 111 323
rect 21 287 111 303
rect 363 320 513 336
rect 363 300 463 320
rect 81 222 111 287
rect 345 286 463 300
rect 497 286 513 320
rect 345 270 513 286
rect 555 320 681 336
rect 555 286 620 320
rect 654 286 681 320
rect 555 270 681 286
rect 345 255 375 270
rect 475 222 505 270
rect 561 222 591 270
rect 647 222 677 270
rect 345 81 375 107
rect 81 48 111 74
rect 475 48 505 74
rect 561 48 591 74
rect 647 48 677 74
<< polycont >>
rect 37 303 71 337
rect 463 286 497 320
rect 620 286 654 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 123 581 369 615
rect 123 580 179 581
rect 123 546 139 580
rect 173 546 179 580
rect 313 580 369 581
rect 123 510 179 546
rect 123 476 139 510
rect 173 476 179 510
rect 123 440 179 476
rect 123 406 139 440
rect 173 406 179 440
rect 123 390 179 406
rect 213 513 229 547
rect 263 513 279 547
rect 213 479 279 513
rect 213 445 229 479
rect 263 445 279 479
rect 313 546 319 580
rect 353 546 369 580
rect 313 508 369 546
rect 409 578 461 649
rect 409 544 410 578
rect 444 544 461 578
rect 409 526 461 544
rect 495 580 561 596
rect 495 546 511 580
rect 545 546 561 580
rect 313 474 319 508
rect 353 492 369 508
rect 495 508 561 546
rect 601 578 635 649
rect 601 526 635 544
rect 675 580 741 596
rect 675 546 691 580
rect 725 546 741 580
rect 495 492 511 508
rect 353 474 511 492
rect 545 492 561 508
rect 675 508 741 546
rect 675 492 691 508
rect 545 474 691 492
rect 725 474 741 508
rect 313 458 741 474
rect 213 411 279 445
rect 213 377 229 411
rect 263 377 279 411
rect 213 356 279 377
rect 21 337 87 356
rect 21 303 37 337
rect 71 303 87 337
rect 21 287 87 303
rect 121 310 279 356
rect 313 390 738 424
rect 20 210 86 226
rect 20 176 36 210
rect 70 176 86 210
rect 20 120 86 176
rect 20 86 36 120
rect 70 86 86 120
rect 20 17 86 86
rect 121 210 172 310
rect 313 252 355 390
rect 272 218 288 252
rect 322 218 355 252
rect 409 320 551 356
rect 409 286 463 320
rect 497 286 551 320
rect 409 236 551 286
rect 601 320 670 356
rect 601 286 620 320
rect 654 286 670 320
rect 601 270 670 286
rect 704 226 738 390
rect 121 176 122 210
rect 156 184 172 210
rect 586 205 636 226
rect 586 184 602 205
rect 156 176 602 184
rect 121 171 602 176
rect 121 150 636 171
rect 672 210 738 226
rect 672 176 688 210
rect 722 176 738 210
rect 121 120 172 150
rect 121 86 122 120
rect 156 86 172 120
rect 672 120 738 176
rect 672 116 688 120
rect 121 70 172 86
rect 400 82 416 116
rect 450 82 466 116
rect 400 17 466 82
rect 500 82 516 116
rect 550 86 688 116
rect 722 86 738 120
rect 550 82 738 86
rect 500 66 738 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a21oi_2
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 2542230
string GDS_START 2535304
<< end >>
