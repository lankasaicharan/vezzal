magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2546 1975
<< nwell >>
rect -38 331 1286 704
<< pwell >>
rect 3 49 1247 243
rect 0 0 1248 49
<< scnmos >>
rect 82 49 112 217
rect 168 49 198 217
rect 254 49 284 217
rect 340 49 370 217
rect 426 49 456 217
rect 512 49 542 217
rect 598 49 628 217
rect 684 49 714 217
rect 876 49 906 217
rect 962 49 992 217
rect 1048 49 1078 217
rect 1134 49 1164 217
<< scpmoshvt >>
rect 82 367 112 619
rect 168 367 198 619
rect 254 367 284 619
rect 340 367 370 619
rect 426 367 456 619
rect 512 367 542 619
rect 598 367 628 619
rect 684 367 714 619
rect 876 367 906 619
rect 962 367 992 619
rect 1048 367 1078 619
rect 1134 367 1164 619
<< ndiff >>
rect 29 182 82 217
rect 29 148 37 182
rect 71 148 82 182
rect 29 114 82 148
rect 29 80 37 114
rect 71 80 82 114
rect 29 49 82 80
rect 112 187 168 217
rect 112 153 123 187
rect 157 153 168 187
rect 112 113 168 153
rect 112 79 123 113
rect 157 79 168 113
rect 112 49 168 79
rect 198 159 254 217
rect 198 125 209 159
rect 243 125 254 159
rect 198 91 254 125
rect 198 57 209 91
rect 243 57 254 91
rect 198 49 254 57
rect 284 187 340 217
rect 284 153 295 187
rect 329 153 340 187
rect 284 113 340 153
rect 284 79 295 113
rect 329 79 340 113
rect 284 49 340 79
rect 370 159 426 217
rect 370 125 381 159
rect 415 125 426 159
rect 370 91 426 125
rect 370 57 381 91
rect 415 57 426 91
rect 370 49 426 57
rect 456 187 512 217
rect 456 153 467 187
rect 501 153 512 187
rect 456 113 512 153
rect 456 79 467 113
rect 501 79 512 113
rect 456 49 512 79
rect 542 159 598 217
rect 542 125 553 159
rect 587 125 598 159
rect 542 91 598 125
rect 542 57 553 91
rect 587 57 598 91
rect 542 49 598 57
rect 628 187 684 217
rect 628 153 639 187
rect 673 153 684 187
rect 628 113 684 153
rect 628 79 639 113
rect 673 79 684 113
rect 628 49 684 79
rect 714 187 767 217
rect 714 153 725 187
rect 759 153 767 187
rect 714 113 767 153
rect 714 79 725 113
rect 759 79 767 113
rect 714 49 767 79
rect 821 187 876 217
rect 821 153 829 187
rect 863 153 876 187
rect 821 113 876 153
rect 821 79 829 113
rect 863 79 876 113
rect 821 49 876 79
rect 906 169 962 217
rect 906 135 917 169
rect 951 135 962 169
rect 906 101 962 135
rect 906 67 917 101
rect 951 67 962 101
rect 906 49 962 67
rect 992 187 1048 217
rect 992 153 1003 187
rect 1037 153 1048 187
rect 992 113 1048 153
rect 992 79 1003 113
rect 1037 79 1048 113
rect 992 49 1048 79
rect 1078 124 1134 217
rect 1078 90 1089 124
rect 1123 90 1134 124
rect 1078 49 1134 90
rect 1164 187 1221 217
rect 1164 153 1179 187
rect 1213 153 1221 187
rect 1164 113 1221 153
rect 1164 79 1179 113
rect 1213 79 1221 113
rect 1164 49 1221 79
<< pdiff >>
rect 29 605 82 619
rect 29 571 37 605
rect 71 571 82 605
rect 29 537 82 571
rect 29 503 37 537
rect 71 503 82 537
rect 29 469 82 503
rect 29 435 37 469
rect 71 435 82 469
rect 29 367 82 435
rect 112 585 168 619
rect 112 551 123 585
rect 157 551 168 585
rect 112 506 168 551
rect 112 472 123 506
rect 157 472 168 506
rect 112 427 168 472
rect 112 393 123 427
rect 157 393 168 427
rect 112 367 168 393
rect 198 605 254 619
rect 198 571 209 605
rect 243 571 254 605
rect 198 537 254 571
rect 198 503 209 537
rect 243 503 254 537
rect 198 469 254 503
rect 198 435 209 469
rect 243 435 254 469
rect 198 367 254 435
rect 284 585 340 619
rect 284 551 295 585
rect 329 551 340 585
rect 284 506 340 551
rect 284 472 295 506
rect 329 472 340 506
rect 284 427 340 472
rect 284 393 295 427
rect 329 393 340 427
rect 284 367 340 393
rect 370 605 426 619
rect 370 571 381 605
rect 415 571 426 605
rect 370 537 426 571
rect 370 503 381 537
rect 415 503 426 537
rect 370 469 426 503
rect 370 435 381 469
rect 415 435 426 469
rect 370 367 426 435
rect 456 585 512 619
rect 456 551 467 585
rect 501 551 512 585
rect 456 506 512 551
rect 456 472 467 506
rect 501 472 512 506
rect 456 427 512 472
rect 456 393 467 427
rect 501 393 512 427
rect 456 367 512 393
rect 542 605 598 619
rect 542 571 553 605
rect 587 571 598 605
rect 542 537 598 571
rect 542 503 553 537
rect 587 503 598 537
rect 542 469 598 503
rect 542 435 553 469
rect 587 435 598 469
rect 542 367 598 435
rect 628 585 684 619
rect 628 551 639 585
rect 673 551 684 585
rect 628 506 684 551
rect 628 472 639 506
rect 673 472 684 506
rect 628 427 684 472
rect 628 393 639 427
rect 673 393 684 427
rect 628 367 684 393
rect 714 585 767 619
rect 714 551 725 585
rect 759 551 767 585
rect 714 506 767 551
rect 714 472 725 506
rect 759 472 767 506
rect 714 427 767 472
rect 714 393 725 427
rect 759 393 767 427
rect 714 367 767 393
rect 823 585 876 619
rect 823 551 831 585
rect 865 551 876 585
rect 823 506 876 551
rect 823 472 831 506
rect 865 472 876 506
rect 823 427 876 472
rect 823 393 831 427
rect 865 393 876 427
rect 823 367 876 393
rect 906 605 962 619
rect 906 571 917 605
rect 951 571 962 605
rect 906 537 962 571
rect 906 503 917 537
rect 951 503 962 537
rect 906 469 962 503
rect 906 435 917 469
rect 951 435 962 469
rect 906 367 962 435
rect 992 585 1048 619
rect 992 551 1003 585
rect 1037 551 1048 585
rect 992 506 1048 551
rect 992 472 1003 506
rect 1037 472 1048 506
rect 992 427 1048 472
rect 992 393 1003 427
rect 1037 393 1048 427
rect 992 367 1048 393
rect 1078 575 1134 619
rect 1078 541 1089 575
rect 1123 541 1134 575
rect 1078 504 1134 541
rect 1078 470 1089 504
rect 1123 470 1134 504
rect 1078 367 1134 470
rect 1164 580 1217 619
rect 1164 546 1175 580
rect 1209 546 1217 580
rect 1164 512 1217 546
rect 1164 478 1175 512
rect 1209 478 1217 512
rect 1164 444 1217 478
rect 1164 410 1175 444
rect 1209 410 1217 444
rect 1164 367 1217 410
<< ndiffc >>
rect 37 148 71 182
rect 37 80 71 114
rect 123 153 157 187
rect 123 79 157 113
rect 209 125 243 159
rect 209 57 243 91
rect 295 153 329 187
rect 295 79 329 113
rect 381 125 415 159
rect 381 57 415 91
rect 467 153 501 187
rect 467 79 501 113
rect 553 125 587 159
rect 553 57 587 91
rect 639 153 673 187
rect 639 79 673 113
rect 725 153 759 187
rect 725 79 759 113
rect 829 153 863 187
rect 829 79 863 113
rect 917 135 951 169
rect 917 67 951 101
rect 1003 153 1037 187
rect 1003 79 1037 113
rect 1089 90 1123 124
rect 1179 153 1213 187
rect 1179 79 1213 113
<< pdiffc >>
rect 37 571 71 605
rect 37 503 71 537
rect 37 435 71 469
rect 123 551 157 585
rect 123 472 157 506
rect 123 393 157 427
rect 209 571 243 605
rect 209 503 243 537
rect 209 435 243 469
rect 295 551 329 585
rect 295 472 329 506
rect 295 393 329 427
rect 381 571 415 605
rect 381 503 415 537
rect 381 435 415 469
rect 467 551 501 585
rect 467 472 501 506
rect 467 393 501 427
rect 553 571 587 605
rect 553 503 587 537
rect 553 435 587 469
rect 639 551 673 585
rect 639 472 673 506
rect 639 393 673 427
rect 725 551 759 585
rect 725 472 759 506
rect 725 393 759 427
rect 831 551 865 585
rect 831 472 865 506
rect 831 393 865 427
rect 917 571 951 605
rect 917 503 951 537
rect 917 435 951 469
rect 1003 551 1037 585
rect 1003 472 1037 506
rect 1003 393 1037 427
rect 1089 541 1123 575
rect 1089 470 1123 504
rect 1175 546 1209 580
rect 1175 478 1209 512
rect 1175 410 1209 444
<< poly >>
rect 82 619 112 645
rect 168 619 198 645
rect 254 619 284 645
rect 340 619 370 645
rect 426 619 456 645
rect 512 619 542 645
rect 598 619 628 645
rect 684 619 714 645
rect 876 619 906 645
rect 962 619 992 645
rect 1048 619 1078 645
rect 1134 619 1164 645
rect 82 331 112 367
rect 168 331 198 367
rect 254 331 284 367
rect 340 331 370 367
rect 426 331 456 367
rect 512 331 542 367
rect 598 331 628 367
rect 684 331 714 367
rect 876 331 906 367
rect 962 331 992 367
rect 1048 331 1078 367
rect 82 315 807 331
rect 82 281 213 315
rect 247 281 281 315
rect 315 281 349 315
rect 383 281 417 315
rect 451 281 485 315
rect 519 281 553 315
rect 587 281 621 315
rect 655 281 689 315
rect 723 281 757 315
rect 791 281 807 315
rect 82 265 807 281
rect 876 315 1078 331
rect 876 281 892 315
rect 926 281 960 315
rect 994 281 1028 315
rect 1062 281 1078 315
rect 876 265 1078 281
rect 82 217 112 265
rect 168 217 198 265
rect 254 217 284 265
rect 340 217 370 265
rect 426 217 456 265
rect 512 217 542 265
rect 598 217 628 265
rect 684 217 714 265
rect 876 217 906 265
rect 962 217 992 265
rect 1048 217 1078 265
rect 1134 308 1164 367
rect 1134 292 1200 308
rect 1134 258 1150 292
rect 1184 258 1200 292
rect 1134 242 1200 258
rect 1134 217 1164 242
rect 82 23 112 49
rect 168 23 198 49
rect 254 23 284 49
rect 340 23 370 49
rect 426 23 456 49
rect 512 23 542 49
rect 598 23 628 49
rect 684 23 714 49
rect 876 23 906 49
rect 962 23 992 49
rect 1048 23 1078 49
rect 1134 23 1164 49
<< polycont >>
rect 213 281 247 315
rect 281 281 315 315
rect 349 281 383 315
rect 417 281 451 315
rect 485 281 519 315
rect 553 281 587 315
rect 621 281 655 315
rect 689 281 723 315
rect 757 281 791 315
rect 892 281 926 315
rect 960 281 994 315
rect 1028 281 1062 315
rect 1150 258 1184 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 21 605 80 649
rect 21 571 37 605
rect 71 571 80 605
rect 21 537 80 571
rect 21 503 37 537
rect 71 503 80 537
rect 21 469 80 503
rect 21 435 37 469
rect 71 435 80 469
rect 21 419 80 435
rect 114 585 166 611
rect 114 551 123 585
rect 157 551 166 585
rect 114 506 166 551
rect 114 472 123 506
rect 157 472 166 506
rect 114 427 166 472
rect 114 393 123 427
rect 157 393 166 427
rect 200 605 252 649
rect 200 571 209 605
rect 243 571 252 605
rect 200 537 252 571
rect 200 503 209 537
rect 243 503 252 537
rect 200 469 252 503
rect 200 435 209 469
rect 243 435 252 469
rect 200 419 252 435
rect 286 585 338 611
rect 286 551 295 585
rect 329 551 338 585
rect 286 506 338 551
rect 286 472 295 506
rect 329 472 338 506
rect 286 427 338 472
rect 114 385 166 393
rect 286 393 295 427
rect 329 393 338 427
rect 372 605 424 649
rect 372 571 381 605
rect 415 571 424 605
rect 372 537 424 571
rect 372 503 381 537
rect 415 503 424 537
rect 372 469 424 503
rect 372 435 381 469
rect 415 435 424 469
rect 372 419 424 435
rect 458 585 510 611
rect 458 551 467 585
rect 501 551 510 585
rect 458 506 510 551
rect 458 472 467 506
rect 501 472 510 506
rect 458 427 510 472
rect 286 385 338 393
rect 458 393 467 427
rect 501 393 510 427
rect 544 605 596 649
rect 544 571 553 605
rect 587 571 596 605
rect 544 537 596 571
rect 544 503 553 537
rect 587 503 596 537
rect 544 469 596 503
rect 544 435 553 469
rect 587 435 596 469
rect 544 419 596 435
rect 630 585 682 611
rect 630 551 639 585
rect 673 551 682 585
rect 630 506 682 551
rect 630 472 639 506
rect 673 472 682 506
rect 630 427 682 472
rect 458 385 510 393
rect 630 393 639 427
rect 673 393 682 427
rect 630 385 682 393
rect 19 351 682 385
rect 716 585 774 649
rect 716 551 725 585
rect 759 551 774 585
rect 716 506 774 551
rect 716 472 725 506
rect 759 472 774 506
rect 716 427 774 472
rect 716 393 725 427
rect 759 393 774 427
rect 716 368 774 393
rect 808 585 875 611
rect 808 551 831 585
rect 865 551 875 585
rect 808 506 875 551
rect 808 472 831 506
rect 865 472 875 506
rect 808 427 875 472
rect 808 393 831 427
rect 865 393 875 427
rect 909 605 960 649
rect 909 571 917 605
rect 951 571 960 605
rect 909 537 960 571
rect 909 503 917 537
rect 951 503 960 537
rect 909 469 960 503
rect 909 435 917 469
rect 951 435 960 469
rect 909 419 960 435
rect 994 585 1039 611
rect 994 551 1003 585
rect 1037 551 1039 585
rect 994 506 1039 551
rect 994 472 1003 506
rect 1037 472 1039 506
rect 994 427 1039 472
rect 1073 575 1139 649
rect 1073 541 1089 575
rect 1123 541 1139 575
rect 1073 504 1139 541
rect 1073 470 1089 504
rect 1123 470 1139 504
rect 1073 462 1139 470
rect 1173 580 1225 611
rect 1173 546 1175 580
rect 1209 546 1225 580
rect 1173 512 1225 546
rect 1173 478 1175 512
rect 1209 478 1225 512
rect 1173 444 1225 478
rect 1173 428 1175 444
rect 808 385 875 393
rect 994 393 1003 427
rect 1037 393 1039 427
rect 994 385 1039 393
rect 808 351 1039 385
rect 1077 410 1175 428
rect 1209 410 1225 444
rect 1077 394 1225 410
rect 19 245 163 351
rect 808 317 842 351
rect 1077 317 1111 394
rect 197 315 842 317
rect 197 281 213 315
rect 247 281 281 315
rect 315 281 349 315
rect 383 281 417 315
rect 451 281 485 315
rect 519 281 553 315
rect 587 281 621 315
rect 655 281 689 315
rect 723 281 757 315
rect 791 281 842 315
rect 197 279 842 281
rect 876 315 1111 317
rect 876 281 892 315
rect 926 281 960 315
rect 994 281 1028 315
rect 1062 281 1111 315
rect 876 279 1111 281
rect 806 245 842 279
rect 19 232 682 245
rect 114 211 682 232
rect 21 182 80 198
rect 21 148 37 182
rect 71 148 80 182
rect 21 114 80 148
rect 21 80 37 114
rect 71 80 80 114
rect 21 17 80 80
rect 114 187 166 211
rect 114 153 123 187
rect 157 153 166 187
rect 286 187 338 211
rect 114 113 166 153
rect 114 79 123 113
rect 157 79 166 113
rect 114 51 166 79
rect 200 159 252 177
rect 200 125 209 159
rect 243 125 252 159
rect 200 91 252 125
rect 200 57 209 91
rect 243 57 252 91
rect 200 17 252 57
rect 286 153 295 187
rect 329 153 338 187
rect 458 187 510 211
rect 286 113 338 153
rect 286 79 295 113
rect 329 79 338 113
rect 286 51 338 79
rect 372 159 424 177
rect 372 125 381 159
rect 415 125 424 159
rect 372 91 424 125
rect 372 57 381 91
rect 415 57 424 91
rect 372 17 424 57
rect 458 153 467 187
rect 501 153 510 187
rect 630 187 682 211
rect 458 113 510 153
rect 458 79 467 113
rect 501 79 510 113
rect 458 51 510 79
rect 544 159 596 177
rect 544 125 553 159
rect 587 125 596 159
rect 544 91 596 125
rect 544 57 553 91
rect 587 57 596 91
rect 544 17 596 57
rect 630 153 639 187
rect 673 153 682 187
rect 630 113 682 153
rect 630 79 639 113
rect 673 79 682 113
rect 630 51 682 79
rect 716 187 772 214
rect 716 153 725 187
rect 759 153 772 187
rect 716 113 772 153
rect 716 79 725 113
rect 759 79 772 113
rect 716 17 772 79
rect 806 211 1039 245
rect 806 187 867 211
rect 806 153 829 187
rect 863 153 867 187
rect 1001 187 1039 211
rect 806 113 867 153
rect 806 79 829 113
rect 863 79 867 113
rect 806 51 867 79
rect 901 169 967 177
rect 901 135 917 169
rect 951 135 967 169
rect 901 101 967 135
rect 901 67 917 101
rect 951 67 967 101
rect 901 17 967 67
rect 1001 153 1003 187
rect 1037 153 1039 187
rect 1077 208 1111 279
rect 1150 292 1231 360
rect 1184 258 1231 292
rect 1150 242 1231 258
rect 1077 187 1229 208
rect 1077 174 1179 187
rect 1001 113 1039 153
rect 1173 153 1179 174
rect 1213 153 1229 187
rect 1001 79 1003 113
rect 1037 79 1039 113
rect 1001 51 1039 79
rect 1073 124 1139 140
rect 1073 90 1089 124
rect 1123 90 1139 124
rect 1073 17 1139 90
rect 1173 113 1229 153
rect 1173 79 1179 113
rect 1213 79 1229 113
rect 1173 51 1229 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
<< metal1 >>
rect 0 683 1248 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1248 683
rect 0 617 1248 649
rect 0 17 1248 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1248 17
rect 0 -49 1248 -17
<< labels >>
flabel pwell s 0 0 1248 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1248 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 bufinv_8
flabel metal1 s 0 617 1248 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1248 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1248 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1623856
string GDS_START 1612638
<< end >>
