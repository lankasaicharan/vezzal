magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 32 230 217 241
rect 32 191 220 230
rect 764 191 976 275
rect 32 189 976 191
rect 1155 189 1343 241
rect 32 49 1343 189
rect 0 0 1344 49
<< scnmos >>
rect 111 47 141 215
rect 847 165 877 249
rect 249 81 279 165
rect 321 81 351 165
rect 407 81 437 165
rect 501 81 531 165
rect 609 81 639 165
rect 972 79 1002 163
rect 1044 79 1074 163
rect 1234 47 1264 215
<< scpmoshvt >>
rect 80 367 110 619
rect 243 480 273 608
rect 315 480 345 608
rect 423 480 453 564
rect 495 480 525 564
rect 639 395 669 523
rect 898 367 928 495
rect 1016 367 1046 495
rect 1102 367 1132 495
rect 1234 367 1264 619
<< ndiff >>
rect 58 203 111 215
rect 58 169 66 203
rect 100 169 111 203
rect 58 101 111 169
rect 58 67 66 101
rect 100 67 111 101
rect 58 47 111 67
rect 141 204 191 215
rect 141 165 194 204
rect 790 241 847 249
rect 790 207 802 241
rect 836 207 847 241
rect 790 165 847 207
rect 877 165 950 249
rect 141 124 249 165
rect 141 90 165 124
rect 199 90 249 124
rect 141 81 249 90
rect 279 81 321 165
rect 351 157 407 165
rect 351 123 362 157
rect 396 123 407 157
rect 351 81 407 123
rect 437 81 501 165
rect 531 140 609 165
rect 531 106 559 140
rect 593 106 609 140
rect 531 81 609 106
rect 639 139 692 165
rect 892 163 950 165
rect 639 105 650 139
rect 684 105 692 139
rect 639 81 692 105
rect 892 101 972 163
rect 141 47 194 81
rect 892 67 904 101
rect 938 79 972 101
rect 1002 79 1044 163
rect 1074 138 1127 163
rect 1074 104 1085 138
rect 1119 104 1127 138
rect 1074 79 1127 104
rect 1181 93 1234 215
rect 938 67 950 79
rect 892 59 950 67
rect 1181 59 1189 93
rect 1223 59 1234 93
rect 1181 47 1234 59
rect 1264 203 1317 215
rect 1264 169 1275 203
rect 1309 169 1317 203
rect 1264 101 1317 169
rect 1264 67 1275 101
rect 1309 67 1317 101
rect 1264 47 1317 67
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 505 80 565
rect 27 471 35 505
rect 69 471 80 505
rect 27 413 80 471
rect 27 379 35 413
rect 69 379 80 413
rect 27 367 80 379
rect 110 608 175 619
rect 110 607 243 608
rect 110 573 127 607
rect 161 573 243 607
rect 110 498 243 573
rect 110 464 121 498
rect 155 480 243 498
rect 273 480 315 608
rect 345 564 398 608
rect 547 566 624 593
rect 547 564 559 566
rect 345 539 423 564
rect 345 505 364 539
rect 398 505 423 539
rect 345 480 423 505
rect 453 480 495 564
rect 525 532 559 564
rect 593 532 624 566
rect 943 619 1001 627
rect 943 585 955 619
rect 989 585 1001 619
rect 525 523 624 532
rect 525 480 639 523
rect 155 464 163 480
rect 110 367 163 464
rect 547 395 639 480
rect 669 441 755 523
rect 943 495 1001 585
rect 1177 611 1234 619
rect 1177 577 1189 611
rect 1223 577 1234 611
rect 1177 543 1234 577
rect 1177 509 1189 543
rect 1223 509 1234 543
rect 1177 495 1234 509
rect 669 407 713 441
rect 747 407 755 441
rect 669 395 755 407
rect 821 409 898 495
rect 821 375 833 409
rect 867 375 898 409
rect 821 367 898 375
rect 928 367 1016 495
rect 1046 483 1102 495
rect 1046 449 1057 483
rect 1091 449 1102 483
rect 1046 409 1102 449
rect 1046 375 1057 409
rect 1091 375 1102 409
rect 1046 367 1102 375
rect 1132 477 1234 495
rect 1132 443 1143 477
rect 1177 443 1234 477
rect 1132 409 1234 443
rect 1132 375 1143 409
rect 1177 375 1234 409
rect 1132 367 1234 375
rect 1264 599 1317 619
rect 1264 565 1275 599
rect 1309 565 1317 599
rect 1264 503 1317 565
rect 1264 469 1275 503
rect 1309 469 1317 503
rect 1264 413 1317 469
rect 1264 379 1275 413
rect 1309 379 1317 413
rect 1264 367 1317 379
<< ndiffc >>
rect 66 169 100 203
rect 66 67 100 101
rect 802 207 836 241
rect 165 90 199 124
rect 362 123 396 157
rect 559 106 593 140
rect 650 105 684 139
rect 904 67 938 101
rect 1085 104 1119 138
rect 1189 59 1223 93
rect 1275 169 1309 203
rect 1275 67 1309 101
<< pdiffc >>
rect 35 565 69 599
rect 35 471 69 505
rect 35 379 69 413
rect 127 573 161 607
rect 121 464 155 498
rect 364 505 398 539
rect 559 532 593 566
rect 955 585 989 619
rect 1189 577 1223 611
rect 1189 509 1223 543
rect 713 407 747 441
rect 833 375 867 409
rect 1057 449 1091 483
rect 1057 375 1091 409
rect 1143 443 1177 477
rect 1143 375 1177 409
rect 1275 565 1309 599
rect 1275 469 1309 503
rect 1275 379 1309 413
<< poly >>
rect 80 619 110 645
rect 243 608 273 634
rect 315 608 345 634
rect 495 608 783 638
rect 423 564 453 590
rect 495 564 525 608
rect 717 605 783 608
rect 717 571 733 605
rect 767 571 783 605
rect 717 555 783 571
rect 1234 619 1264 645
rect 639 523 669 549
rect 80 335 110 367
rect 80 319 159 335
rect 80 285 109 319
rect 143 285 159 319
rect 243 292 273 480
rect 315 448 345 480
rect 315 432 381 448
rect 315 398 331 432
rect 365 398 381 432
rect 315 382 381 398
rect 423 373 453 480
rect 495 454 525 480
rect 898 495 928 521
rect 1016 495 1046 521
rect 1102 495 1132 521
rect 639 373 669 395
rect 423 353 669 373
rect 423 337 469 353
rect 321 319 469 337
rect 503 350 669 353
rect 503 334 675 350
rect 503 319 625 334
rect 321 301 625 319
rect 80 269 159 285
rect 213 276 279 292
rect 111 215 141 269
rect 213 242 229 276
rect 263 242 279 276
rect 213 226 279 242
rect 249 165 279 226
rect 321 165 351 301
rect 609 300 625 301
rect 659 300 675 334
rect 393 243 459 259
rect 609 257 675 300
rect 723 345 789 350
rect 898 345 928 367
rect 1016 345 1046 367
rect 723 334 1046 345
rect 723 300 739 334
rect 773 315 1046 334
rect 773 300 789 315
rect 723 284 789 300
rect 393 209 409 243
rect 443 209 459 243
rect 393 193 459 209
rect 501 237 567 253
rect 501 203 517 237
rect 551 203 567 237
rect 407 165 437 193
rect 501 187 567 203
rect 609 223 625 257
rect 659 223 675 257
rect 847 249 877 315
rect 609 207 675 223
rect 501 165 531 187
rect 609 165 639 207
rect 847 139 877 165
rect 972 163 1002 315
rect 1102 267 1132 367
rect 1234 333 1264 367
rect 1189 317 1264 333
rect 1189 283 1205 317
rect 1239 283 1264 317
rect 1189 267 1264 283
rect 1069 251 1135 267
rect 1069 231 1085 251
rect 1044 217 1085 231
rect 1119 217 1135 251
rect 1044 201 1135 217
rect 1234 215 1264 267
rect 1044 163 1074 201
rect 249 55 279 81
rect 321 55 351 81
rect 407 55 437 81
rect 501 55 531 81
rect 609 55 639 81
rect 972 53 1002 79
rect 1044 53 1074 79
rect 111 21 141 47
rect 1234 21 1264 47
<< polycont >>
rect 733 571 767 605
rect 109 285 143 319
rect 331 398 365 432
rect 469 319 503 353
rect 229 242 263 276
rect 625 300 659 334
rect 739 300 773 334
rect 409 209 443 243
rect 517 203 551 237
rect 625 223 659 257
rect 1205 283 1239 317
rect 1085 217 1119 251
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 19 599 85 615
rect 19 565 35 599
rect 69 565 85 599
rect 19 505 85 565
rect 19 471 35 505
rect 69 471 85 505
rect 19 414 85 471
rect 121 607 161 649
rect 121 573 127 607
rect 121 498 161 573
rect 155 464 161 498
rect 121 448 161 464
rect 195 581 489 615
rect 195 414 229 581
rect 19 413 229 414
rect 19 379 35 413
rect 69 380 229 413
rect 263 539 414 547
rect 263 505 364 539
rect 398 505 414 539
rect 263 497 414 505
rect 69 379 73 380
rect 19 219 73 379
rect 263 348 297 497
rect 455 489 489 581
rect 543 566 609 649
rect 939 619 1005 649
rect 543 532 559 566
rect 593 532 609 566
rect 717 605 783 615
rect 717 571 733 605
rect 767 571 783 605
rect 939 585 955 619
rect 989 585 1005 619
rect 939 581 1005 585
rect 1127 611 1239 649
rect 717 549 783 571
rect 543 523 609 532
rect 645 547 783 549
rect 1127 577 1189 611
rect 1223 577 1239 611
rect 645 513 1019 547
rect 645 489 679 513
rect 455 455 679 489
rect 331 432 419 448
rect 365 421 419 432
rect 713 445 951 479
rect 713 441 765 445
rect 365 407 713 421
rect 747 407 765 441
rect 365 398 765 407
rect 331 387 765 398
rect 817 409 883 411
rect 331 382 419 387
rect 263 346 351 348
rect 107 319 351 346
rect 107 285 109 319
rect 143 312 351 319
rect 143 285 159 312
rect 107 269 159 285
rect 195 276 283 278
rect 195 242 229 276
rect 263 242 283 276
rect 195 232 283 242
rect 19 203 116 219
rect 19 169 66 203
rect 100 198 116 203
rect 100 169 283 198
rect 19 164 283 169
rect 19 101 115 164
rect 19 67 66 101
rect 100 67 115 101
rect 19 51 115 67
rect 149 124 215 130
rect 149 90 165 124
rect 199 90 215 124
rect 149 17 215 90
rect 249 85 283 164
rect 317 159 351 312
rect 385 259 419 382
rect 817 375 833 409
rect 867 375 883 409
rect 453 319 469 353
rect 503 334 659 353
rect 503 319 625 334
rect 453 301 625 319
rect 609 300 625 301
rect 385 243 456 259
rect 609 257 659 300
rect 693 334 783 353
rect 693 300 739 334
rect 773 300 783 334
rect 693 284 783 300
rect 385 209 409 243
rect 443 209 456 243
rect 385 193 456 209
rect 490 237 567 253
rect 490 203 517 237
rect 551 203 567 237
rect 609 223 625 257
rect 817 250 883 375
rect 659 241 883 250
rect 659 223 802 241
rect 609 207 802 223
rect 836 207 883 241
rect 609 205 883 207
rect 490 190 567 203
rect 317 157 412 159
rect 317 123 362 157
rect 396 123 412 157
rect 317 119 412 123
rect 490 85 524 190
rect 917 171 951 445
rect 985 265 1019 513
rect 1127 543 1239 577
rect 1127 509 1189 543
rect 1223 509 1239 543
rect 1053 483 1093 499
rect 1053 449 1057 483
rect 1091 449 1093 483
rect 1053 409 1093 449
rect 1053 375 1057 409
rect 1091 375 1093 409
rect 1053 333 1093 375
rect 1127 477 1239 509
rect 1127 443 1143 477
rect 1177 443 1239 477
rect 1127 409 1239 443
rect 1127 375 1143 409
rect 1177 375 1239 409
rect 1127 367 1239 375
rect 1273 599 1325 615
rect 1273 565 1275 599
rect 1309 565 1325 599
rect 1273 503 1325 565
rect 1273 469 1275 503
rect 1309 469 1325 503
rect 1273 413 1325 469
rect 1273 379 1275 413
rect 1309 379 1325 413
rect 1053 317 1239 333
rect 1053 299 1205 317
rect 1189 283 1205 299
rect 985 251 1135 265
rect 985 217 1085 251
rect 1119 217 1135 251
rect 985 201 1135 217
rect 249 51 524 85
rect 558 140 608 156
rect 558 106 559 140
rect 593 106 608 140
rect 558 17 608 106
rect 642 139 951 171
rect 1189 167 1239 283
rect 642 105 650 139
rect 684 137 951 139
rect 1069 138 1239 167
rect 684 105 700 137
rect 642 89 700 105
rect 1069 104 1085 138
rect 1119 133 1239 138
rect 1273 203 1325 379
rect 1273 169 1275 203
rect 1309 169 1325 203
rect 1119 104 1135 133
rect 888 101 954 103
rect 888 67 904 101
rect 938 67 954 101
rect 1069 88 1135 104
rect 1273 101 1325 169
rect 1173 93 1239 99
rect 888 17 954 67
rect 1173 59 1189 93
rect 1223 59 1239 93
rect 1173 17 1239 59
rect 1273 67 1275 101
rect 1309 67 1325 101
rect 1273 51 1325 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dlclkp_1
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1279 390 1313 424 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1279 464 1313 498 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1279 538 1313 572 0 FreeSans 340 0 0 0 GCLK
port 7 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3567902
string GDS_START 3557472
<< end >>
