magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 5426 1975
<< nwell >>
rect -38 397 4166 704
rect -38 331 1668 397
rect 1922 331 4166 397
<< pwell >>
rect 1712 279 1818 355
rect 328 246 436 275
rect 194 230 701 246
rect 903 230 1230 275
rect 1712 273 2108 279
rect 194 229 1230 230
rect 1498 235 2108 273
rect 1498 229 2359 235
rect 194 220 2807 229
rect 1 49 2807 220
rect 3199 183 3581 207
rect 3935 183 4127 251
rect 3199 49 4127 183
rect 0 0 4128 49
<< scnmos >>
rect 82 110 112 194
rect 302 136 332 220
rect 432 136 462 220
rect 504 136 534 220
rect 590 136 620 220
rect 784 120 814 204
rect 1020 165 1050 249
rect 1120 165 1150 249
rect 1313 119 1343 203
rect 1385 119 1415 203
rect 1579 119 1609 247
rect 1686 163 1716 247
rect 1901 125 1931 253
rect 1973 125 2003 253
rect 2104 125 2134 209
rect 2176 125 2206 209
rect 2248 125 2278 209
rect 2442 119 2472 203
rect 2514 119 2544 203
rect 2600 119 2630 203
rect 2694 119 2724 203
rect 3305 97 3335 181
rect 3377 97 3407 181
rect 3449 97 3479 181
rect 3664 73 3694 157
rect 3736 73 3766 157
rect 3822 73 3852 157
rect 4016 57 4046 225
<< scpmoshvt >>
rect 98 466 128 594
rect 283 466 313 594
rect 361 466 391 594
rect 522 466 552 594
rect 624 466 654 594
rect 860 466 890 594
rect 969 424 999 508
rect 1098 424 1128 508
rect 1176 424 1206 508
rect 1308 424 1338 508
rect 1529 373 1559 541
rect 1654 433 1684 561
rect 2039 397 2069 565
rect 2111 397 2141 565
rect 2786 390 2836 590
rect 2884 390 2934 590
rect 3013 390 3063 590
rect 3105 390 3155 590
rect 3211 390 3261 590
rect 3340 390 3370 518
rect 3432 390 3462 518
rect 3564 390 3614 590
rect 3808 367 3838 495
rect 3974 367 4004 619
<< ndiff >>
rect 354 237 410 249
rect 354 220 366 237
rect 27 169 82 194
rect 27 135 37 169
rect 71 135 82 169
rect 27 110 82 135
rect 112 169 166 194
rect 112 135 123 169
rect 157 135 166 169
rect 220 182 302 220
rect 220 148 230 182
rect 264 148 302 182
rect 220 136 302 148
rect 332 203 366 220
rect 400 220 410 237
rect 400 203 432 220
rect 332 136 432 203
rect 462 136 504 220
rect 534 195 590 220
rect 534 161 545 195
rect 579 161 590 195
rect 534 136 590 161
rect 620 187 675 220
rect 620 153 631 187
rect 665 153 675 187
rect 620 136 675 153
rect 729 179 784 204
rect 729 145 739 179
rect 773 145 784 179
rect 112 110 166 135
rect 729 120 784 145
rect 814 179 869 204
rect 814 145 825 179
rect 859 145 869 179
rect 814 120 869 145
rect 929 199 1020 249
rect 929 165 939 199
rect 973 165 1020 199
rect 1050 237 1120 249
rect 1050 203 1075 237
rect 1109 203 1120 237
rect 1050 165 1120 203
rect 1150 224 1204 249
rect 1150 190 1161 224
rect 1195 190 1204 224
rect 1738 317 1792 329
rect 1738 283 1748 317
rect 1782 283 1792 317
rect 1738 247 1792 283
rect 1150 165 1204 190
rect 1258 166 1313 203
rect 929 152 985 165
rect 1258 132 1268 166
rect 1302 132 1313 166
rect 1258 119 1313 132
rect 1343 119 1385 203
rect 1415 166 1470 203
rect 1415 132 1426 166
rect 1460 132 1470 166
rect 1415 119 1470 132
rect 1524 192 1579 247
rect 1524 158 1534 192
rect 1568 158 1579 192
rect 1524 119 1579 158
rect 1609 165 1686 247
rect 1609 131 1620 165
rect 1654 163 1686 165
rect 1716 163 1792 247
rect 1846 241 1901 253
rect 1846 207 1856 241
rect 1890 207 1901 241
rect 1846 171 1901 207
rect 1654 131 1664 163
rect 1846 137 1856 171
rect 1890 137 1901 171
rect 1609 119 1664 131
rect 1846 125 1901 137
rect 1931 125 1973 253
rect 2003 241 2082 253
rect 2003 207 2038 241
rect 2072 209 2082 241
rect 2072 207 2104 209
rect 2003 171 2104 207
rect 2003 137 2038 171
rect 2072 137 2104 171
rect 2003 125 2104 137
rect 2134 125 2176 209
rect 2206 125 2248 209
rect 2278 176 2333 209
rect 2278 142 2289 176
rect 2323 142 2333 176
rect 2278 125 2333 142
rect 2387 178 2442 203
rect 2387 144 2397 178
rect 2431 144 2442 178
rect 2387 119 2442 144
rect 2472 119 2514 203
rect 2544 178 2600 203
rect 2544 144 2555 178
rect 2589 144 2600 178
rect 2544 119 2600 144
rect 2630 162 2694 203
rect 2630 128 2641 162
rect 2675 128 2694 162
rect 2630 119 2694 128
rect 2724 178 2781 203
rect 2724 144 2735 178
rect 2769 144 2781 178
rect 2724 119 2781 144
rect 3225 169 3305 181
rect 3225 135 3237 169
rect 3271 135 3305 169
rect 3225 97 3305 135
rect 3335 97 3377 181
rect 3407 97 3449 181
rect 3479 103 3555 181
rect 3961 213 4016 225
rect 3961 179 3971 213
rect 4005 179 4016 213
rect 3479 97 3511 103
rect 3501 69 3511 97
rect 3545 69 3555 103
rect 3609 132 3664 157
rect 3609 98 3619 132
rect 3653 98 3664 132
rect 3609 73 3664 98
rect 3694 73 3736 157
rect 3766 132 3822 157
rect 3766 98 3777 132
rect 3811 98 3822 132
rect 3766 73 3822 98
rect 3852 132 3907 157
rect 3852 98 3863 132
rect 3897 98 3907 132
rect 3852 73 3907 98
rect 3961 103 4016 179
rect 3501 54 3555 69
rect 3961 69 3971 103
rect 4005 69 4016 103
rect 3961 57 4016 69
rect 4046 213 4101 225
rect 4046 179 4057 213
rect 4091 179 4101 213
rect 4046 103 4101 179
rect 4046 69 4057 103
rect 4091 69 4101 103
rect 4046 57 4101 69
<< pdiff >>
rect 41 582 98 594
rect 41 548 53 582
rect 87 548 98 582
rect 41 512 98 548
rect 41 478 53 512
rect 87 478 98 512
rect 41 466 98 478
rect 128 550 283 594
rect 128 516 140 550
rect 174 516 283 550
rect 128 466 283 516
rect 313 466 361 594
rect 391 582 522 594
rect 391 548 477 582
rect 511 548 522 582
rect 391 512 522 548
rect 391 478 477 512
rect 511 478 522 512
rect 391 466 522 478
rect 552 466 624 594
rect 654 560 860 594
rect 654 526 665 560
rect 699 526 860 560
rect 654 466 860 526
rect 890 582 947 594
rect 890 548 901 582
rect 935 548 947 582
rect 890 512 947 548
rect 890 478 901 512
rect 935 508 947 512
rect 1228 588 1286 600
rect 1228 554 1240 588
rect 1274 554 1286 588
rect 1574 571 1632 583
rect 1228 508 1286 554
rect 1574 541 1586 571
rect 935 478 969 508
rect 890 466 969 478
rect 919 424 969 466
rect 999 470 1098 508
rect 999 436 1053 470
rect 1087 436 1098 470
rect 999 424 1098 436
rect 1128 424 1176 508
rect 1206 424 1308 508
rect 1338 436 1418 508
rect 1338 424 1372 436
rect 1360 402 1372 424
rect 1406 402 1418 436
rect 1360 390 1418 402
rect 1472 419 1529 541
rect 1472 385 1484 419
rect 1518 385 1529 419
rect 1472 373 1529 385
rect 1559 537 1586 541
rect 1620 561 1632 571
rect 1620 537 1654 561
rect 1559 433 1654 537
rect 1684 549 1741 561
rect 1684 515 1695 549
rect 1729 515 1741 549
rect 1684 479 1741 515
rect 1684 445 1695 479
rect 1729 445 1741 479
rect 1684 433 1741 445
rect 1982 531 2039 565
rect 1982 497 1994 531
rect 2028 497 2039 531
rect 1982 443 2039 497
rect 1559 373 1632 433
rect 1982 409 1994 443
rect 2028 409 2039 443
rect 1982 397 2039 409
rect 2069 397 2111 565
rect 2141 453 2198 565
rect 2141 419 2152 453
rect 2186 419 2198 453
rect 2141 397 2198 419
rect 3484 590 3542 601
rect 3903 607 3974 619
rect 2729 549 2786 590
rect 2729 515 2741 549
rect 2775 515 2786 549
rect 2729 390 2786 515
rect 2836 390 2884 590
rect 2934 575 3013 590
rect 2934 541 2945 575
rect 2979 541 3013 575
rect 2934 390 3013 541
rect 3063 390 3105 590
rect 3155 436 3211 590
rect 3155 402 3166 436
rect 3200 402 3211 436
rect 3155 390 3211 402
rect 3261 575 3318 590
rect 3261 541 3272 575
rect 3306 541 3318 575
rect 3484 588 3564 590
rect 3484 554 3496 588
rect 3530 554 3564 588
rect 3261 518 3318 541
rect 3484 518 3564 554
rect 3261 390 3340 518
rect 3370 436 3432 518
rect 3370 402 3387 436
rect 3421 402 3432 436
rect 3370 390 3432 402
rect 3462 390 3564 518
rect 3614 420 3694 590
rect 3903 573 3915 607
rect 3949 573 3974 607
rect 3903 510 3974 573
rect 3903 495 3915 510
rect 3614 390 3648 420
rect 3636 386 3648 390
rect 3682 386 3694 420
rect 3636 374 3694 386
rect 3751 416 3808 495
rect 3751 382 3763 416
rect 3797 382 3808 416
rect 3751 367 3808 382
rect 3838 476 3915 495
rect 3949 476 3974 510
rect 3838 413 3974 476
rect 3838 379 3915 413
rect 3949 379 3974 413
rect 3838 367 3974 379
rect 4004 599 4061 619
rect 4004 565 4015 599
rect 4049 565 4061 599
rect 4004 506 4061 565
rect 4004 472 4015 506
rect 4049 472 4061 506
rect 4004 413 4061 472
rect 4004 379 4015 413
rect 4049 379 4061 413
rect 4004 367 4061 379
<< ndiffc >>
rect 37 135 71 169
rect 123 135 157 169
rect 230 148 264 182
rect 366 203 400 237
rect 545 161 579 195
rect 631 153 665 187
rect 739 145 773 179
rect 825 145 859 179
rect 939 165 973 199
rect 1075 203 1109 237
rect 1161 190 1195 224
rect 1748 283 1782 317
rect 1268 132 1302 166
rect 1426 132 1460 166
rect 1534 158 1568 192
rect 1620 131 1654 165
rect 1856 207 1890 241
rect 1856 137 1890 171
rect 2038 207 2072 241
rect 2038 137 2072 171
rect 2289 142 2323 176
rect 2397 144 2431 178
rect 2555 144 2589 178
rect 2641 128 2675 162
rect 2735 144 2769 178
rect 3237 135 3271 169
rect 3971 179 4005 213
rect 3511 69 3545 103
rect 3619 98 3653 132
rect 3777 98 3811 132
rect 3863 98 3897 132
rect 3971 69 4005 103
rect 4057 179 4091 213
rect 4057 69 4091 103
<< pdiffc >>
rect 53 548 87 582
rect 53 478 87 512
rect 140 516 174 550
rect 477 548 511 582
rect 477 478 511 512
rect 665 526 699 560
rect 901 548 935 582
rect 901 478 935 512
rect 1240 554 1274 588
rect 1053 436 1087 470
rect 1372 402 1406 436
rect 1484 385 1518 419
rect 1586 537 1620 571
rect 1695 515 1729 549
rect 1695 445 1729 479
rect 1994 497 2028 531
rect 1994 409 2028 443
rect 2152 419 2186 453
rect 2741 515 2775 549
rect 2945 541 2979 575
rect 3166 402 3200 436
rect 3272 541 3306 575
rect 3496 554 3530 588
rect 3387 402 3421 436
rect 3915 573 3949 607
rect 3648 386 3682 420
rect 3763 382 3797 416
rect 3915 476 3949 510
rect 3915 379 3949 413
rect 4015 565 4049 599
rect 4015 472 4049 506
rect 4015 379 4049 413
<< poly >>
rect 98 594 128 620
rect 283 594 313 620
rect 361 594 391 620
rect 522 594 552 620
rect 624 594 654 620
rect 860 594 890 620
rect 1098 615 2358 645
rect 969 508 999 534
rect 1098 508 1128 615
rect 1176 508 1206 534
rect 1529 541 1559 567
rect 1308 508 1338 534
rect 98 434 128 466
rect 283 434 313 466
rect 98 418 313 434
rect 98 384 137 418
rect 171 404 313 418
rect 361 434 391 466
rect 361 418 427 434
rect 171 384 190 404
rect 98 350 190 384
rect 361 384 377 418
rect 411 398 427 418
rect 411 384 462 398
rect 522 386 552 466
rect 361 368 462 384
rect 98 320 137 350
rect 82 316 137 320
rect 171 320 190 350
rect 171 316 332 320
rect 82 290 332 316
rect 82 194 112 290
rect 302 220 332 290
rect 432 220 462 368
rect 504 370 576 386
rect 504 336 526 370
rect 560 336 576 370
rect 504 320 576 336
rect 624 376 654 466
rect 860 376 890 466
rect 624 360 736 376
rect 624 326 686 360
rect 720 326 736 360
rect 504 220 534 320
rect 624 310 736 326
rect 784 360 890 376
rect 784 326 800 360
rect 834 340 890 360
rect 969 384 999 424
rect 969 368 1050 384
rect 834 326 914 340
rect 784 310 914 326
rect 969 334 993 368
rect 1027 334 1050 368
rect 969 318 1050 334
rect 624 272 654 310
rect 590 242 654 272
rect 590 220 620 242
rect 784 204 814 310
rect 302 110 332 136
rect 432 110 462 136
rect 504 110 534 136
rect 590 110 620 136
rect 82 84 112 110
rect 784 94 814 120
rect 884 51 914 310
rect 1020 249 1050 318
rect 1098 301 1128 424
rect 1176 379 1206 424
rect 1176 349 1258 379
rect 1192 315 1208 349
rect 1242 315 1258 349
rect 1308 375 1338 424
rect 1308 345 1421 375
rect 1654 561 1684 615
rect 2039 565 2069 615
rect 2111 565 2141 615
rect 1654 411 1684 433
rect 1654 381 1716 411
rect 1098 271 1150 301
rect 1120 249 1150 271
rect 1192 297 1258 315
rect 1192 281 1343 297
rect 1192 267 1272 281
rect 1256 247 1272 267
rect 1306 247 1343 281
rect 1391 255 1421 345
rect 1529 335 1559 373
rect 1493 319 1559 335
rect 1493 285 1509 319
rect 1543 299 1559 319
rect 1543 285 1609 299
rect 1493 269 1609 285
rect 1256 231 1343 247
rect 1313 203 1343 231
rect 1385 225 1421 255
rect 1579 247 1609 269
rect 1686 247 1716 381
rect 2039 375 2069 397
rect 2111 375 2141 397
rect 1842 349 1931 365
rect 1842 315 1858 349
rect 1892 315 1931 349
rect 2039 345 2141 375
rect 2328 368 2358 615
rect 2625 612 2836 642
rect 3974 619 4004 645
rect 2625 599 2691 612
rect 2625 565 2641 599
rect 2675 565 2691 599
rect 2786 590 2836 612
rect 2884 590 2934 616
rect 3013 590 3063 616
rect 3105 590 3155 616
rect 3211 590 3261 616
rect 3564 590 3614 616
rect 2625 549 2691 565
rect 2442 520 2508 536
rect 2442 486 2458 520
rect 2492 500 2508 520
rect 2492 486 2544 500
rect 2442 470 2544 486
rect 2220 349 2286 365
rect 1842 303 1931 315
rect 1842 299 2003 303
rect 1901 273 2003 299
rect 1901 253 1931 273
rect 1973 253 2003 273
rect 1385 203 1415 225
rect 1020 139 1050 165
rect 1120 139 1150 165
rect 1686 137 1716 163
rect 2104 209 2134 345
rect 2220 315 2236 349
rect 2270 315 2286 349
rect 2220 281 2286 315
rect 2328 352 2394 368
rect 2328 318 2344 352
rect 2378 318 2394 352
rect 2328 302 2394 318
rect 2220 261 2236 281
rect 2176 247 2236 261
rect 2270 247 2286 281
rect 2176 231 2286 247
rect 2176 209 2206 231
rect 2248 209 2278 231
rect 2442 203 2472 470
rect 2514 203 2544 470
rect 3340 518 3370 544
rect 3432 518 3462 544
rect 3808 495 3838 521
rect 2786 364 2836 390
rect 2884 322 2934 390
rect 3013 364 3063 390
rect 2586 299 2652 315
rect 2586 265 2602 299
rect 2636 265 2652 299
rect 2586 249 2652 265
rect 2884 306 2991 322
rect 2884 272 2941 306
rect 2975 272 2991 306
rect 2884 256 2991 272
rect 2600 203 2630 249
rect 2694 203 2724 229
rect 1313 93 1343 119
rect 1385 51 1415 119
rect 1579 93 1609 119
rect 1901 99 1931 125
rect 1973 99 2003 125
rect 2104 99 2134 125
rect 2176 99 2206 125
rect 2248 99 2278 125
rect 3033 159 3063 364
rect 3105 207 3155 390
rect 3211 348 3261 390
rect 3340 358 3370 390
rect 3197 332 3263 348
rect 3197 298 3213 332
rect 3247 298 3263 332
rect 3197 282 3263 298
rect 3305 342 3384 358
rect 3305 308 3334 342
rect 3368 308 3384 342
rect 3305 292 3384 308
rect 2997 143 3063 159
rect 2442 93 2472 119
rect 2514 93 2544 119
rect 2600 93 2630 119
rect 2694 51 2724 119
rect 2997 109 3013 143
rect 3047 109 3063 143
rect 2997 93 3063 109
rect 3125 51 3155 207
rect 3305 181 3335 292
rect 3432 290 3462 390
rect 3564 338 3614 390
rect 3564 290 3594 338
rect 3808 329 3838 367
rect 3974 329 4004 367
rect 3808 313 3875 329
rect 3432 274 3713 290
rect 3432 260 3663 274
rect 3432 233 3479 260
rect 3377 203 3479 233
rect 3647 240 3663 260
rect 3697 240 3713 274
rect 3808 279 3825 313
rect 3859 279 3875 313
rect 3808 263 3875 279
rect 3938 313 4004 329
rect 3938 279 3954 313
rect 3988 293 4004 313
rect 3988 279 4046 293
rect 3938 263 4046 279
rect 3647 224 3713 240
rect 3377 181 3407 203
rect 3449 181 3479 203
rect 3664 215 3713 224
rect 3664 185 3766 215
rect 3664 157 3694 185
rect 3736 157 3766 185
rect 3822 157 3852 263
rect 4016 225 4046 263
rect 3305 71 3335 97
rect 3377 71 3407 97
rect 3449 71 3479 97
rect 884 21 3155 51
rect 3664 47 3694 73
rect 3736 47 3766 73
rect 3822 47 3852 73
rect 4016 31 4046 57
<< polycont >>
rect 137 384 171 418
rect 377 384 411 418
rect 137 316 171 350
rect 526 336 560 370
rect 686 326 720 360
rect 800 326 834 360
rect 993 334 1027 368
rect 1208 315 1242 349
rect 1272 247 1306 281
rect 1509 285 1543 319
rect 1858 315 1892 349
rect 2641 565 2675 599
rect 2458 486 2492 520
rect 2236 315 2270 349
rect 2344 318 2378 352
rect 2236 247 2270 281
rect 2602 265 2636 299
rect 2941 272 2975 306
rect 3213 298 3247 332
rect 3334 308 3368 342
rect 3013 109 3047 143
rect 3663 240 3697 274
rect 3825 279 3859 313
rect 3954 279 3988 313
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3775 683
rect 3809 649 3871 683
rect 3905 649 3967 683
rect 4001 649 4063 683
rect 4097 649 4128 683
rect 21 582 87 598
rect 21 548 53 582
rect 21 512 87 548
rect 21 478 53 512
rect 21 266 87 478
rect 124 550 190 649
rect 124 516 140 550
rect 174 516 190 550
rect 124 468 190 516
rect 461 582 527 598
rect 461 548 477 582
rect 511 548 527 582
rect 461 512 527 548
rect 461 502 477 512
rect 245 478 477 502
rect 511 478 527 512
rect 649 560 715 649
rect 649 526 665 560
rect 699 526 715 560
rect 649 488 715 526
rect 885 582 951 598
rect 885 548 901 582
rect 935 548 951 582
rect 1224 588 1290 649
rect 1224 554 1240 588
rect 1274 554 1290 588
rect 1570 571 1636 649
rect 885 512 951 548
rect 245 468 527 478
rect 121 418 187 434
rect 121 384 137 418
rect 171 384 187 418
rect 121 350 187 384
rect 121 316 137 350
rect 171 316 187 350
rect 121 300 187 316
rect 245 334 279 468
rect 461 454 527 468
rect 885 478 901 512
rect 935 478 951 512
rect 885 454 951 478
rect 313 418 427 434
rect 461 420 951 454
rect 985 520 1190 554
rect 1570 537 1586 571
rect 1620 537 1636 571
rect 1711 599 2691 615
rect 3899 607 3965 649
rect 1711 581 2641 599
rect 1711 565 1745 581
rect 1570 521 1636 537
rect 1679 549 1745 565
rect 2625 565 2641 581
rect 2675 565 2691 599
rect 2625 549 2691 565
rect 2725 549 2791 594
rect 313 384 377 418
rect 411 384 427 418
rect 313 368 427 384
rect 461 370 576 386
rect 461 336 526 370
rect 560 336 576 370
rect 245 300 416 334
rect 21 232 332 266
rect 21 169 71 232
rect 21 135 37 169
rect 21 106 71 135
rect 107 169 173 198
rect 107 135 123 169
rect 157 135 173 169
rect 107 17 173 135
rect 214 182 264 198
rect 214 148 230 182
rect 214 85 264 148
rect 298 153 332 232
rect 366 237 416 300
rect 400 203 416 237
rect 366 187 416 203
rect 461 320 576 336
rect 670 360 743 376
rect 670 326 686 360
rect 720 326 743 360
rect 461 153 495 320
rect 670 310 743 326
rect 784 360 850 376
rect 784 326 800 360
rect 834 326 850 360
rect 784 310 850 326
rect 909 284 943 420
rect 985 384 1019 520
rect 1156 487 1536 520
rect 1679 515 1695 549
rect 1729 515 1745 549
rect 1679 487 1745 515
rect 1156 486 1745 487
rect 1053 470 1111 486
rect 1087 452 1111 470
rect 1502 479 1745 486
rect 1502 453 1695 479
rect 1087 436 1422 452
rect 1053 418 1372 436
rect 977 368 1043 384
rect 977 334 993 368
rect 1027 334 1043 368
rect 977 318 1043 334
rect 298 119 495 153
rect 529 242 875 276
rect 909 250 1041 284
rect 1077 253 1111 418
rect 1356 402 1372 418
rect 1406 402 1422 436
rect 1679 445 1695 453
rect 1729 445 1745 479
rect 1192 349 1258 365
rect 1192 315 1208 349
rect 1242 321 1258 349
rect 1356 335 1422 402
rect 1468 385 1484 419
rect 1518 385 1627 419
rect 1468 369 1627 385
rect 1242 315 1322 321
rect 1192 287 1322 315
rect 1256 281 1322 287
rect 529 195 595 242
rect 529 161 545 195
rect 579 161 595 195
rect 529 148 595 161
rect 631 187 681 208
rect 665 153 681 187
rect 631 85 681 153
rect 214 51 681 85
rect 723 179 773 208
rect 723 145 739 179
rect 723 17 773 145
rect 809 179 875 242
rect 809 145 825 179
rect 859 145 875 179
rect 809 116 875 145
rect 923 199 973 216
rect 923 165 939 199
rect 923 85 973 165
rect 1007 153 1041 250
rect 1075 237 1111 253
rect 1109 203 1111 237
rect 1075 187 1111 203
rect 1145 224 1211 253
rect 1145 190 1161 224
rect 1195 190 1211 224
rect 1256 247 1272 281
rect 1306 247 1322 281
rect 1356 319 1559 335
rect 1356 285 1509 319
rect 1543 285 1559 319
rect 1356 269 1559 285
rect 1256 235 1322 247
rect 1593 235 1627 369
rect 1679 333 1745 445
rect 1978 531 2508 547
rect 1978 497 1994 531
rect 2028 520 2508 531
rect 2028 513 2458 520
rect 2028 497 2100 513
rect 1978 443 2100 497
rect 2442 486 2458 513
rect 2492 504 2508 520
rect 2725 515 2741 549
rect 2775 515 2791 549
rect 2905 581 2995 594
rect 2905 547 2911 581
rect 2945 575 2995 581
rect 2905 541 2945 547
rect 2979 541 2995 575
rect 2905 538 2995 541
rect 3256 581 3335 594
rect 3256 575 3295 581
rect 3256 541 3272 575
rect 3329 547 3335 581
rect 3306 541 3335 547
rect 3256 538 3335 541
rect 3385 588 3546 605
rect 3385 581 3496 588
rect 3385 547 3391 581
rect 3425 554 3496 581
rect 3530 554 3546 588
rect 3425 547 3546 554
rect 3385 538 3546 547
rect 3899 573 3915 607
rect 3949 573 3965 607
rect 2725 504 2791 515
rect 3899 510 3965 573
rect 2492 486 3865 504
rect 1978 409 1994 443
rect 2028 409 2100 443
rect 1978 408 2100 409
rect 1842 349 1908 365
rect 1842 333 1858 349
rect 1679 317 1858 333
rect 1679 283 1748 317
rect 1782 315 1858 317
rect 1892 315 1908 349
rect 1782 299 1908 315
rect 1782 283 1798 299
rect 1679 267 1798 283
rect 1256 233 1627 235
rect 1840 241 1906 257
rect 1840 233 1856 241
rect 1256 207 1856 233
rect 1890 207 1906 241
rect 1256 201 1906 207
rect 1145 153 1211 190
rect 1518 199 1906 201
rect 1518 192 1568 199
rect 1007 119 1211 153
rect 1252 166 1318 167
rect 1252 132 1268 166
rect 1302 132 1318 166
rect 1252 85 1318 132
rect 923 51 1318 85
rect 1410 166 1476 167
rect 1410 132 1426 166
rect 1460 132 1476 166
rect 1410 17 1476 132
rect 1518 158 1534 192
rect 1840 171 1906 199
rect 1518 115 1568 158
rect 1604 131 1620 165
rect 1654 131 1670 165
rect 1604 17 1670 131
rect 1840 137 1856 171
rect 1890 137 1906 171
rect 1840 87 1906 137
rect 2038 241 2100 408
rect 2072 207 2100 241
rect 2038 171 2100 207
rect 2072 137 2100 171
rect 2038 121 2100 137
rect 2136 453 2186 479
rect 2442 470 3865 486
rect 2136 419 2152 453
rect 2136 87 2186 419
rect 2220 402 2991 436
rect 2220 349 2286 402
rect 2220 315 2236 349
rect 2270 315 2286 349
rect 2220 281 2286 315
rect 2328 352 2905 368
rect 2328 318 2344 352
rect 2378 334 2905 352
rect 2378 318 2394 334
rect 2328 302 2394 318
rect 2220 247 2236 281
rect 2270 265 2286 281
rect 2586 299 2837 300
rect 2586 265 2602 299
rect 2636 265 2837 299
rect 2270 247 2447 265
rect 2586 264 2837 265
rect 2220 231 2447 247
rect 1840 53 2186 87
rect 2273 176 2339 197
rect 2273 142 2289 176
rect 2323 142 2339 176
rect 2273 17 2339 142
rect 2381 178 2447 231
rect 2381 144 2397 178
rect 2431 144 2447 178
rect 2381 115 2447 144
rect 2539 196 2769 230
rect 2539 178 2589 196
rect 2539 144 2555 178
rect 2735 178 2769 196
rect 2539 115 2589 144
rect 2625 128 2641 162
rect 2675 128 2691 162
rect 2625 17 2691 128
rect 2735 115 2769 144
rect 2803 154 2837 264
rect 2871 222 2905 334
rect 2939 322 2991 402
rect 3129 402 3166 436
rect 3200 402 3216 436
rect 3129 386 3216 402
rect 3129 322 3163 386
rect 3250 348 3284 470
rect 3371 402 3387 436
rect 3421 402 3499 436
rect 2939 306 3163 322
rect 2939 272 2941 306
rect 2975 288 3163 306
rect 3197 332 3284 348
rect 3197 298 3213 332
rect 3247 298 3284 332
rect 2975 272 2991 288
rect 3197 282 3284 298
rect 3318 342 3431 358
rect 3318 308 3334 342
rect 3368 308 3431 342
rect 3318 292 3431 308
rect 2939 256 2991 272
rect 3465 258 3499 402
rect 3318 224 3499 258
rect 3579 420 3698 436
rect 3579 386 3648 420
rect 3682 386 3698 420
rect 3579 370 3698 386
rect 3747 416 3797 436
rect 3747 382 3763 416
rect 3221 222 3352 224
rect 2871 190 3352 222
rect 3579 190 3613 370
rect 3747 363 3797 382
rect 3647 274 3713 290
rect 3647 240 3663 274
rect 3697 240 3713 274
rect 3647 224 3713 240
rect 3747 229 3781 363
rect 3831 329 3865 470
rect 3899 476 3915 510
rect 3949 476 3965 510
rect 3899 413 3965 476
rect 3899 379 3915 413
rect 3949 379 3965 413
rect 3899 363 3965 379
rect 3999 599 4065 615
rect 3999 565 4015 599
rect 4049 565 4065 599
rect 3999 506 4065 565
rect 3999 472 4015 506
rect 4049 472 4065 506
rect 3999 430 4065 472
rect 3999 413 4107 430
rect 3999 379 4015 413
rect 4049 379 4107 413
rect 3999 363 4107 379
rect 3815 313 3869 329
rect 3815 279 3825 313
rect 3859 279 3869 313
rect 3815 263 3869 279
rect 3903 313 4004 329
rect 3903 279 3954 313
rect 3988 279 4004 313
rect 3903 263 4004 279
rect 3903 229 3937 263
rect 3747 195 3937 229
rect 2871 188 3287 190
rect 3221 169 3287 188
rect 2803 143 3063 154
rect 2803 120 3013 143
rect 2997 109 3013 120
rect 3047 109 3063 143
rect 3221 135 3237 169
rect 3271 135 3287 169
rect 3221 119 3287 135
rect 3386 156 3669 190
rect 2997 85 3063 109
rect 3386 85 3420 156
rect 3603 132 3669 156
rect 2997 51 3420 85
rect 3495 103 3561 122
rect 3495 69 3511 103
rect 3545 69 3561 103
rect 3603 98 3619 132
rect 3653 98 3669 132
rect 3603 69 3669 98
rect 3761 132 3811 161
rect 3761 98 3777 132
rect 3495 17 3561 69
rect 3761 17 3811 98
rect 3847 132 3937 195
rect 3847 98 3863 132
rect 3897 98 3937 132
rect 3847 69 3937 98
rect 3971 213 4005 229
rect 3971 103 4005 179
rect 3971 17 4005 69
rect 4041 213 4107 363
rect 4041 179 4057 213
rect 4091 179 4107 213
rect 4041 103 4107 179
rect 4041 69 4057 103
rect 4091 69 4107 103
rect 4041 53 4107 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4128 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 3583 649 3617 683
rect 3679 649 3713 683
rect 3775 649 3809 683
rect 3871 649 3905 683
rect 3967 649 4001 683
rect 4063 649 4097 683
rect 2911 547 2945 581
rect 3295 575 3329 581
rect 3295 547 3306 575
rect 3306 547 3329 575
rect 3391 547 3425 581
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
rect 4063 -17 4097 17
<< metal1 >>
rect 0 683 4128 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3775 683
rect 3809 649 3871 683
rect 3905 649 3967 683
rect 4001 649 4063 683
rect 4097 649 4128 683
rect 0 617 4128 649
rect 14 581 4114 589
rect 14 547 2911 581
rect 2945 547 3295 581
rect 3329 547 3391 581
rect 3425 547 4114 581
rect 14 535 4114 547
rect 0 17 4128 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4128 17
rect 0 -49 4128 -17
<< labels >>
flabel pwell s 0 0 4128 49 0 FreeSans 200 0 0 0 VNB
port 9 nsew ground bidirectional
flabel nwell s 0 617 4128 666 0 FreeSans 200 0 0 0 VPB
port 10 nsew power bidirectional
rlabel comment s 0 0 0 0 4 srsdfrtp_1
flabel metal1 s 14 535 4114 589 0 FreeSans 340 0 0 0 KAPWR
port 7 nsew power bidirectional
flabel metal1 s 0 617 4128 666 0 FreeSans 340 0 0 0 VPWR
port 11 nsew power bidirectional
flabel metal1 s 0 0 4128 49 0 FreeSans 340 0 0 0 VGND
port 8 nsew ground bidirectional
flabel locali s 3679 242 3713 276 0 FreeSans 340 0 0 0 SLEEP_B
port 6 nsew signal input
flabel locali s 3391 316 3425 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 4063 94 4097 128 0 FreeSans 340 0 0 0 Q
port 12 nsew signal output
flabel locali s 4063 168 4097 202 0 FreeSans 340 0 0 0 Q
port 12 nsew signal output
flabel locali s 4063 242 4097 276 0 FreeSans 340 0 0 0 Q
port 12 nsew signal output
flabel locali s 4063 316 4097 350 0 FreeSans 340 0 0 0 Q
port 12 nsew signal output
flabel locali s 4063 390 4097 424 0 FreeSans 340 0 0 0 Q
port 12 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 4128 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5771440
string GDS_START 5747634
<< end >>
