magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 34 49 824 243
rect 0 0 864 49
<< scnmos >>
rect 113 49 143 217
rect 287 49 317 217
rect 373 49 403 217
rect 481 49 511 217
rect 643 49 673 217
rect 715 49 745 217
<< scpmoshvt >>
rect 105 367 135 619
rect 295 367 325 619
rect 373 367 403 619
rect 481 367 511 619
rect 635 367 665 619
rect 721 367 751 619
<< ndiff >>
rect 60 205 113 217
rect 60 171 68 205
rect 102 171 113 205
rect 60 101 113 171
rect 60 67 68 101
rect 102 67 113 101
rect 60 49 113 67
rect 143 159 287 217
rect 143 125 154 159
rect 188 125 242 159
rect 276 125 287 159
rect 143 91 287 125
rect 143 57 154 91
rect 188 57 242 91
rect 276 57 287 91
rect 143 49 287 57
rect 317 205 373 217
rect 317 171 328 205
rect 362 171 373 205
rect 317 101 373 171
rect 317 67 328 101
rect 362 67 373 101
rect 317 49 373 67
rect 403 165 481 217
rect 403 131 422 165
rect 456 131 481 165
rect 403 91 481 131
rect 403 57 422 91
rect 456 57 481 91
rect 403 49 481 57
rect 511 205 643 217
rect 511 171 522 205
rect 556 171 598 205
rect 632 171 643 205
rect 511 101 643 171
rect 511 67 522 101
rect 556 67 598 101
rect 632 67 643 101
rect 511 49 643 67
rect 673 49 715 217
rect 745 205 798 217
rect 745 171 756 205
rect 790 171 798 205
rect 745 95 798 171
rect 745 61 756 95
rect 790 61 798 95
rect 745 49 798 61
<< pdiff >>
rect 52 599 105 619
rect 52 565 60 599
rect 94 565 105 599
rect 52 504 105 565
rect 52 470 60 504
rect 94 470 105 504
rect 52 413 105 470
rect 52 379 60 413
rect 94 379 105 413
rect 52 367 105 379
rect 135 607 188 619
rect 135 573 146 607
rect 180 573 188 607
rect 135 490 188 573
rect 135 456 146 490
rect 180 456 188 490
rect 135 367 188 456
rect 242 599 295 619
rect 242 565 250 599
rect 284 565 295 599
rect 242 518 295 565
rect 242 484 250 518
rect 284 484 295 518
rect 242 436 295 484
rect 242 402 250 436
rect 284 402 295 436
rect 242 367 295 402
rect 325 367 373 619
rect 403 367 481 619
rect 511 599 635 619
rect 511 565 522 599
rect 556 565 590 599
rect 624 565 635 599
rect 511 512 635 565
rect 511 478 522 512
rect 556 478 590 512
rect 624 478 635 512
rect 511 420 635 478
rect 511 386 522 420
rect 556 386 590 420
rect 624 386 635 420
rect 511 367 635 386
rect 665 611 721 619
rect 665 577 676 611
rect 710 577 721 611
rect 665 492 721 577
rect 665 458 676 492
rect 710 458 721 492
rect 665 367 721 458
rect 751 599 804 619
rect 751 565 762 599
rect 796 565 804 599
rect 751 512 804 565
rect 751 478 762 512
rect 796 478 804 512
rect 751 420 804 478
rect 751 386 762 420
rect 796 386 804 420
rect 751 367 804 386
<< ndiffc >>
rect 68 171 102 205
rect 68 67 102 101
rect 154 125 188 159
rect 242 125 276 159
rect 154 57 188 91
rect 242 57 276 91
rect 328 171 362 205
rect 328 67 362 101
rect 422 131 456 165
rect 422 57 456 91
rect 522 171 556 205
rect 598 171 632 205
rect 522 67 556 101
rect 598 67 632 101
rect 756 171 790 205
rect 756 61 790 95
<< pdiffc >>
rect 60 565 94 599
rect 60 470 94 504
rect 60 379 94 413
rect 146 573 180 607
rect 146 456 180 490
rect 250 565 284 599
rect 250 484 284 518
rect 250 402 284 436
rect 522 565 556 599
rect 590 565 624 599
rect 522 478 556 512
rect 590 478 624 512
rect 522 386 556 420
rect 590 386 624 420
rect 676 577 710 611
rect 676 458 710 492
rect 762 565 796 599
rect 762 478 796 512
rect 762 386 796 420
<< poly >>
rect 105 619 135 645
rect 295 619 325 645
rect 373 619 403 645
rect 481 619 511 645
rect 635 619 665 645
rect 721 619 751 645
rect 105 305 135 367
rect 295 335 325 367
rect 259 319 325 335
rect 105 289 192 305
rect 105 255 142 289
rect 176 255 192 289
rect 259 285 275 319
rect 309 285 325 319
rect 259 269 325 285
rect 373 335 403 367
rect 481 335 511 367
rect 373 319 439 335
rect 373 285 389 319
rect 423 285 439 319
rect 373 269 439 285
rect 481 319 559 335
rect 481 285 503 319
rect 537 285 559 319
rect 635 308 665 367
rect 721 308 751 367
rect 481 269 559 285
rect 601 292 673 308
rect 105 239 192 255
rect 113 217 143 239
rect 287 217 317 269
rect 373 217 403 269
rect 481 217 511 269
rect 601 258 623 292
rect 657 258 673 292
rect 601 242 673 258
rect 643 217 673 242
rect 715 292 823 308
rect 715 258 773 292
rect 807 258 823 292
rect 715 242 823 258
rect 715 217 745 242
rect 113 23 143 49
rect 287 23 317 49
rect 373 23 403 49
rect 481 23 511 49
rect 643 23 673 49
rect 715 23 745 49
<< polycont >>
rect 142 255 176 289
rect 275 285 309 319
rect 389 285 423 319
rect 503 285 537 319
rect 623 258 657 292
rect 773 258 807 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 17 599 96 615
rect 17 565 60 599
rect 94 565 96 599
rect 17 504 96 565
rect 17 470 60 504
rect 94 470 96 504
rect 17 413 96 470
rect 130 607 196 649
rect 130 573 146 607
rect 180 573 196 607
rect 130 490 196 573
rect 130 456 146 490
rect 180 456 196 490
rect 130 452 196 456
rect 234 599 300 615
rect 234 565 250 599
rect 284 565 300 599
rect 506 599 626 615
rect 234 518 300 565
rect 234 484 250 518
rect 284 484 300 518
rect 234 436 300 484
rect 234 418 250 436
rect 17 379 60 413
rect 94 379 96 413
rect 17 355 96 379
rect 138 402 250 418
rect 284 402 300 436
rect 138 384 300 402
rect 17 205 104 355
rect 17 171 68 205
rect 102 171 104 205
rect 138 289 181 384
rect 138 255 142 289
rect 176 255 181 289
rect 215 319 355 350
rect 215 285 275 319
rect 309 285 355 319
rect 215 267 355 285
rect 389 319 453 592
rect 506 565 522 599
rect 556 565 590 599
rect 624 565 626 599
rect 506 512 626 565
rect 506 478 522 512
rect 556 478 590 512
rect 624 478 626 512
rect 506 420 626 478
rect 660 611 726 649
rect 660 577 676 611
rect 710 577 726 611
rect 660 492 726 577
rect 660 458 676 492
rect 710 458 726 492
rect 660 454 726 458
rect 760 599 812 615
rect 760 565 762 599
rect 796 565 812 599
rect 760 512 812 565
rect 760 478 762 512
rect 796 478 812 512
rect 760 420 812 478
rect 506 386 522 420
rect 556 386 590 420
rect 624 386 762 420
rect 796 386 812 420
rect 423 285 453 319
rect 389 267 453 285
rect 487 319 564 350
rect 487 285 503 319
rect 537 285 564 319
rect 487 267 564 285
rect 598 292 739 352
rect 138 233 181 255
rect 598 258 623 292
rect 657 258 739 292
rect 598 242 739 258
rect 773 292 847 352
rect 807 258 847 292
rect 773 242 847 258
rect 138 208 564 233
rect 138 205 648 208
rect 138 199 328 205
rect 17 101 104 171
rect 326 171 328 199
rect 362 199 522 205
rect 362 171 372 199
rect 17 67 68 101
rect 102 67 104 101
rect 17 51 104 67
rect 138 159 292 165
rect 138 125 154 159
rect 188 125 242 159
rect 276 125 292 159
rect 138 91 292 125
rect 138 57 154 91
rect 188 57 242 91
rect 276 57 292 91
rect 138 17 292 57
rect 326 101 372 171
rect 506 171 522 199
rect 556 171 598 205
rect 632 171 648 205
rect 326 67 328 101
rect 362 67 372 101
rect 326 51 372 67
rect 406 131 422 165
rect 456 131 472 165
rect 406 91 472 131
rect 406 57 422 91
rect 456 57 472 91
rect 406 17 472 57
rect 506 101 648 171
rect 506 67 522 101
rect 556 67 598 101
rect 632 67 648 101
rect 506 51 648 67
rect 740 205 806 208
rect 740 171 756 205
rect 790 171 806 205
rect 740 95 806 171
rect 740 61 756 95
rect 790 61 806 95
rect 740 17 806 61
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2111o_1
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1095350
string GDS_START 1085984
<< end >>
