magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2930 1975
<< nwell >>
rect -38 331 1670 704
rect 874 309 1168 331
<< pwell >>
rect 2 241 448 243
rect 2 49 1616 241
rect 0 0 1632 49
<< scnmos >>
rect 81 49 111 217
rect 167 49 197 217
rect 253 49 283 217
rect 339 49 369 217
rect 529 47 559 215
rect 615 47 645 215
rect 701 47 731 215
rect 787 47 817 215
rect 977 47 1007 215
rect 1163 47 1193 215
rect 1249 47 1279 215
rect 1335 47 1365 215
rect 1421 47 1451 215
rect 1507 47 1537 215
<< scpmoshvt >>
rect 156 367 186 619
rect 242 367 272 619
rect 328 367 358 619
rect 414 367 444 619
rect 500 367 530 619
rect 586 367 616 619
rect 687 367 717 619
rect 773 367 803 619
rect 963 345 993 597
rect 1049 345 1079 597
rect 1249 367 1279 619
rect 1335 367 1365 619
rect 1421 367 1451 619
rect 1507 367 1537 619
<< ndiff >>
rect 28 173 81 217
rect 28 139 36 173
rect 70 139 81 173
rect 28 95 81 139
rect 28 61 36 95
rect 70 61 81 95
rect 28 49 81 61
rect 111 205 167 217
rect 111 171 122 205
rect 156 171 167 205
rect 111 101 167 171
rect 111 67 122 101
rect 156 67 167 101
rect 111 49 167 67
rect 197 175 253 217
rect 197 141 208 175
rect 242 141 253 175
rect 197 91 253 141
rect 197 57 208 91
rect 242 57 253 91
rect 197 49 253 57
rect 283 205 339 217
rect 283 171 294 205
rect 328 171 339 205
rect 283 101 339 171
rect 283 67 294 101
rect 328 67 339 101
rect 283 49 339 67
rect 369 205 422 217
rect 369 171 380 205
rect 414 171 422 205
rect 369 95 422 171
rect 369 61 380 95
rect 414 61 422 95
rect 369 49 422 61
rect 476 101 529 215
rect 476 67 484 101
rect 518 67 529 101
rect 476 47 529 67
rect 559 193 615 215
rect 559 159 570 193
rect 604 159 615 193
rect 559 47 615 159
rect 645 189 701 215
rect 645 155 656 189
rect 690 155 701 189
rect 645 101 701 155
rect 645 67 656 101
rect 690 67 701 101
rect 645 47 701 67
rect 731 169 787 215
rect 731 135 742 169
rect 776 135 787 169
rect 731 47 787 135
rect 817 121 870 215
rect 817 87 828 121
rect 862 87 870 121
rect 817 47 870 87
rect 924 192 977 215
rect 924 158 932 192
rect 966 158 977 192
rect 924 101 977 158
rect 924 67 932 101
rect 966 67 977 101
rect 924 47 977 67
rect 1007 130 1163 215
rect 1007 96 1018 130
rect 1052 96 1118 130
rect 1152 96 1163 130
rect 1007 47 1163 96
rect 1193 203 1249 215
rect 1193 169 1204 203
rect 1238 169 1249 203
rect 1193 101 1249 169
rect 1193 67 1204 101
rect 1238 67 1249 101
rect 1193 47 1249 67
rect 1279 183 1335 215
rect 1279 149 1290 183
rect 1324 149 1335 183
rect 1279 93 1335 149
rect 1279 59 1290 93
rect 1324 59 1335 93
rect 1279 47 1335 59
rect 1365 203 1421 215
rect 1365 169 1376 203
rect 1410 169 1421 203
rect 1365 101 1421 169
rect 1365 67 1376 101
rect 1410 67 1421 101
rect 1365 47 1421 67
rect 1451 183 1507 215
rect 1451 149 1462 183
rect 1496 149 1507 183
rect 1451 93 1507 149
rect 1451 59 1462 93
rect 1496 59 1507 93
rect 1451 47 1507 59
rect 1537 203 1590 215
rect 1537 169 1548 203
rect 1582 169 1590 203
rect 1537 101 1590 169
rect 1537 67 1548 101
rect 1582 67 1590 101
rect 1537 47 1590 67
<< pdiff >>
rect 103 607 156 619
rect 103 573 111 607
rect 145 573 156 607
rect 103 528 156 573
rect 103 494 111 528
rect 145 494 156 528
rect 103 453 156 494
rect 103 419 111 453
rect 145 419 156 453
rect 103 367 156 419
rect 186 599 242 619
rect 186 565 197 599
rect 231 565 242 599
rect 186 506 242 565
rect 186 472 197 506
rect 231 472 242 506
rect 186 413 242 472
rect 186 379 197 413
rect 231 379 242 413
rect 186 367 242 379
rect 272 607 328 619
rect 272 573 283 607
rect 317 573 328 607
rect 272 528 328 573
rect 272 494 283 528
rect 317 494 328 528
rect 272 455 328 494
rect 272 421 283 455
rect 317 421 328 455
rect 272 367 328 421
rect 358 599 414 619
rect 358 565 369 599
rect 403 565 414 599
rect 358 506 414 565
rect 358 472 369 506
rect 403 472 414 506
rect 358 413 414 472
rect 358 379 369 413
rect 403 379 414 413
rect 358 367 414 379
rect 444 607 500 619
rect 444 573 455 607
rect 489 573 500 607
rect 444 525 500 573
rect 444 491 455 525
rect 489 491 500 525
rect 444 443 500 491
rect 444 409 455 443
rect 489 409 500 443
rect 444 367 500 409
rect 530 599 586 619
rect 530 565 541 599
rect 575 565 586 599
rect 530 506 586 565
rect 530 472 541 506
rect 575 472 586 506
rect 530 413 586 472
rect 530 379 541 413
rect 575 379 586 413
rect 530 367 586 379
rect 616 607 687 619
rect 616 573 635 607
rect 669 573 687 607
rect 616 525 687 573
rect 616 491 635 525
rect 669 491 687 525
rect 616 443 687 491
rect 616 409 635 443
rect 669 409 687 443
rect 616 367 687 409
rect 717 599 773 619
rect 717 565 728 599
rect 762 565 773 599
rect 717 506 773 565
rect 717 472 728 506
rect 762 472 773 506
rect 717 413 773 472
rect 717 379 728 413
rect 762 379 773 413
rect 717 367 773 379
rect 803 607 856 619
rect 803 573 814 607
rect 848 573 856 607
rect 803 525 856 573
rect 803 491 814 525
rect 848 491 856 525
rect 803 443 856 491
rect 803 409 814 443
rect 848 409 856 443
rect 803 367 856 409
rect 910 585 963 597
rect 910 551 918 585
rect 952 551 963 585
rect 910 517 963 551
rect 910 483 918 517
rect 952 483 963 517
rect 910 443 963 483
rect 910 409 918 443
rect 952 409 963 443
rect 910 345 963 409
rect 993 531 1049 597
rect 993 497 1004 531
rect 1038 497 1049 531
rect 993 463 1049 497
rect 993 429 1004 463
rect 1038 429 1049 463
rect 993 391 1049 429
rect 993 357 1004 391
rect 1038 357 1049 391
rect 993 345 1049 357
rect 1079 585 1132 597
rect 1079 551 1090 585
rect 1124 551 1132 585
rect 1079 484 1132 551
rect 1079 450 1090 484
rect 1124 450 1132 484
rect 1079 391 1132 450
rect 1079 357 1090 391
rect 1124 357 1132 391
rect 1196 531 1249 619
rect 1196 497 1204 531
rect 1238 497 1249 531
rect 1196 420 1249 497
rect 1196 386 1204 420
rect 1238 386 1249 420
rect 1196 367 1249 386
rect 1279 599 1335 619
rect 1279 565 1290 599
rect 1324 565 1335 599
rect 1279 495 1335 565
rect 1279 461 1290 495
rect 1324 461 1335 495
rect 1279 367 1335 461
rect 1365 599 1421 619
rect 1365 565 1376 599
rect 1410 565 1421 599
rect 1365 504 1421 565
rect 1365 470 1376 504
rect 1410 470 1421 504
rect 1365 420 1421 470
rect 1365 386 1376 420
rect 1410 386 1421 420
rect 1365 367 1421 386
rect 1451 607 1507 619
rect 1451 573 1462 607
rect 1496 573 1507 607
rect 1451 495 1507 573
rect 1451 461 1462 495
rect 1496 461 1507 495
rect 1451 367 1507 461
rect 1537 599 1590 619
rect 1537 565 1548 599
rect 1582 565 1590 599
rect 1537 507 1590 565
rect 1537 473 1548 507
rect 1582 473 1590 507
rect 1537 420 1590 473
rect 1537 386 1548 420
rect 1582 386 1590 420
rect 1537 367 1590 386
rect 1079 345 1132 357
<< ndiffc >>
rect 36 139 70 173
rect 36 61 70 95
rect 122 171 156 205
rect 122 67 156 101
rect 208 141 242 175
rect 208 57 242 91
rect 294 171 328 205
rect 294 67 328 101
rect 380 171 414 205
rect 380 61 414 95
rect 484 67 518 101
rect 570 159 604 193
rect 656 155 690 189
rect 656 67 690 101
rect 742 135 776 169
rect 828 87 862 121
rect 932 158 966 192
rect 932 67 966 101
rect 1018 96 1052 130
rect 1118 96 1152 130
rect 1204 169 1238 203
rect 1204 67 1238 101
rect 1290 149 1324 183
rect 1290 59 1324 93
rect 1376 169 1410 203
rect 1376 67 1410 101
rect 1462 149 1496 183
rect 1462 59 1496 93
rect 1548 169 1582 203
rect 1548 67 1582 101
<< pdiffc >>
rect 111 573 145 607
rect 111 494 145 528
rect 111 419 145 453
rect 197 565 231 599
rect 197 472 231 506
rect 197 379 231 413
rect 283 573 317 607
rect 283 494 317 528
rect 283 421 317 455
rect 369 565 403 599
rect 369 472 403 506
rect 369 379 403 413
rect 455 573 489 607
rect 455 491 489 525
rect 455 409 489 443
rect 541 565 575 599
rect 541 472 575 506
rect 541 379 575 413
rect 635 573 669 607
rect 635 491 669 525
rect 635 409 669 443
rect 728 565 762 599
rect 728 472 762 506
rect 728 379 762 413
rect 814 573 848 607
rect 814 491 848 525
rect 814 409 848 443
rect 918 551 952 585
rect 918 483 952 517
rect 918 409 952 443
rect 1004 497 1038 531
rect 1004 429 1038 463
rect 1004 357 1038 391
rect 1090 551 1124 585
rect 1090 450 1124 484
rect 1090 357 1124 391
rect 1204 497 1238 531
rect 1204 386 1238 420
rect 1290 565 1324 599
rect 1290 461 1324 495
rect 1376 565 1410 599
rect 1376 470 1410 504
rect 1376 386 1410 420
rect 1462 573 1496 607
rect 1462 461 1496 495
rect 1548 565 1582 599
rect 1548 473 1582 507
rect 1548 386 1582 420
<< poly >>
rect 156 619 186 645
rect 242 619 272 645
rect 328 619 358 645
rect 414 619 444 645
rect 500 619 530 645
rect 586 619 616 645
rect 687 619 717 645
rect 773 619 803 645
rect 963 597 993 623
rect 1049 597 1079 623
rect 1249 619 1279 645
rect 1335 619 1365 645
rect 1421 619 1451 645
rect 1507 619 1537 645
rect 156 331 186 367
rect 242 331 272 367
rect 328 331 358 367
rect 414 331 444 367
rect 81 315 444 331
rect 81 281 122 315
rect 156 281 190 315
rect 224 281 258 315
rect 292 281 326 315
rect 360 281 394 315
rect 428 281 444 315
rect 81 265 444 281
rect 500 305 530 367
rect 586 305 616 367
rect 687 315 717 367
rect 773 315 803 367
rect 500 289 645 305
rect 500 275 595 289
rect 81 217 111 265
rect 167 217 197 265
rect 253 217 283 265
rect 339 217 369 265
rect 529 255 595 275
rect 629 255 645 289
rect 529 237 645 255
rect 687 289 817 315
rect 687 255 703 289
rect 737 255 817 289
rect 687 239 817 255
rect 529 215 559 237
rect 615 215 645 237
rect 701 215 731 239
rect 787 215 817 239
rect 963 303 993 345
rect 1049 303 1079 345
rect 1249 335 1279 367
rect 1335 335 1365 367
rect 1249 319 1365 335
rect 963 287 1193 303
rect 963 253 979 287
rect 1013 253 1065 287
rect 1099 253 1193 287
rect 963 237 1193 253
rect 977 215 1007 237
rect 1163 215 1193 237
rect 1249 285 1265 319
rect 1299 285 1365 319
rect 1249 269 1365 285
rect 1249 215 1279 269
rect 1335 215 1365 269
rect 1421 335 1451 367
rect 1507 335 1537 367
rect 1421 319 1537 335
rect 1421 285 1487 319
rect 1521 285 1537 319
rect 1421 269 1537 285
rect 1421 215 1451 269
rect 1507 215 1537 269
rect 81 23 111 49
rect 167 23 197 49
rect 253 23 283 49
rect 339 23 369 49
rect 529 21 559 47
rect 615 21 645 47
rect 701 21 731 47
rect 787 21 817 47
rect 977 21 1007 47
rect 1163 21 1193 47
rect 1249 21 1279 47
rect 1335 21 1365 47
rect 1421 21 1451 47
rect 1507 21 1537 47
<< polycont >>
rect 122 281 156 315
rect 190 281 224 315
rect 258 281 292 315
rect 326 281 360 315
rect 394 281 428 315
rect 595 255 629 289
rect 703 255 737 289
rect 979 253 1013 287
rect 1065 253 1099 287
rect 1265 285 1299 319
rect 1487 285 1521 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 95 607 161 649
rect 95 573 111 607
rect 145 573 161 607
rect 95 528 161 573
rect 95 494 111 528
rect 145 494 161 528
rect 95 453 161 494
rect 95 419 111 453
rect 145 419 161 453
rect 195 599 233 615
rect 195 565 197 599
rect 231 565 233 599
rect 195 506 233 565
rect 195 472 197 506
rect 231 472 233 506
rect 195 413 233 472
rect 267 607 333 649
rect 267 573 283 607
rect 317 573 333 607
rect 267 528 333 573
rect 267 494 283 528
rect 317 494 333 528
rect 267 455 333 494
rect 267 421 283 455
rect 317 421 333 455
rect 367 599 405 615
rect 367 565 369 599
rect 403 565 405 599
rect 367 506 405 565
rect 367 472 369 506
rect 403 472 405 506
rect 195 385 197 413
rect 17 379 197 385
rect 231 385 233 413
rect 367 413 405 472
rect 367 385 369 413
rect 231 379 369 385
rect 403 379 405 413
rect 439 607 505 649
rect 439 573 455 607
rect 489 573 505 607
rect 439 525 505 573
rect 439 491 455 525
rect 489 491 505 525
rect 439 443 505 491
rect 439 409 455 443
rect 489 409 505 443
rect 539 599 585 615
rect 539 565 541 599
rect 575 565 585 599
rect 539 506 585 565
rect 539 472 541 506
rect 575 472 585 506
rect 539 413 585 472
rect 17 351 405 379
rect 539 379 541 413
rect 575 379 585 413
rect 619 607 685 649
rect 619 573 635 607
rect 669 573 685 607
rect 619 525 685 573
rect 619 491 635 525
rect 669 491 685 525
rect 619 443 685 491
rect 619 409 635 443
rect 669 409 685 443
rect 719 599 764 615
rect 719 565 728 599
rect 762 565 764 599
rect 719 506 764 565
rect 719 472 728 506
rect 762 472 764 506
rect 719 413 764 472
rect 539 375 585 379
rect 719 379 728 413
rect 762 379 764 413
rect 798 607 864 649
rect 798 573 814 607
rect 848 573 864 607
rect 798 525 864 573
rect 798 491 814 525
rect 848 491 864 525
rect 798 443 864 491
rect 798 409 814 443
rect 848 409 864 443
rect 902 599 1340 615
rect 902 585 1290 599
rect 902 551 918 585
rect 952 581 1090 585
rect 952 551 968 581
rect 902 517 968 551
rect 1081 551 1090 581
rect 1124 581 1290 585
rect 1124 551 1136 581
rect 902 483 918 517
rect 952 483 968 517
rect 902 443 968 483
rect 902 409 918 443
rect 952 409 968 443
rect 1002 531 1047 547
rect 1002 497 1004 531
rect 1038 497 1047 531
rect 1002 463 1047 497
rect 1002 429 1004 463
rect 1038 429 1047 463
rect 719 375 764 379
rect 1002 391 1047 429
rect 1002 375 1004 391
rect 439 357 1004 375
rect 1038 357 1047 391
rect 17 247 72 351
rect 439 341 1047 357
rect 1081 484 1136 551
rect 1274 565 1290 581
rect 1324 565 1340 599
rect 1081 450 1090 484
rect 1124 450 1136 484
rect 1081 391 1136 450
rect 1081 357 1090 391
rect 1124 357 1136 391
rect 1188 531 1240 547
rect 1188 497 1204 531
rect 1238 497 1240 531
rect 1188 420 1240 497
rect 1274 495 1340 565
rect 1274 461 1290 495
rect 1324 461 1340 495
rect 1274 454 1340 461
rect 1374 599 1412 615
rect 1374 565 1376 599
rect 1410 565 1412 599
rect 1374 504 1412 565
rect 1374 470 1376 504
rect 1410 470 1412 504
rect 1374 420 1412 470
rect 1446 607 1512 649
rect 1446 573 1462 607
rect 1496 573 1512 607
rect 1446 495 1512 573
rect 1446 461 1462 495
rect 1496 461 1512 495
rect 1446 454 1512 461
rect 1546 599 1598 615
rect 1546 565 1548 599
rect 1582 565 1598 599
rect 1546 507 1598 565
rect 1546 473 1548 507
rect 1582 473 1598 507
rect 1546 420 1598 473
rect 1188 386 1204 420
rect 1238 386 1376 420
rect 1410 386 1548 420
rect 1582 386 1598 420
rect 1081 341 1136 357
rect 439 317 559 341
rect 106 315 559 317
rect 106 281 122 315
rect 156 281 190 315
rect 224 281 258 315
rect 292 281 326 315
rect 360 281 394 315
rect 428 281 559 315
rect 1170 319 1423 352
rect 17 213 338 247
rect 17 211 158 213
rect 120 205 158 211
rect 20 173 86 177
rect 20 139 36 173
rect 70 139 86 173
rect 20 95 86 139
rect 20 61 36 95
rect 70 61 86 95
rect 20 17 86 61
rect 120 171 122 205
rect 156 171 158 205
rect 292 205 338 213
rect 120 101 158 171
rect 120 67 122 101
rect 156 67 158 101
rect 120 51 158 67
rect 192 175 258 179
rect 192 141 208 175
rect 242 141 258 175
rect 192 91 258 141
rect 192 57 208 91
rect 242 57 258 91
rect 192 17 258 57
rect 292 171 294 205
rect 328 171 338 205
rect 292 101 338 171
rect 292 67 294 101
rect 328 67 338 101
rect 292 51 338 67
rect 372 205 430 221
rect 372 171 380 205
rect 414 171 430 205
rect 372 95 430 171
rect 464 203 559 281
rect 593 289 653 305
rect 593 255 595 289
rect 629 255 653 289
rect 593 239 653 255
rect 687 289 757 305
rect 687 255 703 289
rect 737 255 757 289
rect 687 239 757 255
rect 791 287 1136 303
rect 791 253 979 287
rect 1013 253 1065 287
rect 1099 253 1136 287
rect 1170 285 1265 319
rect 1299 285 1423 319
rect 1457 319 1615 352
rect 1457 285 1487 319
rect 1521 285 1615 319
rect 791 242 1136 253
rect 1200 217 1598 251
rect 1200 208 1240 217
rect 791 205 1240 208
rect 464 193 620 203
rect 464 159 570 193
rect 604 159 620 193
rect 464 153 620 159
rect 654 189 692 205
rect 654 155 656 189
rect 690 155 692 189
rect 654 119 692 155
rect 726 203 1240 205
rect 726 192 1204 203
rect 726 171 932 192
rect 726 169 792 171
rect 726 135 742 169
rect 776 135 792 169
rect 916 158 932 171
rect 966 174 1204 192
rect 966 158 968 174
rect 726 123 792 135
rect 372 61 380 95
rect 414 61 430 95
rect 372 17 430 61
rect 468 101 692 119
rect 468 67 484 101
rect 518 67 656 101
rect 690 87 692 101
rect 826 121 878 137
rect 826 87 828 121
rect 862 87 878 121
rect 690 67 878 87
rect 468 51 878 67
rect 916 101 968 158
rect 1202 169 1204 174
rect 1238 169 1240 203
rect 1374 203 1412 217
rect 916 67 932 101
rect 966 67 968 101
rect 916 51 968 67
rect 1002 130 1168 140
rect 1002 96 1018 130
rect 1052 96 1118 130
rect 1152 96 1168 130
rect 1002 17 1168 96
rect 1202 101 1240 169
rect 1202 67 1204 101
rect 1238 67 1240 101
rect 1202 51 1240 67
rect 1274 149 1290 183
rect 1324 149 1340 183
rect 1274 93 1340 149
rect 1274 59 1290 93
rect 1324 59 1340 93
rect 1274 17 1340 59
rect 1374 169 1376 203
rect 1410 169 1412 203
rect 1546 203 1598 217
rect 1374 101 1412 169
rect 1374 67 1376 101
rect 1410 67 1412 101
rect 1374 51 1412 67
rect 1446 149 1462 183
rect 1496 149 1512 183
rect 1446 93 1512 149
rect 1446 59 1462 93
rect 1496 59 1512 93
rect 1446 17 1512 59
rect 1546 169 1548 203
rect 1582 169 1598 203
rect 1546 101 1598 169
rect 1546 67 1548 101
rect 1582 67 1598 101
rect 1546 51 1598 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 683 1632 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1632 683
rect 0 617 1632 649
rect 0 17 1632 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -49 1632 -17
<< labels >>
flabel pwell s 0 0 1632 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 1632 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o311a_4
flabel metal1 s 0 617 1632 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 1632 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1632 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4392476
string GDS_START 4378248
<< end >>
