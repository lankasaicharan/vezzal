magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 18 261 296 263
rect 18 241 1179 261
rect 18 49 2015 241
rect 0 0 2016 49
<< scnmos >>
rect 101 69 131 237
rect 187 69 217 237
rect 404 67 434 235
rect 490 67 520 235
rect 608 67 638 235
rect 694 67 724 235
rect 812 67 842 235
rect 898 67 928 235
rect 984 67 1014 235
rect 1070 67 1100 235
rect 1304 47 1334 215
rect 1390 47 1420 215
rect 1476 47 1506 215
rect 1562 47 1592 215
rect 1648 47 1678 215
rect 1734 47 1764 215
rect 1820 47 1850 215
rect 1906 47 1936 215
<< scpmoshvt >>
rect 101 367 131 619
rect 187 367 217 619
rect 430 367 460 619
rect 516 367 546 619
rect 602 367 632 619
rect 688 367 718 619
rect 774 367 804 619
rect 860 367 890 619
rect 946 367 976 619
rect 1032 367 1062 619
rect 1298 367 1328 619
rect 1384 367 1414 619
rect 1470 367 1500 619
rect 1556 367 1586 619
rect 1642 367 1672 619
rect 1728 367 1758 619
rect 1814 367 1844 619
rect 1900 367 1930 619
<< ndiff >>
rect 44 192 101 237
rect 44 158 52 192
rect 86 158 101 192
rect 44 115 101 158
rect 44 81 52 115
rect 86 81 101 115
rect 44 69 101 81
rect 131 208 187 237
rect 131 174 142 208
rect 176 174 187 208
rect 131 111 187 174
rect 131 77 142 111
rect 176 77 187 111
rect 131 69 187 77
rect 217 192 270 237
rect 217 158 228 192
rect 262 158 270 192
rect 217 115 270 158
rect 217 81 228 115
rect 262 81 270 115
rect 217 69 270 81
rect 324 87 404 235
rect 324 53 336 87
rect 370 67 404 87
rect 434 227 490 235
rect 434 193 445 227
rect 479 193 490 227
rect 434 67 490 193
rect 520 87 608 235
rect 520 67 547 87
rect 370 53 382 67
rect 324 45 382 53
rect 535 53 547 67
rect 581 67 608 87
rect 638 227 694 235
rect 638 193 649 227
rect 683 193 694 227
rect 638 67 694 193
rect 724 87 812 235
rect 724 67 751 87
rect 581 53 593 67
rect 535 45 593 53
rect 739 53 751 67
rect 785 67 812 87
rect 842 227 898 235
rect 842 193 853 227
rect 887 193 898 227
rect 842 67 898 193
rect 928 177 984 235
rect 928 143 939 177
rect 973 143 984 177
rect 928 109 984 143
rect 928 75 939 109
rect 973 75 984 109
rect 928 67 984 75
rect 1014 222 1070 235
rect 1014 188 1025 222
rect 1059 188 1070 222
rect 1014 67 1070 188
rect 1100 142 1153 235
rect 1100 108 1111 142
rect 1145 108 1153 142
rect 1100 67 1153 108
rect 1251 190 1304 215
rect 1251 156 1259 190
rect 1293 156 1304 190
rect 785 53 797 67
rect 739 45 797 53
rect 1251 47 1304 156
rect 1334 100 1390 215
rect 1334 66 1345 100
rect 1379 66 1390 100
rect 1334 47 1390 66
rect 1420 190 1476 215
rect 1420 156 1431 190
rect 1465 156 1476 190
rect 1420 47 1476 156
rect 1506 112 1562 215
rect 1506 78 1517 112
rect 1551 78 1562 112
rect 1506 47 1562 78
rect 1592 190 1648 215
rect 1592 156 1603 190
rect 1637 156 1648 190
rect 1592 101 1648 156
rect 1592 67 1603 101
rect 1637 67 1648 101
rect 1592 47 1648 67
rect 1678 122 1734 215
rect 1678 88 1689 122
rect 1723 88 1734 122
rect 1678 47 1734 88
rect 1764 190 1820 215
rect 1764 156 1775 190
rect 1809 156 1820 190
rect 1764 101 1820 156
rect 1764 67 1775 101
rect 1809 67 1820 101
rect 1764 47 1820 67
rect 1850 122 1906 215
rect 1850 88 1861 122
rect 1895 88 1906 122
rect 1850 47 1906 88
rect 1936 190 1989 215
rect 1936 156 1947 190
rect 1981 156 1989 190
rect 1936 101 1989 156
rect 1936 67 1947 101
rect 1981 67 1989 101
rect 1936 47 1989 67
<< pdiff >>
rect 48 572 101 619
rect 48 538 56 572
rect 90 538 101 572
rect 48 504 101 538
rect 48 470 56 504
rect 90 470 101 504
rect 48 436 101 470
rect 48 402 56 436
rect 90 402 101 436
rect 48 367 101 402
rect 131 586 187 619
rect 131 552 142 586
rect 176 552 187 586
rect 131 367 187 552
rect 217 426 270 619
rect 217 392 228 426
rect 262 392 270 426
rect 217 367 270 392
rect 377 586 430 619
rect 377 552 385 586
rect 419 552 430 586
rect 377 367 430 552
rect 460 599 516 619
rect 460 565 471 599
rect 505 565 516 599
rect 460 506 516 565
rect 460 472 471 506
rect 505 472 516 506
rect 460 409 516 472
rect 460 375 471 409
rect 505 375 516 409
rect 460 367 516 375
rect 546 611 602 619
rect 546 577 557 611
rect 591 577 602 611
rect 546 536 602 577
rect 546 502 557 536
rect 591 502 602 536
rect 546 457 602 502
rect 546 423 557 457
rect 591 423 602 457
rect 546 367 602 423
rect 632 599 688 619
rect 632 565 643 599
rect 677 565 688 599
rect 632 506 688 565
rect 632 472 643 506
rect 677 472 688 506
rect 632 409 688 472
rect 632 375 643 409
rect 677 375 688 409
rect 632 367 688 375
rect 718 611 774 619
rect 718 577 729 611
rect 763 577 774 611
rect 718 543 774 577
rect 718 509 729 543
rect 763 509 774 543
rect 718 473 774 509
rect 718 439 729 473
rect 763 439 774 473
rect 718 367 774 439
rect 804 599 860 619
rect 804 565 815 599
rect 849 565 860 599
rect 804 506 860 565
rect 804 472 815 506
rect 849 472 860 506
rect 804 409 860 472
rect 804 375 815 409
rect 849 375 860 409
rect 804 367 860 375
rect 890 611 946 619
rect 890 577 901 611
rect 935 577 946 611
rect 890 492 946 577
rect 890 458 901 492
rect 935 458 946 492
rect 890 367 946 458
rect 976 599 1032 619
rect 976 565 987 599
rect 1021 565 1032 599
rect 976 506 1032 565
rect 976 472 987 506
rect 1021 472 1032 506
rect 976 409 1032 472
rect 976 375 987 409
rect 1021 375 1032 409
rect 976 367 1032 375
rect 1062 611 1298 619
rect 1062 577 1073 611
rect 1107 577 1160 611
rect 1194 577 1253 611
rect 1287 577 1298 611
rect 1062 543 1298 577
rect 1062 509 1253 543
rect 1287 509 1298 543
rect 1062 500 1298 509
rect 1062 466 1073 500
rect 1107 466 1160 500
rect 1194 475 1298 500
rect 1194 466 1253 475
rect 1062 441 1253 466
rect 1287 441 1298 475
rect 1062 367 1298 441
rect 1328 599 1384 619
rect 1328 565 1339 599
rect 1373 565 1384 599
rect 1328 506 1384 565
rect 1328 472 1339 506
rect 1373 472 1384 506
rect 1328 409 1384 472
rect 1328 375 1339 409
rect 1373 375 1384 409
rect 1328 367 1384 375
rect 1414 611 1470 619
rect 1414 577 1425 611
rect 1459 577 1470 611
rect 1414 533 1470 577
rect 1414 499 1425 533
rect 1459 499 1470 533
rect 1414 457 1470 499
rect 1414 423 1425 457
rect 1459 423 1470 457
rect 1414 367 1470 423
rect 1500 599 1556 619
rect 1500 565 1511 599
rect 1545 565 1556 599
rect 1500 506 1556 565
rect 1500 472 1511 506
rect 1545 472 1556 506
rect 1500 409 1556 472
rect 1500 375 1511 409
rect 1545 375 1556 409
rect 1500 367 1556 375
rect 1586 611 1642 619
rect 1586 577 1597 611
rect 1631 577 1642 611
rect 1586 533 1642 577
rect 1586 499 1597 533
rect 1631 499 1642 533
rect 1586 457 1642 499
rect 1586 423 1597 457
rect 1631 423 1642 457
rect 1586 367 1642 423
rect 1672 599 1728 619
rect 1672 565 1683 599
rect 1717 565 1728 599
rect 1672 506 1728 565
rect 1672 472 1683 506
rect 1717 472 1728 506
rect 1672 409 1728 472
rect 1672 375 1683 409
rect 1717 375 1728 409
rect 1672 367 1728 375
rect 1758 611 1814 619
rect 1758 577 1769 611
rect 1803 577 1814 611
rect 1758 533 1814 577
rect 1758 499 1769 533
rect 1803 499 1814 533
rect 1758 457 1814 499
rect 1758 423 1769 457
rect 1803 423 1814 457
rect 1758 367 1814 423
rect 1844 599 1900 619
rect 1844 565 1855 599
rect 1889 565 1900 599
rect 1844 506 1900 565
rect 1844 472 1855 506
rect 1889 472 1900 506
rect 1844 409 1900 472
rect 1844 375 1855 409
rect 1889 375 1900 409
rect 1844 367 1900 375
rect 1930 607 1983 619
rect 1930 573 1941 607
rect 1975 573 1983 607
rect 1930 506 1983 573
rect 1930 472 1941 506
rect 1975 472 1983 506
rect 1930 413 1983 472
rect 1930 379 1941 413
rect 1975 379 1983 413
rect 1930 367 1983 379
<< ndiffc >>
rect 52 158 86 192
rect 52 81 86 115
rect 142 174 176 208
rect 142 77 176 111
rect 228 158 262 192
rect 228 81 262 115
rect 336 53 370 87
rect 445 193 479 227
rect 547 53 581 87
rect 649 193 683 227
rect 751 53 785 87
rect 853 193 887 227
rect 939 143 973 177
rect 939 75 973 109
rect 1025 188 1059 222
rect 1111 108 1145 142
rect 1259 156 1293 190
rect 1345 66 1379 100
rect 1431 156 1465 190
rect 1517 78 1551 112
rect 1603 156 1637 190
rect 1603 67 1637 101
rect 1689 88 1723 122
rect 1775 156 1809 190
rect 1775 67 1809 101
rect 1861 88 1895 122
rect 1947 156 1981 190
rect 1947 67 1981 101
<< pdiffc >>
rect 56 538 90 572
rect 56 470 90 504
rect 56 402 90 436
rect 142 552 176 586
rect 228 392 262 426
rect 385 552 419 586
rect 471 565 505 599
rect 471 472 505 506
rect 471 375 505 409
rect 557 577 591 611
rect 557 502 591 536
rect 557 423 591 457
rect 643 565 677 599
rect 643 472 677 506
rect 643 375 677 409
rect 729 577 763 611
rect 729 509 763 543
rect 729 439 763 473
rect 815 565 849 599
rect 815 472 849 506
rect 815 375 849 409
rect 901 577 935 611
rect 901 458 935 492
rect 987 565 1021 599
rect 987 472 1021 506
rect 987 375 1021 409
rect 1073 577 1107 611
rect 1160 577 1194 611
rect 1253 577 1287 611
rect 1253 509 1287 543
rect 1073 466 1107 500
rect 1160 466 1194 500
rect 1253 441 1287 475
rect 1339 565 1373 599
rect 1339 472 1373 506
rect 1339 375 1373 409
rect 1425 577 1459 611
rect 1425 499 1459 533
rect 1425 423 1459 457
rect 1511 565 1545 599
rect 1511 472 1545 506
rect 1511 375 1545 409
rect 1597 577 1631 611
rect 1597 499 1631 533
rect 1597 423 1631 457
rect 1683 565 1717 599
rect 1683 472 1717 506
rect 1683 375 1717 409
rect 1769 577 1803 611
rect 1769 499 1803 533
rect 1769 423 1803 457
rect 1855 565 1889 599
rect 1855 472 1889 506
rect 1855 375 1889 409
rect 1941 573 1975 607
rect 1941 472 1975 506
rect 1941 379 1975 413
<< poly >>
rect 101 619 131 645
rect 187 619 217 645
rect 430 619 460 645
rect 516 619 546 645
rect 602 619 632 645
rect 688 619 718 645
rect 774 619 804 645
rect 860 619 890 645
rect 946 619 976 645
rect 1032 619 1062 645
rect 1298 619 1328 645
rect 1384 619 1414 645
rect 1470 619 1500 645
rect 1556 619 1586 645
rect 1642 619 1672 645
rect 1728 619 1758 645
rect 1814 619 1844 645
rect 1900 619 1930 645
rect 101 325 131 367
rect 187 325 217 367
rect 430 335 460 367
rect 516 335 546 367
rect 602 335 632 367
rect 688 335 718 367
rect 73 309 139 325
rect 73 275 89 309
rect 123 275 139 309
rect 73 259 139 275
rect 187 309 273 325
rect 187 275 223 309
rect 257 275 273 309
rect 187 259 273 275
rect 398 319 718 335
rect 398 285 414 319
rect 448 285 482 319
rect 516 285 550 319
rect 584 285 618 319
rect 652 299 718 319
rect 774 333 804 367
rect 860 333 890 367
rect 946 333 976 367
rect 1032 333 1062 367
rect 774 317 1180 333
rect 652 285 724 299
rect 398 269 724 285
rect 101 237 131 259
rect 187 237 217 259
rect 404 235 434 269
rect 490 235 520 269
rect 608 235 638 269
rect 694 235 724 269
rect 774 283 790 317
rect 824 283 858 317
rect 892 283 926 317
rect 960 283 994 317
rect 1028 283 1062 317
rect 1096 283 1130 317
rect 1164 283 1180 317
rect 1298 303 1328 367
rect 1384 303 1414 367
rect 1470 303 1500 367
rect 1556 303 1586 367
rect 1642 303 1672 367
rect 1728 303 1758 367
rect 1814 303 1844 367
rect 1900 303 1930 367
rect 774 267 1180 283
rect 1254 287 1592 303
rect 812 235 842 267
rect 898 235 928 267
rect 984 235 1014 267
rect 1070 235 1100 267
rect 1254 253 1270 287
rect 1304 253 1338 287
rect 1372 253 1406 287
rect 1440 253 1474 287
rect 1508 253 1542 287
rect 1576 253 1592 287
rect 1254 237 1592 253
rect 1642 287 1980 303
rect 1642 253 1658 287
rect 1692 253 1726 287
rect 1760 253 1794 287
rect 1828 253 1862 287
rect 1896 253 1930 287
rect 1964 253 1980 287
rect 1642 237 1980 253
rect 101 43 131 69
rect 187 43 217 69
rect 404 41 434 67
rect 490 41 520 67
rect 608 41 638 67
rect 694 41 724 67
rect 1304 215 1334 237
rect 1390 215 1420 237
rect 1476 215 1506 237
rect 1562 215 1592 237
rect 1648 215 1678 237
rect 1734 215 1764 237
rect 1820 215 1850 237
rect 1906 215 1936 237
rect 812 41 842 67
rect 898 41 928 67
rect 984 41 1014 67
rect 1070 41 1100 67
rect 1304 21 1334 47
rect 1390 21 1420 47
rect 1476 21 1506 47
rect 1562 21 1592 47
rect 1648 21 1678 47
rect 1734 21 1764 47
rect 1820 21 1850 47
rect 1906 21 1936 47
<< polycont >>
rect 89 275 123 309
rect 223 275 257 309
rect 414 285 448 319
rect 482 285 516 319
rect 550 285 584 319
rect 618 285 652 319
rect 790 283 824 317
rect 858 283 892 317
rect 926 283 960 317
rect 994 283 1028 317
rect 1062 283 1096 317
rect 1130 283 1164 317
rect 1270 253 1304 287
rect 1338 253 1372 287
rect 1406 253 1440 287
rect 1474 253 1508 287
rect 1542 253 1576 287
rect 1658 253 1692 287
rect 1726 253 1760 287
rect 1794 253 1828 287
rect 1862 253 1896 287
rect 1930 253 1964 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 17 572 90 588
rect 17 538 56 572
rect 17 504 90 538
rect 126 586 192 649
rect 126 552 142 586
rect 176 552 192 586
rect 126 536 192 552
rect 369 586 435 649
rect 369 552 385 586
rect 419 552 435 586
rect 369 536 435 552
rect 469 599 507 615
rect 469 565 471 599
rect 505 565 507 599
rect 17 470 56 504
rect 469 506 507 565
rect 90 470 404 502
rect 17 468 404 470
rect 17 436 90 468
rect 17 402 56 436
rect 17 386 90 402
rect 212 426 336 434
rect 212 392 228 426
rect 262 392 336 426
rect 17 208 55 386
rect 212 384 336 392
rect 89 309 173 350
rect 123 275 173 309
rect 89 242 173 275
rect 207 309 257 350
rect 207 275 223 309
rect 207 242 257 275
rect 17 192 92 208
rect 17 158 52 192
rect 86 158 92 192
rect 17 115 92 158
rect 17 81 52 115
rect 86 81 92 115
rect 17 65 92 81
rect 126 174 142 208
rect 176 174 192 208
rect 126 111 192 174
rect 126 77 142 111
rect 176 77 192 111
rect 126 17 192 77
rect 226 192 266 208
rect 226 158 228 192
rect 262 158 266 192
rect 226 157 266 158
rect 300 157 336 384
rect 370 321 404 468
rect 469 472 471 506
rect 505 472 507 506
rect 469 409 507 472
rect 541 611 607 649
rect 541 577 557 611
rect 591 577 607 611
rect 541 536 607 577
rect 541 502 557 536
rect 591 502 607 536
rect 541 457 607 502
rect 541 423 557 457
rect 591 423 607 457
rect 641 599 685 615
rect 641 565 643 599
rect 677 565 685 599
rect 641 506 685 565
rect 641 472 643 506
rect 677 472 685 506
rect 469 375 471 409
rect 505 389 507 409
rect 641 409 685 472
rect 719 611 765 649
rect 719 577 729 611
rect 763 577 765 611
rect 719 543 765 577
rect 719 509 729 543
rect 763 509 765 543
rect 719 473 765 509
rect 719 439 729 473
rect 763 439 765 473
rect 719 423 765 439
rect 799 599 851 615
rect 799 565 815 599
rect 849 565 851 599
rect 799 506 851 565
rect 799 472 815 506
rect 849 472 851 506
rect 799 424 851 472
rect 885 611 951 649
rect 885 577 901 611
rect 935 577 951 611
rect 885 492 951 577
rect 885 458 901 492
rect 935 458 951 492
rect 985 599 1023 615
rect 985 565 987 599
rect 1021 565 1023 599
rect 985 506 1023 565
rect 985 472 987 506
rect 1021 472 1023 506
rect 985 432 1023 472
rect 1057 611 1295 649
rect 1057 577 1073 611
rect 1107 577 1160 611
rect 1194 577 1253 611
rect 1287 577 1295 611
rect 1057 543 1295 577
rect 1057 509 1253 543
rect 1287 509 1295 543
rect 1057 500 1295 509
rect 1057 466 1073 500
rect 1107 466 1160 500
rect 1194 475 1295 500
rect 1194 466 1253 475
rect 1251 441 1253 466
rect 1287 441 1295 475
rect 985 424 1217 432
rect 1251 425 1295 441
rect 1329 599 1375 615
rect 1329 565 1339 599
rect 1373 565 1375 599
rect 1329 506 1375 565
rect 1329 472 1339 506
rect 1373 472 1375 506
rect 641 389 643 409
rect 505 375 643 389
rect 677 389 685 409
rect 799 409 1217 424
rect 799 389 815 409
rect 677 375 815 389
rect 849 375 987 409
rect 1021 389 1217 409
rect 1329 409 1375 472
rect 1409 611 1475 649
rect 1409 577 1425 611
rect 1459 577 1475 611
rect 1409 533 1475 577
rect 1409 499 1425 533
rect 1459 499 1475 533
rect 1409 457 1475 499
rect 1409 423 1425 457
rect 1459 423 1475 457
rect 1509 599 1547 615
rect 1509 565 1511 599
rect 1545 565 1547 599
rect 1509 506 1547 565
rect 1509 472 1511 506
rect 1545 472 1547 506
rect 1329 389 1339 409
rect 1021 375 1339 389
rect 1373 389 1375 409
rect 1509 409 1547 472
rect 1581 611 1647 649
rect 1581 577 1597 611
rect 1631 577 1647 611
rect 1581 533 1647 577
rect 1581 499 1597 533
rect 1631 499 1647 533
rect 1581 457 1647 499
rect 1581 423 1597 457
rect 1631 423 1647 457
rect 1681 599 1719 615
rect 1681 565 1683 599
rect 1717 565 1719 599
rect 1681 506 1719 565
rect 1681 472 1683 506
rect 1717 472 1719 506
rect 1509 389 1511 409
rect 1373 375 1511 389
rect 1545 389 1547 409
rect 1681 409 1719 472
rect 1753 611 1819 649
rect 1753 577 1769 611
rect 1803 577 1819 611
rect 1753 533 1819 577
rect 1753 499 1769 533
rect 1803 499 1819 533
rect 1753 457 1819 499
rect 1753 423 1769 457
rect 1803 423 1819 457
rect 1853 599 1897 615
rect 1853 565 1855 599
rect 1889 565 1897 599
rect 1853 506 1897 565
rect 1853 472 1855 506
rect 1889 472 1897 506
rect 1681 389 1683 409
rect 1545 375 1683 389
rect 1717 389 1719 409
rect 1853 409 1897 472
rect 1853 389 1855 409
rect 1717 375 1855 389
rect 1889 375 1897 409
rect 469 355 1897 375
rect 1931 607 1991 649
rect 1931 573 1941 607
rect 1975 573 1991 607
rect 1931 506 1991 573
rect 1931 472 1941 506
rect 1975 472 1991 506
rect 1931 413 1991 472
rect 1931 379 1941 413
rect 1975 379 1991 413
rect 1931 363 1991 379
rect 370 319 668 321
rect 370 285 414 319
rect 448 285 482 319
rect 516 285 550 319
rect 584 285 618 319
rect 652 285 668 319
rect 370 277 668 285
rect 704 243 738 355
rect 1251 337 1897 355
rect 429 227 738 243
rect 429 193 445 227
rect 479 193 649 227
rect 683 193 738 227
rect 429 191 738 193
rect 774 317 1180 321
rect 774 283 790 317
rect 824 283 858 317
rect 892 283 926 317
rect 960 283 994 317
rect 1028 283 1062 317
rect 1096 283 1130 317
rect 1164 283 1180 317
rect 1254 287 1601 303
rect 774 157 808 283
rect 1254 253 1270 287
rect 1304 253 1338 287
rect 1372 253 1406 287
rect 1440 253 1474 287
rect 1508 253 1542 287
rect 1576 253 1601 287
rect 849 227 1220 249
rect 1254 240 1601 253
rect 1642 287 1985 303
rect 1642 253 1658 287
rect 1692 253 1726 287
rect 1760 253 1794 287
rect 1828 253 1862 287
rect 1896 253 1930 287
rect 1964 253 1985 287
rect 1642 240 1985 253
rect 849 193 853 227
rect 887 222 1220 227
rect 887 211 1025 222
rect 887 193 889 211
rect 849 177 889 193
rect 1023 188 1025 211
rect 1059 192 1220 222
rect 1059 188 1061 192
rect 226 123 808 157
rect 923 143 939 177
rect 973 143 989 177
rect 1023 172 1061 188
rect 226 115 266 123
rect 226 81 228 115
rect 262 81 266 115
rect 923 109 989 143
rect 923 89 939 109
rect 226 65 266 81
rect 320 87 939 89
rect 320 53 336 87
rect 370 53 547 87
rect 581 53 751 87
rect 785 75 939 87
rect 973 85 989 109
rect 1095 142 1152 158
rect 1095 108 1111 142
rect 1145 108 1152 142
rect 1095 85 1152 108
rect 973 75 1152 85
rect 785 53 1152 75
rect 1186 104 1220 192
rect 1256 190 1985 206
rect 1256 156 1259 190
rect 1293 156 1431 190
rect 1465 172 1603 190
rect 1465 156 1469 172
rect 1256 140 1469 156
rect 1599 156 1603 172
rect 1637 172 1775 190
rect 1637 156 1639 172
rect 1503 112 1555 138
rect 1503 104 1517 112
rect 1186 100 1517 104
rect 1186 66 1345 100
rect 1379 78 1517 100
rect 1551 78 1555 112
rect 1379 66 1555 78
rect 1186 62 1555 66
rect 1599 101 1639 156
rect 1773 156 1775 172
rect 1809 172 1947 190
rect 1599 67 1603 101
rect 1637 67 1639 101
rect 320 51 1152 53
rect 1599 51 1639 67
rect 1673 122 1739 138
rect 1673 88 1689 122
rect 1723 88 1739 122
rect 1673 17 1739 88
rect 1773 101 1809 156
rect 1945 156 1947 172
rect 1981 156 1985 190
rect 1773 67 1775 101
rect 1773 51 1809 67
rect 1845 122 1911 138
rect 1845 88 1861 122
rect 1895 88 1911 122
rect 1845 17 1911 88
rect 1945 101 1985 156
rect 1945 67 1947 101
rect 1981 67 1985 101
rect 1945 51 1985 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nand4bb_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1567 242 1601 276 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1663 242 1697 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 1759 242 1793 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 1855 242 1889 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 D
port 4 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A_N
port 1 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B_N
port 2 nsew signal input
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1087 390 1121 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 1183 390 1217 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 5667884
string GDS_START 5651126
<< end >>
