magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2258 1975
<< nwell >>
rect -38 332 998 704
<< pwell >>
rect 770 228 959 248
rect 6 49 959 228
rect 0 0 960 49
<< scnmos >>
rect 89 74 119 202
rect 167 74 197 202
rect 356 74 386 202
rect 434 74 464 202
rect 621 74 651 202
rect 699 74 729 202
rect 846 74 876 222
<< scpmoshvt >>
rect 86 390 116 590
rect 207 390 237 590
rect 307 390 337 590
rect 425 390 455 590
rect 637 383 667 583
rect 727 383 757 583
rect 844 368 874 592
<< ndiff >>
rect 796 202 846 222
rect 32 188 89 202
rect 32 154 44 188
rect 78 154 89 188
rect 32 120 89 154
rect 32 86 44 120
rect 78 86 89 120
rect 32 74 89 86
rect 119 74 167 202
rect 197 120 356 202
rect 197 86 208 120
rect 242 86 311 120
rect 345 86 356 120
rect 197 74 356 86
rect 386 74 434 202
rect 464 184 621 202
rect 464 150 475 184
rect 509 150 576 184
rect 610 150 621 184
rect 464 116 621 150
rect 464 82 475 116
rect 509 82 576 116
rect 610 82 621 116
rect 464 74 621 82
rect 651 74 699 202
rect 729 120 846 202
rect 729 86 763 120
rect 797 86 846 120
rect 729 74 846 86
rect 876 210 933 222
rect 876 176 887 210
rect 921 176 933 210
rect 876 120 933 176
rect 876 86 887 120
rect 921 86 933 120
rect 876 74 933 86
<< pdiff >>
rect 27 578 86 590
rect 27 544 39 578
rect 73 544 86 578
rect 27 510 86 544
rect 27 476 39 510
rect 73 476 86 510
rect 27 442 86 476
rect 27 408 39 442
rect 73 408 86 442
rect 27 390 86 408
rect 116 531 207 590
rect 116 497 160 531
rect 194 497 207 531
rect 116 436 207 497
rect 116 402 160 436
rect 194 402 207 436
rect 116 390 207 402
rect 237 578 307 590
rect 237 544 260 578
rect 294 544 307 578
rect 237 507 307 544
rect 237 473 260 507
rect 294 473 307 507
rect 237 436 307 473
rect 237 402 260 436
rect 294 402 307 436
rect 237 390 307 402
rect 337 531 425 590
rect 337 497 360 531
rect 394 497 425 531
rect 337 436 425 497
rect 337 402 360 436
rect 394 402 425 436
rect 337 390 425 402
rect 455 578 514 590
rect 775 583 844 592
rect 455 544 468 578
rect 502 544 514 578
rect 455 510 514 544
rect 455 476 468 510
rect 502 476 514 510
rect 455 390 514 476
rect 568 570 637 583
rect 568 536 580 570
rect 614 536 637 570
rect 568 494 637 536
rect 568 460 580 494
rect 614 460 637 494
rect 568 383 637 460
rect 667 571 727 583
rect 667 537 680 571
rect 714 537 727 571
rect 667 500 727 537
rect 667 466 680 500
rect 714 466 727 500
rect 667 429 727 466
rect 667 395 680 429
rect 714 395 727 429
rect 667 383 727 395
rect 757 580 844 583
rect 757 546 787 580
rect 821 546 844 580
rect 757 504 844 546
rect 757 470 787 504
rect 821 470 844 504
rect 757 429 844 470
rect 757 395 787 429
rect 821 395 844 429
rect 757 383 844 395
rect 791 368 844 383
rect 874 580 933 592
rect 874 546 887 580
rect 921 546 933 580
rect 874 497 933 546
rect 874 463 887 497
rect 921 463 933 497
rect 874 414 933 463
rect 874 380 887 414
rect 921 380 933 414
rect 874 368 933 380
<< ndiffc >>
rect 44 154 78 188
rect 44 86 78 120
rect 208 86 242 120
rect 311 86 345 120
rect 475 150 509 184
rect 576 150 610 184
rect 475 82 509 116
rect 576 82 610 116
rect 763 86 797 120
rect 887 176 921 210
rect 887 86 921 120
<< pdiffc >>
rect 39 544 73 578
rect 39 476 73 510
rect 39 408 73 442
rect 160 497 194 531
rect 160 402 194 436
rect 260 544 294 578
rect 260 473 294 507
rect 260 402 294 436
rect 360 497 394 531
rect 360 402 394 436
rect 468 544 502 578
rect 468 476 502 510
rect 580 536 614 570
rect 580 460 614 494
rect 680 537 714 571
rect 680 466 714 500
rect 680 395 714 429
rect 787 546 821 580
rect 787 470 821 504
rect 787 395 821 429
rect 887 546 921 580
rect 887 463 921 497
rect 887 380 921 414
<< poly >>
rect 86 590 116 616
rect 207 590 237 616
rect 307 590 337 616
rect 425 590 455 616
rect 637 583 667 609
rect 727 583 757 609
rect 844 592 874 618
rect 86 375 116 390
rect 207 375 237 390
rect 307 375 337 390
rect 425 375 455 390
rect 83 290 119 375
rect 44 274 119 290
rect 44 240 60 274
rect 94 240 119 274
rect 204 290 240 375
rect 304 368 340 375
rect 304 338 350 368
rect 425 358 458 375
rect 637 368 667 383
rect 727 368 757 383
rect 320 302 350 338
rect 204 274 278 290
rect 204 254 228 274
rect 44 224 119 240
rect 89 202 119 224
rect 167 240 228 254
rect 262 240 278 274
rect 167 224 278 240
rect 320 286 386 302
rect 320 252 336 286
rect 370 252 386 286
rect 320 236 386 252
rect 167 202 197 224
rect 356 202 386 236
rect 428 290 458 358
rect 621 338 670 368
rect 621 290 651 338
rect 724 290 760 368
rect 844 353 874 368
rect 841 326 877 353
rect 808 310 877 326
rect 428 274 510 290
rect 428 240 460 274
rect 494 240 510 274
rect 428 224 510 240
rect 585 274 651 290
rect 585 240 601 274
rect 635 240 651 274
rect 585 224 651 240
rect 434 202 464 224
rect 621 202 651 224
rect 699 274 765 290
rect 699 240 715 274
rect 749 240 765 274
rect 808 276 824 310
rect 858 276 877 310
rect 808 260 877 276
rect 699 224 765 240
rect 699 202 729 224
rect 846 222 876 260
rect 89 48 119 74
rect 167 48 197 74
rect 356 48 386 74
rect 434 48 464 74
rect 621 48 651 74
rect 699 48 729 74
rect 846 48 876 74
<< polycont >>
rect 60 240 94 274
rect 228 240 262 274
rect 336 252 370 286
rect 460 240 494 274
rect 601 240 635 274
rect 715 240 749 274
rect 824 276 858 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 23 581 518 615
rect 23 578 89 581
rect 23 544 39 578
rect 73 544 89 578
rect 244 578 310 581
rect 23 510 89 544
rect 23 476 39 510
rect 73 476 89 510
rect 23 442 89 476
rect 23 408 39 442
rect 73 408 89 442
rect 23 392 89 408
rect 144 531 210 547
rect 144 497 160 531
rect 194 497 210 531
rect 144 436 210 497
rect 144 402 160 436
rect 194 402 210 436
rect 144 386 210 402
rect 244 544 260 578
rect 294 544 310 578
rect 452 578 518 581
rect 244 507 310 544
rect 244 473 260 507
rect 294 473 310 507
rect 244 436 310 473
rect 244 402 260 436
rect 294 402 310 436
rect 244 386 310 402
rect 344 531 410 547
rect 344 497 360 531
rect 394 497 410 531
rect 344 436 410 497
rect 452 544 468 578
rect 502 544 518 578
rect 452 510 518 544
rect 452 476 468 510
rect 502 476 518 510
rect 452 460 518 476
rect 564 570 630 649
rect 564 536 580 570
rect 614 536 630 570
rect 564 494 630 536
rect 564 460 580 494
rect 614 460 630 494
rect 664 571 730 587
rect 664 537 680 571
rect 714 537 730 571
rect 664 500 730 537
rect 664 466 680 500
rect 714 466 730 500
rect 344 402 360 436
rect 394 426 410 436
rect 664 429 730 466
rect 664 426 680 429
rect 394 402 680 426
rect 344 395 680 402
rect 714 395 730 429
rect 344 392 730 395
rect 344 386 410 392
rect 25 274 110 358
rect 25 240 60 274
rect 94 240 110 274
rect 25 224 110 240
rect 144 190 178 386
rect 664 379 730 392
rect 771 580 837 649
rect 771 546 787 580
rect 821 546 837 580
rect 771 504 837 546
rect 771 470 787 504
rect 821 470 837 504
rect 771 429 837 470
rect 771 395 787 429
rect 821 395 837 429
rect 771 379 837 395
rect 871 580 942 596
rect 871 546 887 580
rect 921 546 942 580
rect 871 497 942 546
rect 871 463 887 497
rect 921 463 942 497
rect 871 414 942 463
rect 871 380 887 414
rect 921 380 942 414
rect 871 364 942 380
rect 212 274 278 352
rect 212 240 228 274
rect 262 240 278 274
rect 212 224 278 240
rect 313 286 386 352
rect 313 252 336 286
rect 370 252 386 286
rect 313 236 386 252
rect 444 274 551 358
rect 803 310 874 326
rect 444 240 460 274
rect 494 240 551 274
rect 444 224 551 240
rect 585 274 651 304
rect 585 240 601 274
rect 635 240 651 274
rect 585 224 651 240
rect 697 274 765 309
rect 697 240 715 274
rect 749 240 765 274
rect 697 224 765 240
rect 803 276 824 310
rect 858 276 874 310
rect 803 260 874 276
rect 803 190 837 260
rect 908 226 942 364
rect 28 188 837 190
rect 28 154 44 188
rect 78 184 837 188
rect 78 156 475 184
rect 78 154 94 156
rect 28 120 94 154
rect 459 150 475 156
rect 509 150 576 184
rect 610 156 837 184
rect 871 210 942 226
rect 871 176 887 210
rect 921 176 942 210
rect 610 150 626 156
rect 28 86 44 120
rect 78 86 94 120
rect 28 70 94 86
rect 192 86 208 120
rect 242 86 311 120
rect 345 86 361 120
rect 192 17 361 86
rect 459 116 626 150
rect 459 82 475 116
rect 509 82 576 116
rect 610 82 626 116
rect 459 66 626 82
rect 724 120 837 122
rect 724 86 763 120
rect 797 86 837 120
rect 724 17 837 86
rect 871 120 942 176
rect 871 86 887 120
rect 921 86 942 120
rect 871 70 942 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
<< metal1 >>
rect 0 683 960 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 960 683
rect 0 617 960 649
rect 0 17 960 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 960 17
rect 0 -49 960 -17
<< labels >>
rlabel comment s 0 0 0 0 4 a222o_1
flabel pwell s 0 0 960 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 960 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
flabel metal1 s 0 617 960 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional abutment
flabel metal1 s 0 0 960 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional abutment
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 C2
port 6 nsew signal input
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 895 464 929 498 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 895 538 929 572 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 B2
port 4 nsew signal input
flabel locali s 703 242 737 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 960 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 127338
string GDS_START 118370
<< end >>
