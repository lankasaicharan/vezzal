magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 9 49 667 241
rect 0 0 672 49
<< scnmos >>
rect 88 47 118 215
rect 264 47 294 215
rect 342 47 372 215
rect 456 47 486 215
rect 558 47 588 215
<< scpmoshvt >>
rect 80 367 110 619
rect 270 367 300 619
rect 372 367 402 619
rect 474 367 504 619
rect 558 367 588 619
<< ndiff >>
rect 35 203 88 215
rect 35 169 43 203
rect 77 169 88 203
rect 35 101 88 169
rect 35 67 43 101
rect 77 67 88 101
rect 35 47 88 67
rect 118 129 264 215
rect 118 95 133 129
rect 167 95 219 129
rect 253 95 264 129
rect 118 47 264 95
rect 294 47 342 215
rect 372 205 456 215
rect 372 171 397 205
rect 431 171 456 205
rect 372 92 456 171
rect 372 58 397 92
rect 431 58 456 92
rect 372 47 456 58
rect 486 129 558 215
rect 486 95 505 129
rect 539 95 558 129
rect 486 47 558 95
rect 588 187 641 215
rect 588 153 599 187
rect 633 153 641 187
rect 588 101 641 153
rect 588 67 599 101
rect 633 67 641 101
rect 588 47 641 67
<< pdiff >>
rect 27 599 80 619
rect 27 565 35 599
rect 69 565 80 599
rect 27 504 80 565
rect 27 470 35 504
rect 69 470 80 504
rect 27 420 80 470
rect 27 386 35 420
rect 69 386 80 420
rect 27 367 80 386
rect 110 607 163 619
rect 110 573 121 607
rect 155 573 163 607
rect 110 534 163 573
rect 110 500 121 534
rect 155 500 163 534
rect 110 459 163 500
rect 110 425 121 459
rect 155 425 163 459
rect 110 367 163 425
rect 217 599 270 619
rect 217 565 225 599
rect 259 565 270 599
rect 217 529 270 565
rect 217 495 225 529
rect 259 495 270 529
rect 217 441 270 495
rect 217 407 225 441
rect 259 407 270 441
rect 217 367 270 407
rect 300 607 372 619
rect 300 573 319 607
rect 353 573 372 607
rect 300 517 372 573
rect 300 483 319 517
rect 353 483 372 517
rect 300 367 372 483
rect 402 605 474 619
rect 402 571 422 605
rect 456 571 474 605
rect 402 529 474 571
rect 402 495 422 529
rect 456 495 474 529
rect 402 441 474 495
rect 402 407 422 441
rect 456 407 474 441
rect 402 367 474 407
rect 504 367 558 619
rect 588 599 641 619
rect 588 565 599 599
rect 633 565 641 599
rect 588 509 641 565
rect 588 475 599 509
rect 633 475 641 509
rect 588 413 641 475
rect 588 379 599 413
rect 633 379 641 413
rect 588 367 641 379
<< ndiffc >>
rect 43 169 77 203
rect 43 67 77 101
rect 133 95 167 129
rect 219 95 253 129
rect 397 171 431 205
rect 397 58 431 92
rect 505 95 539 129
rect 599 153 633 187
rect 599 67 633 101
<< pdiffc >>
rect 35 565 69 599
rect 35 470 69 504
rect 35 386 69 420
rect 121 573 155 607
rect 121 500 155 534
rect 121 425 155 459
rect 225 565 259 599
rect 225 495 259 529
rect 225 407 259 441
rect 319 573 353 607
rect 319 483 353 517
rect 422 571 456 605
rect 422 495 456 529
rect 422 407 456 441
rect 599 565 633 599
rect 599 475 633 509
rect 599 379 633 413
<< poly >>
rect 80 619 110 645
rect 270 619 300 645
rect 372 619 402 645
rect 474 619 504 645
rect 558 619 588 645
rect 80 303 110 367
rect 270 305 300 367
rect 80 287 183 303
rect 80 253 133 287
rect 167 253 183 287
rect 80 237 183 253
rect 228 289 300 305
rect 372 303 402 367
rect 474 303 504 367
rect 558 303 588 367
rect 228 255 244 289
rect 278 275 300 289
rect 342 287 408 303
rect 278 255 294 275
rect 228 239 294 255
rect 88 215 118 237
rect 264 215 294 239
rect 342 253 358 287
rect 392 253 408 287
rect 342 237 408 253
rect 450 287 516 303
rect 450 253 466 287
rect 500 253 516 287
rect 450 237 516 253
rect 558 287 647 303
rect 558 253 597 287
rect 631 253 647 287
rect 558 237 647 253
rect 342 215 372 237
rect 456 215 486 237
rect 558 215 588 237
rect 88 21 118 47
rect 264 21 294 47
rect 342 21 372 47
rect 456 21 486 47
rect 558 21 588 47
<< polycont >>
rect 133 253 167 287
rect 244 255 278 289
rect 358 253 392 287
rect 466 253 500 287
rect 597 253 631 287
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 19 599 81 615
rect 19 565 35 599
rect 69 565 81 599
rect 19 504 81 565
rect 19 470 35 504
rect 69 470 81 504
rect 19 420 81 470
rect 19 386 35 420
rect 69 386 81 420
rect 115 607 171 649
rect 115 573 121 607
rect 155 573 171 607
rect 115 534 171 573
rect 115 500 121 534
rect 155 500 171 534
rect 115 459 171 500
rect 115 425 121 459
rect 155 425 171 459
rect 115 409 171 425
rect 209 599 269 615
rect 209 565 225 599
rect 259 565 269 599
rect 209 529 269 565
rect 209 495 225 529
rect 259 495 269 529
rect 209 441 269 495
rect 303 607 369 649
rect 303 573 319 607
rect 353 573 369 607
rect 303 517 369 573
rect 303 483 319 517
rect 353 483 369 517
rect 303 475 369 483
rect 406 605 472 615
rect 406 571 422 605
rect 456 571 472 605
rect 406 529 472 571
rect 406 495 422 529
rect 456 495 472 529
rect 406 441 472 495
rect 209 407 225 441
rect 259 407 422 441
rect 456 407 472 441
rect 583 599 649 615
rect 583 565 599 599
rect 633 565 649 599
rect 583 509 649 565
rect 583 475 599 509
rect 633 475 649 509
rect 583 413 649 475
rect 19 203 81 386
rect 583 379 599 413
rect 633 379 649 413
rect 583 373 649 379
rect 19 169 43 203
rect 77 169 81 203
rect 117 339 649 373
rect 117 287 183 339
rect 117 253 133 287
rect 167 253 183 287
rect 117 205 183 253
rect 217 289 278 305
rect 217 255 244 289
rect 217 239 278 255
rect 312 287 408 305
rect 312 253 358 287
rect 392 253 408 287
rect 312 242 408 253
rect 450 287 547 305
rect 450 253 466 287
rect 500 253 547 287
rect 450 242 547 253
rect 581 287 647 305
rect 581 253 597 287
rect 631 253 647 287
rect 581 242 647 253
rect 117 171 397 205
rect 431 187 649 205
rect 431 171 599 187
rect 19 101 81 169
rect 19 67 43 101
rect 77 67 81 101
rect 19 51 81 67
rect 115 129 269 137
rect 115 95 133 129
rect 167 95 219 129
rect 253 95 269 129
rect 115 17 269 95
rect 381 92 447 171
rect 589 153 599 171
rect 633 153 649 187
rect 381 58 397 92
rect 431 58 447 92
rect 381 51 447 58
rect 489 129 555 137
rect 489 95 505 129
rect 539 95 555 129
rect 489 17 555 95
rect 589 101 649 153
rect 589 67 599 101
rect 633 67 649 101
rect 589 51 649 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a211o_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1954138
string GDS_START 1947106
<< end >>
