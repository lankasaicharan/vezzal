magic
tech sky130A
magscale 1 2
timestamp 1627202626
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 332 902 704
<< pwell >>
rect 6 49 863 248
rect 0 0 864 49
<< scpmos >>
rect 108 368 138 568
rect 222 368 252 568
rect 330 368 360 592
rect 414 368 444 592
rect 522 368 552 592
rect 639 368 669 592
rect 729 368 759 592
<< nmoslvt >>
rect 105 74 135 222
rect 189 74 219 222
rect 297 74 327 222
rect 441 74 471 222
rect 527 74 557 222
rect 646 74 676 222
rect 732 74 762 222
<< ndiff >>
rect 32 196 105 222
rect 32 162 60 196
rect 94 162 105 196
rect 32 120 105 162
rect 32 86 60 120
rect 94 86 105 120
rect 32 74 105 86
rect 135 74 189 222
rect 219 136 297 222
rect 219 102 252 136
rect 286 102 297 136
rect 219 74 297 102
rect 327 84 441 222
rect 327 74 367 84
rect 342 50 367 74
rect 401 74 441 84
rect 471 136 527 222
rect 471 102 482 136
rect 516 102 527 136
rect 471 74 527 102
rect 557 136 646 222
rect 557 102 582 136
rect 616 102 646 136
rect 557 74 646 102
rect 676 194 732 222
rect 676 160 687 194
rect 721 160 732 194
rect 676 120 732 160
rect 676 86 687 120
rect 721 86 732 120
rect 676 74 732 86
rect 762 120 837 222
rect 762 86 789 120
rect 823 86 837 120
rect 762 74 837 86
rect 401 50 426 74
rect 342 38 426 50
<< pdiff >>
rect 271 580 330 592
rect 271 568 283 580
rect 49 556 108 568
rect 49 522 61 556
rect 95 522 108 556
rect 49 485 108 522
rect 49 451 61 485
rect 95 451 108 485
rect 49 414 108 451
rect 49 380 61 414
rect 95 380 108 414
rect 49 368 108 380
rect 138 560 222 568
rect 138 526 171 560
rect 205 526 222 560
rect 138 492 222 526
rect 138 458 171 492
rect 205 458 222 492
rect 138 368 222 458
rect 252 546 283 568
rect 317 546 330 580
rect 252 510 330 546
rect 252 476 283 510
rect 317 476 330 510
rect 252 440 330 476
rect 252 406 283 440
rect 317 406 330 440
rect 252 368 330 406
rect 360 368 414 592
rect 444 368 522 592
rect 552 580 639 592
rect 552 546 565 580
rect 599 546 639 580
rect 552 510 639 546
rect 552 476 565 510
rect 599 476 639 510
rect 552 440 639 476
rect 552 406 565 440
rect 599 406 639 440
rect 552 368 639 406
rect 669 580 729 592
rect 669 546 682 580
rect 716 546 729 580
rect 669 497 729 546
rect 669 463 682 497
rect 716 463 729 497
rect 669 414 729 463
rect 669 380 682 414
rect 716 380 729 414
rect 669 368 729 380
rect 759 582 828 592
rect 759 548 782 582
rect 816 548 828 582
rect 759 514 828 548
rect 759 480 782 514
rect 816 480 828 514
rect 759 446 828 480
rect 759 412 782 446
rect 816 412 828 446
rect 759 368 828 412
<< ndiffc >>
rect 60 162 94 196
rect 60 86 94 120
rect 252 102 286 136
rect 367 50 401 84
rect 482 102 516 136
rect 582 102 616 136
rect 687 160 721 194
rect 687 86 721 120
rect 789 86 823 120
<< pdiffc >>
rect 61 522 95 556
rect 61 451 95 485
rect 61 380 95 414
rect 171 526 205 560
rect 171 458 205 492
rect 283 546 317 580
rect 283 476 317 510
rect 283 406 317 440
rect 565 546 599 580
rect 565 476 599 510
rect 565 406 599 440
rect 682 546 716 580
rect 682 463 716 497
rect 682 380 716 414
rect 782 548 816 582
rect 782 480 816 514
rect 782 412 816 446
<< poly >>
rect 108 568 138 594
rect 222 568 252 594
rect 330 592 360 618
rect 414 592 444 618
rect 522 592 552 618
rect 639 592 669 618
rect 729 592 759 618
rect 108 353 138 368
rect 222 353 252 368
rect 330 353 360 368
rect 414 353 444 368
rect 522 353 552 368
rect 639 353 669 368
rect 729 353 759 368
rect 105 310 141 353
rect 219 336 255 353
rect 327 336 363 353
rect 411 336 447 353
rect 519 336 555 353
rect 21 294 141 310
rect 21 260 37 294
rect 71 260 141 294
rect 21 244 141 260
rect 189 320 255 336
rect 189 286 205 320
rect 239 286 255 320
rect 189 270 255 286
rect 297 320 363 336
rect 297 286 313 320
rect 347 286 363 320
rect 297 270 363 286
rect 405 320 471 336
rect 405 286 421 320
rect 455 286 471 320
rect 405 270 471 286
rect 519 320 585 336
rect 519 286 535 320
rect 569 286 585 320
rect 519 270 585 286
rect 636 310 672 353
rect 726 310 762 353
rect 636 294 762 310
rect 105 222 135 244
rect 189 222 219 270
rect 297 222 327 270
rect 441 222 471 270
rect 527 222 557 270
rect 636 260 652 294
rect 686 260 762 294
rect 636 244 762 260
rect 646 222 676 244
rect 732 222 762 244
rect 105 48 135 74
rect 189 48 219 74
rect 297 48 327 74
rect 441 48 471 74
rect 527 48 557 74
rect 646 48 676 74
rect 732 48 762 74
<< polycont >>
rect 37 260 71 294
rect 205 286 239 320
rect 313 286 347 320
rect 421 286 455 320
rect 535 286 569 320
rect 652 260 686 294
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 45 556 121 572
rect 45 522 61 556
rect 95 522 121 556
rect 45 485 121 522
rect 45 451 61 485
rect 95 451 121 485
rect 155 560 221 649
rect 155 526 171 560
rect 205 526 221 560
rect 155 492 221 526
rect 155 458 171 492
rect 205 458 221 492
rect 267 580 333 596
rect 267 546 283 580
rect 317 546 333 580
rect 549 580 615 649
rect 267 510 333 546
rect 267 476 283 510
rect 317 476 333 510
rect 45 424 121 451
rect 267 440 333 476
rect 267 424 283 440
rect 45 414 283 424
rect 45 380 61 414
rect 95 406 283 414
rect 317 406 333 440
rect 95 390 333 406
rect 95 380 155 390
rect 45 364 155 380
rect 21 294 87 310
rect 21 260 37 294
rect 71 260 87 294
rect 21 236 87 260
rect 121 236 155 364
rect 189 320 263 356
rect 189 286 205 320
rect 239 286 263 320
rect 189 270 263 286
rect 297 320 363 356
rect 297 286 313 320
rect 347 286 363 320
rect 297 270 363 286
rect 405 320 471 578
rect 549 546 565 580
rect 599 546 615 580
rect 549 510 615 546
rect 549 476 565 510
rect 599 476 615 510
rect 549 440 615 476
rect 549 406 565 440
rect 599 406 615 440
rect 549 390 615 406
rect 666 580 732 596
rect 666 546 682 580
rect 716 546 732 580
rect 666 497 732 546
rect 666 463 682 497
rect 716 463 732 497
rect 666 414 732 463
rect 666 380 682 414
rect 716 380 732 414
rect 766 582 832 649
rect 766 548 782 582
rect 816 548 832 582
rect 766 514 832 548
rect 766 480 782 514
rect 816 480 832 514
rect 766 446 832 480
rect 766 412 782 446
rect 816 412 832 446
rect 666 378 732 380
rect 405 286 421 320
rect 455 286 471 320
rect 405 270 471 286
rect 505 320 585 356
rect 666 344 839 378
rect 505 286 535 320
rect 569 286 585 320
rect 505 270 585 286
rect 619 294 702 310
rect 619 260 652 294
rect 686 260 702 294
rect 619 244 702 260
rect 619 236 653 244
rect 121 202 653 236
rect 793 210 839 344
rect 41 196 155 202
rect 41 162 60 196
rect 94 162 155 196
rect 687 194 839 210
rect 41 120 155 162
rect 41 86 60 120
rect 94 86 155 120
rect 41 70 155 86
rect 236 136 532 168
rect 236 102 252 136
rect 286 134 482 136
rect 286 102 302 134
rect 236 70 302 102
rect 466 102 482 134
rect 516 102 532 136
rect 338 84 430 100
rect 338 50 367 84
rect 401 50 430 84
rect 466 70 532 102
rect 566 136 632 168
rect 566 102 582 136
rect 616 102 632 136
rect 338 17 430 50
rect 566 17 632 102
rect 721 162 839 194
rect 721 160 737 162
rect 687 120 737 160
rect 721 86 737 120
rect 687 70 737 86
rect 771 86 789 120
rect 823 86 841 120
rect 771 17 841 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o311a_2
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 C1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hs/gds/sky130_fd_sc_hs.gds
string LEFsymmetry X Y
string GDS_END 2445826
string GDS_START 2437850
<< end >>
