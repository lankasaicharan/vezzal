magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 331 1382 704
<< pwell >>
rect 48 49 1326 241
rect 0 0 1344 49
<< scnmos >>
rect 127 47 157 215
rect 229 47 259 215
rect 315 47 345 215
rect 417 47 447 215
rect 503 47 533 215
rect 589 47 619 215
rect 675 47 705 215
rect 761 47 791 215
rect 847 47 877 215
rect 959 47 989 215
rect 1045 47 1075 215
rect 1131 47 1161 215
rect 1217 47 1247 215
<< scpmoshvt >>
rect 95 367 125 619
rect 181 367 211 619
rect 267 367 297 619
rect 353 367 383 619
rect 439 367 469 619
rect 629 367 659 619
rect 715 367 745 619
rect 801 367 831 619
rect 887 367 917 619
rect 973 367 1003 619
rect 1059 367 1089 619
rect 1145 367 1175 619
rect 1231 367 1261 619
<< ndiff >>
rect 74 187 127 215
rect 74 153 82 187
rect 116 153 127 187
rect 74 101 127 153
rect 74 67 82 101
rect 116 67 127 101
rect 74 47 127 67
rect 157 198 229 215
rect 157 164 177 198
rect 211 164 229 198
rect 157 93 229 164
rect 157 59 177 93
rect 211 59 229 93
rect 157 47 229 59
rect 259 187 315 215
rect 259 153 270 187
rect 304 153 315 187
rect 259 101 315 153
rect 259 67 270 101
rect 304 67 315 101
rect 259 47 315 67
rect 345 126 417 215
rect 345 92 364 126
rect 398 92 417 126
rect 345 47 417 92
rect 447 203 503 215
rect 447 169 458 203
rect 492 169 503 203
rect 447 101 503 169
rect 447 67 458 101
rect 492 67 503 101
rect 447 47 503 67
rect 533 163 589 215
rect 533 129 544 163
rect 578 129 589 163
rect 533 89 589 129
rect 533 55 544 89
rect 578 55 589 89
rect 533 47 589 55
rect 619 203 675 215
rect 619 169 630 203
rect 664 169 675 203
rect 619 101 675 169
rect 619 67 630 101
rect 664 67 675 101
rect 619 47 675 67
rect 705 163 761 215
rect 705 129 716 163
rect 750 129 761 163
rect 705 89 761 129
rect 705 55 716 89
rect 750 55 761 89
rect 705 47 761 55
rect 791 203 847 215
rect 791 169 802 203
rect 836 169 847 203
rect 791 101 847 169
rect 791 67 802 101
rect 836 67 847 101
rect 791 47 847 67
rect 877 129 959 215
rect 877 95 901 129
rect 935 95 959 129
rect 877 47 959 95
rect 989 192 1045 215
rect 989 158 1000 192
rect 1034 158 1045 192
rect 989 101 1045 158
rect 989 67 1000 101
rect 1034 67 1045 101
rect 989 47 1045 67
rect 1075 129 1131 215
rect 1075 95 1086 129
rect 1120 95 1131 129
rect 1075 47 1131 95
rect 1161 203 1217 215
rect 1161 169 1172 203
rect 1206 169 1217 203
rect 1161 101 1217 169
rect 1161 67 1172 101
rect 1206 67 1217 101
rect 1161 47 1217 67
rect 1247 163 1300 215
rect 1247 129 1258 163
rect 1292 129 1300 163
rect 1247 93 1300 129
rect 1247 59 1258 93
rect 1292 59 1300 93
rect 1247 47 1300 59
<< pdiff >>
rect 38 599 95 619
rect 38 565 46 599
rect 80 565 95 599
rect 38 507 95 565
rect 38 473 46 507
rect 80 473 95 507
rect 38 413 95 473
rect 38 379 46 413
rect 80 379 95 413
rect 38 367 95 379
rect 125 607 181 619
rect 125 573 136 607
rect 170 573 181 607
rect 125 529 181 573
rect 125 495 136 529
rect 170 495 181 529
rect 125 455 181 495
rect 125 421 136 455
rect 170 421 181 455
rect 125 367 181 421
rect 211 597 267 619
rect 211 563 222 597
rect 256 563 267 597
rect 211 529 267 563
rect 211 495 222 529
rect 256 495 267 529
rect 211 459 267 495
rect 211 425 222 459
rect 256 425 267 459
rect 211 367 267 425
rect 297 607 353 619
rect 297 573 308 607
rect 342 573 353 607
rect 297 521 353 573
rect 297 487 308 521
rect 342 487 353 521
rect 297 367 353 487
rect 383 597 439 619
rect 383 563 394 597
rect 428 563 439 597
rect 383 529 439 563
rect 383 495 394 529
rect 428 495 439 529
rect 383 461 439 495
rect 383 427 394 461
rect 428 427 439 461
rect 383 367 439 427
rect 469 583 522 619
rect 469 549 480 583
rect 514 549 522 583
rect 469 367 522 549
rect 576 583 629 619
rect 576 549 584 583
rect 618 549 629 583
rect 576 367 629 549
rect 659 413 715 619
rect 659 379 670 413
rect 704 379 715 413
rect 659 367 715 379
rect 745 583 801 619
rect 745 549 756 583
rect 790 549 801 583
rect 745 367 801 549
rect 831 413 887 619
rect 831 379 842 413
rect 876 379 887 413
rect 831 367 887 379
rect 917 611 973 619
rect 917 577 928 611
rect 962 577 973 611
rect 917 367 973 577
rect 1003 541 1059 619
rect 1003 507 1014 541
rect 1048 507 1059 541
rect 1003 439 1059 507
rect 1003 405 1014 439
rect 1048 405 1059 439
rect 1003 367 1059 405
rect 1089 599 1145 619
rect 1089 565 1100 599
rect 1134 565 1145 599
rect 1089 525 1145 565
rect 1089 491 1100 525
rect 1134 491 1145 525
rect 1089 367 1145 491
rect 1175 541 1231 619
rect 1175 507 1186 541
rect 1220 507 1231 541
rect 1175 439 1231 507
rect 1175 405 1186 439
rect 1220 405 1231 439
rect 1175 367 1231 405
rect 1261 599 1314 619
rect 1261 565 1272 599
rect 1306 565 1314 599
rect 1261 527 1314 565
rect 1261 493 1272 527
rect 1306 493 1314 527
rect 1261 455 1314 493
rect 1261 421 1272 455
rect 1306 421 1314 455
rect 1261 367 1314 421
<< ndiffc >>
rect 82 153 116 187
rect 82 67 116 101
rect 177 164 211 198
rect 177 59 211 93
rect 270 153 304 187
rect 270 67 304 101
rect 364 92 398 126
rect 458 169 492 203
rect 458 67 492 101
rect 544 129 578 163
rect 544 55 578 89
rect 630 169 664 203
rect 630 67 664 101
rect 716 129 750 163
rect 716 55 750 89
rect 802 169 836 203
rect 802 67 836 101
rect 901 95 935 129
rect 1000 158 1034 192
rect 1000 67 1034 101
rect 1086 95 1120 129
rect 1172 169 1206 203
rect 1172 67 1206 101
rect 1258 129 1292 163
rect 1258 59 1292 93
<< pdiffc >>
rect 46 565 80 599
rect 46 473 80 507
rect 46 379 80 413
rect 136 573 170 607
rect 136 495 170 529
rect 136 421 170 455
rect 222 563 256 597
rect 222 495 256 529
rect 222 425 256 459
rect 308 573 342 607
rect 308 487 342 521
rect 394 563 428 597
rect 394 495 428 529
rect 394 427 428 461
rect 480 549 514 583
rect 584 549 618 583
rect 670 379 704 413
rect 756 549 790 583
rect 842 379 876 413
rect 928 577 962 611
rect 1014 507 1048 541
rect 1014 405 1048 439
rect 1100 565 1134 599
rect 1100 491 1134 525
rect 1186 507 1220 541
rect 1186 405 1220 439
rect 1272 565 1306 599
rect 1272 493 1306 527
rect 1272 421 1306 455
<< poly >>
rect 95 619 125 645
rect 181 619 211 645
rect 267 619 297 645
rect 353 619 383 645
rect 439 619 469 645
rect 629 619 659 645
rect 715 619 745 645
rect 801 619 831 645
rect 887 619 917 645
rect 973 619 1003 645
rect 1059 619 1089 645
rect 1145 619 1175 645
rect 1231 619 1261 645
rect 95 303 125 367
rect 181 345 211 367
rect 267 345 297 367
rect 353 345 383 367
rect 439 345 469 367
rect 629 345 659 367
rect 715 345 745 367
rect 801 345 831 367
rect 887 345 917 367
rect 181 315 537 345
rect 629 317 917 345
rect 973 317 1003 367
rect 1059 317 1089 367
rect 1145 317 1175 367
rect 1231 317 1261 367
rect 199 305 537 315
rect 73 287 139 303
rect 73 253 89 287
rect 123 267 139 287
rect 199 271 215 305
rect 249 271 283 305
rect 317 271 351 305
rect 385 271 419 305
rect 453 271 487 305
rect 521 271 537 305
rect 123 253 157 267
rect 199 255 537 271
rect 579 301 917 317
rect 579 267 595 301
rect 629 267 663 301
rect 697 267 731 301
rect 765 267 799 301
rect 833 267 867 301
rect 901 267 917 301
rect 73 237 157 253
rect 127 215 157 237
rect 229 215 259 255
rect 315 215 345 255
rect 417 215 447 255
rect 503 215 533 255
rect 579 251 917 267
rect 959 301 1261 317
rect 959 267 989 301
rect 1023 267 1057 301
rect 1091 267 1125 301
rect 1159 267 1193 301
rect 1227 267 1261 301
rect 959 251 1261 267
rect 589 215 619 251
rect 675 215 705 251
rect 761 215 791 251
rect 847 215 877 251
rect 959 215 989 251
rect 1045 215 1075 251
rect 1131 215 1161 251
rect 1217 215 1247 251
rect 127 21 157 47
rect 229 21 259 47
rect 315 21 345 47
rect 417 21 447 47
rect 503 21 533 47
rect 589 21 619 47
rect 675 21 705 47
rect 761 21 791 47
rect 847 21 877 47
rect 959 21 989 47
rect 1045 21 1075 47
rect 1131 21 1161 47
rect 1217 21 1247 47
<< polycont >>
rect 89 253 123 287
rect 215 271 249 305
rect 283 271 317 305
rect 351 271 385 305
rect 419 271 453 305
rect 487 271 521 305
rect 595 267 629 301
rect 663 267 697 301
rect 731 267 765 301
rect 799 267 833 301
rect 867 267 901 301
rect 989 267 1023 301
rect 1057 267 1091 301
rect 1125 267 1159 301
rect 1193 267 1227 301
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 19 599 84 615
rect 19 565 46 599
rect 80 565 84 599
rect 19 507 84 565
rect 19 473 46 507
rect 80 473 84 507
rect 19 413 84 473
rect 120 607 186 649
rect 120 573 136 607
rect 170 573 186 607
rect 120 529 186 573
rect 120 495 136 529
rect 170 495 186 529
rect 120 455 186 495
rect 120 421 136 455
rect 170 421 186 455
rect 220 597 258 613
rect 220 563 222 597
rect 256 563 258 597
rect 220 529 258 563
rect 220 495 222 529
rect 256 495 258 529
rect 220 459 258 495
rect 292 607 358 649
rect 292 573 308 607
rect 342 573 358 607
rect 292 521 358 573
rect 292 487 308 521
rect 342 487 358 521
rect 292 479 358 487
rect 392 597 430 613
rect 392 563 394 597
rect 428 563 430 597
rect 392 529 430 563
rect 464 583 530 649
rect 464 549 480 583
rect 514 549 530 583
rect 464 533 530 549
rect 580 611 1322 615
rect 580 583 928 611
rect 580 549 584 583
rect 618 549 756 583
rect 790 577 928 583
rect 962 599 1322 611
rect 962 577 1100 599
rect 790 575 1100 577
rect 790 549 806 575
rect 580 533 806 549
rect 1098 565 1100 575
rect 1134 577 1272 599
rect 1134 565 1136 577
rect 392 495 394 529
rect 428 499 430 529
rect 998 507 1014 541
rect 1048 507 1064 541
rect 998 499 1064 507
rect 428 495 1064 499
rect 220 425 222 459
rect 256 445 258 459
rect 392 465 1064 495
rect 1098 525 1136 565
rect 1270 565 1272 577
rect 1306 565 1322 599
rect 1098 491 1100 525
rect 1134 491 1136 525
rect 1098 475 1136 491
rect 1170 507 1186 541
rect 1220 507 1236 541
rect 392 461 444 465
rect 392 445 394 461
rect 256 427 394 445
rect 428 427 444 461
rect 998 441 1064 465
rect 1170 441 1236 507
rect 998 439 1236 441
rect 256 425 444 427
rect 19 379 46 413
rect 80 379 84 413
rect 220 409 444 425
rect 666 413 880 429
rect 19 375 84 379
rect 666 379 670 413
rect 704 379 842 413
rect 876 379 880 413
rect 998 405 1014 439
rect 1048 405 1186 439
rect 1220 405 1236 439
rect 1270 527 1322 565
rect 1270 493 1272 527
rect 1306 493 1322 527
rect 1270 455 1322 493
rect 1270 421 1272 455
rect 1306 421 1322 455
rect 1270 405 1322 421
rect 19 341 613 375
rect 19 203 55 341
rect 89 287 165 303
rect 123 253 165 287
rect 199 271 215 305
rect 249 271 283 305
rect 317 271 351 305
rect 385 271 419 305
rect 453 271 487 305
rect 521 271 537 305
rect 89 237 165 253
rect 223 265 537 271
rect 579 301 613 341
rect 666 371 880 379
rect 666 335 1327 371
rect 579 267 595 301
rect 629 267 663 301
rect 697 267 731 301
rect 765 267 799 301
rect 833 267 867 301
rect 901 267 917 301
rect 579 265 917 267
rect 973 267 989 301
rect 1023 267 1057 301
rect 1091 267 1125 301
rect 1159 267 1193 301
rect 1227 267 1243 301
rect 223 237 391 265
rect 973 242 1134 267
rect 1277 231 1327 335
rect 442 208 852 231
rect 1168 208 1327 231
rect 442 203 1327 208
rect 19 187 116 203
rect 19 153 82 187
rect 19 101 116 153
rect 19 67 82 101
rect 19 51 116 67
rect 161 198 227 203
rect 161 164 177 198
rect 211 164 227 198
rect 161 93 227 164
rect 161 59 177 93
rect 211 59 227 93
rect 161 17 227 59
rect 261 187 458 203
rect 261 153 270 187
rect 304 169 458 187
rect 492 197 630 203
rect 492 169 494 197
rect 304 153 314 169
rect 261 101 314 153
rect 261 67 270 101
rect 304 67 314 101
rect 261 51 314 67
rect 348 126 414 135
rect 348 92 364 126
rect 398 92 414 126
rect 348 17 414 92
rect 448 101 494 169
rect 628 169 630 197
rect 664 197 802 203
rect 664 169 666 197
rect 448 67 458 101
rect 492 67 494 101
rect 448 51 494 67
rect 528 129 544 163
rect 578 129 594 163
rect 528 89 594 129
rect 528 55 544 89
rect 578 55 594 89
rect 528 17 594 55
rect 628 101 666 169
rect 800 169 802 197
rect 836 192 1172 203
rect 836 174 1000 192
rect 836 169 851 174
rect 628 67 630 101
rect 664 67 666 101
rect 628 51 666 67
rect 700 129 716 163
rect 750 129 766 163
rect 700 89 766 129
rect 700 55 716 89
rect 750 55 766 89
rect 700 17 766 55
rect 800 101 851 169
rect 985 158 1000 174
rect 1034 174 1172 192
rect 1034 158 1036 174
rect 800 67 802 101
rect 836 67 851 101
rect 800 51 851 67
rect 885 129 951 140
rect 885 95 901 129
rect 935 95 951 129
rect 885 17 951 95
rect 985 101 1036 158
rect 1170 169 1172 174
rect 1206 197 1327 203
rect 1206 169 1208 197
rect 985 67 1000 101
rect 1034 67 1036 101
rect 985 51 1036 67
rect 1070 129 1136 140
rect 1070 95 1086 129
rect 1120 95 1136 129
rect 1070 17 1136 95
rect 1170 101 1208 169
rect 1170 67 1172 101
rect 1206 67 1208 101
rect 1170 51 1208 67
rect 1242 129 1258 163
rect 1292 129 1308 163
rect 1242 93 1308 129
rect 1242 59 1258 93
rect 1292 59 1308 93
rect 1242 17 1308 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor3b_4
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 C_N
port 3 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1174280
string GDS_START 1163396
<< end >>
