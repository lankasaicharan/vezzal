magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2066 1975
<< nwell >>
rect -38 331 806 704
<< pwell >>
rect 5 199 217 211
rect 5 49 767 199
rect 0 0 768 49
<< scnmos >>
rect 104 101 134 185
rect 206 89 236 173
rect 292 89 322 173
rect 410 89 440 173
rect 496 89 526 173
rect 582 89 612 173
rect 654 89 684 173
<< scpmoshvt >>
rect 101 419 151 619
rect 199 419 249 619
rect 326 419 376 619
rect 424 419 474 619
rect 522 419 572 619
rect 630 419 680 619
<< ndiff >>
rect 31 160 104 185
rect 31 126 43 160
rect 77 126 104 160
rect 31 101 104 126
rect 134 173 191 185
rect 134 139 145 173
rect 179 139 206 173
rect 134 101 206 139
rect 156 89 206 101
rect 236 139 292 173
rect 236 105 247 139
rect 281 105 292 139
rect 236 89 292 105
rect 322 89 410 173
rect 440 139 496 173
rect 440 105 451 139
rect 485 105 496 139
rect 440 89 496 105
rect 526 139 582 173
rect 526 105 537 139
rect 571 105 582 139
rect 526 89 582 105
rect 612 89 654 173
rect 684 148 741 173
rect 684 114 695 148
rect 729 114 741 148
rect 684 89 741 114
rect 337 74 395 89
rect 337 40 349 74
rect 383 40 395 74
rect 337 28 395 40
<< pdiff >>
rect 41 607 101 619
rect 41 573 53 607
rect 87 573 101 607
rect 41 536 101 573
rect 41 502 53 536
rect 87 502 101 536
rect 41 465 101 502
rect 41 431 53 465
rect 87 431 101 465
rect 41 419 101 431
rect 151 419 199 619
rect 249 597 326 619
rect 249 563 281 597
rect 315 563 326 597
rect 249 465 326 563
rect 249 431 281 465
rect 315 431 326 465
rect 249 419 326 431
rect 376 419 424 619
rect 474 419 522 619
rect 572 607 630 619
rect 572 573 583 607
rect 617 573 630 607
rect 572 512 630 573
rect 572 478 583 512
rect 617 478 630 512
rect 572 419 630 478
rect 680 597 737 619
rect 680 563 691 597
rect 725 563 737 597
rect 680 465 737 563
rect 680 431 691 465
rect 725 431 737 465
rect 680 419 737 431
<< ndiffc >>
rect 43 126 77 160
rect 145 139 179 173
rect 247 105 281 139
rect 451 105 485 139
rect 537 105 571 139
rect 695 114 729 148
rect 349 40 383 74
<< pdiffc >>
rect 53 573 87 607
rect 53 502 87 536
rect 53 431 87 465
rect 281 563 315 597
rect 281 431 315 465
rect 583 573 617 607
rect 583 478 617 512
rect 691 563 725 597
rect 691 431 725 465
<< poly >>
rect 101 619 151 645
rect 199 619 249 645
rect 326 619 376 645
rect 424 619 474 645
rect 522 619 572 645
rect 630 619 680 645
rect 101 393 151 419
rect 199 393 249 419
rect 326 404 376 419
rect 101 302 131 393
rect 199 351 229 393
rect 323 374 376 404
rect 424 393 474 419
rect 21 286 131 302
rect 21 252 37 286
rect 71 252 131 286
rect 179 335 245 351
rect 323 345 353 374
rect 179 301 195 335
rect 229 301 245 335
rect 179 285 245 301
rect 287 329 353 345
rect 424 332 454 393
rect 522 390 572 419
rect 522 345 552 390
rect 630 348 680 419
rect 287 295 303 329
rect 337 295 353 329
rect 21 236 131 252
rect 101 230 131 236
rect 101 200 134 230
rect 104 185 134 200
rect 206 173 236 285
rect 287 279 353 295
rect 395 316 461 332
rect 395 282 411 316
rect 445 282 461 316
rect 292 173 322 279
rect 395 266 461 282
rect 503 329 569 345
rect 503 295 519 329
rect 553 295 569 329
rect 503 279 569 295
rect 611 332 684 348
rect 611 298 627 332
rect 661 298 684 332
rect 410 173 440 266
rect 509 218 539 279
rect 611 264 684 298
rect 611 230 627 264
rect 661 230 684 264
rect 611 218 684 230
rect 496 188 539 218
rect 582 188 684 218
rect 496 173 526 188
rect 582 173 612 188
rect 654 173 684 188
rect 104 75 134 101
rect 206 63 236 89
rect 292 63 322 89
rect 410 63 440 89
rect 496 63 526 89
rect 582 63 612 89
rect 654 63 684 89
<< polycont >>
rect 37 252 71 286
rect 195 301 229 335
rect 303 295 337 329
rect 411 282 445 316
rect 519 295 553 329
rect 627 298 661 332
rect 627 230 661 264
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 37 607 87 649
rect 37 573 53 607
rect 281 597 331 613
rect 37 536 87 573
rect 37 502 53 536
rect 37 465 87 502
rect 37 431 53 465
rect 37 415 87 431
rect 21 286 87 356
rect 21 252 37 286
rect 71 252 87 286
rect 123 335 245 578
rect 315 563 331 597
rect 281 465 331 563
rect 315 431 331 465
rect 567 607 633 649
rect 567 573 583 607
rect 617 573 633 607
rect 567 512 633 573
rect 567 478 583 512
rect 617 478 633 512
rect 567 462 633 478
rect 675 597 747 613
rect 675 563 691 597
rect 725 563 747 597
rect 675 465 747 563
rect 281 426 331 431
rect 675 431 691 465
rect 725 431 747 465
rect 281 392 639 426
rect 123 301 195 335
rect 229 301 245 335
rect 123 285 245 301
rect 287 329 359 356
rect 287 295 303 329
rect 337 295 359 329
rect 287 279 359 295
rect 395 316 461 356
rect 395 282 411 316
rect 445 282 461 316
rect 395 266 461 282
rect 503 329 569 356
rect 503 295 519 329
rect 553 295 569 329
rect 503 279 569 295
rect 605 348 639 392
rect 675 384 747 431
rect 605 332 677 348
rect 605 298 627 332
rect 661 298 677 332
rect 21 236 87 252
rect 605 264 677 298
rect 605 230 627 264
rect 661 230 677 264
rect 129 214 677 230
rect 129 196 639 214
rect 27 160 93 189
rect 27 126 43 160
rect 77 126 93 160
rect 27 87 93 126
rect 129 173 195 196
rect 713 177 747 384
rect 129 139 145 173
rect 179 139 195 173
rect 129 123 195 139
rect 231 139 485 160
rect 231 105 247 139
rect 281 126 451 139
rect 281 105 297 126
rect 231 87 297 105
rect 435 105 451 126
rect 27 53 297 87
rect 333 74 399 90
rect 435 85 485 105
rect 521 139 587 160
rect 521 105 537 139
rect 571 105 587 139
rect 333 40 349 74
rect 383 40 399 74
rect 333 17 399 40
rect 521 17 587 105
rect 679 148 747 177
rect 679 114 695 148
rect 729 114 747 148
rect 679 85 747 114
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 683 768 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 768 683
rect 0 617 768 649
rect 0 17 768 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -49 768 -17
<< labels >>
flabel pwell s 0 0 768 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 768 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o32a_lp
flabel metal1 s 0 617 768 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 768 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 768 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1765314
string GDS_START 1757820
<< end >>
