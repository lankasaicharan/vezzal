magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 3410 1975
<< nwell >>
rect -38 332 2150 704
<< pwell >>
rect 1 49 2111 248
rect 0 0 2112 49
<< scpmos >>
rect 84 368 120 592
rect 183 368 219 592
rect 273 368 309 592
rect 363 368 399 592
rect 463 368 499 592
rect 563 368 599 592
rect 663 368 699 592
rect 763 368 799 592
rect 891 368 927 592
rect 991 368 1027 592
rect 1081 368 1117 592
rect 1191 368 1227 592
rect 1283 368 1319 592
rect 1391 368 1427 592
rect 1481 368 1517 592
rect 1581 368 1617 592
rect 1681 368 1717 592
rect 1781 368 1817 592
rect 1881 368 1917 592
rect 1992 368 2028 592
<< nmoslvt >>
rect 84 74 114 222
rect 184 74 214 222
rect 270 74 300 222
rect 369 74 399 222
rect 455 74 485 222
rect 541 74 571 222
rect 641 74 671 222
rect 727 74 757 222
rect 925 74 955 222
rect 1025 74 1055 222
rect 1111 74 1141 222
rect 1197 74 1227 222
rect 1283 74 1313 222
rect 1369 74 1399 222
rect 1456 74 1486 222
rect 1542 74 1572 222
rect 1740 74 1770 222
rect 1826 74 1856 222
rect 1912 74 1942 222
rect 1998 74 2028 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 136 184 222
rect 114 102 139 136
rect 173 102 184 136
rect 114 74 184 102
rect 214 210 270 222
rect 214 176 225 210
rect 259 176 270 210
rect 214 120 270 176
rect 214 86 225 120
rect 259 86 270 120
rect 214 74 270 86
rect 300 136 369 222
rect 300 102 311 136
rect 345 102 369 136
rect 300 74 369 102
rect 399 210 455 222
rect 399 176 410 210
rect 444 176 455 210
rect 399 120 455 176
rect 399 86 410 120
rect 444 86 455 120
rect 399 74 455 86
rect 485 189 541 222
rect 485 155 496 189
rect 530 155 541 189
rect 485 74 541 155
rect 571 123 641 222
rect 571 89 596 123
rect 630 89 641 123
rect 571 74 641 89
rect 671 210 727 222
rect 671 176 682 210
rect 716 176 727 210
rect 671 74 727 176
rect 757 123 814 222
rect 757 89 768 123
rect 802 89 814 123
rect 757 74 814 89
rect 868 136 925 222
rect 868 102 880 136
rect 914 102 925 136
rect 868 74 925 102
rect 955 207 1025 222
rect 955 173 980 207
rect 1014 173 1025 207
rect 955 74 1025 173
rect 1055 120 1111 222
rect 1055 86 1066 120
rect 1100 86 1111 120
rect 1055 74 1111 86
rect 1141 207 1197 222
rect 1141 173 1152 207
rect 1186 173 1197 207
rect 1141 74 1197 173
rect 1227 120 1283 222
rect 1227 86 1238 120
rect 1272 86 1283 120
rect 1227 74 1283 86
rect 1313 207 1369 222
rect 1313 173 1324 207
rect 1358 173 1369 207
rect 1313 74 1369 173
rect 1399 120 1456 222
rect 1399 86 1410 120
rect 1444 86 1456 120
rect 1399 74 1456 86
rect 1486 207 1542 222
rect 1486 173 1497 207
rect 1531 173 1542 207
rect 1486 74 1542 173
rect 1572 120 1629 222
rect 1572 86 1583 120
rect 1617 86 1629 120
rect 1572 74 1629 86
rect 1683 136 1740 222
rect 1683 102 1695 136
rect 1729 102 1740 136
rect 1683 74 1740 102
rect 1770 210 1826 222
rect 1770 176 1781 210
rect 1815 176 1826 210
rect 1770 120 1826 176
rect 1770 86 1781 120
rect 1815 86 1826 120
rect 1770 74 1826 86
rect 1856 136 1912 222
rect 1856 102 1867 136
rect 1901 102 1912 136
rect 1856 74 1912 102
rect 1942 210 1998 222
rect 1942 176 1953 210
rect 1987 176 1998 210
rect 1942 120 1998 176
rect 1942 86 1953 120
rect 1987 86 1998 120
rect 1942 74 1998 86
rect 2028 210 2085 222
rect 2028 176 2039 210
rect 2073 176 2085 210
rect 2028 120 2085 176
rect 2028 86 2039 120
rect 2073 86 2085 120
rect 2028 74 2085 86
<< pdiff >>
rect 27 580 84 592
rect 27 546 39 580
rect 73 546 84 580
rect 27 510 84 546
rect 27 476 39 510
rect 73 476 84 510
rect 27 440 84 476
rect 27 406 39 440
rect 73 406 84 440
rect 27 368 84 406
rect 120 531 183 592
rect 120 497 139 531
rect 173 497 183 531
rect 120 440 183 497
rect 120 406 139 440
rect 173 406 183 440
rect 120 368 183 406
rect 219 580 273 592
rect 219 546 229 580
rect 263 546 273 580
rect 219 508 273 546
rect 219 474 229 508
rect 263 474 273 508
rect 219 368 273 474
rect 309 531 363 592
rect 309 497 319 531
rect 353 497 363 531
rect 309 440 363 497
rect 309 406 319 440
rect 353 406 363 440
rect 309 368 363 406
rect 399 580 463 592
rect 399 546 419 580
rect 453 546 463 580
rect 399 508 463 546
rect 399 474 419 508
rect 453 474 463 508
rect 399 368 463 474
rect 499 531 563 592
rect 499 497 519 531
rect 553 497 563 531
rect 499 440 563 497
rect 499 406 519 440
rect 553 406 563 440
rect 499 368 563 406
rect 599 580 663 592
rect 599 546 619 580
rect 653 546 663 580
rect 599 508 663 546
rect 599 474 619 508
rect 653 474 663 508
rect 599 368 663 474
rect 699 531 763 592
rect 699 497 719 531
rect 753 497 763 531
rect 699 440 763 497
rect 699 406 719 440
rect 753 406 763 440
rect 699 368 763 406
rect 799 580 891 592
rect 799 546 819 580
rect 853 546 891 580
rect 799 508 891 546
rect 799 474 819 508
rect 853 474 891 508
rect 799 368 891 474
rect 927 578 991 592
rect 927 544 937 578
rect 971 544 991 578
rect 927 368 991 544
rect 1027 580 1081 592
rect 1027 546 1037 580
rect 1071 546 1081 580
rect 1027 508 1081 546
rect 1027 474 1037 508
rect 1071 474 1081 508
rect 1027 368 1081 474
rect 1117 578 1191 592
rect 1117 544 1137 578
rect 1171 544 1191 578
rect 1117 368 1191 544
rect 1227 580 1283 592
rect 1227 546 1237 580
rect 1271 546 1283 580
rect 1227 508 1283 546
rect 1227 474 1237 508
rect 1271 474 1283 508
rect 1227 368 1283 474
rect 1319 578 1391 592
rect 1319 544 1337 578
rect 1371 544 1391 578
rect 1319 368 1391 544
rect 1427 580 1481 592
rect 1427 546 1437 580
rect 1471 546 1481 580
rect 1427 510 1481 546
rect 1427 476 1437 510
rect 1471 476 1481 510
rect 1427 440 1481 476
rect 1427 406 1437 440
rect 1471 406 1481 440
rect 1427 368 1481 406
rect 1517 580 1581 592
rect 1517 546 1537 580
rect 1571 546 1581 580
rect 1517 508 1581 546
rect 1517 474 1537 508
rect 1571 474 1581 508
rect 1517 368 1581 474
rect 1617 580 1681 592
rect 1617 546 1637 580
rect 1671 546 1681 580
rect 1617 510 1681 546
rect 1617 476 1637 510
rect 1671 476 1681 510
rect 1617 440 1681 476
rect 1617 406 1637 440
rect 1671 406 1681 440
rect 1617 368 1681 406
rect 1717 580 1781 592
rect 1717 546 1737 580
rect 1771 546 1781 580
rect 1717 508 1781 546
rect 1717 474 1737 508
rect 1771 474 1781 508
rect 1717 368 1781 474
rect 1817 580 1881 592
rect 1817 546 1837 580
rect 1871 546 1881 580
rect 1817 510 1881 546
rect 1817 476 1837 510
rect 1871 476 1881 510
rect 1817 440 1881 476
rect 1817 406 1837 440
rect 1871 406 1881 440
rect 1817 368 1881 406
rect 1917 580 1992 592
rect 1917 546 1937 580
rect 1971 546 1992 580
rect 1917 508 1992 546
rect 1917 474 1937 508
rect 1971 474 1992 508
rect 1917 368 1992 474
rect 2028 580 2084 592
rect 2028 546 2038 580
rect 2072 546 2084 580
rect 2028 510 2084 546
rect 2028 476 2038 510
rect 2072 476 2084 510
rect 2028 440 2084 476
rect 2028 406 2038 440
rect 2072 406 2084 440
rect 2028 368 2084 406
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 139 102 173 136
rect 225 176 259 210
rect 225 86 259 120
rect 311 102 345 136
rect 410 176 444 210
rect 410 86 444 120
rect 496 155 530 189
rect 596 89 630 123
rect 682 176 716 210
rect 768 89 802 123
rect 880 102 914 136
rect 980 173 1014 207
rect 1066 86 1100 120
rect 1152 173 1186 207
rect 1238 86 1272 120
rect 1324 173 1358 207
rect 1410 86 1444 120
rect 1497 173 1531 207
rect 1583 86 1617 120
rect 1695 102 1729 136
rect 1781 176 1815 210
rect 1781 86 1815 120
rect 1867 102 1901 136
rect 1953 176 1987 210
rect 1953 86 1987 120
rect 2039 176 2073 210
rect 2039 86 2073 120
<< pdiffc >>
rect 39 546 73 580
rect 39 476 73 510
rect 39 406 73 440
rect 139 497 173 531
rect 139 406 173 440
rect 229 546 263 580
rect 229 474 263 508
rect 319 497 353 531
rect 319 406 353 440
rect 419 546 453 580
rect 419 474 453 508
rect 519 497 553 531
rect 519 406 553 440
rect 619 546 653 580
rect 619 474 653 508
rect 719 497 753 531
rect 719 406 753 440
rect 819 546 853 580
rect 819 474 853 508
rect 937 544 971 578
rect 1037 546 1071 580
rect 1037 474 1071 508
rect 1137 544 1171 578
rect 1237 546 1271 580
rect 1237 474 1271 508
rect 1337 544 1371 578
rect 1437 546 1471 580
rect 1437 476 1471 510
rect 1437 406 1471 440
rect 1537 546 1571 580
rect 1537 474 1571 508
rect 1637 546 1671 580
rect 1637 476 1671 510
rect 1637 406 1671 440
rect 1737 546 1771 580
rect 1737 474 1771 508
rect 1837 546 1871 580
rect 1837 476 1871 510
rect 1837 406 1871 440
rect 1937 546 1971 580
rect 1937 474 1971 508
rect 2038 546 2072 580
rect 2038 476 2072 510
rect 2038 406 2072 440
<< poly >>
rect 84 592 120 618
rect 183 592 219 618
rect 273 592 309 618
rect 363 592 399 618
rect 463 592 499 618
rect 563 592 599 618
rect 663 592 699 618
rect 763 592 799 618
rect 891 592 927 618
rect 991 592 1027 618
rect 1081 592 1117 618
rect 1191 592 1227 618
rect 1283 592 1319 618
rect 1391 592 1427 618
rect 1481 592 1517 618
rect 1581 592 1617 618
rect 1681 592 1717 618
rect 1781 592 1817 618
rect 1881 592 1917 618
rect 1992 592 2028 618
rect 84 336 120 368
rect 183 336 219 368
rect 273 336 309 368
rect 363 336 399 368
rect 463 336 499 368
rect 563 336 599 368
rect 663 336 699 368
rect 763 336 799 368
rect 84 320 399 336
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 304 320
rect 338 286 399 320
rect 84 270 399 286
rect 84 222 114 270
rect 184 222 214 270
rect 270 222 300 270
rect 369 222 399 270
rect 455 320 799 336
rect 455 286 471 320
rect 505 286 539 320
rect 573 286 607 320
rect 641 286 675 320
rect 709 286 743 320
rect 777 286 799 320
rect 455 270 799 286
rect 891 336 927 368
rect 991 336 1027 368
rect 1081 336 1117 368
rect 1191 336 1227 368
rect 891 320 1227 336
rect 891 286 907 320
rect 941 286 975 320
rect 1009 286 1043 320
rect 1077 286 1111 320
rect 1145 286 1227 320
rect 891 270 1227 286
rect 455 222 485 270
rect 541 222 571 270
rect 641 222 671 270
rect 727 222 757 270
rect 925 222 955 270
rect 1025 222 1055 270
rect 1111 222 1141 270
rect 1197 222 1227 270
rect 1283 336 1319 368
rect 1391 336 1427 368
rect 1481 336 1517 368
rect 1581 336 1617 368
rect 1283 320 1617 336
rect 1283 286 1363 320
rect 1397 286 1431 320
rect 1465 286 1499 320
rect 1533 286 1567 320
rect 1601 286 1617 320
rect 1681 336 1717 368
rect 1781 336 1817 368
rect 1881 336 1917 368
rect 1992 336 2028 368
rect 1681 320 2028 336
rect 1681 306 1769 320
rect 1283 270 1617 286
rect 1740 286 1769 306
rect 1803 286 1837 320
rect 1871 286 1905 320
rect 1939 286 1973 320
rect 2007 286 2028 320
rect 1740 270 2028 286
rect 1283 222 1313 270
rect 1369 222 1399 270
rect 1456 222 1486 270
rect 1542 222 1572 270
rect 1740 222 1770 270
rect 1826 222 1856 270
rect 1912 222 1942 270
rect 1998 222 2028 270
rect 84 48 114 74
rect 184 48 214 74
rect 270 48 300 74
rect 369 48 399 74
rect 455 48 485 74
rect 541 48 571 74
rect 641 48 671 74
rect 727 48 757 74
rect 925 48 955 74
rect 1025 48 1055 74
rect 1111 48 1141 74
rect 1197 48 1227 74
rect 1283 48 1313 74
rect 1369 48 1399 74
rect 1456 48 1486 74
rect 1542 48 1572 74
rect 1740 48 1770 74
rect 1826 48 1856 74
rect 1912 48 1942 74
rect 1998 48 2028 74
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 236 286 270 320
rect 304 286 338 320
rect 471 286 505 320
rect 539 286 573 320
rect 607 286 641 320
rect 675 286 709 320
rect 743 286 777 320
rect 907 286 941 320
rect 975 286 1009 320
rect 1043 286 1077 320
rect 1111 286 1145 320
rect 1363 286 1397 320
rect 1431 286 1465 320
rect 1499 286 1533 320
rect 1567 286 1601 320
rect 1769 286 1803 320
rect 1837 286 1871 320
rect 1905 286 1939 320
rect 1973 286 2007 320
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 23 581 869 615
rect 23 580 89 581
rect 23 546 39 580
rect 73 546 89 580
rect 229 580 263 581
rect 23 510 89 546
rect 23 476 39 510
rect 73 476 89 510
rect 23 440 89 476
rect 23 406 39 440
rect 73 406 89 440
rect 23 390 89 406
rect 123 531 189 547
rect 123 497 139 531
rect 173 497 189 531
rect 123 440 189 497
rect 403 580 469 581
rect 229 508 263 546
rect 229 458 263 474
rect 303 531 369 547
rect 303 497 319 531
rect 353 497 369 531
rect 123 406 139 440
rect 173 424 189 440
rect 303 440 369 497
rect 403 546 419 580
rect 453 546 469 580
rect 603 580 669 581
rect 403 508 469 546
rect 403 474 419 508
rect 453 474 469 508
rect 403 458 469 474
rect 503 531 569 547
rect 503 497 519 531
rect 553 497 569 531
rect 303 424 319 440
rect 173 406 319 424
rect 353 424 369 440
rect 503 440 569 497
rect 603 546 619 580
rect 653 546 669 580
rect 803 580 869 581
rect 603 508 669 546
rect 603 474 619 508
rect 653 474 669 508
rect 603 458 669 474
rect 703 531 769 547
rect 703 497 719 531
rect 753 497 769 531
rect 503 424 519 440
rect 353 406 519 424
rect 553 424 569 440
rect 703 440 769 497
rect 803 546 819 580
rect 853 546 869 580
rect 803 508 869 546
rect 921 578 987 649
rect 921 544 937 578
rect 971 544 987 578
rect 921 526 987 544
rect 1021 580 1087 596
rect 1021 546 1037 580
rect 1071 546 1087 580
rect 803 474 819 508
rect 853 492 869 508
rect 1021 508 1087 546
rect 1121 578 1187 649
rect 1121 544 1137 578
rect 1171 544 1187 578
rect 1121 526 1187 544
rect 1221 580 1287 596
rect 1221 546 1237 580
rect 1271 546 1287 580
rect 1021 492 1037 508
rect 853 474 1037 492
rect 1071 492 1087 508
rect 1221 508 1287 546
rect 1321 578 1387 649
rect 1321 544 1337 578
rect 1371 544 1387 578
rect 1321 526 1387 544
rect 1421 580 1487 596
rect 1421 546 1437 580
rect 1471 546 1487 580
rect 1221 492 1237 508
rect 1071 474 1237 492
rect 1271 492 1287 508
rect 1421 510 1487 546
rect 1421 492 1437 510
rect 1271 476 1437 492
rect 1471 476 1487 510
rect 1271 474 1487 476
rect 803 458 1487 474
rect 1521 580 1587 649
rect 1521 546 1537 580
rect 1571 546 1587 580
rect 1521 508 1587 546
rect 1521 474 1537 508
rect 1571 474 1587 508
rect 1521 458 1587 474
rect 1621 580 1687 596
rect 1621 546 1637 580
rect 1671 546 1687 580
rect 1621 510 1687 546
rect 1621 476 1637 510
rect 1671 476 1687 510
rect 703 424 719 440
rect 553 406 719 424
rect 753 424 769 440
rect 1421 440 1487 458
rect 753 406 1270 424
rect 123 390 1270 406
rect 1421 406 1437 440
rect 1471 424 1487 440
rect 1621 440 1687 476
rect 1721 580 1787 649
rect 1721 546 1737 580
rect 1771 546 1787 580
rect 1721 508 1787 546
rect 1721 474 1737 508
rect 1771 474 1787 508
rect 1721 458 1787 474
rect 1821 580 1887 596
rect 1821 546 1837 580
rect 1871 546 1887 580
rect 1821 510 1887 546
rect 1821 476 1837 510
rect 1871 476 1887 510
rect 1621 424 1637 440
rect 1471 406 1637 424
rect 1671 424 1687 440
rect 1821 440 1887 476
rect 1921 580 1987 649
rect 1921 546 1937 580
rect 1971 546 1987 580
rect 1921 508 1987 546
rect 1921 474 1937 508
rect 1971 474 1987 508
rect 1921 458 1987 474
rect 2022 580 2088 596
rect 2022 546 2038 580
rect 2072 546 2088 580
rect 2022 510 2088 546
rect 2022 476 2038 510
rect 2072 476 2088 510
rect 1821 424 1837 440
rect 1671 406 1837 424
rect 1871 424 1887 440
rect 2022 440 2088 476
rect 2022 424 2038 440
rect 1871 406 2038 424
rect 2072 406 2088 440
rect 1421 390 2088 406
rect 25 320 359 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 304 320
rect 338 286 359 320
rect 25 270 359 286
rect 409 320 839 356
rect 409 286 471 320
rect 505 286 539 320
rect 573 286 607 320
rect 641 286 675 320
rect 709 286 743 320
rect 777 286 839 320
rect 409 270 839 286
rect 889 320 1161 356
rect 889 286 907 320
rect 941 286 975 320
rect 1009 286 1043 320
rect 1077 286 1111 320
rect 1145 286 1161 320
rect 889 270 1161 286
rect 23 210 444 236
rect 23 176 39 210
rect 73 202 225 210
rect 73 176 89 202
rect 23 120 89 176
rect 259 202 410 210
rect 23 86 39 120
rect 73 86 89 120
rect 23 70 89 86
rect 123 136 189 168
rect 123 102 139 136
rect 173 102 189 136
rect 123 17 189 102
rect 225 120 259 176
rect 225 70 259 86
rect 295 136 361 168
rect 295 102 311 136
rect 345 102 361 136
rect 295 17 361 102
rect 410 120 444 176
rect 480 226 1030 236
rect 1236 226 1270 390
rect 1347 320 1703 356
rect 1347 286 1363 320
rect 1397 286 1431 320
rect 1465 286 1499 320
rect 1533 286 1567 320
rect 1601 286 1703 320
rect 1347 270 1703 286
rect 1753 320 2087 356
rect 1753 286 1769 320
rect 1803 286 1837 320
rect 1871 286 1905 320
rect 1939 286 1973 320
rect 2007 286 2087 320
rect 1753 270 2087 286
rect 480 210 1270 226
rect 480 189 682 210
rect 480 155 496 189
rect 530 176 682 189
rect 716 207 1270 210
rect 716 202 980 207
rect 716 176 732 202
rect 530 155 546 176
rect 964 173 980 202
rect 1014 173 1152 207
rect 1186 173 1270 207
rect 480 119 546 155
rect 580 123 646 142
rect 410 85 444 86
rect 580 89 596 123
rect 630 89 646 123
rect 580 85 646 89
rect 752 123 818 142
rect 752 89 768 123
rect 802 89 818 123
rect 752 85 818 89
rect 410 51 818 85
rect 864 136 930 168
rect 964 154 1270 173
rect 1308 210 1987 236
rect 1308 207 1781 210
rect 1308 173 1324 207
rect 1358 173 1497 207
rect 1531 202 1781 207
rect 1531 173 1547 202
rect 1308 170 1547 173
rect 1815 202 1953 210
rect 1308 154 1374 170
rect 1679 136 1745 168
rect 864 102 880 136
rect 914 120 930 136
rect 1567 120 1633 136
rect 914 102 1066 120
rect 864 86 1066 102
rect 1100 86 1238 120
rect 1272 86 1410 120
rect 1444 86 1583 120
rect 1617 86 1633 120
rect 864 70 1633 86
rect 1679 102 1695 136
rect 1729 102 1745 136
rect 1679 17 1745 102
rect 1781 120 1815 176
rect 1781 70 1815 86
rect 1851 136 1917 168
rect 1851 102 1867 136
rect 1901 102 1917 136
rect 1851 17 1917 102
rect 1953 120 1987 176
rect 1953 70 1987 86
rect 2023 210 2089 226
rect 2023 176 2039 210
rect 2073 176 2089 210
rect 2023 120 2089 176
rect 2023 86 2039 120
rect 2073 86 2089 120
rect 2023 17 2089 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
<< metal1 >>
rect 0 683 2112 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2112 683
rect 0 617 2112 649
rect 0 17 2112 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2112 17
rect 0 -49 2112 -17
<< labels >>
flabel pwell s 0 0 2112 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2112 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a32oi_4
flabel metal1 s 0 617 2112 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2112 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 1759 316 1793 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1855 316 1889 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 2047 316 2081 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1471 316 1505 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 991 168 1025 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1087 168 1121 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1183 168 1217 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2112 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 67956
string GDS_START 51380
<< end >>
