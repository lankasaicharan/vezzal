magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 23 49 639 160
rect 0 0 672 49
<< scnmos >>
rect 106 50 136 134
rect 242 50 272 134
rect 331 50 361 134
rect 422 50 452 134
rect 530 50 560 134
<< scpmoshvt >>
rect 150 483 180 611
rect 236 483 266 611
rect 322 483 352 611
rect 408 483 438 611
rect 494 483 524 611
<< ndiff >>
rect 49 92 106 134
rect 49 58 61 92
rect 95 58 106 92
rect 49 50 106 58
rect 136 92 242 134
rect 136 58 163 92
rect 197 58 242 92
rect 136 50 242 58
rect 272 50 331 134
rect 361 50 422 134
rect 452 109 530 134
rect 452 75 471 109
rect 505 75 530 109
rect 452 50 530 75
rect 560 109 613 134
rect 560 75 571 109
rect 605 75 613 109
rect 560 50 613 75
<< pdiff >>
rect 97 599 150 611
rect 97 565 105 599
rect 139 565 150 599
rect 97 529 150 565
rect 97 495 105 529
rect 139 495 150 529
rect 97 483 150 495
rect 180 599 236 611
rect 180 565 191 599
rect 225 565 236 599
rect 180 529 236 565
rect 180 495 191 529
rect 225 495 236 529
rect 180 483 236 495
rect 266 599 322 611
rect 266 565 277 599
rect 311 565 322 599
rect 266 529 322 565
rect 266 495 277 529
rect 311 495 322 529
rect 266 483 322 495
rect 352 599 408 611
rect 352 565 363 599
rect 397 565 408 599
rect 352 529 408 565
rect 352 495 363 529
rect 397 495 408 529
rect 352 483 408 495
rect 438 599 494 611
rect 438 565 449 599
rect 483 565 494 599
rect 438 529 494 565
rect 438 495 449 529
rect 483 495 494 529
rect 438 483 494 495
rect 524 599 577 611
rect 524 565 535 599
rect 569 565 577 599
rect 524 529 577 565
rect 524 495 535 529
rect 569 495 577 529
rect 524 483 577 495
<< ndiffc >>
rect 61 58 95 92
rect 163 58 197 92
rect 471 75 505 109
rect 571 75 605 109
<< pdiffc >>
rect 105 565 139 599
rect 105 495 139 529
rect 191 565 225 599
rect 191 495 225 529
rect 277 565 311 599
rect 277 495 311 529
rect 363 565 397 599
rect 363 495 397 529
rect 449 565 483 599
rect 449 495 483 529
rect 535 565 569 599
rect 535 495 569 529
<< poly >>
rect 150 611 180 637
rect 236 611 266 637
rect 322 611 352 637
rect 408 611 438 637
rect 494 611 524 637
rect 150 398 180 483
rect 86 368 180 398
rect 86 359 152 368
rect 86 325 102 359
rect 136 325 152 359
rect 86 291 152 325
rect 236 320 266 483
rect 86 257 102 291
rect 136 257 152 291
rect 86 241 152 257
rect 200 304 272 320
rect 200 270 216 304
rect 250 270 272 304
rect 322 302 352 483
rect 408 380 438 483
rect 494 458 524 483
rect 494 428 572 458
rect 408 350 458 380
rect 422 302 458 350
rect 530 302 572 428
rect 106 134 136 241
rect 200 236 272 270
rect 200 202 216 236
rect 250 202 272 236
rect 200 186 272 202
rect 242 134 272 186
rect 314 286 380 302
rect 314 252 330 286
rect 364 252 380 286
rect 314 218 380 252
rect 314 184 330 218
rect 364 184 380 218
rect 314 168 380 184
rect 422 286 488 302
rect 422 252 438 286
rect 472 252 488 286
rect 422 218 488 252
rect 422 184 438 218
rect 472 184 488 218
rect 422 168 488 184
rect 530 286 651 302
rect 530 252 601 286
rect 635 252 651 286
rect 530 218 651 252
rect 530 184 601 218
rect 635 184 651 218
rect 530 168 651 184
rect 331 134 361 168
rect 422 134 452 168
rect 530 134 560 168
rect 106 24 136 50
rect 242 24 272 50
rect 331 24 361 50
rect 422 24 452 50
rect 530 24 560 50
<< polycont >>
rect 102 325 136 359
rect 102 257 136 291
rect 216 270 250 304
rect 216 202 250 236
rect 330 252 364 286
rect 330 184 364 218
rect 438 252 472 286
rect 438 184 472 218
rect 601 252 635 286
rect 601 184 635 218
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 17 599 148 615
rect 17 565 105 599
rect 139 565 148 599
rect 17 529 148 565
rect 17 495 105 529
rect 139 495 148 529
rect 17 479 148 495
rect 182 599 234 649
rect 182 565 191 599
rect 225 565 234 599
rect 182 529 234 565
rect 182 495 191 529
rect 225 495 234 529
rect 182 479 234 495
rect 268 599 321 615
rect 268 565 277 599
rect 311 565 321 599
rect 268 529 321 565
rect 268 495 277 529
rect 311 495 321 529
rect 17 100 68 479
rect 268 445 321 495
rect 355 599 405 649
rect 355 565 363 599
rect 397 565 405 599
rect 355 529 405 565
rect 355 495 363 529
rect 397 495 405 529
rect 355 479 405 495
rect 439 599 491 615
rect 439 565 449 599
rect 483 565 491 599
rect 439 529 491 565
rect 439 495 449 529
rect 483 495 491 529
rect 439 445 491 495
rect 268 411 491 445
rect 525 599 585 615
rect 525 565 535 599
rect 569 565 585 599
rect 525 529 585 565
rect 525 495 535 529
rect 569 495 585 529
rect 525 479 585 495
rect 525 375 565 479
rect 102 359 565 375
rect 136 341 565 359
rect 136 325 152 341
rect 102 291 152 325
rect 136 257 152 291
rect 102 168 152 257
rect 200 270 216 304
rect 250 270 272 304
rect 200 236 272 270
rect 200 202 216 236
rect 250 202 272 236
rect 315 286 368 302
rect 315 252 330 286
rect 364 252 368 286
rect 315 218 368 252
rect 315 184 330 218
rect 364 184 368 218
rect 102 134 281 168
rect 315 159 368 184
rect 402 286 478 302
rect 402 252 438 286
rect 472 252 478 286
rect 402 218 478 252
rect 402 184 438 218
rect 472 184 478 218
rect 402 159 478 184
rect 599 286 655 368
rect 599 252 601 286
rect 635 252 655 286
rect 599 218 655 252
rect 599 184 601 218
rect 635 184 655 218
rect 599 159 655 184
rect 247 125 281 134
rect 247 109 521 125
rect 17 92 111 100
rect 17 58 61 92
rect 95 58 111 92
rect 17 54 111 58
rect 147 92 213 100
rect 147 58 163 92
rect 197 58 213 92
rect 247 75 471 109
rect 505 75 521 109
rect 247 59 521 75
rect 555 109 621 125
rect 555 75 571 109
rect 605 75 621 109
rect 147 17 213 58
rect 555 17 621 75
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a31o_0
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 415 168 449 202 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 31 94 65 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 168 65 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 464 65 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 31 538 65 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2646686
string GDS_START 2639328
<< end >>
