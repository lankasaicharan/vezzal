magic
tech sky130A
magscale 1 2
timestamp 1627201311
<< checkpaint >>
rect -1288 -1260 1388 2749
use sky130_fd_pr__hvdfm1sd__example_55959141808163  sky130_fd_pr__hvdfm1sd__example_55959141808163_0
timestamp 1627201311
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808163  sky130_fd_pr__hvdfm1sd__example_55959141808163_1
timestamp 1627201311
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 1489 128 1489 0 FreeSans 300 0 0 0 D
flabel comment s -28 1489 -28 1489 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 39926742
string GDS_START 39925688
<< end >>
