magic
tech sky130A
magscale 1 2
timestamp 1627202631
<< checkpaint >>
rect -1298 -1309 2642 1975
<< nwell >>
rect -38 332 1382 704
<< pwell >>
rect 466 248 1338 279
rect 7 49 1338 248
rect 0 0 1344 49
<< scnmos >>
rect 90 74 120 222
rect 176 74 206 222
rect 265 74 295 222
rect 351 74 381 222
rect 553 125 583 253
rect 649 125 679 253
rect 767 125 797 253
rect 853 125 883 253
rect 939 125 969 253
rect 1025 125 1055 253
rect 1125 125 1155 253
rect 1225 125 1255 253
<< scpmoshvt >>
rect 89 368 119 592
rect 179 368 209 592
rect 269 368 299 592
rect 359 368 389 592
rect 466 392 496 592
rect 556 392 586 592
rect 758 392 788 592
rect 848 392 878 592
rect 938 392 968 592
rect 1028 392 1058 592
rect 1128 392 1158 592
rect 1226 392 1256 592
<< ndiff >>
rect 33 210 90 222
rect 33 176 45 210
rect 79 176 90 210
rect 33 120 90 176
rect 33 86 45 120
rect 79 86 90 120
rect 33 74 90 86
rect 120 210 176 222
rect 120 176 131 210
rect 165 176 176 210
rect 120 120 176 176
rect 120 86 131 120
rect 165 86 176 120
rect 120 74 176 86
rect 206 131 265 222
rect 206 97 217 131
rect 251 97 265 131
rect 206 74 265 97
rect 295 210 351 222
rect 295 176 306 210
rect 340 176 351 210
rect 295 120 351 176
rect 295 86 306 120
rect 340 86 351 120
rect 295 74 351 86
rect 381 210 438 222
rect 381 176 392 210
rect 426 176 438 210
rect 381 120 438 176
rect 492 173 553 253
rect 492 139 504 173
rect 538 139 553 173
rect 492 125 553 139
rect 583 241 649 253
rect 583 207 604 241
rect 638 207 649 241
rect 583 171 649 207
rect 583 137 604 171
rect 638 137 649 171
rect 583 125 649 137
rect 679 241 767 253
rect 679 207 706 241
rect 740 207 767 241
rect 679 171 767 207
rect 679 137 706 171
rect 740 137 767 171
rect 679 125 767 137
rect 797 172 853 253
rect 797 138 808 172
rect 842 138 853 172
rect 797 125 853 138
rect 883 241 939 253
rect 883 207 894 241
rect 928 207 939 241
rect 883 171 939 207
rect 883 137 894 171
rect 928 137 939 171
rect 883 125 939 137
rect 969 172 1025 253
rect 969 138 980 172
rect 1014 138 1025 172
rect 969 125 1025 138
rect 1055 241 1125 253
rect 1055 207 1080 241
rect 1114 207 1125 241
rect 1055 171 1125 207
rect 1055 137 1080 171
rect 1114 137 1125 171
rect 1055 125 1125 137
rect 1155 172 1225 253
rect 1155 138 1166 172
rect 1200 138 1225 172
rect 1155 125 1225 138
rect 1255 241 1312 253
rect 1255 207 1266 241
rect 1300 207 1312 241
rect 1255 171 1312 207
rect 1255 137 1266 171
rect 1300 137 1312 171
rect 1255 125 1312 137
rect 381 86 392 120
rect 426 86 438 120
rect 381 74 438 86
<< pdiff >>
rect 30 580 89 592
rect 30 546 42 580
rect 76 546 89 580
rect 30 497 89 546
rect 30 463 42 497
rect 76 463 89 497
rect 30 414 89 463
rect 30 380 42 414
rect 76 380 89 414
rect 30 368 89 380
rect 119 580 179 592
rect 119 546 132 580
rect 166 546 179 580
rect 119 497 179 546
rect 119 463 132 497
rect 166 463 179 497
rect 119 414 179 463
rect 119 380 132 414
rect 166 380 179 414
rect 119 368 179 380
rect 209 580 269 592
rect 209 546 222 580
rect 256 546 269 580
rect 209 478 269 546
rect 209 444 222 478
rect 256 444 269 478
rect 209 368 269 444
rect 299 580 359 592
rect 299 546 312 580
rect 346 546 359 580
rect 299 497 359 546
rect 299 463 312 497
rect 346 463 359 497
rect 299 414 359 463
rect 299 380 312 414
rect 346 380 359 414
rect 299 368 359 380
rect 389 580 466 592
rect 389 546 402 580
rect 436 546 466 580
rect 389 497 466 546
rect 389 463 402 497
rect 436 463 466 497
rect 389 414 466 463
rect 389 380 402 414
rect 436 392 466 414
rect 496 580 556 592
rect 496 546 509 580
rect 543 546 556 580
rect 496 509 556 546
rect 496 475 509 509
rect 543 475 556 509
rect 496 438 556 475
rect 496 404 509 438
rect 543 404 556 438
rect 496 392 556 404
rect 586 578 645 592
rect 586 544 599 578
rect 633 544 645 578
rect 586 392 645 544
rect 699 441 758 592
rect 699 407 711 441
rect 745 407 758 441
rect 699 392 758 407
rect 788 580 848 592
rect 788 546 801 580
rect 835 546 848 580
rect 788 509 848 546
rect 788 475 801 509
rect 835 475 848 509
rect 788 392 848 475
rect 878 580 938 592
rect 878 546 891 580
rect 925 546 938 580
rect 878 512 938 546
rect 878 478 891 512
rect 925 478 938 512
rect 878 441 938 478
rect 878 407 891 441
rect 925 407 938 441
rect 878 392 938 407
rect 968 580 1028 592
rect 968 546 981 580
rect 1015 546 1028 580
rect 968 493 1028 546
rect 968 459 981 493
rect 1015 459 1028 493
rect 968 392 1028 459
rect 1058 577 1128 592
rect 1058 543 1071 577
rect 1105 543 1128 577
rect 1058 392 1128 543
rect 1158 580 1226 592
rect 1158 546 1171 580
rect 1205 546 1226 580
rect 1158 493 1226 546
rect 1158 459 1171 493
rect 1205 459 1226 493
rect 1158 392 1226 459
rect 1256 580 1317 592
rect 1256 546 1271 580
rect 1305 546 1317 580
rect 1256 510 1317 546
rect 1256 476 1271 510
rect 1305 476 1317 510
rect 1256 441 1317 476
rect 1256 407 1271 441
rect 1305 407 1317 441
rect 1256 392 1317 407
rect 436 380 448 392
rect 389 368 448 380
<< ndiffc >>
rect 45 176 79 210
rect 45 86 79 120
rect 131 176 165 210
rect 131 86 165 120
rect 217 97 251 131
rect 306 176 340 210
rect 306 86 340 120
rect 392 176 426 210
rect 504 139 538 173
rect 604 207 638 241
rect 604 137 638 171
rect 706 207 740 241
rect 706 137 740 171
rect 808 138 842 172
rect 894 207 928 241
rect 894 137 928 171
rect 980 138 1014 172
rect 1080 207 1114 241
rect 1080 137 1114 171
rect 1166 138 1200 172
rect 1266 207 1300 241
rect 1266 137 1300 171
rect 392 86 426 120
<< pdiffc >>
rect 42 546 76 580
rect 42 463 76 497
rect 42 380 76 414
rect 132 546 166 580
rect 132 463 166 497
rect 132 380 166 414
rect 222 546 256 580
rect 222 444 256 478
rect 312 546 346 580
rect 312 463 346 497
rect 312 380 346 414
rect 402 546 436 580
rect 402 463 436 497
rect 402 380 436 414
rect 509 546 543 580
rect 509 475 543 509
rect 509 404 543 438
rect 599 544 633 578
rect 711 407 745 441
rect 801 546 835 580
rect 801 475 835 509
rect 891 546 925 580
rect 891 478 925 512
rect 891 407 925 441
rect 981 546 1015 580
rect 981 459 1015 493
rect 1071 543 1105 577
rect 1171 546 1205 580
rect 1171 459 1205 493
rect 1271 546 1305 580
rect 1271 476 1305 510
rect 1271 407 1305 441
<< poly >>
rect 89 592 119 618
rect 179 592 209 618
rect 269 592 299 618
rect 359 592 389 618
rect 466 592 496 618
rect 556 592 586 618
rect 758 592 788 618
rect 848 592 878 618
rect 938 592 968 618
rect 1028 592 1058 618
rect 1128 592 1158 618
rect 1226 592 1256 618
rect 466 377 496 392
rect 556 377 586 392
rect 758 377 788 392
rect 848 377 878 392
rect 938 377 968 392
rect 1028 377 1058 392
rect 1128 377 1158 392
rect 1226 377 1256 392
rect 89 353 119 368
rect 179 353 209 368
rect 269 353 299 368
rect 359 353 389 368
rect 86 308 122 353
rect 176 326 212 353
rect 266 326 302 353
rect 356 326 392 353
rect 176 310 403 326
rect 176 308 217 310
rect 86 276 217 308
rect 251 276 285 310
rect 319 276 353 310
rect 387 276 403 310
rect 463 324 499 377
rect 553 360 589 377
rect 553 344 679 360
rect 755 357 791 377
rect 845 357 881 377
rect 553 324 597 344
rect 463 310 597 324
rect 631 310 679 344
rect 463 294 679 310
rect 86 260 403 276
rect 90 222 120 260
rect 176 222 206 260
rect 265 222 295 260
rect 351 222 381 260
rect 553 253 583 294
rect 649 253 679 294
rect 747 341 881 357
rect 747 307 763 341
rect 797 307 831 341
rect 865 321 881 341
rect 865 307 883 321
rect 747 291 883 307
rect 767 253 797 291
rect 853 253 883 291
rect 935 268 971 377
rect 1025 357 1061 377
rect 1125 357 1161 377
rect 1223 357 1259 377
rect 1025 341 1175 357
rect 1025 307 1125 341
rect 1159 307 1175 341
rect 1025 291 1175 307
rect 1223 341 1289 357
rect 1223 307 1239 341
rect 1273 307 1289 341
rect 1223 291 1289 307
rect 939 253 969 268
rect 1025 253 1055 291
rect 1125 253 1155 291
rect 1225 253 1255 291
rect 553 99 583 125
rect 649 99 679 125
rect 767 99 797 125
rect 853 99 883 125
rect 90 48 120 74
rect 176 48 206 74
rect 265 48 295 74
rect 351 48 381 74
rect 939 51 969 125
rect 1025 99 1055 125
rect 1125 99 1155 125
rect 1225 51 1255 125
rect 939 21 1255 51
<< polycont >>
rect 217 276 251 310
rect 285 276 319 310
rect 353 276 387 310
rect 597 310 631 344
rect 763 307 797 341
rect 831 307 865 341
rect 1125 307 1159 341
rect 1239 307 1273 341
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 26 580 76 649
rect 26 546 42 580
rect 26 497 76 546
rect 26 463 42 497
rect 26 414 76 463
rect 26 380 42 414
rect 26 364 76 380
rect 115 580 167 596
rect 115 546 132 580
rect 166 546 167 580
rect 115 497 167 546
rect 115 463 132 497
rect 166 463 167 497
rect 115 414 167 463
rect 206 580 256 649
rect 206 546 222 580
rect 206 478 256 546
rect 206 444 222 478
rect 206 428 256 444
rect 296 580 362 596
rect 296 546 312 580
rect 346 546 362 580
rect 296 497 362 546
rect 296 463 312 497
rect 346 463 362 497
rect 115 380 132 414
rect 166 394 167 414
rect 296 414 362 463
rect 296 394 312 414
rect 166 380 312 394
rect 346 380 362 414
rect 115 360 362 380
rect 402 580 452 649
rect 436 546 452 580
rect 402 497 452 546
rect 436 463 452 497
rect 402 414 452 463
rect 436 380 452 414
rect 402 364 452 380
rect 493 580 543 596
rect 493 546 509 580
rect 493 509 543 546
rect 583 578 649 649
rect 583 544 599 578
rect 633 544 649 578
rect 583 543 649 544
rect 785 580 851 596
rect 785 546 801 580
rect 835 546 851 580
rect 785 509 851 546
rect 493 475 509 509
rect 543 475 801 509
rect 835 475 851 509
rect 887 580 929 596
rect 887 546 891 580
rect 925 546 929 580
rect 887 512 929 546
rect 887 478 891 512
rect 925 478 929 512
rect 493 438 543 475
rect 887 441 929 478
rect 965 580 1015 596
rect 965 546 981 580
rect 965 493 1015 546
rect 1055 577 1121 649
rect 1055 543 1071 577
rect 1105 543 1121 577
rect 1055 527 1121 543
rect 1155 580 1221 596
rect 1155 546 1171 580
rect 1205 546 1221 580
rect 1155 493 1221 546
rect 965 459 981 493
rect 1015 459 1171 493
rect 1205 459 1221 493
rect 1255 580 1321 596
rect 1255 546 1271 580
rect 1305 546 1321 580
rect 1255 510 1321 546
rect 1255 476 1271 510
rect 1305 476 1321 510
rect 493 404 509 438
rect 115 226 167 360
rect 493 326 543 404
rect 201 310 543 326
rect 201 276 217 310
rect 251 276 285 310
rect 319 276 353 310
rect 387 276 543 310
rect 581 344 647 430
rect 695 407 711 441
rect 745 407 891 441
rect 925 425 929 441
rect 1255 441 1321 476
rect 1255 425 1271 441
rect 925 407 1271 425
rect 1305 407 1321 441
rect 695 391 1321 407
rect 581 310 597 344
rect 631 310 647 344
rect 581 294 647 310
rect 697 341 1031 357
rect 697 307 763 341
rect 797 307 831 341
rect 865 307 1031 341
rect 697 291 1031 307
rect 1081 341 1175 357
rect 1081 307 1125 341
rect 1159 307 1175 341
rect 1081 291 1175 307
rect 1223 341 1319 357
rect 1223 307 1239 341
rect 1273 307 1319 341
rect 1223 291 1319 307
rect 201 260 543 276
rect 509 241 654 260
rect 509 226 604 241
rect 29 210 79 226
rect 29 176 45 210
rect 29 120 79 176
rect 29 86 45 120
rect 29 17 79 86
rect 115 210 340 226
rect 115 176 131 210
rect 165 192 306 210
rect 165 176 181 192
rect 115 120 181 176
rect 290 176 306 192
rect 115 86 131 120
rect 165 86 181 120
rect 115 70 181 86
rect 217 131 251 158
rect 217 17 251 97
rect 290 120 340 176
rect 290 86 306 120
rect 290 70 340 86
rect 376 210 442 226
rect 376 176 392 210
rect 426 176 442 210
rect 588 207 604 226
rect 638 207 654 241
rect 376 120 442 176
rect 376 86 392 120
rect 426 86 442 120
rect 376 17 442 86
rect 488 173 554 192
rect 488 139 504 173
rect 538 139 554 173
rect 488 87 554 139
rect 588 171 654 207
rect 588 137 604 171
rect 638 137 654 171
rect 588 121 654 137
rect 690 241 1316 257
rect 690 207 706 241
rect 740 223 894 241
rect 740 207 756 223
rect 690 171 756 207
rect 878 207 894 223
rect 928 223 1080 241
rect 690 137 706 171
rect 740 137 756 171
rect 690 87 756 137
rect 488 53 756 87
rect 792 172 842 189
rect 792 138 808 172
rect 792 17 842 138
rect 878 171 928 207
rect 1064 207 1080 223
rect 1114 223 1266 241
rect 878 137 894 171
rect 878 121 928 137
rect 964 172 1030 189
rect 964 138 980 172
rect 1014 138 1030 172
rect 964 17 1030 138
rect 1064 171 1114 207
rect 1250 207 1266 223
rect 1300 207 1316 241
rect 1064 137 1080 171
rect 1064 121 1114 137
rect 1150 172 1216 189
rect 1150 138 1166 172
rect 1200 138 1216 172
rect 1150 17 1216 138
rect 1250 171 1316 207
rect 1250 137 1266 171
rect 1300 137 1316 171
rect 1250 121 1316 137
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
<< metal1 >>
rect 0 683 1344 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1344 683
rect 0 617 1344 649
rect 0 17 1344 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1344 17
rect 0 -49 1344 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o31a_4
flabel pwell s 0 0 1344 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 1344 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 0 617 1344 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 0 0 1344 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1344 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ls/gds/sky130_fd_sc_ls.gds
string LEFsymmetry X Y
string GDS_END 553920
string GDS_START 541666
<< end >>
