magic
tech sky130A
magscale 1 2
timestamp 1627202617
<< checkpaint >>
rect -1298 -1308 2402 1852
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 8 67 1103 203
rect 29 -17 63 67
rect 285 21 1103 67
<< scnmos >>
rect 86 93 116 177
rect 175 93 205 177
rect 363 47 393 177
rect 469 47 499 177
rect 553 47 583 177
rect 637 47 667 177
rect 743 47 773 177
rect 827 47 857 177
rect 911 47 941 177
rect 995 47 1025 177
<< scpmoshvt >>
rect 79 410 109 494
rect 176 297 206 381
rect 367 297 397 497
rect 469 297 499 497
rect 553 297 583 497
rect 637 297 667 497
rect 743 297 773 497
rect 827 297 857 497
rect 911 297 941 497
rect 995 297 1025 497
<< ndiff >>
rect 34 149 86 177
rect 34 115 42 149
rect 76 115 86 149
rect 34 93 86 115
rect 116 149 175 177
rect 116 115 131 149
rect 165 115 175 149
rect 116 93 175 115
rect 205 149 257 177
rect 205 115 215 149
rect 249 115 257 149
rect 205 93 257 115
rect 311 96 363 177
rect 311 62 319 96
rect 353 62 363 96
rect 311 47 363 62
rect 393 115 469 177
rect 393 81 419 115
rect 453 81 469 115
rect 393 47 469 81
rect 499 97 553 177
rect 499 63 509 97
rect 543 63 553 97
rect 499 47 553 63
rect 583 115 637 177
rect 583 81 593 115
rect 627 81 637 115
rect 583 47 637 81
rect 667 97 743 177
rect 667 63 697 97
rect 731 63 743 97
rect 667 47 743 63
rect 773 114 827 177
rect 773 80 783 114
rect 817 80 827 114
rect 773 47 827 80
rect 857 95 911 177
rect 857 61 867 95
rect 901 61 911 95
rect 857 47 911 61
rect 941 163 995 177
rect 941 129 951 163
rect 985 129 995 163
rect 941 95 995 129
rect 941 61 951 95
rect 985 61 995 95
rect 941 47 995 61
rect 1025 95 1077 177
rect 1025 61 1035 95
rect 1069 61 1077 95
rect 1025 47 1077 61
<< pdiff >>
rect 27 475 79 494
rect 27 441 35 475
rect 69 441 79 475
rect 27 410 79 441
rect 109 475 161 494
rect 109 441 119 475
rect 153 441 161 475
rect 109 410 161 441
rect 124 381 161 410
rect 315 425 367 497
rect 315 391 323 425
rect 357 391 367 425
rect 124 297 176 381
rect 206 350 256 381
rect 315 380 367 391
rect 206 339 262 350
rect 206 305 216 339
rect 250 305 262 339
rect 206 297 262 305
rect 316 297 367 380
rect 397 297 469 497
rect 499 297 553 497
rect 583 297 637 497
rect 667 477 743 497
rect 667 443 688 477
rect 722 443 743 477
rect 667 409 743 443
rect 667 375 688 409
rect 722 375 743 409
rect 667 297 743 375
rect 773 477 827 497
rect 773 443 783 477
rect 817 443 827 477
rect 773 409 827 443
rect 773 375 783 409
rect 817 375 827 409
rect 773 341 827 375
rect 773 307 783 341
rect 817 307 827 341
rect 773 297 827 307
rect 857 477 911 497
rect 857 443 867 477
rect 901 443 911 477
rect 857 409 911 443
rect 857 375 867 409
rect 901 375 911 409
rect 857 297 911 375
rect 941 477 995 497
rect 941 443 951 477
rect 985 443 995 477
rect 941 409 995 443
rect 941 375 951 409
rect 985 375 995 409
rect 941 341 995 375
rect 941 307 951 341
rect 985 307 995 341
rect 941 297 995 307
rect 1025 477 1077 497
rect 1025 443 1035 477
rect 1069 443 1077 477
rect 1025 409 1077 443
rect 1025 375 1035 409
rect 1069 375 1077 409
rect 1025 297 1077 375
<< ndiffc >>
rect 42 115 76 149
rect 131 115 165 149
rect 215 115 249 149
rect 319 62 353 96
rect 419 81 453 115
rect 509 63 543 97
rect 593 81 627 115
rect 697 63 731 97
rect 783 80 817 114
rect 867 61 901 95
rect 951 129 985 163
rect 951 61 985 95
rect 1035 61 1069 95
<< pdiffc >>
rect 35 441 69 475
rect 119 441 153 475
rect 323 391 357 425
rect 216 305 250 339
rect 688 443 722 477
rect 688 375 722 409
rect 783 443 817 477
rect 783 375 817 409
rect 783 307 817 341
rect 867 443 901 477
rect 867 375 901 409
rect 951 443 985 477
rect 951 375 985 409
rect 951 307 985 341
rect 1035 443 1069 477
rect 1035 375 1069 409
<< poly >>
rect 79 494 109 520
rect 367 497 397 523
rect 469 497 499 523
rect 553 497 583 523
rect 637 497 667 523
rect 743 497 773 523
rect 827 497 857 523
rect 911 497 941 523
rect 995 497 1025 523
rect 79 265 109 410
rect 176 381 206 407
rect 176 265 206 297
rect 367 265 397 297
rect 469 265 499 297
rect 553 265 583 297
rect 637 265 667 297
rect 743 265 773 297
rect 827 265 857 297
rect 911 265 941 297
rect 995 265 1025 297
rect 75 249 129 265
rect 75 215 85 249
rect 119 215 129 249
rect 75 199 129 215
rect 173 249 239 265
rect 173 215 189 249
rect 223 215 239 249
rect 173 199 239 215
rect 295 249 397 265
rect 295 215 305 249
rect 339 215 397 249
rect 295 199 397 215
rect 445 249 499 265
rect 445 215 455 249
rect 489 215 499 249
rect 445 199 499 215
rect 541 249 595 265
rect 541 215 551 249
rect 585 215 595 249
rect 541 199 595 215
rect 637 249 691 265
rect 637 215 647 249
rect 681 215 691 249
rect 637 199 691 215
rect 743 249 1025 265
rect 743 215 753 249
rect 787 215 821 249
rect 855 215 889 249
rect 923 215 957 249
rect 991 215 1025 249
rect 743 199 1025 215
rect 86 177 116 199
rect 175 177 205 199
rect 363 177 393 199
rect 469 177 499 199
rect 553 177 583 199
rect 637 177 667 199
rect 743 177 773 199
rect 827 177 857 199
rect 911 177 941 199
rect 995 177 1025 199
rect 86 67 116 93
rect 175 67 205 93
rect 363 21 393 47
rect 469 21 499 47
rect 553 21 583 47
rect 637 21 667 47
rect 743 21 773 47
rect 827 21 857 47
rect 911 21 941 47
rect 995 21 1025 47
<< polycont >>
rect 85 215 119 249
rect 189 215 223 249
rect 305 215 339 249
rect 455 215 489 249
rect 551 215 585 249
rect 647 215 681 249
rect 753 215 787 249
rect 821 215 855 249
rect 889 215 923 249
rect 957 215 991 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 17 475 69 491
rect 17 441 35 475
rect 103 475 169 527
rect 103 441 119 475
rect 153 441 169 475
rect 225 459 489 493
rect 680 477 730 527
rect 17 407 69 441
rect 225 407 259 459
rect 17 373 259 407
rect 302 391 323 425
rect 357 391 421 425
rect 17 165 51 373
rect 85 249 155 339
rect 198 305 216 339
rect 250 305 319 339
rect 281 265 319 305
rect 119 215 155 249
rect 85 199 155 215
rect 189 249 247 265
rect 223 215 247 249
rect 189 199 247 215
rect 281 249 339 265
rect 281 215 305 249
rect 281 199 339 215
rect 281 165 319 199
rect 17 149 80 165
rect 17 115 42 149
rect 76 115 80 149
rect 17 90 80 115
rect 131 149 165 165
rect 131 17 165 115
rect 215 149 319 165
rect 249 131 319 149
rect 387 165 421 391
rect 455 249 489 459
rect 559 357 623 475
rect 680 443 688 477
rect 722 443 730 477
rect 680 409 730 443
rect 680 375 688 409
rect 722 375 730 409
rect 680 359 730 375
rect 775 477 825 493
rect 775 443 783 477
rect 817 443 825 477
rect 775 409 825 443
rect 775 375 783 409
rect 817 375 825 409
rect 559 290 601 357
rect 775 341 825 375
rect 859 477 909 527
rect 859 443 867 477
rect 901 443 909 477
rect 859 409 909 443
rect 859 375 867 409
rect 901 375 909 409
rect 859 359 909 375
rect 943 477 993 493
rect 943 443 951 477
rect 985 443 993 477
rect 943 409 993 443
rect 943 375 951 409
rect 985 375 993 409
rect 455 199 489 215
rect 535 249 601 290
rect 535 215 551 249
rect 585 215 601 249
rect 535 199 601 215
rect 647 289 734 323
rect 775 307 783 341
rect 817 325 825 341
rect 943 341 993 375
rect 1027 477 1077 527
rect 1027 443 1035 477
rect 1069 443 1077 477
rect 1027 409 1077 443
rect 1027 375 1035 409
rect 1069 375 1077 409
rect 1027 359 1077 375
rect 943 325 951 341
rect 817 307 951 325
rect 985 325 993 341
rect 985 307 1087 325
rect 775 291 1087 307
rect 647 249 681 289
rect 647 199 681 215
rect 715 215 753 249
rect 787 215 821 249
rect 855 215 889 249
rect 923 215 957 249
rect 991 215 1007 249
rect 715 165 749 215
rect 1041 181 1087 291
rect 387 131 749 165
rect 783 163 1087 181
rect 783 145 951 163
rect 215 90 249 115
rect 419 115 453 131
rect 303 62 319 96
rect 353 62 369 96
rect 303 17 369 62
rect 593 115 627 131
rect 419 61 453 81
rect 493 63 509 97
rect 543 63 559 97
rect 493 17 559 63
rect 783 114 833 145
rect 593 61 627 81
rect 671 63 697 97
rect 731 63 747 97
rect 671 17 747 63
rect 817 80 833 114
rect 935 129 951 145
rect 985 145 1087 163
rect 985 129 1001 145
rect 783 51 833 80
rect 867 95 901 111
rect 867 17 901 61
rect 935 95 1001 129
rect 935 61 951 95
rect 985 61 1001 95
rect 935 51 1001 61
rect 1035 95 1069 111
rect 1035 17 1069 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 585 425 619 459 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 585 357 619 391 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 677 289 711 323 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel locali s 1045 153 1079 187 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 or4bb_4
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 3880124
string GDS_START 3871366
string path 0.000 0.000 27.600 0.000 
<< end >>
