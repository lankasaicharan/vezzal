magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 2126 1852
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 157 618 203
rect 1 67 827 157
rect 29 21 827 67
rect 29 -17 63 21
<< scnmos >>
rect 79 93 109 177
rect 188 47 218 177
rect 304 47 334 177
rect 404 47 434 177
rect 500 47 530 177
rect 698 47 728 131
<< scpmoshvt >>
rect 81 413 117 497
rect 190 297 226 497
rect 306 297 342 497
rect 406 297 442 497
rect 502 297 538 497
rect 700 413 736 497
<< ndiff >>
rect 27 139 79 177
rect 27 105 35 139
rect 69 105 79 139
rect 27 93 79 105
rect 109 93 188 177
rect 134 59 142 93
rect 176 59 188 93
rect 134 47 188 59
rect 218 47 304 177
rect 334 47 404 177
rect 434 47 500 177
rect 530 161 592 177
rect 530 127 550 161
rect 584 127 592 161
rect 530 93 592 127
rect 530 59 550 93
rect 584 59 592 93
rect 530 47 592 59
rect 646 93 698 131
rect 646 59 654 93
rect 688 59 698 93
rect 646 47 698 59
rect 728 93 801 131
rect 728 59 758 93
rect 792 59 801 93
rect 728 47 801 59
<< pdiff >>
rect 27 485 81 497
rect 27 451 35 485
rect 69 451 81 485
rect 27 413 81 451
rect 117 485 190 497
rect 117 451 142 485
rect 176 451 190 485
rect 117 417 190 451
rect 117 413 142 417
rect 134 383 142 413
rect 176 383 190 417
rect 134 297 190 383
rect 226 485 306 497
rect 226 451 247 485
rect 281 451 306 485
rect 226 417 306 451
rect 226 383 247 417
rect 281 383 306 417
rect 226 349 306 383
rect 226 315 247 349
rect 281 315 306 349
rect 226 297 306 315
rect 342 485 406 497
rect 342 451 355 485
rect 389 451 406 485
rect 342 417 406 451
rect 342 383 355 417
rect 389 383 406 417
rect 342 297 406 383
rect 442 485 502 497
rect 442 451 454 485
rect 488 451 502 485
rect 442 417 502 451
rect 442 383 454 417
rect 488 383 502 417
rect 442 349 502 383
rect 442 315 454 349
rect 488 315 502 349
rect 442 297 502 315
rect 538 485 700 497
rect 538 451 550 485
rect 584 451 654 485
rect 688 451 700 485
rect 538 413 700 451
rect 736 477 801 497
rect 736 443 748 477
rect 782 443 801 477
rect 736 413 801 443
rect 538 297 592 413
<< ndiffc >>
rect 35 105 69 139
rect 142 59 176 93
rect 550 127 584 161
rect 550 59 584 93
rect 654 59 688 93
rect 758 59 792 93
<< pdiffc >>
rect 35 451 69 485
rect 142 451 176 485
rect 142 383 176 417
rect 247 451 281 485
rect 247 383 281 417
rect 247 315 281 349
rect 355 451 389 485
rect 355 383 389 417
rect 454 451 488 485
rect 454 383 488 417
rect 454 315 488 349
rect 550 451 584 485
rect 654 451 688 485
rect 748 443 782 477
<< poly >>
rect 81 497 117 523
rect 190 497 226 523
rect 306 497 342 523
rect 406 497 442 523
rect 502 497 538 523
rect 700 497 736 523
rect 81 398 117 413
rect 79 265 119 398
rect 700 398 736 413
rect 190 282 226 297
rect 306 282 342 297
rect 406 282 442 297
rect 502 282 538 297
rect 188 265 228 282
rect 304 265 344 282
rect 404 265 444 282
rect 500 265 540 282
rect 79 249 146 265
rect 79 215 102 249
rect 136 215 146 249
rect 79 199 146 215
rect 188 249 262 265
rect 188 215 215 249
rect 249 215 262 249
rect 188 199 262 215
rect 304 249 362 265
rect 304 215 318 249
rect 352 215 362 249
rect 304 199 362 215
rect 404 249 458 265
rect 404 215 414 249
rect 448 215 458 249
rect 404 199 458 215
rect 500 249 614 265
rect 500 215 570 249
rect 604 215 614 249
rect 500 199 614 215
rect 698 264 738 398
rect 698 248 762 264
rect 698 214 708 248
rect 742 214 762 248
rect 79 177 109 199
rect 188 177 218 199
rect 304 177 334 199
rect 404 177 434 199
rect 500 177 530 199
rect 698 198 762 214
rect 79 67 109 93
rect 698 131 728 198
rect 188 21 218 47
rect 304 21 334 47
rect 404 21 434 47
rect 500 21 530 47
rect 698 21 728 47
<< polycont >>
rect 102 215 136 249
rect 215 215 249 249
rect 318 215 352 249
rect 414 215 448 249
rect 570 215 604 249
rect 708 214 742 248
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 485 85 493
rect 17 451 35 485
rect 69 451 85 485
rect 17 413 85 451
rect 129 485 195 527
rect 129 451 142 485
rect 176 451 195 485
rect 129 417 195 451
rect 17 181 52 413
rect 129 383 142 417
rect 176 383 195 417
rect 129 367 195 383
rect 231 485 297 493
rect 231 451 247 485
rect 281 451 297 485
rect 231 417 297 451
rect 231 383 247 417
rect 281 383 297 417
rect 231 349 297 383
rect 339 485 403 527
rect 339 451 355 485
rect 389 451 403 485
rect 339 417 403 451
rect 339 383 355 417
rect 389 383 403 417
rect 339 367 403 383
rect 438 485 516 493
rect 438 451 454 485
rect 488 451 516 485
rect 438 417 516 451
rect 550 485 704 527
rect 584 451 654 485
rect 688 451 704 485
rect 550 435 704 451
rect 748 477 811 493
rect 782 443 811 477
rect 438 383 454 417
rect 488 401 516 417
rect 748 401 811 443
rect 488 383 536 401
rect 86 249 165 331
rect 231 315 247 349
rect 281 333 297 349
rect 438 349 536 383
rect 438 333 454 349
rect 281 315 454 333
rect 488 315 536 349
rect 231 299 536 315
rect 86 215 102 249
rect 136 215 165 249
rect 199 249 265 265
rect 199 215 215 249
rect 249 215 265 249
rect 299 249 352 265
rect 299 215 318 249
rect 17 143 244 181
rect 299 147 352 215
rect 398 249 448 265
rect 398 215 414 249
rect 17 139 85 143
rect 17 105 35 139
rect 69 105 85 139
rect 210 111 244 143
rect 398 111 448 215
rect 17 97 85 105
rect 129 93 176 109
rect 129 59 142 93
rect 210 73 448 111
rect 482 165 536 299
rect 570 367 811 401
rect 570 249 625 367
rect 604 215 625 249
rect 570 199 625 215
rect 660 248 742 323
rect 660 214 708 248
rect 482 161 600 165
rect 482 127 550 161
rect 584 127 600 161
rect 660 145 742 214
rect 482 93 600 127
rect 777 109 811 367
rect 129 17 176 59
rect 482 59 550 93
rect 584 59 600 93
rect 482 51 600 59
rect 638 93 708 109
rect 638 59 654 93
rect 688 59 708 93
rect 638 17 708 59
rect 742 93 811 109
rect 742 59 758 93
rect 792 59 811 93
rect 742 51 811 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 318 221 352 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 220 221 254 255 0 FreeSans 250 0 0 0 D
port 4 nsew signal input
flabel locali s 692 289 726 323 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel locali s 692 221 726 255 0 FreeSans 250 0 0 0 A_N
port 1 nsew signal input
flabel locali s 490 289 524 323 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 490 221 524 255 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 490 153 524 187 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 113 221 147 255 0 FreeSans 250 0 0 0 B_N
port 2 nsew signal input
flabel locali s 490 85 524 119 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 nand4bb_1
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 2284458
string GDS_START 2277126
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
