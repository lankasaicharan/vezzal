magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 2162 1975
<< nwell >>
rect -38 331 902 704
<< pwell >>
rect 6 49 837 241
rect 0 0 864 49
<< scnmos >>
rect 85 47 115 215
rect 171 47 201 215
rect 311 47 341 215
rect 397 47 427 215
rect 541 47 571 215
rect 627 47 657 215
rect 721 47 751 215
<< scpmoshvt >>
rect 85 367 115 619
rect 171 367 201 619
rect 325 367 355 619
rect 397 367 427 619
rect 505 367 535 619
rect 613 367 643 619
rect 721 367 751 619
<< ndiff >>
rect 32 202 85 215
rect 32 168 40 202
rect 74 168 85 202
rect 32 93 85 168
rect 32 59 40 93
rect 74 59 85 93
rect 32 47 85 59
rect 115 203 171 215
rect 115 169 126 203
rect 160 169 171 203
rect 115 101 171 169
rect 115 67 126 101
rect 160 67 171 101
rect 115 47 171 67
rect 201 203 311 215
rect 201 169 238 203
rect 272 169 311 203
rect 201 93 311 169
rect 201 59 238 93
rect 272 59 311 93
rect 201 47 311 59
rect 341 192 397 215
rect 341 158 352 192
rect 386 158 397 192
rect 341 101 397 158
rect 341 67 352 101
rect 386 67 397 101
rect 341 47 397 67
rect 427 132 541 215
rect 427 98 466 132
rect 500 98 541 132
rect 427 47 541 98
rect 571 192 627 215
rect 571 158 582 192
rect 616 158 627 192
rect 571 101 627 158
rect 571 67 582 101
rect 616 67 627 101
rect 571 47 627 67
rect 657 169 721 215
rect 657 135 676 169
rect 710 135 721 169
rect 657 47 721 135
rect 751 192 811 215
rect 751 158 765 192
rect 799 158 811 192
rect 751 101 811 158
rect 751 67 765 101
rect 799 67 811 101
rect 751 47 811 67
<< pdiff >>
rect 32 607 85 619
rect 32 573 40 607
rect 74 573 85 607
rect 32 506 85 573
rect 32 472 40 506
rect 74 472 85 506
rect 32 413 85 472
rect 32 379 40 413
rect 74 379 85 413
rect 32 367 85 379
rect 115 599 171 619
rect 115 565 126 599
rect 160 565 171 599
rect 115 504 171 565
rect 115 470 126 504
rect 160 470 171 504
rect 115 420 171 470
rect 115 386 126 420
rect 160 386 171 420
rect 115 367 171 386
rect 201 607 325 619
rect 201 573 212 607
rect 246 573 280 607
rect 314 573 325 607
rect 201 525 325 573
rect 201 491 212 525
rect 246 491 280 525
rect 314 491 325 525
rect 201 439 325 491
rect 201 405 212 439
rect 246 405 280 439
rect 314 405 325 439
rect 201 367 325 405
rect 355 367 397 619
rect 427 367 505 619
rect 535 599 613 619
rect 535 565 556 599
rect 590 565 613 599
rect 535 511 613 565
rect 535 477 556 511
rect 590 477 613 511
rect 535 413 613 477
rect 535 379 556 413
rect 590 379 613 413
rect 535 367 613 379
rect 643 367 721 619
rect 751 607 804 619
rect 751 573 762 607
rect 796 573 804 607
rect 751 524 804 573
rect 751 490 762 524
rect 796 490 804 524
rect 751 450 804 490
rect 751 416 762 450
rect 796 416 804 450
rect 751 367 804 416
<< ndiffc >>
rect 40 168 74 202
rect 40 59 74 93
rect 126 169 160 203
rect 126 67 160 101
rect 238 169 272 203
rect 238 59 272 93
rect 352 158 386 192
rect 352 67 386 101
rect 466 98 500 132
rect 582 158 616 192
rect 582 67 616 101
rect 676 135 710 169
rect 765 158 799 192
rect 765 67 799 101
<< pdiffc >>
rect 40 573 74 607
rect 40 472 74 506
rect 40 379 74 413
rect 126 565 160 599
rect 126 470 160 504
rect 126 386 160 420
rect 212 573 246 607
rect 280 573 314 607
rect 212 491 246 525
rect 280 491 314 525
rect 212 405 246 439
rect 280 405 314 439
rect 556 565 590 599
rect 556 477 590 511
rect 556 379 590 413
rect 762 573 796 607
rect 762 490 796 524
rect 762 416 796 450
<< poly >>
rect 85 619 115 645
rect 171 619 201 645
rect 325 619 355 645
rect 397 619 427 645
rect 505 619 535 645
rect 613 619 643 645
rect 721 619 751 645
rect 85 334 115 367
rect 171 334 201 367
rect 85 318 247 334
rect 85 284 197 318
rect 231 284 247 318
rect 325 303 355 367
rect 85 268 247 284
rect 289 287 355 303
rect 85 215 115 268
rect 171 215 201 268
rect 289 253 305 287
rect 339 253 355 287
rect 289 237 355 253
rect 397 303 427 367
rect 505 303 535 367
rect 613 308 643 367
rect 721 308 751 367
rect 397 287 463 303
rect 397 253 413 287
rect 447 253 463 287
rect 397 237 463 253
rect 505 287 571 303
rect 505 253 521 287
rect 555 253 571 287
rect 505 237 571 253
rect 613 292 679 308
rect 613 258 629 292
rect 663 258 679 292
rect 613 242 679 258
rect 721 292 819 308
rect 721 258 769 292
rect 803 258 819 292
rect 721 242 819 258
rect 311 215 341 237
rect 397 215 427 237
rect 541 215 571 237
rect 627 215 657 242
rect 721 215 751 242
rect 85 21 115 47
rect 171 21 201 47
rect 311 21 341 47
rect 397 21 427 47
rect 541 21 571 47
rect 627 21 657 47
rect 721 21 751 47
<< polycont >>
rect 197 284 231 318
rect 305 253 339 287
rect 413 253 447 287
rect 521 253 555 287
rect 629 258 663 292
rect 769 258 803 292
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 24 607 83 649
rect 24 573 40 607
rect 74 573 83 607
rect 24 506 83 573
rect 24 472 40 506
rect 74 472 83 506
rect 24 413 83 472
rect 24 379 40 413
rect 74 379 83 413
rect 24 363 83 379
rect 117 599 162 615
rect 117 565 126 599
rect 160 565 162 599
rect 117 504 162 565
rect 117 470 126 504
rect 160 470 162 504
rect 117 420 162 470
rect 117 386 126 420
rect 160 386 162 420
rect 196 607 330 649
rect 196 573 212 607
rect 246 573 280 607
rect 314 573 330 607
rect 196 525 330 573
rect 196 491 212 525
rect 246 491 280 525
rect 314 491 330 525
rect 196 439 330 491
rect 196 405 212 439
rect 246 405 280 439
rect 314 405 330 439
rect 540 599 606 615
rect 540 565 556 599
rect 590 565 606 599
rect 540 511 606 565
rect 540 477 556 511
rect 590 477 606 511
rect 540 413 606 477
rect 24 202 83 218
rect 24 168 40 202
rect 74 168 83 202
rect 24 93 83 168
rect 24 59 40 93
rect 74 59 83 93
rect 24 17 83 59
rect 117 203 162 386
rect 540 379 556 413
rect 590 385 606 413
rect 762 607 812 649
rect 796 573 812 607
rect 762 524 812 573
rect 796 490 812 524
rect 762 450 812 490
rect 796 416 812 450
rect 762 400 812 416
rect 590 379 731 385
rect 540 371 731 379
rect 235 342 731 371
rect 235 337 583 342
rect 235 334 269 337
rect 197 318 269 334
rect 231 284 269 318
rect 197 268 269 284
rect 305 287 363 303
rect 339 253 363 287
rect 305 237 363 253
rect 397 287 463 303
rect 397 253 413 287
rect 447 253 463 287
rect 397 242 463 253
rect 497 287 571 303
rect 497 253 521 287
rect 555 253 571 287
rect 497 242 571 253
rect 605 292 663 308
rect 605 258 629 292
rect 605 242 663 258
rect 117 169 126 203
rect 160 169 162 203
rect 117 101 162 169
rect 117 67 126 101
rect 160 67 162 101
rect 117 51 162 67
rect 222 203 288 207
rect 382 203 626 208
rect 222 169 238 203
rect 272 169 288 203
rect 222 93 288 169
rect 222 59 238 93
rect 272 59 288 93
rect 222 17 288 59
rect 336 192 626 203
rect 336 158 352 192
rect 386 174 582 192
rect 386 158 402 174
rect 336 101 402 158
rect 566 158 582 174
rect 616 158 626 192
rect 697 187 731 342
rect 769 292 847 366
rect 803 258 847 292
rect 769 242 847 258
rect 336 67 352 101
rect 386 67 402 101
rect 336 51 402 67
rect 450 132 516 140
rect 450 98 466 132
rect 500 98 516 132
rect 450 17 516 98
rect 566 101 626 158
rect 660 169 731 187
rect 660 135 676 169
rect 710 135 731 169
rect 660 119 731 135
rect 765 192 819 208
rect 799 158 819 192
rect 566 67 582 101
rect 616 85 626 101
rect 765 101 819 158
rect 616 67 765 85
rect 799 67 819 101
rect 566 51 819 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
<< metal1 >>
rect 0 683 864 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 864 683
rect 0 617 864 649
rect 0 17 864 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 864 17
rect 0 -49 864 -17
<< labels >>
flabel pwell s 0 0 864 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 864 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 o32a_2
flabel metal1 s 0 617 864 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 864 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 127 94 161 128 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 168 161 202 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 390 161 424 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 127 538 161 572 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A3
port 3 nsew signal input
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 4 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 B2
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 864 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1740974
string GDS_START 1732668
<< end >>
