magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3218 1975
<< nwell >>
rect -38 331 1958 704
<< pwell >>
rect 1 241 875 263
rect 1 49 1871 241
rect 0 0 1920 49
<< scnmos >>
rect 80 69 110 237
rect 166 69 196 237
rect 268 69 298 237
rect 354 69 384 237
rect 440 69 470 237
rect 558 69 588 237
rect 644 69 674 237
rect 762 69 792 237
rect 1074 47 1104 215
rect 1160 47 1190 215
rect 1246 47 1276 215
rect 1332 47 1362 215
rect 1418 47 1448 215
rect 1504 47 1534 215
rect 1590 47 1620 215
rect 1676 47 1706 215
rect 1762 47 1792 215
<< scpmoshvt >>
rect 96 367 126 619
rect 182 367 212 619
rect 268 367 298 619
rect 354 367 384 619
rect 440 367 470 619
rect 526 367 556 619
rect 612 367 642 619
rect 698 367 728 619
rect 1072 367 1102 619
rect 1158 367 1188 619
rect 1244 367 1274 619
rect 1334 367 1364 619
rect 1420 367 1450 619
rect 1506 367 1536 619
rect 1624 367 1654 619
rect 1710 367 1740 619
rect 1800 367 1830 619
<< ndiff >>
rect 27 225 80 237
rect 27 191 35 225
rect 69 191 80 225
rect 27 115 80 191
rect 27 81 35 115
rect 69 81 80 115
rect 27 69 80 81
rect 110 179 166 237
rect 110 145 121 179
rect 155 145 166 179
rect 110 111 166 145
rect 110 77 121 111
rect 155 77 166 111
rect 110 69 166 77
rect 196 229 268 237
rect 196 195 223 229
rect 257 195 268 229
rect 196 161 268 195
rect 196 127 223 161
rect 257 127 268 161
rect 196 69 268 127
rect 298 143 354 237
rect 298 109 309 143
rect 343 109 354 143
rect 298 69 354 109
rect 384 229 440 237
rect 384 195 395 229
rect 429 195 440 229
rect 384 69 440 195
rect 470 89 558 237
rect 470 69 497 89
rect 485 55 497 69
rect 531 69 558 89
rect 588 229 644 237
rect 588 195 599 229
rect 633 195 644 229
rect 588 69 644 195
rect 674 89 762 237
rect 674 69 701 89
rect 531 55 543 69
rect 485 47 543 55
rect 689 55 701 69
rect 735 69 762 89
rect 792 229 849 237
rect 792 195 803 229
rect 837 195 849 229
rect 792 69 849 195
rect 1021 97 1074 215
rect 735 55 747 69
rect 689 47 747 55
rect 1021 63 1029 97
rect 1063 63 1074 97
rect 1021 47 1074 63
rect 1104 178 1160 215
rect 1104 144 1115 178
rect 1149 144 1160 178
rect 1104 107 1160 144
rect 1104 73 1115 107
rect 1149 73 1160 107
rect 1104 47 1160 73
rect 1190 97 1246 215
rect 1190 63 1201 97
rect 1235 63 1246 97
rect 1190 47 1246 63
rect 1276 178 1332 215
rect 1276 144 1287 178
rect 1321 144 1332 178
rect 1276 101 1332 144
rect 1276 67 1287 101
rect 1321 67 1332 101
rect 1276 47 1332 67
rect 1362 165 1418 215
rect 1362 131 1373 165
rect 1407 131 1418 165
rect 1362 89 1418 131
rect 1362 55 1373 89
rect 1407 55 1418 89
rect 1362 47 1418 55
rect 1448 207 1504 215
rect 1448 173 1459 207
rect 1493 173 1504 207
rect 1448 101 1504 173
rect 1448 67 1459 101
rect 1493 67 1504 101
rect 1448 47 1504 67
rect 1534 157 1590 215
rect 1534 123 1545 157
rect 1579 123 1590 157
rect 1534 89 1590 123
rect 1534 55 1545 89
rect 1579 55 1590 89
rect 1534 47 1590 55
rect 1620 207 1676 215
rect 1620 173 1631 207
rect 1665 173 1676 207
rect 1620 101 1676 173
rect 1620 67 1631 101
rect 1665 67 1676 101
rect 1620 47 1676 67
rect 1706 161 1762 215
rect 1706 127 1717 161
rect 1751 127 1762 161
rect 1706 89 1762 127
rect 1706 55 1717 89
rect 1751 55 1762 89
rect 1706 47 1762 55
rect 1792 203 1845 215
rect 1792 169 1803 203
rect 1837 169 1845 203
rect 1792 101 1845 169
rect 1792 67 1803 101
rect 1837 67 1845 101
rect 1792 47 1845 67
<< pdiff >>
rect 992 630 1050 638
rect 43 572 96 619
rect 43 538 51 572
rect 85 538 96 572
rect 43 504 96 538
rect 43 470 51 504
rect 85 470 96 504
rect 43 436 96 470
rect 43 402 51 436
rect 85 402 96 436
rect 43 367 96 402
rect 126 574 182 619
rect 126 540 137 574
rect 171 540 182 574
rect 126 506 182 540
rect 126 472 137 506
rect 171 472 182 506
rect 126 367 182 472
rect 212 504 268 619
rect 212 470 223 504
rect 257 470 268 504
rect 212 436 268 470
rect 212 402 223 436
rect 257 402 268 436
rect 212 367 268 402
rect 298 574 354 619
rect 298 540 309 574
rect 343 540 354 574
rect 298 506 354 540
rect 298 472 309 506
rect 343 472 354 506
rect 298 367 354 472
rect 384 420 440 619
rect 384 386 395 420
rect 429 386 440 420
rect 384 367 440 386
rect 470 576 526 619
rect 470 542 481 576
rect 515 542 526 576
rect 470 367 526 542
rect 556 420 612 619
rect 556 386 567 420
rect 601 386 612 420
rect 556 367 612 386
rect 642 576 698 619
rect 642 542 653 576
rect 687 542 698 576
rect 642 367 698 542
rect 728 420 781 619
rect 728 386 739 420
rect 773 386 781 420
rect 728 367 781 386
rect 992 596 1004 630
rect 1038 619 1050 630
rect 1038 596 1072 619
rect 992 367 1072 596
rect 1102 451 1158 619
rect 1102 417 1113 451
rect 1147 417 1158 451
rect 1102 367 1158 417
rect 1188 609 1244 619
rect 1188 575 1199 609
rect 1233 575 1244 609
rect 1188 367 1244 575
rect 1274 451 1334 619
rect 1274 417 1285 451
rect 1319 417 1334 451
rect 1274 367 1334 417
rect 1364 606 1420 619
rect 1364 572 1375 606
rect 1409 572 1420 606
rect 1364 367 1420 572
rect 1450 597 1506 619
rect 1450 563 1461 597
rect 1495 563 1506 597
rect 1450 527 1506 563
rect 1450 493 1461 527
rect 1495 493 1506 527
rect 1450 457 1506 493
rect 1450 423 1461 457
rect 1495 423 1506 457
rect 1450 367 1506 423
rect 1536 605 1624 619
rect 1536 571 1563 605
rect 1597 571 1624 605
rect 1536 525 1624 571
rect 1536 491 1563 525
rect 1597 491 1624 525
rect 1536 367 1624 491
rect 1654 609 1710 619
rect 1654 575 1665 609
rect 1699 575 1710 609
rect 1654 541 1710 575
rect 1654 507 1665 541
rect 1699 507 1710 541
rect 1654 473 1710 507
rect 1654 439 1665 473
rect 1699 439 1710 473
rect 1654 367 1710 439
rect 1740 611 1800 619
rect 1740 577 1755 611
rect 1789 577 1800 611
rect 1740 543 1800 577
rect 1740 509 1755 543
rect 1789 509 1800 543
rect 1740 475 1800 509
rect 1740 441 1755 475
rect 1789 441 1800 475
rect 1740 367 1800 441
rect 1830 599 1883 619
rect 1830 565 1841 599
rect 1875 565 1883 599
rect 1830 512 1883 565
rect 1830 478 1841 512
rect 1875 478 1883 512
rect 1830 419 1883 478
rect 1830 385 1841 419
rect 1875 385 1883 419
rect 1830 367 1883 385
<< ndiffc >>
rect 35 191 69 225
rect 35 81 69 115
rect 121 145 155 179
rect 121 77 155 111
rect 223 195 257 229
rect 223 127 257 161
rect 309 109 343 143
rect 395 195 429 229
rect 497 55 531 89
rect 599 195 633 229
rect 701 55 735 89
rect 803 195 837 229
rect 1029 63 1063 97
rect 1115 144 1149 178
rect 1115 73 1149 107
rect 1201 63 1235 97
rect 1287 144 1321 178
rect 1287 67 1321 101
rect 1373 131 1407 165
rect 1373 55 1407 89
rect 1459 173 1493 207
rect 1459 67 1493 101
rect 1545 123 1579 157
rect 1545 55 1579 89
rect 1631 173 1665 207
rect 1631 67 1665 101
rect 1717 127 1751 161
rect 1717 55 1751 89
rect 1803 169 1837 203
rect 1803 67 1837 101
<< pdiffc >>
rect 51 538 85 572
rect 51 470 85 504
rect 51 402 85 436
rect 137 540 171 574
rect 137 472 171 506
rect 223 470 257 504
rect 223 402 257 436
rect 309 540 343 574
rect 309 472 343 506
rect 395 386 429 420
rect 481 542 515 576
rect 567 386 601 420
rect 653 542 687 576
rect 739 386 773 420
rect 1004 596 1038 630
rect 1113 417 1147 451
rect 1199 575 1233 609
rect 1285 417 1319 451
rect 1375 572 1409 606
rect 1461 563 1495 597
rect 1461 493 1495 527
rect 1461 423 1495 457
rect 1563 571 1597 605
rect 1563 491 1597 525
rect 1665 575 1699 609
rect 1665 507 1699 541
rect 1665 439 1699 473
rect 1755 577 1789 611
rect 1755 509 1789 543
rect 1755 441 1789 475
rect 1841 565 1875 599
rect 1841 478 1875 512
rect 1841 385 1875 419
<< poly >>
rect 96 619 126 645
rect 182 619 212 645
rect 268 619 298 645
rect 354 619 384 645
rect 440 619 470 645
rect 526 619 556 645
rect 612 619 642 645
rect 698 619 728 645
rect 1072 619 1102 645
rect 1158 619 1188 645
rect 1244 619 1274 645
rect 1334 619 1364 645
rect 1420 619 1450 645
rect 1506 619 1536 645
rect 1624 619 1654 645
rect 1710 619 1740 645
rect 1800 619 1830 645
rect 96 335 126 367
rect 182 335 212 367
rect 268 335 298 367
rect 354 335 384 367
rect 73 319 384 335
rect 73 285 89 319
rect 123 285 157 319
rect 191 285 225 319
rect 259 285 293 319
rect 327 285 384 319
rect 73 269 384 285
rect 80 237 110 269
rect 166 237 196 269
rect 268 237 298 269
rect 354 237 384 269
rect 440 335 470 367
rect 526 335 556 367
rect 612 335 642 367
rect 698 335 728 367
rect 1072 335 1102 367
rect 1158 335 1188 367
rect 1244 335 1274 367
rect 1334 335 1364 367
rect 440 319 792 335
rect 440 285 501 319
rect 535 285 569 319
rect 603 285 637 319
rect 671 285 705 319
rect 739 285 792 319
rect 1072 319 1364 335
rect 1072 305 1090 319
rect 440 269 792 285
rect 440 237 470 269
rect 558 237 588 269
rect 644 237 674 269
rect 762 237 792 269
rect 1074 285 1090 305
rect 1124 285 1158 319
rect 1192 285 1226 319
rect 1260 285 1294 319
rect 1328 305 1364 319
rect 1420 345 1450 367
rect 1506 345 1536 367
rect 1624 345 1654 367
rect 1710 345 1740 367
rect 1420 319 1740 345
rect 1800 333 1830 367
rect 1328 285 1362 305
rect 1420 299 1461 319
rect 1074 269 1362 285
rect 80 43 110 69
rect 166 43 196 69
rect 268 43 298 69
rect 354 43 384 69
rect 440 43 470 69
rect 558 43 588 69
rect 644 43 674 69
rect 1074 215 1104 269
rect 1160 215 1190 269
rect 1246 215 1276 269
rect 1332 215 1362 269
rect 1418 285 1461 299
rect 1495 285 1529 319
rect 1563 285 1597 319
rect 1631 285 1665 319
rect 1699 315 1740 319
rect 1782 317 1848 333
rect 1699 285 1715 315
rect 1418 269 1715 285
rect 1782 283 1798 317
rect 1832 283 1848 317
rect 1418 215 1448 269
rect 1504 215 1534 269
rect 1590 215 1620 269
rect 1676 215 1706 269
rect 1782 267 1848 283
rect 1762 237 1848 267
rect 1762 215 1792 237
rect 762 43 792 69
rect 1074 21 1104 47
rect 1160 21 1190 47
rect 1246 21 1276 47
rect 1332 21 1362 47
rect 1418 21 1448 47
rect 1504 21 1534 47
rect 1590 21 1620 47
rect 1676 21 1706 47
rect 1762 21 1792 47
<< polycont >>
rect 89 285 123 319
rect 157 285 191 319
rect 225 285 259 319
rect 293 285 327 319
rect 501 285 535 319
rect 569 285 603 319
rect 637 285 671 319
rect 705 285 739 319
rect 1090 285 1124 319
rect 1158 285 1192 319
rect 1226 285 1260 319
rect 1294 285 1328 319
rect 1461 285 1495 319
rect 1529 285 1563 319
rect 1597 285 1631 319
rect 1665 285 1699 319
rect 1798 283 1832 317
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 988 630 1054 649
rect 47 572 85 588
rect 47 538 51 572
rect 47 504 85 538
rect 47 470 51 504
rect 47 436 85 470
rect 133 574 347 590
rect 133 540 137 574
rect 171 556 309 574
rect 171 540 175 556
rect 133 506 175 540
rect 305 540 309 556
rect 343 540 347 574
rect 133 472 137 506
rect 171 472 175 506
rect 133 456 175 472
rect 223 504 257 520
rect 47 402 51 436
rect 223 436 257 470
rect 305 506 347 540
rect 477 576 691 615
rect 988 596 1004 630
rect 1038 596 1054 630
rect 988 594 1054 596
rect 1183 609 1249 649
rect 477 542 481 576
rect 515 542 653 576
rect 687 560 691 576
rect 1183 575 1199 609
rect 1233 575 1249 609
rect 1183 569 1249 575
rect 1359 606 1425 649
rect 1359 572 1375 606
rect 1409 572 1425 606
rect 1359 569 1425 572
rect 1459 597 1513 613
rect 1459 563 1461 597
rect 1495 563 1513 597
rect 687 542 993 560
rect 477 535 993 542
rect 1459 535 1513 563
rect 477 527 1513 535
rect 477 526 1461 527
rect 305 472 309 506
rect 343 492 347 506
rect 959 501 1461 526
rect 1376 493 1461 501
rect 1495 493 1513 527
rect 343 472 923 492
rect 305 467 923 472
rect 305 456 1323 467
rect 85 402 223 420
rect 889 451 1323 456
rect 257 420 853 422
rect 257 402 395 420
rect 47 386 395 402
rect 429 386 567 420
rect 601 386 739 420
rect 773 386 853 420
rect 889 417 1113 451
rect 1147 417 1285 451
rect 1319 417 1323 451
rect 1376 457 1513 493
rect 1547 605 1613 649
rect 1547 571 1563 605
rect 1597 571 1613 605
rect 1547 525 1613 571
rect 1547 491 1563 525
rect 1597 491 1613 525
rect 1647 609 1715 613
rect 1647 575 1665 609
rect 1699 575 1715 609
rect 1647 541 1715 575
rect 1647 507 1665 541
rect 1699 507 1715 541
rect 1647 473 1715 507
rect 1647 457 1665 473
rect 1376 423 1461 457
rect 1495 439 1665 457
rect 1699 439 1715 473
rect 1495 423 1715 439
rect 1749 611 1805 649
rect 1749 577 1755 611
rect 1789 577 1805 611
rect 1749 543 1805 577
rect 1749 509 1755 543
rect 1789 509 1805 543
rect 1749 475 1805 509
rect 1749 441 1755 475
rect 1789 441 1805 475
rect 1749 425 1805 441
rect 1839 599 1902 615
rect 1839 565 1841 599
rect 1875 565 1902 599
rect 1839 512 1902 565
rect 1839 478 1841 512
rect 1875 478 1902 512
rect 889 401 1323 417
rect 1839 419 1902 478
rect 31 319 343 350
rect 31 285 89 319
rect 123 285 157 319
rect 191 285 225 319
rect 259 285 293 319
rect 327 285 343 319
rect 485 319 755 352
rect 379 249 451 294
rect 485 285 501 319
rect 535 285 569 319
rect 603 285 637 319
rect 671 285 705 319
rect 739 285 755 319
rect 485 267 755 285
rect 31 233 451 249
rect 819 233 853 386
rect 1375 367 1805 389
rect 1839 385 1841 419
rect 1875 385 1902 419
rect 1839 369 1902 385
rect 887 355 1805 367
rect 887 319 1409 355
rect 1771 333 1805 355
rect 887 285 1090 319
rect 1124 285 1158 319
rect 1192 285 1226 319
rect 1260 285 1294 319
rect 1328 285 1409 319
rect 887 283 1409 285
rect 1445 319 1735 321
rect 1445 285 1461 319
rect 1495 285 1529 319
rect 1563 285 1597 319
rect 1631 285 1665 319
rect 1699 285 1735 319
rect 1445 283 1735 285
rect 31 229 853 233
rect 31 225 223 229
rect 31 191 35 225
rect 69 215 223 225
rect 31 115 69 191
rect 207 195 223 215
rect 257 195 395 229
rect 429 195 599 229
rect 633 195 803 229
rect 837 195 853 229
rect 207 193 853 195
rect 889 215 1667 249
rect 31 81 35 115
rect 31 65 69 81
rect 105 179 171 181
rect 105 145 121 179
rect 155 145 171 179
rect 105 111 171 145
rect 207 161 273 193
rect 207 127 223 161
rect 257 127 273 161
rect 889 159 923 215
rect 1457 207 1495 215
rect 307 143 923 159
rect 105 77 121 111
rect 155 91 171 111
rect 307 109 309 143
rect 343 125 923 143
rect 959 178 1337 181
rect 959 147 1115 178
rect 343 109 359 125
rect 307 91 359 109
rect 959 91 993 147
rect 1099 144 1115 147
rect 1149 147 1287 178
rect 1149 144 1165 147
rect 155 77 359 91
rect 105 51 359 77
rect 481 89 993 91
rect 481 55 497 89
rect 531 55 701 89
rect 735 55 993 89
rect 481 51 993 55
rect 1027 97 1065 113
rect 1027 63 1029 97
rect 1063 63 1065 97
rect 1099 107 1165 144
rect 1271 144 1287 147
rect 1321 144 1337 178
rect 1099 73 1115 107
rect 1149 73 1165 107
rect 1099 69 1165 73
rect 1199 97 1237 113
rect 1027 17 1065 63
rect 1199 63 1201 97
rect 1235 63 1237 97
rect 1199 17 1237 63
rect 1271 101 1337 144
rect 1271 67 1287 101
rect 1321 67 1337 101
rect 1271 51 1337 67
rect 1371 165 1423 181
rect 1371 131 1373 165
rect 1407 131 1423 165
rect 1371 89 1423 131
rect 1371 55 1373 89
rect 1407 55 1423 89
rect 1371 17 1423 55
rect 1457 173 1459 207
rect 1493 173 1495 207
rect 1457 101 1495 173
rect 1629 207 1667 215
rect 1629 173 1631 207
rect 1665 173 1667 207
rect 1701 233 1735 283
rect 1771 317 1834 333
rect 1771 283 1798 317
rect 1832 283 1834 317
rect 1771 267 1834 283
rect 1868 233 1902 369
rect 1701 203 1902 233
rect 1701 197 1803 203
rect 1457 67 1459 101
rect 1493 67 1495 101
rect 1457 51 1495 67
rect 1529 157 1595 161
rect 1529 123 1545 157
rect 1579 123 1595 157
rect 1529 89 1595 123
rect 1529 55 1545 89
rect 1579 55 1595 89
rect 1529 17 1595 55
rect 1629 101 1667 173
rect 1801 169 1803 197
rect 1837 197 1902 203
rect 1837 169 1841 197
rect 1629 67 1631 101
rect 1665 67 1667 101
rect 1629 51 1667 67
rect 1701 161 1767 163
rect 1701 127 1717 161
rect 1751 127 1767 161
rect 1701 89 1767 127
rect 1701 55 1717 89
rect 1751 55 1767 89
rect 1701 17 1767 55
rect 1801 101 1841 169
rect 1801 67 1803 101
rect 1837 67 1841 101
rect 1801 51 1841 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
<< metal1 >>
rect 0 683 1920 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1920 683
rect 0 617 1920 649
rect 0 17 1920 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1920 17
rect 0 -49 1920 -17
<< labels >>
flabel pwell s 0 0 1920 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 1920 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux2i_4
flabel metal1 s 0 617 1920 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 1920 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 1183 316 1217 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 1279 316 1313 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 S
port 3 nsew signal input
flabel locali s 415 242 449 276 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1920 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3863264
string GDS_START 3849196
<< end >>
