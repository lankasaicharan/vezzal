magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 1970 1975
<< nwell >>
rect -38 331 710 704
<< pwell >>
rect 54 49 638 241
rect 0 0 672 49
<< scnmos >>
rect 133 131 163 215
rect 241 47 271 215
rect 336 47 366 215
rect 443 47 473 215
rect 529 47 559 215
<< scpmoshvt >>
rect 133 367 163 451
rect 241 367 271 619
rect 313 367 343 619
rect 421 367 451 619
rect 529 367 559 619
<< ndiff >>
rect 80 190 133 215
rect 80 156 88 190
rect 122 156 133 190
rect 80 131 133 156
rect 163 182 241 215
rect 163 148 174 182
rect 208 148 241 182
rect 163 131 241 148
rect 188 93 241 131
rect 188 59 196 93
rect 230 59 241 93
rect 188 47 241 59
rect 271 203 336 215
rect 271 169 291 203
rect 325 169 336 203
rect 271 101 336 169
rect 271 67 291 101
rect 325 67 336 101
rect 271 47 336 67
rect 366 165 443 215
rect 366 131 387 165
rect 421 131 443 165
rect 366 93 443 131
rect 366 59 387 93
rect 421 59 443 93
rect 366 47 443 59
rect 473 203 529 215
rect 473 169 484 203
rect 518 169 529 203
rect 473 101 529 169
rect 473 67 484 101
rect 518 67 529 101
rect 473 47 529 67
rect 559 163 612 215
rect 559 129 570 163
rect 604 129 612 163
rect 559 93 612 129
rect 559 59 570 93
rect 604 59 612 93
rect 559 47 612 59
<< pdiff >>
rect 188 607 241 619
rect 188 573 196 607
rect 230 573 241 607
rect 188 502 241 573
rect 188 468 196 502
rect 230 468 241 502
rect 188 451 241 468
rect 80 424 133 451
rect 80 390 88 424
rect 122 390 133 424
rect 80 367 133 390
rect 163 367 241 451
rect 271 367 313 619
rect 343 367 421 619
rect 451 367 529 619
rect 559 599 619 619
rect 559 565 577 599
rect 611 565 619 599
rect 559 506 619 565
rect 559 472 577 506
rect 611 472 619 506
rect 559 419 619 472
rect 559 385 577 419
rect 611 385 619 419
rect 559 367 619 385
<< ndiffc >>
rect 88 156 122 190
rect 174 148 208 182
rect 196 59 230 93
rect 291 169 325 203
rect 291 67 325 101
rect 387 131 421 165
rect 387 59 421 93
rect 484 169 518 203
rect 484 67 518 101
rect 570 129 604 163
rect 570 59 604 93
<< pdiffc >>
rect 196 573 230 607
rect 196 468 230 502
rect 88 390 122 424
rect 577 565 611 599
rect 577 472 611 506
rect 577 385 611 419
<< poly >>
rect 241 619 271 645
rect 313 619 343 645
rect 421 619 451 645
rect 529 619 559 645
rect 133 451 163 477
rect 133 335 163 367
rect 49 319 163 335
rect 49 285 69 319
rect 103 285 163 319
rect 241 303 271 367
rect 49 269 163 285
rect 133 215 163 269
rect 205 287 271 303
rect 205 253 221 287
rect 255 253 271 287
rect 205 237 271 253
rect 313 317 343 367
rect 421 345 451 367
rect 421 319 487 345
rect 313 301 379 317
rect 313 267 329 301
rect 363 267 379 301
rect 421 285 437 319
rect 471 285 487 319
rect 421 269 487 285
rect 529 335 559 367
rect 529 319 595 335
rect 529 285 545 319
rect 579 285 595 319
rect 529 269 595 285
rect 313 237 379 267
rect 241 215 271 237
rect 336 215 366 237
rect 443 215 473 269
rect 529 215 559 269
rect 133 105 163 131
rect 241 21 271 47
rect 336 21 366 47
rect 443 21 473 47
rect 529 21 559 47
<< polycont >>
rect 69 285 103 319
rect 221 253 255 287
rect 329 267 363 301
rect 437 285 471 319
rect 545 285 579 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 180 607 246 649
rect 180 573 196 607
rect 230 573 246 607
rect 180 502 246 573
rect 180 468 196 502
rect 230 468 246 502
rect 180 462 246 468
rect 573 599 655 615
rect 573 565 577 599
rect 611 565 655 599
rect 573 506 655 565
rect 573 472 577 506
rect 611 472 655 506
rect 72 424 539 428
rect 72 390 88 424
rect 122 394 539 424
rect 122 390 187 394
rect 72 386 187 390
rect 17 319 119 352
rect 17 285 69 319
rect 103 285 119 319
rect 153 251 187 386
rect 72 217 187 251
rect 221 287 257 360
rect 255 253 257 287
rect 313 301 379 360
rect 313 267 329 301
rect 363 267 379 301
rect 413 319 471 360
rect 413 285 437 319
rect 413 269 471 285
rect 505 335 539 394
rect 573 419 655 472
rect 573 385 577 419
rect 611 385 655 419
rect 573 369 655 385
rect 505 319 579 335
rect 505 285 545 319
rect 505 269 579 285
rect 221 219 257 253
rect 613 233 655 369
rect 72 190 124 217
rect 72 156 88 190
rect 122 156 124 190
rect 291 203 655 233
rect 72 140 124 156
rect 158 182 248 183
rect 158 148 174 182
rect 208 148 248 182
rect 158 93 248 148
rect 158 59 196 93
rect 230 59 248 93
rect 158 17 248 59
rect 325 199 484 203
rect 325 169 337 199
rect 291 101 337 169
rect 471 169 484 199
rect 518 197 655 203
rect 518 169 520 197
rect 325 67 337 101
rect 291 51 337 67
rect 371 131 387 165
rect 421 131 437 165
rect 371 93 437 131
rect 371 59 387 93
rect 421 59 437 93
rect 371 17 437 59
rect 471 101 520 169
rect 471 67 484 101
rect 518 67 520 101
rect 471 51 520 67
rect 554 129 570 163
rect 604 129 620 163
rect 554 93 620 129
rect 554 59 570 93
rect 604 59 620 93
rect 554 17 620 59
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 683 672 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 672 683
rect 0 617 672 649
rect 0 17 672 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -49 672 -17
<< labels >>
flabel pwell s 0 0 672 49 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 0 617 672 666 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 nor4b_1
flabel metal1 s 0 617 672 666 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 0 672 49 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D_N
port 4 nsew signal input
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 672 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1815216
string GDS_START 1809184
<< end >>
