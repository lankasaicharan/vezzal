magic
tech sky130A
magscale 1 2
timestamp 1627202621
<< checkpaint >>
rect -1298 -1308 3138 1852
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 1 201 1431 203
rect 1 23 1835 201
rect 1 21 207 23
rect 695 21 905 23
rect 1346 21 1835 23
rect 29 -17 63 21
<< scnmos >>
rect 83 47 113 177
rect 196 93 226 177
rect 439 49 469 177
rect 537 49 567 177
rect 799 47 829 177
rect 995 49 1025 177
rect 1156 49 1186 133
rect 1315 49 1345 177
rect 1454 47 1484 167
rect 1565 47 1595 175
rect 1722 47 1752 175
<< scpmoshvt >>
rect 85 297 121 497
rect 198 297 234 425
rect 418 325 454 493
rect 525 297 561 465
rect 747 297 783 497
rect 987 297 1023 465
rect 1148 297 1184 425
rect 1333 329 1369 457
rect 1446 329 1482 497
rect 1557 297 1593 497
rect 1714 297 1750 497
<< ndiff >>
rect 27 129 83 177
rect 27 95 35 129
rect 69 95 83 129
rect 27 47 83 95
rect 113 93 196 177
rect 226 169 321 177
rect 226 135 275 169
rect 309 135 321 169
rect 226 93 321 135
rect 375 165 439 177
rect 375 131 385 165
rect 419 131 439 165
rect 113 89 181 93
rect 113 55 129 89
rect 163 55 181 89
rect 113 47 181 55
rect 375 49 439 131
rect 469 91 537 177
rect 469 57 481 91
rect 515 57 537 91
rect 469 49 537 57
rect 567 91 637 177
rect 567 57 591 91
rect 625 57 637 91
rect 567 49 637 57
rect 721 157 799 177
rect 721 123 735 157
rect 769 123 799 157
rect 721 89 799 123
rect 721 55 735 89
rect 769 55 799 89
rect 721 47 799 55
rect 829 165 881 177
rect 829 131 839 165
rect 873 131 881 165
rect 829 124 881 131
rect 829 47 879 124
rect 935 104 995 177
rect 933 97 995 104
rect 933 63 941 97
rect 975 63 995 97
rect 933 49 995 63
rect 1025 133 1125 177
rect 1211 169 1315 177
rect 1211 135 1257 169
rect 1291 135 1315 169
rect 1211 133 1315 135
rect 1025 126 1156 133
rect 1025 92 1035 126
rect 1069 92 1156 126
rect 1025 49 1156 92
rect 1186 49 1315 133
rect 1345 167 1405 177
rect 1505 167 1565 175
rect 1345 93 1454 167
rect 1345 59 1367 93
rect 1401 59 1454 93
rect 1345 49 1454 59
rect 1372 47 1454 49
rect 1484 142 1565 167
rect 1484 108 1511 142
rect 1545 108 1565 142
rect 1484 47 1565 108
rect 1595 97 1722 175
rect 1595 63 1640 97
rect 1674 63 1722 97
rect 1595 47 1722 63
rect 1752 101 1809 175
rect 1752 67 1762 101
rect 1796 67 1809 101
rect 1752 47 1809 67
<< pdiff >>
rect 27 477 85 497
rect 27 443 39 477
rect 73 443 85 477
rect 27 409 85 443
rect 27 375 39 409
rect 73 375 85 409
rect 27 341 85 375
rect 27 307 39 341
rect 73 307 85 341
rect 27 297 85 307
rect 121 477 181 497
rect 121 443 134 477
rect 168 443 181 477
rect 121 425 181 443
rect 121 297 198 425
rect 234 341 292 425
rect 234 307 246 341
rect 280 307 292 341
rect 351 413 418 493
rect 351 379 372 413
rect 406 379 418 413
rect 351 325 418 379
rect 454 481 508 493
rect 454 447 466 481
rect 500 465 508 481
rect 693 481 747 497
rect 500 447 525 465
rect 454 325 525 447
rect 234 297 292 307
rect 473 297 525 325
rect 561 423 639 465
rect 693 447 701 481
rect 735 447 747 481
rect 693 435 747 447
rect 561 339 640 423
rect 561 305 594 339
rect 628 305 640 339
rect 561 297 640 305
rect 694 297 747 435
rect 783 343 847 497
rect 1386 489 1446 497
rect 783 309 795 343
rect 829 309 847 343
rect 783 297 847 309
rect 901 405 987 465
rect 901 371 909 405
rect 943 371 987 405
rect 901 297 987 371
rect 1023 425 1124 465
rect 1386 457 1398 489
rect 1246 425 1333 457
rect 1023 409 1148 425
rect 1023 375 1075 409
rect 1109 375 1148 409
rect 1023 341 1148 375
rect 1023 307 1075 341
rect 1109 307 1148 341
rect 1023 297 1148 307
rect 1184 421 1333 425
rect 1184 387 1287 421
rect 1321 387 1333 421
rect 1184 329 1333 387
rect 1369 455 1398 457
rect 1432 455 1446 489
rect 1369 329 1446 455
rect 1482 341 1557 497
rect 1482 329 1511 341
rect 1184 297 1281 329
rect 1499 307 1511 329
rect 1545 307 1557 341
rect 1499 297 1557 307
rect 1593 489 1714 497
rect 1593 455 1638 489
rect 1672 455 1714 489
rect 1593 297 1714 455
rect 1750 477 1809 497
rect 1750 443 1763 477
rect 1797 443 1809 477
rect 1750 409 1809 443
rect 1750 375 1763 409
rect 1797 375 1809 409
rect 1750 297 1809 375
<< ndiffc >>
rect 35 95 69 129
rect 275 135 309 169
rect 385 131 419 165
rect 129 55 163 89
rect 481 57 515 91
rect 591 57 625 91
rect 735 123 769 157
rect 735 55 769 89
rect 839 131 873 165
rect 941 63 975 97
rect 1257 135 1291 169
rect 1035 92 1069 126
rect 1367 59 1401 93
rect 1511 108 1545 142
rect 1640 63 1674 97
rect 1762 67 1796 101
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 134 443 168 477
rect 246 307 280 341
rect 372 379 406 413
rect 466 447 500 481
rect 701 447 735 481
rect 594 305 628 339
rect 795 309 829 343
rect 909 371 943 405
rect 1075 375 1109 409
rect 1075 307 1109 341
rect 1287 387 1321 421
rect 1398 455 1432 489
rect 1511 307 1545 341
rect 1638 455 1672 489
rect 1763 443 1797 477
rect 1763 375 1797 409
<< poly >>
rect 85 497 121 523
rect 418 493 454 519
rect 196 451 236 483
rect 198 425 234 451
rect 525 465 561 504
rect 747 497 783 523
rect 418 310 454 325
rect 85 282 121 297
rect 198 282 234 297
rect 83 265 123 282
rect 196 265 236 282
rect 416 271 456 310
rect 985 493 1371 523
rect 1446 497 1482 523
rect 1557 497 1593 523
rect 1714 497 1750 523
rect 985 491 1025 493
rect 987 465 1023 491
rect 1331 483 1371 493
rect 1333 457 1369 483
rect 1148 425 1184 451
rect 1333 314 1369 329
rect 1446 314 1482 329
rect 525 282 561 297
rect 747 282 783 297
rect 987 282 1023 297
rect 1148 282 1184 297
rect 416 265 469 271
rect 523 265 563 282
rect 83 249 154 265
rect 83 215 103 249
rect 137 215 154 249
rect 83 199 154 215
rect 196 249 469 265
rect 196 215 386 249
rect 420 215 469 249
rect 196 199 469 215
rect 511 249 575 265
rect 511 215 521 249
rect 555 215 575 249
rect 745 247 785 282
rect 985 247 1025 282
rect 1146 265 1186 282
rect 1331 265 1371 314
rect 745 217 1025 247
rect 511 199 575 215
rect 83 177 113 199
rect 196 177 226 199
rect 439 177 469 199
rect 537 177 567 199
rect 799 177 829 217
rect 995 177 1025 217
rect 1067 249 1186 265
rect 1067 215 1077 249
rect 1111 215 1186 249
rect 1067 199 1186 215
rect 196 67 226 93
rect 83 21 113 47
rect 439 21 469 49
rect 537 21 567 49
rect 1156 133 1186 199
rect 1315 249 1379 265
rect 1444 255 1484 314
rect 1557 282 1593 297
rect 1714 282 1750 297
rect 1555 265 1595 282
rect 1712 265 1752 282
rect 1315 215 1325 249
rect 1359 215 1379 249
rect 1315 199 1379 215
rect 1421 239 1484 255
rect 1421 205 1431 239
rect 1465 205 1484 239
rect 1315 177 1345 199
rect 1421 189 1484 205
rect 1527 249 1595 265
rect 1527 215 1537 249
rect 1571 215 1595 249
rect 1527 199 1595 215
rect 1700 249 1764 265
rect 1700 215 1710 249
rect 1744 215 1764 249
rect 1700 199 1764 215
rect 1454 167 1484 189
rect 1565 175 1595 199
rect 1722 175 1752 199
rect 799 21 829 47
rect 995 21 1025 49
rect 1156 23 1186 49
rect 1315 21 1345 49
rect 1454 21 1484 47
rect 1565 21 1595 47
rect 1722 21 1752 47
<< polycont >>
rect 103 215 137 249
rect 386 215 420 249
rect 521 215 555 249
rect 1077 215 1111 249
rect 1325 215 1359 249
rect 1431 205 1465 239
rect 1537 215 1571 249
rect 1710 215 1744 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 17 477 73 493
rect 17 443 39 477
rect 107 477 184 527
rect 685 481 751 527
rect 1583 489 1719 527
rect 107 443 134 477
rect 168 443 184 477
rect 220 447 466 481
rect 500 447 534 481
rect 685 447 701 481
rect 735 447 751 481
rect 838 455 1398 489
rect 1432 455 1497 489
rect 1583 455 1638 489
rect 1672 455 1719 489
rect 1763 477 1822 493
rect 17 409 73 443
rect 220 409 264 447
rect 838 413 872 455
rect 17 375 39 409
rect 17 341 73 375
rect 17 307 39 341
rect 17 288 73 307
rect 107 375 264 409
rect 332 379 372 413
rect 406 379 872 413
rect 909 405 943 421
rect 17 129 69 288
rect 107 266 151 375
rect 197 307 246 341
rect 280 307 534 341
rect 103 249 151 266
rect 137 215 151 249
rect 103 173 151 215
rect 103 139 241 173
rect 17 95 35 129
rect 17 70 69 95
rect 103 89 163 105
rect 103 55 129 89
rect 103 17 163 55
rect 197 85 241 139
rect 275 169 309 307
rect 500 265 534 307
rect 578 305 594 339
rect 628 323 655 339
rect 599 289 621 305
rect 599 275 655 289
rect 343 249 466 265
rect 343 215 386 249
rect 420 215 466 249
rect 500 249 565 265
rect 500 215 521 249
rect 555 215 565 249
rect 500 199 565 215
rect 275 119 309 135
rect 369 165 445 181
rect 369 131 385 165
rect 419 159 445 165
rect 599 159 633 275
rect 689 241 723 379
rect 769 309 795 343
rect 829 309 873 343
rect 769 289 873 309
rect 419 131 633 159
rect 369 125 633 131
rect 667 207 723 241
rect 667 91 701 207
rect 815 187 873 289
rect 434 85 481 91
rect 197 57 481 85
rect 515 57 531 91
rect 575 57 591 91
rect 625 57 701 91
rect 735 157 769 173
rect 735 89 769 123
rect 197 51 531 57
rect 849 165 873 187
rect 815 131 839 153
rect 815 83 873 131
rect 909 119 943 371
rect 977 178 1011 455
rect 1797 443 1822 477
rect 1763 421 1822 443
rect 1057 375 1075 409
rect 1109 375 1140 409
rect 1057 341 1140 375
rect 1057 307 1075 341
rect 1109 323 1140 341
rect 1257 387 1287 421
rect 1321 409 1822 421
rect 1321 387 1763 409
rect 1109 307 1111 323
rect 1057 289 1111 307
rect 1145 289 1223 323
rect 1060 249 1145 254
rect 1060 215 1077 249
rect 1111 215 1145 249
rect 1060 199 1145 215
rect 1103 187 1145 199
rect 977 165 1029 178
rect 977 144 1069 165
rect 985 131 1069 144
rect 1035 126 1069 131
rect 1103 153 1111 187
rect 1103 126 1145 153
rect 909 85 917 119
rect 735 17 769 55
rect 909 63 941 85
rect 975 63 991 97
rect 1035 64 1069 92
rect 1189 85 1223 289
rect 1257 169 1291 387
rect 1715 375 1763 387
rect 1797 375 1822 409
rect 1325 289 1451 323
rect 1495 307 1511 341
rect 1545 307 1732 341
rect 1495 299 1732 307
rect 1325 249 1369 289
rect 1698 265 1732 299
rect 1359 215 1369 249
rect 1325 199 1369 215
rect 1403 239 1465 255
rect 1403 205 1431 239
rect 1499 249 1643 265
rect 1499 215 1537 249
rect 1571 215 1643 249
rect 1698 249 1754 265
rect 1698 215 1710 249
rect 1744 215 1754 249
rect 1403 189 1465 205
rect 1698 199 1754 215
rect 1403 187 1444 189
rect 1403 153 1407 187
rect 1441 153 1444 187
rect 1698 181 1732 199
rect 1403 146 1444 153
rect 1511 150 1732 181
rect 1503 147 1732 150
rect 1257 119 1291 135
rect 1503 142 1561 147
rect 1503 119 1511 142
rect 1325 85 1367 93
rect 909 53 991 63
rect 1189 59 1367 85
rect 1401 59 1428 93
rect 1503 85 1509 119
rect 1545 108 1561 142
rect 1788 117 1822 375
rect 1543 85 1561 108
rect 1503 59 1561 85
rect 1610 97 1702 113
rect 1610 63 1640 97
rect 1674 63 1702 97
rect 1189 51 1428 59
rect 1610 17 1702 63
rect 1762 101 1822 117
rect 1796 67 1822 101
rect 1762 51 1822 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 621 305 628 323
rect 628 305 655 323
rect 621 289 655 305
rect 815 165 849 187
rect 815 153 839 165
rect 839 153 849 165
rect 1111 289 1145 323
rect 1111 153 1145 187
rect 917 97 951 119
rect 917 85 941 97
rect 941 85 951 97
rect 1407 153 1441 187
rect 1509 108 1511 119
rect 1511 108 1543 119
rect 1509 85 1543 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 609 323 667 329
rect 609 289 621 323
rect 655 320 667 323
rect 1099 323 1157 329
rect 1099 320 1111 323
rect 655 292 1111 320
rect 655 289 667 292
rect 609 283 667 289
rect 1099 289 1111 292
rect 1145 289 1157 323
rect 1099 283 1157 289
rect 803 187 861 193
rect 803 153 815 187
rect 849 184 861 187
rect 1099 187 1157 193
rect 1099 184 1111 187
rect 849 156 1111 184
rect 849 153 861 156
rect 803 147 861 153
rect 1099 153 1111 156
rect 1145 184 1157 187
rect 1395 187 1453 193
rect 1395 184 1407 187
rect 1145 156 1407 184
rect 1145 153 1157 156
rect 1099 147 1157 153
rect 1395 153 1407 156
rect 1441 153 1453 187
rect 1395 147 1453 153
rect 905 119 963 125
rect 905 85 917 119
rect 951 116 963 119
rect 1497 119 1555 125
rect 1497 116 1509 119
rect 951 88 1509 116
rect 951 85 963 88
rect 905 79 963 85
rect 1497 85 1509 88
rect 1543 85 1555 119
rect 1497 79 1555 85
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel locali s 29 357 63 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1325 289 1451 323 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1592 221 1626 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 xnor3_1
rlabel locali s 1325 199 1369 289 1 B
port 2 nsew signal input
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hdll/gds/sky130_fd_sc_hdll.gds
string LEFsymmetry X Y R90
string GDS_END 1275986
string GDS_START 1263724
string LEFproperties maskLayoutSubType "abstract" prCellType "standard" originalViewName "layout"
<< end >>
