magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4850 1975
<< nwell >>
rect -38 331 3590 704
<< pwell >>
rect 1828 273 1937 281
rect 9 160 707 229
rect 1183 214 1395 235
rect 1828 224 2853 273
rect 3062 224 3551 251
rect 1828 214 3551 224
rect 1183 176 3551 214
rect 969 160 3551 176
rect 9 49 3551 160
rect 0 0 3552 49
<< scnmos >>
rect 92 119 122 203
rect 170 119 200 203
rect 284 119 314 203
rect 412 119 442 203
rect 578 119 608 203
rect 808 50 838 134
rect 1054 66 1084 150
rect 1266 125 1296 209
rect 1409 104 1439 188
rect 1523 104 1553 188
rect 1722 60 1752 188
rect 1809 60 1839 188
rect 1926 66 1956 194
rect 2168 119 2198 247
rect 2269 119 2299 247
rect 2371 163 2401 247
rect 2449 163 2479 247
rect 2606 119 2636 247
rect 2724 119 2754 247
rect 2842 70 2872 198
rect 3043 57 3073 141
rect 3145 57 3175 225
rect 3343 57 3373 141
rect 3438 57 3468 225
<< scpmoshvt >>
rect 84 474 114 602
rect 170 474 200 602
rect 242 474 272 602
rect 328 474 358 602
rect 578 411 608 539
rect 858 411 888 539
rect 1054 367 1084 495
rect 1265 379 1295 463
rect 1367 379 1397 463
rect 1445 379 1475 463
rect 1737 379 1767 547
rect 1966 379 1996 547
rect 2044 379 2074 547
rect 2168 379 2198 547
rect 2269 428 2299 596
rect 2371 506 2401 590
rect 2534 506 2564 590
rect 2682 451 2712 619
rect 2768 451 2798 619
rect 2840 451 2870 619
rect 3037 367 3067 495
rect 3139 367 3169 619
rect 3336 367 3366 495
rect 3438 367 3468 619
<< ndiff >>
rect 35 178 92 203
rect 35 144 47 178
rect 81 144 92 178
rect 35 119 92 144
rect 122 119 170 203
rect 200 178 284 203
rect 200 144 212 178
rect 246 144 284 178
rect 200 119 284 144
rect 314 119 412 203
rect 442 174 578 203
rect 442 140 486 174
rect 520 140 578 174
rect 442 119 578 140
rect 608 178 681 203
rect 608 144 635 178
rect 669 144 681 178
rect 608 119 681 144
rect 1209 184 1266 209
rect 1209 150 1221 184
rect 1255 150 1266 184
rect 735 109 808 134
rect 735 75 747 109
rect 781 75 808 109
rect 735 50 808 75
rect 838 112 895 134
rect 838 78 849 112
rect 883 78 895 112
rect 838 50 895 78
rect 995 125 1054 150
rect 995 91 1007 125
rect 1041 91 1054 125
rect 995 66 1054 91
rect 1084 125 1155 150
rect 1209 125 1266 150
rect 1296 188 1369 209
rect 1854 243 1911 255
rect 1854 209 1865 243
rect 1899 209 1911 243
rect 1854 194 1911 209
rect 1854 188 1926 194
rect 1296 173 1409 188
rect 1296 139 1323 173
rect 1357 139 1409 173
rect 1296 125 1409 139
rect 1084 91 1109 125
rect 1143 91 1155 125
rect 1311 104 1409 125
rect 1439 104 1523 188
rect 1553 104 1722 188
rect 1084 66 1155 91
rect 1579 89 1722 104
rect 1579 55 1591 89
rect 1625 60 1722 89
rect 1752 160 1809 188
rect 1752 126 1763 160
rect 1797 126 1809 160
rect 1752 60 1809 126
rect 1839 66 1926 188
rect 1956 158 2013 194
rect 1956 124 1967 158
rect 2001 124 2013 158
rect 1956 66 2013 124
rect 2111 165 2168 247
rect 2111 131 2123 165
rect 2157 131 2168 165
rect 2111 119 2168 131
rect 2198 119 2269 247
rect 2299 191 2371 247
rect 2299 157 2310 191
rect 2344 163 2371 191
rect 2401 163 2449 247
rect 2479 163 2606 247
rect 2344 157 2356 163
rect 2299 119 2356 157
rect 2533 119 2606 163
rect 2636 119 2724 247
rect 2754 204 2827 247
rect 2754 170 2781 204
rect 2815 198 2827 204
rect 2815 170 2842 198
rect 2754 119 2842 170
rect 2533 114 2591 119
rect 2533 80 2545 114
rect 2579 80 2591 114
rect 2651 114 2709 119
rect 2533 68 2591 80
rect 2651 80 2663 114
rect 2697 80 2709 114
rect 2651 68 2709 80
rect 2769 70 2842 119
rect 2872 131 2929 198
rect 3088 213 3145 225
rect 3088 179 3100 213
rect 3134 179 3145 213
rect 3088 141 3145 179
rect 2872 97 2883 131
rect 2917 97 2929 131
rect 2872 70 2929 97
rect 2986 116 3043 141
rect 2986 82 2998 116
rect 3032 82 3043 116
rect 1839 60 1889 66
rect 1625 55 1637 60
rect 1579 43 1637 55
rect 2986 57 3043 82
rect 3073 103 3145 141
rect 3073 69 3100 103
rect 3134 69 3145 103
rect 3073 57 3145 69
rect 3175 213 3232 225
rect 3175 179 3186 213
rect 3220 179 3232 213
rect 3175 103 3232 179
rect 3388 141 3438 225
rect 3175 69 3186 103
rect 3220 69 3232 103
rect 3175 57 3232 69
rect 3286 116 3343 141
rect 3286 82 3298 116
rect 3332 82 3343 116
rect 3286 57 3343 82
rect 3373 116 3438 141
rect 3373 82 3384 116
rect 3418 82 3438 116
rect 3373 57 3438 82
rect 3468 209 3525 225
rect 3468 175 3479 209
rect 3513 175 3525 209
rect 3468 103 3525 175
rect 3468 69 3479 103
rect 3513 69 3525 103
rect 3468 57 3525 69
<< pdiff >>
rect 27 590 84 602
rect 27 556 39 590
rect 73 556 84 590
rect 27 520 84 556
rect 27 486 39 520
rect 73 486 84 520
rect 27 474 84 486
rect 114 561 170 602
rect 114 527 125 561
rect 159 527 170 561
rect 114 474 170 527
rect 200 474 242 602
rect 272 523 328 602
rect 272 489 283 523
rect 317 489 328 523
rect 272 474 328 489
rect 358 590 414 602
rect 358 556 369 590
rect 403 556 414 590
rect 358 520 414 556
rect 358 486 369 520
rect 403 486 414 520
rect 358 474 414 486
rect 468 527 578 539
rect 468 493 479 527
rect 513 493 578 527
rect 468 457 578 493
rect 468 423 479 457
rect 513 423 578 457
rect 468 411 578 423
rect 608 527 665 539
rect 608 493 619 527
rect 653 493 665 527
rect 608 457 665 493
rect 608 423 619 457
rect 653 423 665 457
rect 608 411 665 423
rect 747 495 858 539
rect 747 461 759 495
rect 793 461 858 495
rect 747 411 858 461
rect 888 527 944 539
rect 888 493 899 527
rect 933 493 944 527
rect 1099 585 1155 597
rect 1099 551 1110 585
rect 1144 551 1155 585
rect 1099 495 1155 551
rect 888 457 944 493
rect 888 423 899 457
rect 933 423 944 457
rect 888 411 944 423
rect 998 413 1054 495
rect 998 379 1009 413
rect 1043 379 1054 413
rect 998 367 1054 379
rect 1084 367 1155 495
rect 2219 547 2269 596
rect 1664 521 1737 547
rect 1664 487 1676 521
rect 1710 487 1737 521
rect 1664 463 1737 487
rect 1209 438 1265 463
rect 1209 404 1220 438
rect 1254 404 1265 438
rect 1209 379 1265 404
rect 1295 438 1367 463
rect 1295 404 1322 438
rect 1356 404 1367 438
rect 1295 379 1367 404
rect 1397 379 1445 463
rect 1475 379 1737 463
rect 1767 535 1966 547
rect 1767 501 1921 535
rect 1955 501 1966 535
rect 1767 433 1966 501
rect 1767 399 1921 433
rect 1955 399 1966 433
rect 1767 379 1966 399
rect 1996 379 2044 547
rect 2074 535 2168 547
rect 2074 501 2085 535
rect 2119 501 2168 535
rect 2074 431 2168 501
rect 2074 397 2085 431
rect 2119 397 2168 431
rect 2074 379 2168 397
rect 2198 428 2269 547
rect 2299 590 2349 596
rect 2626 590 2682 619
rect 2299 506 2371 590
rect 2401 506 2534 590
rect 2564 575 2682 590
rect 2564 541 2637 575
rect 2671 541 2682 575
rect 2564 506 2682 541
rect 2299 500 2356 506
rect 2299 466 2310 500
rect 2344 466 2356 500
rect 2299 428 2356 466
rect 2198 379 2248 428
rect 2626 451 2682 506
rect 2712 597 2768 619
rect 2712 563 2723 597
rect 2757 563 2768 597
rect 2712 497 2768 563
rect 2712 463 2723 497
rect 2757 463 2768 497
rect 2712 451 2768 463
rect 2798 451 2840 619
rect 2870 602 2927 619
rect 2870 568 2881 602
rect 2915 568 2927 602
rect 2870 451 2927 568
rect 3082 602 3139 619
rect 3082 568 3094 602
rect 3128 568 3139 602
rect 3082 495 3139 568
rect 2981 442 3037 495
rect 2981 408 2992 442
rect 3026 408 3037 442
rect 2981 367 3037 408
rect 3067 367 3139 495
rect 3169 597 3225 619
rect 3169 563 3180 597
rect 3214 563 3225 597
rect 3169 507 3225 563
rect 3381 607 3438 619
rect 3381 573 3393 607
rect 3427 573 3438 607
rect 3169 473 3180 507
rect 3214 473 3225 507
rect 3381 510 3438 573
rect 3381 495 3393 510
rect 3169 417 3225 473
rect 3169 383 3180 417
rect 3214 383 3225 417
rect 3169 367 3225 383
rect 3279 483 3336 495
rect 3279 449 3291 483
rect 3325 449 3336 483
rect 3279 413 3336 449
rect 3279 379 3291 413
rect 3325 379 3336 413
rect 3279 367 3336 379
rect 3366 476 3393 495
rect 3427 476 3438 510
rect 3366 413 3438 476
rect 3366 379 3393 413
rect 3427 379 3438 413
rect 3366 367 3438 379
rect 3468 597 3525 619
rect 3468 563 3479 597
rect 3513 563 3525 597
rect 3468 505 3525 563
rect 3468 471 3479 505
rect 3513 471 3525 505
rect 3468 413 3525 471
rect 3468 379 3479 413
rect 3513 379 3525 413
rect 3468 367 3525 379
<< ndiffc >>
rect 47 144 81 178
rect 212 144 246 178
rect 486 140 520 174
rect 635 144 669 178
rect 1221 150 1255 184
rect 747 75 781 109
rect 849 78 883 112
rect 1007 91 1041 125
rect 1865 209 1899 243
rect 1323 139 1357 173
rect 1109 91 1143 125
rect 1591 55 1625 89
rect 1763 126 1797 160
rect 1967 124 2001 158
rect 2123 131 2157 165
rect 2310 157 2344 191
rect 2781 170 2815 204
rect 2545 80 2579 114
rect 2663 80 2697 114
rect 3100 179 3134 213
rect 2883 97 2917 131
rect 2998 82 3032 116
rect 3100 69 3134 103
rect 3186 179 3220 213
rect 3186 69 3220 103
rect 3298 82 3332 116
rect 3384 82 3418 116
rect 3479 175 3513 209
rect 3479 69 3513 103
<< pdiffc >>
rect 39 556 73 590
rect 39 486 73 520
rect 125 527 159 561
rect 283 489 317 523
rect 369 556 403 590
rect 369 486 403 520
rect 479 493 513 527
rect 479 423 513 457
rect 619 493 653 527
rect 619 423 653 457
rect 759 461 793 495
rect 899 493 933 527
rect 1110 551 1144 585
rect 899 423 933 457
rect 1009 379 1043 413
rect 1676 487 1710 521
rect 1220 404 1254 438
rect 1322 404 1356 438
rect 1921 501 1955 535
rect 1921 399 1955 433
rect 2085 501 2119 535
rect 2085 397 2119 431
rect 2637 541 2671 575
rect 2310 466 2344 500
rect 2723 563 2757 597
rect 2723 463 2757 497
rect 2881 568 2915 602
rect 3094 568 3128 602
rect 2992 408 3026 442
rect 3180 563 3214 597
rect 3393 573 3427 607
rect 3180 473 3214 507
rect 3180 383 3214 417
rect 3291 449 3325 483
rect 3291 379 3325 413
rect 3393 476 3427 510
rect 3393 379 3427 413
rect 3479 563 3513 597
rect 3479 471 3513 505
rect 3479 379 3513 413
<< poly >>
rect 84 602 114 628
rect 170 602 200 628
rect 242 602 272 628
rect 328 602 358 628
rect 1054 612 1295 642
rect 578 539 608 565
rect 858 539 888 565
rect 84 377 114 474
rect 44 361 122 377
rect 44 327 60 361
rect 94 327 122 361
rect 44 293 122 327
rect 44 259 60 293
rect 94 259 122 293
rect 44 243 122 259
rect 92 203 122 243
rect 170 309 200 474
rect 242 387 272 474
rect 328 459 358 474
rect 328 429 442 459
rect 242 357 364 387
rect 284 348 364 357
rect 284 314 314 348
rect 348 314 364 348
rect 170 293 236 309
rect 170 259 186 293
rect 220 259 236 293
rect 170 243 236 259
rect 284 280 364 314
rect 284 246 314 280
rect 348 246 364 280
rect 170 203 200 243
rect 284 230 364 246
rect 412 301 442 429
rect 1054 495 1084 612
rect 412 285 536 301
rect 412 251 486 285
rect 520 251 536 285
rect 412 235 536 251
rect 284 203 314 230
rect 412 203 442 235
rect 578 203 608 411
rect 858 386 888 411
rect 808 356 888 386
rect 1265 463 1295 612
rect 1367 615 2299 645
rect 2682 619 2712 645
rect 2768 619 2798 645
rect 2840 619 2870 645
rect 3139 619 3169 645
rect 3438 619 3468 645
rect 1367 463 1397 615
rect 2269 596 2299 615
rect 1737 547 1767 573
rect 1966 547 1996 573
rect 2044 547 2074 573
rect 2168 547 2198 573
rect 1445 463 1475 489
rect 2371 590 2401 616
rect 2534 590 2564 616
rect 2371 491 2401 506
rect 2371 461 2486 491
rect 2420 458 2486 461
rect 2534 458 2564 506
rect 2269 413 2299 428
rect 2420 424 2436 458
rect 2470 424 2486 458
rect 2269 383 2378 413
rect 808 308 838 356
rect 1054 308 1084 367
rect 1265 353 1295 379
rect 1367 354 1397 379
rect 772 292 838 308
rect 772 258 788 292
rect 822 258 838 292
rect 772 224 838 258
rect 772 190 788 224
rect 822 190 838 224
rect 772 174 838 190
rect 886 292 1084 308
rect 886 258 902 292
rect 936 258 1084 292
rect 1134 319 1200 335
rect 1134 285 1150 319
rect 1184 299 1200 319
rect 1337 324 1397 354
rect 1445 354 1475 379
rect 1445 331 1621 354
rect 1445 324 1571 331
rect 1337 299 1367 324
rect 1184 285 1367 299
rect 1134 269 1367 285
rect 1523 297 1571 324
rect 1605 297 1621 331
rect 1523 281 1621 297
rect 1737 282 1767 379
rect 1966 347 1996 379
rect 1835 331 1996 347
rect 1835 311 1851 331
rect 886 224 1084 258
rect 886 190 902 224
rect 936 190 1084 224
rect 1266 209 1296 269
rect 1409 260 1475 276
rect 1409 226 1425 260
rect 1459 226 1475 260
rect 1409 210 1475 226
rect 886 174 1084 190
rect 808 134 838 174
rect 1054 150 1084 174
rect 92 93 122 119
rect 170 51 200 119
rect 284 93 314 119
rect 412 93 442 119
rect 578 51 608 119
rect 170 21 608 51
rect 1409 188 1439 210
rect 1523 188 1553 281
rect 1701 266 1767 282
rect 1701 232 1717 266
rect 1751 232 1767 266
rect 1701 216 1767 232
rect 1809 297 1851 311
rect 1885 317 1996 331
rect 1885 297 1901 317
rect 1809 281 1901 297
rect 1722 188 1752 216
rect 1809 188 1839 281
rect 2044 239 2074 379
rect 2168 345 2198 379
rect 2122 329 2198 345
rect 2122 295 2138 329
rect 2172 295 2198 329
rect 2122 279 2198 295
rect 2168 247 2198 279
rect 2240 319 2306 335
rect 2240 285 2256 319
rect 2290 285 2306 319
rect 2240 269 2306 285
rect 2348 292 2378 383
rect 2420 390 2486 424
rect 2420 356 2436 390
rect 2470 356 2486 390
rect 2420 340 2486 356
rect 2528 442 2594 458
rect 3037 495 3067 521
rect 2528 408 2544 442
rect 2578 408 2594 442
rect 2682 425 2712 451
rect 2528 392 2594 408
rect 2636 395 2712 425
rect 2528 292 2558 392
rect 2636 335 2666 395
rect 2768 353 2798 451
rect 2269 247 2299 269
rect 2348 262 2401 292
rect 2371 247 2401 262
rect 2449 262 2558 292
rect 2600 319 2666 335
rect 2600 285 2616 319
rect 2650 285 2666 319
rect 2708 337 2798 353
rect 2708 303 2724 337
rect 2758 323 2798 337
rect 2840 354 2870 451
rect 3336 495 3366 521
rect 2840 338 2946 354
rect 2840 324 2896 338
rect 2758 303 2774 323
rect 2708 287 2774 303
rect 2880 304 2896 324
rect 2930 304 2946 338
rect 3037 335 3067 367
rect 2600 269 2666 285
rect 2449 247 2479 262
rect 2606 247 2636 269
rect 2724 247 2754 287
rect 2880 270 2946 304
rect 2880 250 2896 270
rect 1926 209 2074 239
rect 1926 194 1956 209
rect 1266 99 1296 125
rect 1054 51 1084 66
rect 1409 51 1439 104
rect 1523 78 1553 104
rect 808 24 838 50
rect 1054 21 1439 51
rect 2371 137 2401 163
rect 2449 137 2479 163
rect 2842 236 2896 250
rect 2930 236 2946 270
rect 3007 319 3073 335
rect 3139 331 3169 367
rect 3007 285 3023 319
rect 3057 285 3073 319
rect 3007 269 3073 285
rect 2842 220 2946 236
rect 2842 198 2872 220
rect 2168 93 2198 119
rect 2269 93 2299 119
rect 2606 93 2636 119
rect 2724 93 2754 119
rect 3043 141 3073 269
rect 3115 315 3181 331
rect 3115 281 3131 315
rect 3165 295 3181 315
rect 3336 295 3366 367
rect 3438 327 3468 367
rect 3165 281 3366 295
rect 3115 265 3366 281
rect 3145 225 3175 265
rect 1722 34 1752 60
rect 1809 34 1839 60
rect 1926 51 1956 66
rect 2842 51 2872 70
rect 3336 186 3366 265
rect 3408 311 3474 327
rect 3408 277 3424 311
rect 3458 277 3474 311
rect 3408 261 3474 277
rect 3438 225 3468 261
rect 3336 156 3373 186
rect 3343 141 3373 156
rect 1926 21 2872 51
rect 3043 31 3073 57
rect 3145 31 3175 57
rect 3343 31 3373 57
rect 3438 31 3468 57
<< polycont >>
rect 60 327 94 361
rect 60 259 94 293
rect 314 314 348 348
rect 186 259 220 293
rect 314 246 348 280
rect 486 251 520 285
rect 2436 424 2470 458
rect 788 258 822 292
rect 788 190 822 224
rect 902 258 936 292
rect 1150 285 1184 319
rect 1571 297 1605 331
rect 902 190 936 224
rect 1425 226 1459 260
rect 1717 232 1751 266
rect 1851 297 1885 331
rect 2138 295 2172 329
rect 2256 285 2290 319
rect 2436 356 2470 390
rect 2544 408 2578 442
rect 2616 285 2650 319
rect 2724 303 2758 337
rect 2896 304 2930 338
rect 2896 236 2930 270
rect 3023 285 3057 319
rect 3131 281 3165 315
rect 3424 277 3458 311
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3552 683
rect 23 590 73 606
rect 23 556 39 590
rect 23 520 73 556
rect 23 486 39 520
rect 23 447 73 486
rect 109 561 159 649
rect 109 527 125 561
rect 109 483 159 527
rect 195 590 419 613
rect 195 579 369 590
rect 195 447 229 579
rect 353 556 369 579
rect 403 556 419 590
rect 23 413 229 447
rect 267 523 317 543
rect 267 489 283 523
rect 267 434 317 489
rect 353 520 419 556
rect 353 486 369 520
rect 403 486 419 520
rect 353 470 419 486
rect 479 527 513 649
rect 479 457 513 493
rect 267 400 434 434
rect 479 407 513 423
rect 549 579 723 613
rect 25 361 110 377
rect 400 371 434 400
rect 549 371 583 579
rect 25 327 60 361
rect 94 327 110 361
rect 25 293 110 327
rect 25 259 60 293
rect 94 259 110 293
rect 25 243 110 259
rect 170 293 262 356
rect 170 259 186 293
rect 220 259 262 293
rect 170 243 262 259
rect 298 348 364 364
rect 298 314 314 348
rect 348 314 364 348
rect 298 280 364 314
rect 298 246 314 280
rect 348 246 364 280
rect 31 178 97 207
rect 31 144 47 178
rect 81 144 97 178
rect 31 17 97 144
rect 196 178 262 207
rect 196 144 212 178
rect 246 144 262 178
rect 298 162 364 246
rect 400 337 583 371
rect 619 527 653 543
rect 619 457 653 493
rect 196 126 262 144
rect 400 126 434 337
rect 619 301 653 423
rect 689 378 723 579
rect 759 495 793 649
rect 759 414 793 461
rect 829 579 1058 613
rect 829 378 863 579
rect 689 344 863 378
rect 899 527 952 543
rect 933 493 952 527
rect 899 457 952 493
rect 1024 499 1058 579
rect 1094 585 1160 649
rect 1094 551 1110 585
rect 1144 551 1160 585
rect 1094 535 1160 551
rect 1660 521 1726 649
rect 1024 465 1270 499
rect 1660 487 1676 521
rect 1710 487 1726 521
rect 933 423 952 457
rect 1204 438 1270 465
rect 899 308 952 423
rect 470 285 653 301
rect 470 251 486 285
rect 520 251 653 285
rect 470 235 653 251
rect 619 207 653 235
rect 772 292 839 308
rect 772 258 788 292
rect 822 258 839 292
rect 772 224 839 258
rect 196 92 434 126
rect 470 174 536 199
rect 470 140 486 174
rect 520 140 536 174
rect 470 17 536 140
rect 619 178 685 207
rect 619 144 635 178
rect 669 144 685 178
rect 772 190 788 224
rect 822 190 839 224
rect 772 174 839 190
rect 875 292 952 308
rect 875 258 902 292
rect 936 258 952 292
rect 875 224 952 258
rect 875 190 902 224
rect 936 190 952 224
rect 875 174 952 190
rect 991 413 1059 429
rect 991 379 1009 413
rect 1043 379 1059 413
rect 991 335 1059 379
rect 1204 404 1220 438
rect 1254 404 1270 438
rect 1204 375 1270 404
rect 1306 438 1373 467
rect 1660 458 1726 487
rect 1905 535 1971 551
rect 1905 501 1921 535
rect 1955 501 1971 535
rect 1306 404 1322 438
rect 1356 409 1373 438
rect 1905 433 1971 501
rect 1905 422 1921 433
rect 1356 404 1532 409
rect 1306 375 1532 404
rect 991 319 1200 335
rect 991 285 1150 319
rect 1184 285 1200 319
rect 991 269 1200 285
rect 619 115 685 144
rect 875 138 909 174
rect 731 109 797 138
rect 731 75 747 109
rect 781 75 797 109
rect 731 17 797 75
rect 833 112 909 138
rect 833 78 849 112
rect 883 78 909 112
rect 833 53 909 78
rect 991 125 1057 269
rect 1236 213 1270 375
rect 1205 184 1271 213
rect 991 91 1007 125
rect 1041 91 1057 125
rect 991 62 1057 91
rect 1093 125 1159 154
rect 1093 91 1109 125
rect 1143 91 1159 125
rect 1205 150 1221 184
rect 1255 150 1271 184
rect 1205 121 1271 150
rect 1307 173 1373 375
rect 1307 139 1323 173
rect 1357 139 1373 173
rect 1409 260 1462 276
rect 1409 226 1425 260
rect 1459 226 1462 260
rect 1409 175 1462 226
rect 1498 245 1532 375
rect 1568 399 1921 422
rect 1955 399 1971 433
rect 1568 388 1971 399
rect 1568 331 1608 388
rect 1905 383 1971 388
rect 1568 297 1571 331
rect 1605 297 1608 331
rect 1568 281 1608 297
rect 1644 347 1869 352
rect 1644 331 1901 347
rect 1644 318 1851 331
rect 1644 245 1678 318
rect 1835 297 1851 318
rect 1885 297 1901 331
rect 1498 211 1678 245
rect 1714 276 1799 282
rect 1835 281 1901 297
rect 1937 345 1971 383
rect 2069 535 2135 649
rect 2069 501 2085 535
rect 2119 501 2135 535
rect 2069 431 2135 501
rect 2069 397 2085 431
rect 2119 397 2135 431
rect 2069 381 2135 397
rect 2224 579 2486 613
rect 1937 329 2188 345
rect 1937 295 2138 329
rect 2172 295 2188 329
rect 1937 287 2188 295
rect 2224 335 2258 579
rect 2294 500 2376 543
rect 2294 466 2310 500
rect 2344 466 2376 500
rect 2294 424 2376 466
rect 2224 319 2306 335
rect 1714 266 1759 276
rect 1714 232 1717 266
rect 1751 242 1759 266
rect 1793 242 1799 276
rect 1937 245 1971 287
rect 2224 285 2256 319
rect 2290 285 2306 319
rect 2224 269 2306 285
rect 2224 251 2258 269
rect 1751 232 1799 242
rect 1714 216 1799 232
rect 1849 243 1971 245
rect 1849 209 1865 243
rect 1899 211 1971 243
rect 2053 217 2258 251
rect 2342 233 2376 424
rect 2420 458 2486 579
rect 2621 575 2671 649
rect 2621 541 2637 575
rect 2621 494 2671 541
rect 2707 597 2773 613
rect 2707 563 2723 597
rect 2757 563 2773 597
rect 2865 602 2931 649
rect 2865 568 2881 602
rect 2915 568 2931 602
rect 2865 564 2931 568
rect 3078 602 3144 649
rect 3078 568 3094 602
rect 3128 568 3144 602
rect 3078 564 3144 568
rect 3180 597 3251 613
rect 2707 528 2773 563
rect 3214 563 3251 597
rect 2707 497 3144 528
rect 2707 463 2723 497
rect 2757 494 3144 497
rect 2757 463 2773 494
rect 2707 458 2773 463
rect 2420 424 2436 458
rect 2470 424 2486 458
rect 2420 390 2486 424
rect 2528 442 2773 458
rect 2528 408 2544 442
rect 2578 408 2773 442
rect 2528 392 2773 408
rect 2420 356 2436 390
rect 2470 356 2486 390
rect 2420 340 2486 356
rect 2600 319 2666 356
rect 2600 285 2616 319
rect 2650 285 2666 319
rect 2600 276 2666 285
rect 2600 242 2623 276
rect 2657 242 2666 276
rect 2600 236 2666 242
rect 2708 337 2774 353
rect 2708 303 2724 337
rect 2758 303 2774 337
rect 2708 287 2774 303
rect 1899 209 1915 211
rect 1849 193 1915 209
rect 1409 141 1711 175
rect 1307 100 1373 139
rect 1093 17 1159 91
rect 1575 89 1641 105
rect 1575 55 1591 89
rect 1625 55 1641 89
rect 1575 17 1641 55
rect 1677 87 1711 141
rect 1747 160 1813 180
rect 1747 126 1763 160
rect 1797 157 1813 160
rect 1951 158 2017 175
rect 1951 157 1967 158
rect 1797 126 1967 157
rect 1747 124 1967 126
rect 2001 124 2017 158
rect 1747 123 2017 124
rect 2053 87 2087 217
rect 2294 200 2376 233
rect 2708 200 2742 287
rect 2810 251 2844 494
rect 2294 191 2742 200
rect 1677 53 2087 87
rect 2123 165 2173 181
rect 2157 131 2173 165
rect 2123 17 2173 131
rect 2294 157 2310 191
rect 2344 166 2742 191
rect 2781 217 2844 251
rect 2880 442 3042 458
rect 2880 408 2992 442
rect 3026 408 3042 442
rect 2880 392 3042 408
rect 2880 338 2946 392
rect 2880 304 2896 338
rect 2930 304 2946 338
rect 2880 270 2946 304
rect 2880 236 2896 270
rect 2930 236 2946 270
rect 3001 319 3073 356
rect 3001 285 3023 319
rect 3057 285 3073 319
rect 3001 269 3073 285
rect 3110 331 3144 494
rect 3180 507 3251 563
rect 3214 473 3251 507
rect 3377 607 3427 649
rect 3377 573 3393 607
rect 3377 510 3427 573
rect 3180 417 3251 473
rect 3214 383 3251 417
rect 3180 367 3251 383
rect 3110 315 3181 331
rect 3110 281 3131 315
rect 3165 281 3181 315
rect 3110 265 3181 281
rect 2880 233 2946 236
rect 2781 204 2831 217
rect 2815 170 2831 204
rect 2880 199 3048 233
rect 3217 229 3251 367
rect 2344 157 2376 166
rect 2294 115 2376 157
rect 2529 114 2595 130
rect 2529 80 2545 114
rect 2579 80 2595 114
rect 2529 17 2595 80
rect 2647 114 2713 130
rect 2781 123 2831 170
rect 2867 131 2933 163
rect 2647 80 2663 114
rect 2697 87 2713 114
rect 2867 97 2883 131
rect 2917 97 2933 131
rect 2867 87 2933 97
rect 2697 80 2933 87
rect 2647 53 2933 80
rect 2982 116 3048 199
rect 2982 82 2998 116
rect 3032 82 3048 116
rect 2982 53 3048 82
rect 3084 213 3134 229
rect 3084 179 3100 213
rect 3084 103 3134 179
rect 3084 69 3100 103
rect 3084 17 3134 69
rect 3170 213 3251 229
rect 3170 179 3186 213
rect 3220 179 3251 213
rect 3170 103 3251 179
rect 3170 69 3186 103
rect 3220 69 3251 103
rect 3170 53 3251 69
rect 3291 483 3341 499
rect 3325 449 3341 483
rect 3291 413 3341 449
rect 3325 379 3341 413
rect 3291 327 3341 379
rect 3377 476 3393 510
rect 3377 413 3427 476
rect 3377 379 3393 413
rect 3377 363 3427 379
rect 3463 597 3534 613
rect 3463 563 3479 597
rect 3513 563 3534 597
rect 3463 505 3534 563
rect 3463 471 3479 505
rect 3513 471 3534 505
rect 3463 413 3534 471
rect 3463 379 3479 413
rect 3513 379 3534 413
rect 3463 363 3534 379
rect 3291 311 3464 327
rect 3291 277 3424 311
rect 3458 277 3464 311
rect 3291 261 3464 277
rect 3291 116 3332 261
rect 3500 225 3534 363
rect 3463 209 3534 225
rect 3463 175 3479 209
rect 3513 175 3534 209
rect 3291 82 3298 116
rect 3291 53 3332 82
rect 3368 116 3418 145
rect 3368 82 3384 116
rect 3368 17 3418 82
rect 3463 103 3534 175
rect 3463 69 3479 103
rect 3513 69 3534 103
rect 3463 53 3534 69
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 1759 242 1793 276
rect 2623 242 2657 276
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
<< metal1 >>
rect 0 683 3552 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3552 683
rect 0 617 3552 649
rect 1747 276 1805 282
rect 1747 242 1759 276
rect 1793 273 1805 276
rect 2611 276 2669 282
rect 2611 273 2623 276
rect 1793 245 2623 273
rect 1793 242 1805 245
rect 1747 236 1805 242
rect 2611 242 2623 245
rect 2657 242 2669 276
rect 2611 236 2669 242
rect 0 17 3552 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
rect 0 -49 3552 -17
<< labels >>
flabel pwell s 0 0 3552 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 3552 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 sdfbbn_1
flabel comment s 1064 243 1064 243 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 3552 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 3552 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 3007 316 3041 350 0 FreeSans 340 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 3487 94 3521 128 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 3487 168 3521 202 0 FreeSans 340 0 0 0 Q
port 11 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 3199 390 3233 424 0 FreeSans 340 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 3199 464 3233 498 0 FreeSans 340 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 3199 538 3233 572 0 FreeSans 340 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 SCE
port 5 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 SCD
port 4 nsew signal input
flabel locali s 319 168 353 202 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 2623 316 2657 350 0 FreeSans 340 0 0 0 SET_B
port 6 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 3552 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2990680
string GDS_START 2967988
<< end >>
