magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 1827 259 2015 273
rect 1472 229 2015 259
rect 497 227 682 229
rect 497 224 958 227
rect 494 191 958 224
rect 7 157 958 191
rect 1280 157 2015 229
rect 7 49 2015 157
rect 0 0 2016 49
<< scnmos >>
rect 86 81 116 165
rect 182 81 212 165
rect 254 81 284 165
rect 340 81 370 165
rect 573 119 603 203
rect 763 117 793 201
rect 849 117 879 201
rect 1039 47 1069 131
rect 1141 47 1171 131
rect 1359 119 1389 203
rect 1605 149 1635 233
rect 1691 149 1721 233
rect 1906 79 1936 247
<< scpmoshvt >>
rect 80 519 110 603
rect 166 519 196 603
rect 356 459 386 543
rect 442 459 472 543
rect 638 494 668 578
rect 852 501 882 585
rect 938 501 968 585
rect 1010 501 1040 585
rect 1110 501 1140 585
rect 1359 445 1389 529
rect 1605 367 1635 451
rect 1691 367 1721 451
rect 1906 367 1936 619
<< ndiff >>
rect 523 198 573 203
rect 520 178 573 198
rect 33 140 86 165
rect 33 106 41 140
rect 75 106 86 140
rect 33 81 86 106
rect 116 123 182 165
rect 116 89 127 123
rect 161 89 182 123
rect 116 81 182 89
rect 212 81 254 165
rect 284 157 340 165
rect 284 123 295 157
rect 329 123 340 157
rect 284 81 340 123
rect 370 128 437 165
rect 370 94 395 128
rect 429 94 437 128
rect 520 144 528 178
rect 562 144 573 178
rect 520 119 573 144
rect 603 178 656 203
rect 603 144 614 178
rect 648 144 656 178
rect 603 119 656 144
rect 710 175 763 201
rect 710 141 718 175
rect 752 141 763 175
rect 370 81 437 94
rect 710 117 763 141
rect 793 175 849 201
rect 793 141 804 175
rect 838 141 849 175
rect 793 117 849 141
rect 879 166 932 201
rect 879 132 890 166
rect 924 132 932 166
rect 879 117 932 132
rect 986 93 1039 131
rect 986 59 994 93
rect 1028 59 1039 93
rect 986 47 1039 59
rect 1069 89 1141 131
rect 1069 55 1094 89
rect 1128 55 1141 89
rect 1069 47 1141 55
rect 1171 105 1224 131
rect 1171 71 1182 105
rect 1216 71 1224 105
rect 1171 47 1224 71
rect 1498 208 1605 233
rect 1306 169 1359 203
rect 1306 135 1314 169
rect 1348 135 1359 169
rect 1306 119 1359 135
rect 1389 178 1442 203
rect 1389 144 1400 178
rect 1434 144 1442 178
rect 1498 174 1506 208
rect 1540 174 1605 208
rect 1498 149 1605 174
rect 1635 208 1691 233
rect 1635 174 1646 208
rect 1680 174 1691 208
rect 1635 149 1691 174
rect 1721 208 1774 233
rect 1721 174 1732 208
rect 1766 174 1774 208
rect 1721 149 1774 174
rect 1389 119 1442 144
rect 1853 235 1906 247
rect 1853 201 1861 235
rect 1895 201 1906 235
rect 1853 125 1906 201
rect 1853 91 1861 125
rect 1895 91 1906 125
rect 1853 79 1906 91
rect 1936 235 1989 247
rect 1936 201 1947 235
rect 1981 201 1989 235
rect 1936 125 1989 201
rect 1936 91 1947 125
rect 1981 91 1989 125
rect 1936 79 1989 91
<< pdiff >>
rect 27 578 80 603
rect 27 544 35 578
rect 69 544 80 578
rect 27 519 80 544
rect 110 578 166 603
rect 110 544 121 578
rect 155 544 166 578
rect 110 519 166 544
rect 196 587 249 603
rect 196 553 207 587
rect 241 553 249 587
rect 196 519 249 553
rect 585 553 638 578
rect 303 519 356 543
rect 303 485 311 519
rect 345 485 356 519
rect 303 459 356 485
rect 386 518 442 543
rect 386 484 397 518
rect 431 484 442 518
rect 386 459 442 484
rect 472 518 531 543
rect 472 484 483 518
rect 517 484 531 518
rect 585 519 593 553
rect 627 519 638 553
rect 585 494 638 519
rect 668 553 721 578
rect 668 519 679 553
rect 713 519 721 553
rect 668 494 721 519
rect 799 559 852 585
rect 799 525 807 559
rect 841 525 852 559
rect 799 501 852 525
rect 882 543 938 585
rect 882 509 893 543
rect 927 509 938 543
rect 882 501 938 509
rect 968 501 1010 585
rect 1040 573 1110 585
rect 1040 539 1060 573
rect 1094 539 1110 573
rect 1040 501 1110 539
rect 1140 560 1193 585
rect 1140 526 1151 560
rect 1185 526 1193 560
rect 1140 501 1193 526
rect 472 459 531 484
rect 1853 607 1906 619
rect 1853 573 1861 607
rect 1895 573 1906 607
rect 1290 513 1359 529
rect 1290 479 1300 513
rect 1334 479 1359 513
rect 1290 445 1359 479
rect 1389 513 1442 529
rect 1389 479 1400 513
rect 1434 479 1442 513
rect 1389 445 1442 479
rect 1853 510 1906 573
rect 1853 476 1861 510
rect 1895 476 1906 510
rect 1552 426 1605 451
rect 1552 392 1560 426
rect 1594 392 1605 426
rect 1552 367 1605 392
rect 1635 426 1691 451
rect 1635 392 1646 426
rect 1680 392 1691 426
rect 1635 367 1691 392
rect 1721 426 1774 451
rect 1721 392 1732 426
rect 1766 392 1774 426
rect 1721 367 1774 392
rect 1853 413 1906 476
rect 1853 379 1861 413
rect 1895 379 1906 413
rect 1853 367 1906 379
rect 1936 599 1989 619
rect 1936 565 1947 599
rect 1981 565 1989 599
rect 1936 502 1989 565
rect 1936 468 1947 502
rect 1981 468 1989 502
rect 1936 413 1989 468
rect 1936 379 1947 413
rect 1981 379 1989 413
rect 1936 367 1989 379
<< ndiffc >>
rect 41 106 75 140
rect 127 89 161 123
rect 295 123 329 157
rect 395 94 429 128
rect 528 144 562 178
rect 614 144 648 178
rect 718 141 752 175
rect 804 141 838 175
rect 890 132 924 166
rect 994 59 1028 93
rect 1094 55 1128 89
rect 1182 71 1216 105
rect 1314 135 1348 169
rect 1400 144 1434 178
rect 1506 174 1540 208
rect 1646 174 1680 208
rect 1732 174 1766 208
rect 1861 201 1895 235
rect 1861 91 1895 125
rect 1947 201 1981 235
rect 1947 91 1981 125
<< pdiffc >>
rect 35 544 69 578
rect 121 544 155 578
rect 207 553 241 587
rect 311 485 345 519
rect 397 484 431 518
rect 483 484 517 518
rect 593 519 627 553
rect 679 519 713 553
rect 807 525 841 559
rect 893 509 927 543
rect 1060 539 1094 573
rect 1151 526 1185 560
rect 1861 573 1895 607
rect 1300 479 1334 513
rect 1400 479 1434 513
rect 1861 476 1895 510
rect 1560 392 1594 426
rect 1646 392 1680 426
rect 1732 392 1766 426
rect 1861 379 1895 413
rect 1947 565 1981 599
rect 1947 468 1981 502
rect 1947 379 1981 413
<< poly >>
rect 80 603 110 629
rect 166 603 196 629
rect 638 578 668 604
rect 852 585 882 611
rect 938 585 968 611
rect 1010 585 1040 611
rect 1110 585 1140 611
rect 1245 606 1530 627
rect 1906 619 1936 645
rect 1245 597 1480 606
rect 356 543 386 569
rect 442 543 472 569
rect 80 376 110 519
rect 166 451 196 519
rect 166 435 232 451
rect 166 401 182 435
rect 216 401 232 435
rect 44 360 116 376
rect 44 326 60 360
rect 94 326 116 360
rect 44 292 116 326
rect 166 367 232 401
rect 166 333 182 367
rect 216 333 232 367
rect 166 317 232 333
rect 44 258 60 292
rect 94 258 116 292
rect 44 242 116 258
rect 86 165 116 242
rect 182 165 212 317
rect 356 269 386 459
rect 442 437 472 459
rect 638 437 668 494
rect 852 479 882 501
rect 442 407 668 437
rect 716 449 882 479
rect 435 338 501 354
rect 435 304 451 338
rect 485 304 501 338
rect 435 270 501 304
rect 435 269 451 270
rect 254 239 451 269
rect 254 165 284 239
rect 435 236 451 239
rect 485 236 501 270
rect 435 220 501 236
rect 573 255 603 407
rect 716 359 746 449
rect 938 428 968 501
rect 924 407 968 428
rect 680 343 746 359
rect 680 309 696 343
rect 730 309 746 343
rect 680 275 746 309
rect 680 255 696 275
rect 573 241 696 255
rect 730 255 746 275
rect 835 398 968 407
rect 835 391 954 398
rect 835 357 851 391
rect 885 357 954 391
rect 835 323 954 357
rect 1010 350 1040 501
rect 1110 366 1140 501
rect 1110 350 1176 366
rect 835 289 851 323
rect 885 289 954 323
rect 835 273 954 289
rect 996 334 1062 350
rect 996 300 1012 334
rect 1046 300 1062 334
rect 730 241 793 255
rect 573 225 793 241
rect 573 203 603 225
rect 340 165 370 191
rect 763 201 793 225
rect 849 201 879 273
rect 996 266 1062 300
rect 996 232 1012 266
rect 1046 232 1062 266
rect 1110 316 1126 350
rect 1160 316 1176 350
rect 1110 282 1176 316
rect 1110 248 1126 282
rect 1160 248 1176 282
rect 1110 232 1176 248
rect 1245 359 1275 597
rect 1464 572 1480 597
rect 1514 572 1530 606
rect 1464 556 1530 572
rect 1359 529 1389 555
rect 1605 451 1635 477
rect 1691 451 1721 477
rect 1359 389 1389 445
rect 1359 373 1425 389
rect 1245 343 1311 359
rect 1245 309 1261 343
rect 1295 309 1311 343
rect 1245 275 1311 309
rect 1245 241 1261 275
rect 1295 241 1311 275
rect 996 216 1062 232
rect 573 93 603 119
rect 1032 184 1062 216
rect 1032 154 1069 184
rect 1039 131 1069 154
rect 1141 131 1171 232
rect 1245 225 1311 241
rect 1359 339 1375 373
rect 1409 339 1425 373
rect 1359 305 1425 339
rect 1359 271 1375 305
rect 1409 285 1425 305
rect 1605 285 1635 367
rect 1409 271 1635 285
rect 1359 255 1635 271
rect 86 55 116 81
rect 182 55 212 81
rect 254 55 284 81
rect 340 51 370 81
rect 763 51 793 117
rect 849 91 879 117
rect 340 21 793 51
rect 1245 51 1275 225
rect 1359 203 1389 255
rect 1605 233 1635 255
rect 1691 285 1721 367
rect 1906 335 1936 367
rect 1861 319 1936 335
rect 1861 285 1877 319
rect 1911 285 1936 319
rect 1691 255 1819 285
rect 1861 269 1936 285
rect 1691 233 1721 255
rect 1605 123 1635 149
rect 1691 123 1721 149
rect 1359 93 1389 119
rect 1789 51 1819 255
rect 1906 247 1936 269
rect 1906 53 1936 79
rect 1039 21 1069 47
rect 1141 21 1171 47
rect 1245 21 1819 51
<< polycont >>
rect 182 401 216 435
rect 60 326 94 360
rect 182 333 216 367
rect 60 258 94 292
rect 451 304 485 338
rect 451 236 485 270
rect 696 309 730 343
rect 696 241 730 275
rect 851 357 885 391
rect 851 289 885 323
rect 1012 300 1046 334
rect 1012 232 1046 266
rect 1126 316 1160 350
rect 1126 248 1160 282
rect 1480 572 1514 606
rect 1261 309 1295 343
rect 1261 241 1295 275
rect 1375 339 1409 373
rect 1375 271 1409 305
rect 1877 285 1911 319
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 19 578 71 594
rect 19 544 35 578
rect 69 544 71 578
rect 19 503 71 544
rect 105 578 171 649
rect 105 544 121 578
rect 155 544 171 578
rect 105 537 171 544
rect 205 587 533 607
rect 205 553 207 587
rect 241 573 533 587
rect 241 553 257 573
rect 205 537 257 553
rect 295 519 347 535
rect 295 503 311 519
rect 19 485 311 503
rect 345 485 347 519
rect 19 469 347 485
rect 381 518 447 534
rect 381 484 397 518
rect 431 484 447 518
rect 17 360 110 435
rect 17 326 60 360
rect 94 326 110 360
rect 17 292 110 326
rect 17 258 60 292
rect 94 258 110 292
rect 17 231 110 258
rect 166 401 182 435
rect 216 401 290 435
rect 166 367 290 401
rect 166 333 182 367
rect 216 333 290 367
rect 166 235 290 333
rect 381 434 447 484
rect 481 518 533 573
rect 481 484 483 518
rect 517 484 533 518
rect 481 468 533 484
rect 577 553 635 569
rect 577 519 593 553
rect 627 519 635 553
rect 381 424 461 434
rect 577 429 635 519
rect 669 553 729 649
rect 669 519 679 553
rect 713 519 729 553
rect 669 503 729 519
rect 791 581 1023 615
rect 791 559 841 581
rect 791 525 807 559
rect 791 509 841 525
rect 877 543 955 547
rect 877 509 893 543
rect 927 509 955 543
rect 877 505 955 509
rect 381 390 415 424
rect 449 390 461 424
rect 381 388 461 390
rect 530 395 887 429
rect 381 201 415 388
rect 530 354 564 395
rect 835 391 887 395
rect 451 338 564 354
rect 485 304 564 338
rect 451 270 564 304
rect 485 236 564 270
rect 451 220 564 236
rect 598 343 730 359
rect 598 309 696 343
rect 598 275 730 309
rect 598 241 696 275
rect 835 357 851 391
rect 885 357 887 391
rect 835 323 887 357
rect 835 289 851 323
rect 885 289 887 323
rect 835 273 887 289
rect 921 421 955 505
rect 989 489 1023 581
rect 1057 573 1107 649
rect 1057 539 1060 573
rect 1094 539 1107 573
rect 1057 523 1107 539
rect 1141 560 1201 576
rect 1141 526 1151 560
rect 1185 526 1201 560
rect 1141 489 1201 526
rect 989 455 1201 489
rect 1282 513 1350 649
rect 1282 479 1300 513
rect 1334 479 1350 513
rect 1282 475 1350 479
rect 1384 606 1530 615
rect 1384 572 1480 606
rect 1514 572 1530 606
rect 1384 556 1530 572
rect 1845 607 1911 649
rect 1845 573 1861 607
rect 1895 573 1911 607
rect 1384 513 1450 556
rect 1384 479 1400 513
rect 1434 479 1450 513
rect 1384 475 1450 479
rect 1486 476 1770 522
rect 1486 441 1520 476
rect 1289 421 1520 441
rect 921 407 1520 421
rect 921 387 1323 407
rect 598 225 730 241
rect 921 237 955 387
rect 25 163 245 197
rect 25 140 77 163
rect 25 106 41 140
rect 75 106 77 140
rect 25 90 77 106
rect 111 123 177 129
rect 111 89 127 123
rect 161 89 177 123
rect 111 17 177 89
rect 211 87 245 163
rect 279 167 415 201
rect 512 178 564 220
rect 795 203 955 237
rect 989 334 1046 353
rect 989 300 1012 334
rect 989 266 1046 300
rect 989 232 1012 266
rect 1080 350 1176 353
rect 1080 316 1126 350
rect 1160 316 1176 350
rect 1080 282 1176 316
rect 1080 248 1126 282
rect 1160 248 1176 282
rect 1080 242 1176 248
rect 1245 343 1311 353
rect 1245 309 1261 343
rect 1295 309 1311 343
rect 1245 275 1311 309
rect 989 216 1046 232
rect 1245 241 1261 275
rect 1295 241 1311 275
rect 1359 339 1375 373
rect 1409 339 1425 373
rect 1359 305 1425 339
rect 1359 271 1375 305
rect 1409 271 1425 305
rect 1245 237 1311 241
rect 1245 203 1450 237
rect 279 157 345 167
rect 279 123 295 157
rect 329 123 345 157
rect 512 144 528 178
rect 562 144 564 178
rect 379 128 445 133
rect 512 128 564 144
rect 598 178 664 191
rect 598 144 614 178
rect 648 144 664 178
rect 379 94 395 128
rect 429 94 445 128
rect 379 87 445 94
rect 211 53 445 87
rect 598 17 664 144
rect 702 175 761 191
rect 702 141 718 175
rect 752 141 761 175
rect 702 89 761 141
rect 795 175 840 203
rect 795 141 804 175
rect 838 141 840 175
rect 1400 178 1450 203
rect 795 125 840 141
rect 874 166 1232 169
rect 874 132 890 166
rect 924 132 1232 166
rect 874 129 1232 132
rect 874 123 940 129
rect 1178 105 1232 129
rect 978 93 1044 95
rect 978 89 994 93
rect 702 59 994 89
rect 1028 59 1044 93
rect 702 51 1044 59
rect 1078 89 1144 95
rect 1078 55 1094 89
rect 1128 55 1144 89
rect 1178 71 1182 105
rect 1216 71 1232 105
rect 1178 55 1232 71
rect 1298 135 1314 169
rect 1348 135 1364 169
rect 1078 17 1144 55
rect 1298 17 1364 135
rect 1434 144 1450 178
rect 1486 224 1520 407
rect 1556 426 1610 442
rect 1556 392 1560 426
rect 1594 424 1610 426
rect 1556 390 1567 392
rect 1601 390 1610 424
rect 1556 376 1610 390
rect 1486 208 1542 224
rect 1486 174 1506 208
rect 1540 174 1542 208
rect 1486 158 1542 174
rect 1400 128 1450 144
rect 1576 124 1610 376
rect 1644 426 1688 442
rect 1644 392 1646 426
rect 1680 392 1688 426
rect 1644 335 1688 392
rect 1722 426 1770 476
rect 1722 392 1732 426
rect 1766 392 1770 426
rect 1722 376 1770 392
rect 1845 510 1911 573
rect 1845 476 1861 510
rect 1895 476 1911 510
rect 1845 413 1911 476
rect 1845 379 1861 413
rect 1895 379 1911 413
rect 1845 369 1911 379
rect 1945 599 1999 615
rect 1945 565 1947 599
rect 1981 565 1999 599
rect 1945 502 1999 565
rect 1945 468 1947 502
rect 1981 468 1999 502
rect 1945 413 1999 468
rect 1945 379 1947 413
rect 1981 379 1999 413
rect 1644 319 1911 335
rect 1644 285 1877 319
rect 1644 269 1911 285
rect 1644 208 1689 269
rect 1945 235 1999 379
rect 1644 174 1646 208
rect 1680 174 1689 208
rect 1644 158 1689 174
rect 1723 208 1782 224
rect 1723 174 1732 208
rect 1766 174 1782 208
rect 1723 124 1782 174
rect 1576 78 1782 124
rect 1845 201 1861 235
rect 1895 201 1911 235
rect 1845 125 1911 201
rect 1845 91 1861 125
rect 1895 91 1911 125
rect 1845 17 1911 91
rect 1945 201 1947 235
rect 1981 201 1999 235
rect 1945 125 1999 201
rect 1945 91 1947 125
rect 1981 91 1999 125
rect 1945 75 1999 91
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 415 390 449 424
rect 1567 392 1594 424
rect 1594 392 1601 424
rect 1567 390 1601 392
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 403 424 461 430
rect 403 390 415 424
rect 449 421 461 424
rect 1555 424 1613 430
rect 1555 421 1567 424
rect 449 393 1567 421
rect 449 390 461 393
rect 403 384 461 390
rect 1555 390 1567 393
rect 1601 390 1613 424
rect 1555 384 1613 390
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
rlabel comment s 0 0 0 0 4 mux4_1
flabel comment s 1256 486 1256 486 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 31 390 65 424 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 1087 242 1121 276 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 1951 94 1985 128 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 168 1985 202 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 242 1985 276 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 316 1985 350 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 390 1985 424 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 464 1985 498 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1951 538 1985 572 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 1522152
string GDS_START 1505708
<< end >>
