magic
tech sky130A
magscale 1 2
timestamp 1627202635
<< checkpaint >>
rect -1298 -1309 2450 1975
<< nwell >>
rect -38 332 1190 704
<< pwell >>
rect 1 49 1151 248
rect 0 0 1152 49
<< scpmos >>
rect 84 368 120 592
rect 174 368 210 592
rect 264 368 300 592
rect 354 368 390 592
rect 454 368 490 592
rect 554 368 590 592
rect 644 368 680 592
rect 744 368 780 592
rect 834 368 870 592
rect 931 368 967 592
rect 1024 368 1060 592
<< nmoslvt >>
rect 84 74 114 222
rect 179 74 209 222
rect 265 74 295 222
rect 351 74 381 222
rect 437 74 467 222
rect 537 74 567 222
rect 623 74 653 222
rect 737 74 767 222
rect 823 74 853 222
rect 937 74 967 222
rect 1024 74 1054 222
<< ndiff >>
rect 27 210 84 222
rect 27 176 39 210
rect 73 176 84 210
rect 27 120 84 176
rect 27 86 39 120
rect 73 86 84 120
rect 27 74 84 86
rect 114 152 179 222
rect 114 118 125 152
rect 159 118 179 152
rect 114 74 179 118
rect 209 210 265 222
rect 209 176 220 210
rect 254 176 265 210
rect 209 120 265 176
rect 209 86 220 120
rect 254 86 265 120
rect 209 74 265 86
rect 295 152 351 222
rect 295 118 306 152
rect 340 118 351 152
rect 295 74 351 118
rect 381 210 437 222
rect 381 176 392 210
rect 426 176 437 210
rect 381 120 437 176
rect 381 86 392 120
rect 426 86 437 120
rect 381 74 437 86
rect 467 142 537 222
rect 467 108 478 142
rect 512 108 537 142
rect 467 74 537 108
rect 567 210 623 222
rect 567 176 578 210
rect 612 176 623 210
rect 567 120 623 176
rect 567 86 578 120
rect 612 86 623 120
rect 567 74 623 86
rect 653 142 737 222
rect 653 108 678 142
rect 712 108 737 142
rect 653 74 737 108
rect 767 210 823 222
rect 767 176 778 210
rect 812 176 823 210
rect 767 120 823 176
rect 767 86 778 120
rect 812 86 823 120
rect 767 74 823 86
rect 853 142 937 222
rect 853 108 878 142
rect 912 108 937 142
rect 853 74 937 108
rect 967 210 1024 222
rect 967 176 978 210
rect 1012 176 1024 210
rect 967 120 1024 176
rect 967 86 978 120
rect 1012 86 1024 120
rect 967 74 1024 86
rect 1054 210 1125 222
rect 1054 176 1079 210
rect 1113 176 1125 210
rect 1054 120 1125 176
rect 1054 86 1079 120
rect 1113 86 1125 120
rect 1054 74 1125 86
<< pdiff >>
rect 28 580 84 592
rect 28 546 40 580
rect 74 546 84 580
rect 28 510 84 546
rect 28 476 40 510
rect 74 476 84 510
rect 28 440 84 476
rect 28 406 40 440
rect 74 406 84 440
rect 28 368 84 406
rect 120 580 174 592
rect 120 546 130 580
rect 164 546 174 580
rect 120 508 174 546
rect 120 474 130 508
rect 164 474 174 508
rect 120 368 174 474
rect 210 580 264 592
rect 210 546 220 580
rect 254 546 264 580
rect 210 510 264 546
rect 210 476 220 510
rect 254 476 264 510
rect 210 440 264 476
rect 210 406 220 440
rect 254 406 264 440
rect 210 368 264 406
rect 300 580 354 592
rect 300 546 310 580
rect 344 546 354 580
rect 300 508 354 546
rect 300 474 310 508
rect 344 474 354 508
rect 300 368 354 474
rect 390 580 454 592
rect 390 546 410 580
rect 444 546 454 580
rect 390 497 454 546
rect 390 463 410 497
rect 444 463 454 497
rect 390 414 454 463
rect 390 380 410 414
rect 444 380 454 414
rect 390 368 454 380
rect 490 580 554 592
rect 490 546 500 580
rect 534 546 554 580
rect 490 478 554 546
rect 490 444 500 478
rect 534 444 554 478
rect 490 368 554 444
rect 590 580 644 592
rect 590 546 600 580
rect 634 546 644 580
rect 590 497 644 546
rect 590 463 600 497
rect 634 463 644 497
rect 590 414 644 463
rect 590 380 600 414
rect 634 380 644 414
rect 590 368 644 380
rect 680 580 744 592
rect 680 546 690 580
rect 724 546 744 580
rect 680 478 744 546
rect 680 444 690 478
rect 724 444 744 478
rect 680 368 744 444
rect 780 580 834 592
rect 780 546 790 580
rect 824 546 834 580
rect 780 497 834 546
rect 780 463 790 497
rect 824 463 834 497
rect 780 414 834 463
rect 780 380 790 414
rect 824 380 834 414
rect 780 368 834 380
rect 870 580 931 592
rect 870 546 880 580
rect 914 546 931 580
rect 870 478 931 546
rect 870 444 880 478
rect 914 444 931 478
rect 870 368 931 444
rect 967 580 1024 592
rect 967 546 980 580
rect 1014 546 1024 580
rect 967 497 1024 546
rect 967 463 980 497
rect 1014 463 1024 497
rect 967 414 1024 463
rect 967 380 980 414
rect 1014 380 1024 414
rect 967 368 1024 380
rect 1060 580 1116 592
rect 1060 546 1070 580
rect 1104 546 1116 580
rect 1060 497 1116 546
rect 1060 463 1070 497
rect 1104 463 1116 497
rect 1060 414 1116 463
rect 1060 380 1070 414
rect 1104 380 1116 414
rect 1060 368 1116 380
<< ndiffc >>
rect 39 176 73 210
rect 39 86 73 120
rect 125 118 159 152
rect 220 176 254 210
rect 220 86 254 120
rect 306 118 340 152
rect 392 176 426 210
rect 392 86 426 120
rect 478 108 512 142
rect 578 176 612 210
rect 578 86 612 120
rect 678 108 712 142
rect 778 176 812 210
rect 778 86 812 120
rect 878 108 912 142
rect 978 176 1012 210
rect 978 86 1012 120
rect 1079 176 1113 210
rect 1079 86 1113 120
<< pdiffc >>
rect 40 546 74 580
rect 40 476 74 510
rect 40 406 74 440
rect 130 546 164 580
rect 130 474 164 508
rect 220 546 254 580
rect 220 476 254 510
rect 220 406 254 440
rect 310 546 344 580
rect 310 474 344 508
rect 410 546 444 580
rect 410 463 444 497
rect 410 380 444 414
rect 500 546 534 580
rect 500 444 534 478
rect 600 546 634 580
rect 600 463 634 497
rect 600 380 634 414
rect 690 546 724 580
rect 690 444 724 478
rect 790 546 824 580
rect 790 463 824 497
rect 790 380 824 414
rect 880 546 914 580
rect 880 444 914 478
rect 980 546 1014 580
rect 980 463 1014 497
rect 980 380 1014 414
rect 1070 546 1104 580
rect 1070 463 1104 497
rect 1070 380 1104 414
<< poly >>
rect 84 592 120 618
rect 174 592 210 618
rect 264 592 300 618
rect 354 592 390 618
rect 454 592 490 618
rect 554 592 590 618
rect 644 592 680 618
rect 744 592 780 618
rect 834 592 870 618
rect 931 592 967 618
rect 1024 592 1060 618
rect 84 336 120 368
rect 174 336 210 368
rect 264 336 300 368
rect 84 320 300 336
rect 354 326 390 368
rect 454 326 490 368
rect 554 326 590 368
rect 644 326 680 368
rect 744 326 780 368
rect 834 326 870 368
rect 931 326 967 368
rect 1024 326 1060 368
rect 84 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 300 320
rect 84 270 300 286
rect 351 310 1060 326
rect 351 276 367 310
rect 401 276 435 310
rect 469 276 503 310
rect 537 276 571 310
rect 605 276 639 310
rect 673 276 707 310
rect 741 276 775 310
rect 809 276 843 310
rect 877 276 911 310
rect 945 276 1060 310
rect 84 222 114 270
rect 179 222 209 270
rect 265 222 295 270
rect 351 260 1060 276
rect 351 222 381 260
rect 437 222 467 260
rect 537 222 567 260
rect 623 222 653 260
rect 737 222 767 260
rect 823 222 853 260
rect 937 222 967 260
rect 1024 222 1054 260
rect 84 48 114 74
rect 179 48 209 74
rect 265 48 295 74
rect 351 48 381 74
rect 437 48 467 74
rect 537 48 567 74
rect 623 48 653 74
rect 737 48 767 74
rect 823 48 853 74
rect 937 48 967 74
rect 1024 48 1054 74
<< polycont >>
rect 100 286 134 320
rect 168 286 202 320
rect 236 286 270 320
rect 367 276 401 310
rect 435 276 469 310
rect 503 276 537 310
rect 571 276 605 310
rect 639 276 673 310
rect 707 276 741 310
rect 775 276 809 310
rect 843 276 877 310
rect 911 276 945 310
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 24 580 90 596
rect 24 546 40 580
rect 74 546 90 580
rect 24 510 90 546
rect 24 476 40 510
rect 74 476 90 510
rect 24 440 90 476
rect 130 580 164 649
rect 130 508 164 546
rect 130 458 164 474
rect 204 580 270 596
rect 204 546 220 580
rect 254 546 270 580
rect 204 510 270 546
rect 204 476 220 510
rect 254 476 270 510
rect 24 406 40 440
rect 74 424 90 440
rect 204 440 270 476
rect 310 580 360 649
rect 344 546 360 580
rect 310 508 360 546
rect 344 474 360 508
rect 310 458 360 474
rect 394 580 460 596
rect 394 546 410 580
rect 444 546 460 580
rect 394 497 460 546
rect 394 463 410 497
rect 444 463 460 497
rect 204 424 220 440
rect 74 406 220 424
rect 254 424 270 440
rect 254 406 354 424
rect 24 390 354 406
rect 25 320 286 356
rect 25 286 100 320
rect 134 286 168 320
rect 202 286 236 320
rect 270 286 286 320
rect 25 270 286 286
rect 320 326 354 390
rect 394 414 460 463
rect 500 580 550 649
rect 534 546 550 580
rect 500 478 550 546
rect 534 444 550 478
rect 500 428 550 444
rect 584 580 650 596
rect 584 546 600 580
rect 634 546 650 580
rect 584 497 650 546
rect 584 463 600 497
rect 634 463 650 497
rect 394 380 410 414
rect 444 394 460 414
rect 584 414 650 463
rect 690 580 740 649
rect 724 546 740 580
rect 690 478 740 546
rect 724 444 740 478
rect 690 428 740 444
rect 774 580 840 596
rect 774 546 790 580
rect 824 546 840 580
rect 774 497 840 546
rect 774 463 790 497
rect 824 463 840 497
rect 584 394 600 414
rect 444 380 600 394
rect 634 394 650 414
rect 774 414 840 463
rect 880 580 930 649
rect 914 546 930 580
rect 880 478 930 546
rect 914 444 930 478
rect 880 428 930 444
rect 964 580 1031 596
rect 964 546 980 580
rect 1014 546 1031 580
rect 964 497 1031 546
rect 964 463 980 497
rect 1014 463 1031 497
rect 774 394 790 414
rect 634 380 790 394
rect 824 394 840 414
rect 964 414 1031 463
rect 964 394 980 414
rect 824 380 980 394
rect 1014 380 1031 414
rect 394 360 1031 380
rect 1070 580 1120 649
rect 1104 546 1120 580
rect 1070 497 1120 546
rect 1104 463 1120 497
rect 1070 414 1120 463
rect 1104 380 1120 414
rect 1070 364 1120 380
rect 320 310 961 326
rect 320 276 367 310
rect 401 276 435 310
rect 469 276 503 310
rect 537 276 571 310
rect 605 276 639 310
rect 673 276 707 310
rect 741 276 775 310
rect 809 276 843 310
rect 877 276 911 310
rect 945 276 961 310
rect 320 260 961 276
rect 320 236 354 260
rect 23 210 354 236
rect 995 226 1029 360
rect 23 176 39 210
rect 73 202 220 210
rect 23 120 73 176
rect 254 202 354 210
rect 392 210 1029 226
rect 23 86 39 120
rect 23 70 73 86
rect 109 152 175 168
rect 109 118 125 152
rect 159 118 175 152
rect 109 17 175 118
rect 220 120 254 176
rect 426 192 578 210
rect 220 70 254 86
rect 290 152 356 168
rect 290 118 306 152
rect 340 118 356 152
rect 290 17 356 118
rect 392 120 426 176
rect 562 176 578 192
rect 612 192 778 210
rect 612 176 628 192
rect 392 70 426 86
rect 462 142 528 158
rect 462 108 478 142
rect 512 108 528 142
rect 462 17 528 108
rect 562 120 628 176
rect 762 176 778 192
rect 812 192 978 210
rect 812 176 828 192
rect 562 86 578 120
rect 612 86 628 120
rect 562 70 628 86
rect 662 142 728 158
rect 662 108 678 142
rect 712 108 728 142
rect 662 17 728 108
rect 762 120 828 176
rect 962 176 978 192
rect 1012 176 1029 210
rect 762 86 778 120
rect 812 86 828 120
rect 762 70 828 86
rect 862 142 928 158
rect 862 108 878 142
rect 912 108 928 142
rect 862 17 928 108
rect 962 120 1029 176
rect 962 86 978 120
rect 1012 86 1029 120
rect 962 70 1029 86
rect 1063 210 1129 226
rect 1063 176 1079 210
rect 1113 176 1129 210
rect 1063 120 1129 176
rect 1063 86 1079 120
rect 1113 86 1129 120
rect 1063 17 1129 86
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
<< metal1 >>
rect 0 683 1152 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1152 683
rect 0 617 1152 649
rect 0 17 1152 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1152 17
rect 0 -49 1152 -17
<< labels >>
flabel pwell s 0 0 1152 49 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 0 617 1152 666 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
rlabel comment s 0 0 0 0 4 buf_8
flabel metal1 s 0 617 1152 666 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1152 49 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 464 1025 498 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 538 1025 572 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1152 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_ms/gds/sky130_fd_sc_ms.gds
string LEFsymmetry X Y
string GDS_END 3030600
string GDS_START 3021160
<< end >>
