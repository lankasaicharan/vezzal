magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3122 1975
<< nwell >>
rect -38 331 1862 704
<< pwell >>
rect 89 241 281 263
rect 89 49 1823 241
rect 0 0 1824 49
<< scnmos >>
rect 172 69 202 237
rect 424 47 454 215
rect 510 47 540 215
rect 596 47 626 215
rect 682 47 712 215
rect 768 47 798 215
rect 854 47 884 215
rect 940 47 970 215
rect 1026 47 1056 215
rect 1112 47 1142 215
rect 1198 47 1228 215
rect 1284 47 1314 215
rect 1370 47 1400 215
rect 1456 47 1486 215
rect 1542 47 1572 215
rect 1628 47 1658 215
rect 1714 47 1744 215
<< scpmoshvt >>
rect 152 367 182 619
rect 418 367 448 619
rect 504 367 534 619
rect 590 367 620 619
rect 676 367 706 619
rect 762 367 792 619
rect 848 367 878 619
rect 934 367 964 619
rect 1020 367 1050 619
rect 1106 367 1136 619
rect 1192 367 1222 619
rect 1278 367 1308 619
rect 1364 367 1394 619
rect 1450 367 1480 619
rect 1536 367 1566 619
rect 1622 367 1652 619
rect 1708 367 1738 619
<< ndiff >>
rect 115 192 172 237
rect 115 158 127 192
rect 161 158 172 192
rect 115 115 172 158
rect 115 81 127 115
rect 161 81 172 115
rect 115 69 172 81
rect 202 225 255 237
rect 202 191 213 225
rect 247 191 255 225
rect 202 115 255 191
rect 202 81 213 115
rect 247 81 255 115
rect 202 69 255 81
rect 371 203 424 215
rect 371 169 379 203
rect 413 169 424 203
rect 371 101 424 169
rect 371 67 379 101
rect 413 67 424 101
rect 371 47 424 67
rect 454 207 510 215
rect 454 173 465 207
rect 499 173 510 207
rect 454 93 510 173
rect 454 59 465 93
rect 499 59 510 93
rect 454 47 510 59
rect 540 203 596 215
rect 540 169 551 203
rect 585 169 596 203
rect 540 101 596 169
rect 540 67 551 101
rect 585 67 596 101
rect 540 47 596 67
rect 626 207 682 215
rect 626 173 637 207
rect 671 173 682 207
rect 626 93 682 173
rect 626 59 637 93
rect 671 59 682 93
rect 626 47 682 59
rect 712 203 768 215
rect 712 169 723 203
rect 757 169 768 203
rect 712 101 768 169
rect 712 67 723 101
rect 757 67 768 101
rect 712 47 768 67
rect 798 207 854 215
rect 798 173 809 207
rect 843 173 854 207
rect 798 93 854 173
rect 798 59 809 93
rect 843 59 854 93
rect 798 47 854 59
rect 884 203 940 215
rect 884 169 895 203
rect 929 169 940 203
rect 884 101 940 169
rect 884 67 895 101
rect 929 67 940 101
rect 884 47 940 67
rect 970 192 1026 215
rect 970 158 981 192
rect 1015 158 1026 192
rect 970 89 1026 158
rect 970 55 981 89
rect 1015 55 1026 89
rect 970 47 1026 55
rect 1056 203 1112 215
rect 1056 169 1067 203
rect 1101 169 1112 203
rect 1056 93 1112 169
rect 1056 59 1067 93
rect 1101 59 1112 93
rect 1056 47 1112 59
rect 1142 195 1198 215
rect 1142 161 1153 195
rect 1187 161 1198 195
rect 1142 47 1198 161
rect 1228 105 1284 215
rect 1228 71 1239 105
rect 1273 71 1284 105
rect 1228 47 1284 71
rect 1314 190 1370 215
rect 1314 156 1325 190
rect 1359 156 1370 190
rect 1314 47 1370 156
rect 1400 105 1456 215
rect 1400 71 1411 105
rect 1445 71 1456 105
rect 1400 47 1456 71
rect 1486 195 1542 215
rect 1486 161 1497 195
rect 1531 161 1542 195
rect 1486 47 1542 161
rect 1572 165 1628 215
rect 1572 131 1583 165
rect 1617 131 1628 165
rect 1572 90 1628 131
rect 1572 56 1583 90
rect 1617 56 1628 90
rect 1572 47 1628 56
rect 1658 173 1714 215
rect 1658 139 1669 173
rect 1703 139 1714 173
rect 1658 47 1714 139
rect 1744 203 1797 215
rect 1744 169 1755 203
rect 1789 169 1797 203
rect 1744 105 1797 169
rect 1744 71 1755 105
rect 1789 71 1797 105
rect 1744 47 1797 71
<< pdiff >>
rect 99 607 152 619
rect 99 573 107 607
rect 141 573 152 607
rect 99 520 152 573
rect 99 486 107 520
rect 141 486 152 520
rect 99 434 152 486
rect 99 400 107 434
rect 141 400 152 434
rect 99 367 152 400
rect 182 599 235 619
rect 182 565 193 599
rect 227 565 235 599
rect 182 508 235 565
rect 365 599 418 619
rect 365 565 373 599
rect 407 565 418 599
rect 182 474 193 508
rect 227 474 235 508
rect 182 421 235 474
rect 182 387 193 421
rect 227 387 235 421
rect 182 367 235 387
rect 365 510 418 565
rect 365 476 373 510
rect 407 476 418 510
rect 365 413 418 476
rect 365 379 373 413
rect 407 379 418 413
rect 365 367 418 379
rect 448 607 504 619
rect 448 573 459 607
rect 493 573 504 607
rect 448 516 504 573
rect 448 482 459 516
rect 493 482 504 516
rect 448 428 504 482
rect 448 394 459 428
rect 493 394 504 428
rect 448 367 504 394
rect 534 599 590 619
rect 534 565 545 599
rect 579 565 590 599
rect 534 510 590 565
rect 534 476 545 510
rect 579 476 590 510
rect 534 413 590 476
rect 534 379 545 413
rect 579 379 590 413
rect 534 367 590 379
rect 620 607 676 619
rect 620 573 631 607
rect 665 573 676 607
rect 620 516 676 573
rect 620 482 631 516
rect 665 482 676 516
rect 620 428 676 482
rect 620 394 631 428
rect 665 394 676 428
rect 620 367 676 394
rect 706 599 762 619
rect 706 565 717 599
rect 751 565 762 599
rect 706 510 762 565
rect 706 476 717 510
rect 751 476 762 510
rect 706 413 762 476
rect 706 379 717 413
rect 751 379 762 413
rect 706 367 762 379
rect 792 607 848 619
rect 792 573 803 607
rect 837 573 848 607
rect 792 516 848 573
rect 792 482 803 516
rect 837 482 848 516
rect 792 428 848 482
rect 792 394 803 428
rect 837 394 848 428
rect 792 367 848 394
rect 878 599 934 619
rect 878 565 889 599
rect 923 565 934 599
rect 878 510 934 565
rect 878 476 889 510
rect 923 476 934 510
rect 878 413 934 476
rect 878 379 889 413
rect 923 379 934 413
rect 878 367 934 379
rect 964 607 1020 619
rect 964 573 975 607
rect 1009 573 1020 607
rect 964 516 1020 573
rect 964 482 975 516
rect 1009 482 1020 516
rect 964 428 1020 482
rect 964 394 975 428
rect 1009 394 1020 428
rect 964 367 1020 394
rect 1050 599 1106 619
rect 1050 565 1061 599
rect 1095 565 1106 599
rect 1050 510 1106 565
rect 1050 476 1061 510
rect 1095 476 1106 510
rect 1050 413 1106 476
rect 1050 379 1061 413
rect 1095 379 1106 413
rect 1050 367 1106 379
rect 1136 531 1192 619
rect 1136 497 1147 531
rect 1181 497 1192 531
rect 1136 413 1192 497
rect 1136 379 1147 413
rect 1181 379 1192 413
rect 1136 367 1192 379
rect 1222 597 1278 619
rect 1222 563 1233 597
rect 1267 563 1278 597
rect 1222 526 1278 563
rect 1222 492 1233 526
rect 1267 492 1278 526
rect 1222 455 1278 492
rect 1222 421 1233 455
rect 1267 421 1278 455
rect 1222 367 1278 421
rect 1308 531 1364 619
rect 1308 497 1319 531
rect 1353 497 1364 531
rect 1308 413 1364 497
rect 1308 379 1319 413
rect 1353 379 1364 413
rect 1308 367 1364 379
rect 1394 597 1450 619
rect 1394 563 1405 597
rect 1439 563 1450 597
rect 1394 526 1450 563
rect 1394 492 1405 526
rect 1439 492 1450 526
rect 1394 455 1450 492
rect 1394 421 1405 455
rect 1439 421 1450 455
rect 1394 367 1450 421
rect 1480 531 1536 619
rect 1480 497 1491 531
rect 1525 497 1536 531
rect 1480 413 1536 497
rect 1480 379 1491 413
rect 1525 379 1536 413
rect 1480 367 1536 379
rect 1566 597 1622 619
rect 1566 563 1577 597
rect 1611 563 1622 597
rect 1566 526 1622 563
rect 1566 492 1577 526
rect 1611 492 1622 526
rect 1566 455 1622 492
rect 1566 421 1577 455
rect 1611 421 1622 455
rect 1566 367 1622 421
rect 1652 531 1708 619
rect 1652 497 1663 531
rect 1697 497 1708 531
rect 1652 413 1708 497
rect 1652 379 1663 413
rect 1697 379 1708 413
rect 1652 367 1708 379
rect 1738 599 1791 619
rect 1738 565 1749 599
rect 1783 565 1791 599
rect 1738 506 1791 565
rect 1738 472 1749 506
rect 1783 472 1791 506
rect 1738 413 1791 472
rect 1738 379 1749 413
rect 1783 379 1791 413
rect 1738 367 1791 379
<< ndiffc >>
rect 127 158 161 192
rect 127 81 161 115
rect 213 191 247 225
rect 213 81 247 115
rect 379 169 413 203
rect 379 67 413 101
rect 465 173 499 207
rect 465 59 499 93
rect 551 169 585 203
rect 551 67 585 101
rect 637 173 671 207
rect 637 59 671 93
rect 723 169 757 203
rect 723 67 757 101
rect 809 173 843 207
rect 809 59 843 93
rect 895 169 929 203
rect 895 67 929 101
rect 981 158 1015 192
rect 981 55 1015 89
rect 1067 169 1101 203
rect 1067 59 1101 93
rect 1153 161 1187 195
rect 1239 71 1273 105
rect 1325 156 1359 190
rect 1411 71 1445 105
rect 1497 161 1531 195
rect 1583 131 1617 165
rect 1583 56 1617 90
rect 1669 139 1703 173
rect 1755 169 1789 203
rect 1755 71 1789 105
<< pdiffc >>
rect 107 573 141 607
rect 107 486 141 520
rect 107 400 141 434
rect 193 565 227 599
rect 373 565 407 599
rect 193 474 227 508
rect 193 387 227 421
rect 373 476 407 510
rect 373 379 407 413
rect 459 573 493 607
rect 459 482 493 516
rect 459 394 493 428
rect 545 565 579 599
rect 545 476 579 510
rect 545 379 579 413
rect 631 573 665 607
rect 631 482 665 516
rect 631 394 665 428
rect 717 565 751 599
rect 717 476 751 510
rect 717 379 751 413
rect 803 573 837 607
rect 803 482 837 516
rect 803 394 837 428
rect 889 565 923 599
rect 889 476 923 510
rect 889 379 923 413
rect 975 573 1009 607
rect 975 482 1009 516
rect 975 394 1009 428
rect 1061 565 1095 599
rect 1061 476 1095 510
rect 1061 379 1095 413
rect 1147 497 1181 531
rect 1147 379 1181 413
rect 1233 563 1267 597
rect 1233 492 1267 526
rect 1233 421 1267 455
rect 1319 497 1353 531
rect 1319 379 1353 413
rect 1405 563 1439 597
rect 1405 492 1439 526
rect 1405 421 1439 455
rect 1491 497 1525 531
rect 1491 379 1525 413
rect 1577 563 1611 597
rect 1577 492 1611 526
rect 1577 421 1611 455
rect 1663 497 1697 531
rect 1663 379 1697 413
rect 1749 565 1783 599
rect 1749 472 1783 506
rect 1749 379 1783 413
<< poly >>
rect 152 619 182 645
rect 418 619 448 645
rect 504 619 534 645
rect 590 619 620 645
rect 676 619 706 645
rect 762 619 792 645
rect 848 619 878 645
rect 934 619 964 645
rect 1020 619 1050 645
rect 1106 619 1136 645
rect 1192 619 1222 645
rect 1278 619 1308 645
rect 1364 619 1394 645
rect 1450 619 1480 645
rect 1536 619 1566 645
rect 1622 619 1652 645
rect 1708 619 1738 645
rect 267 504 333 520
rect 267 470 283 504
rect 317 470 333 504
rect 267 436 333 470
rect 267 402 283 436
rect 317 416 333 436
rect 317 402 350 416
rect 267 386 350 402
rect 152 325 182 367
rect 320 352 350 386
rect 418 352 448 367
rect 320 345 448 352
rect 504 345 534 367
rect 590 345 620 367
rect 676 345 706 367
rect 762 345 792 367
rect 848 345 878 367
rect 934 345 964 367
rect 1020 345 1050 367
rect 27 309 202 325
rect 320 322 1050 345
rect 418 315 1050 322
rect 1106 331 1136 367
rect 1192 331 1222 367
rect 1278 331 1308 367
rect 1364 331 1394 367
rect 1450 331 1480 367
rect 1536 331 1566 367
rect 1622 331 1652 367
rect 1708 331 1738 367
rect 1106 315 1744 331
rect 27 275 43 309
rect 77 275 111 309
rect 145 282 202 309
rect 145 275 300 282
rect 27 273 300 275
rect 1106 281 1275 315
rect 1309 281 1343 315
rect 1377 281 1411 315
rect 1445 281 1479 315
rect 1513 281 1547 315
rect 1581 281 1744 315
rect 27 259 1056 273
rect 1106 265 1744 281
rect 172 252 1056 259
rect 172 237 202 252
rect 270 243 1056 252
rect 319 237 1056 243
rect 424 215 454 237
rect 510 215 540 237
rect 596 215 626 237
rect 682 215 712 237
rect 768 215 798 237
rect 854 215 884 237
rect 940 215 970 237
rect 1026 215 1056 237
rect 1112 215 1142 265
rect 1198 215 1228 265
rect 1284 215 1314 265
rect 1370 215 1400 265
rect 1456 215 1486 265
rect 1542 215 1572 265
rect 1628 215 1658 265
rect 1714 215 1744 265
rect 172 43 202 69
rect 424 21 454 47
rect 510 21 540 47
rect 596 21 626 47
rect 682 21 712 47
rect 768 21 798 47
rect 854 21 884 47
rect 940 21 970 47
rect 1026 21 1056 47
rect 1112 21 1142 47
rect 1198 21 1228 47
rect 1284 21 1314 47
rect 1370 21 1400 47
rect 1456 21 1486 47
rect 1542 21 1572 47
rect 1628 21 1658 47
rect 1714 21 1744 47
<< polycont >>
rect 283 470 317 504
rect 283 402 317 436
rect 43 275 77 309
rect 111 275 145 309
rect 1275 281 1309 315
rect 1343 281 1377 315
rect 1411 281 1445 315
rect 1479 281 1513 315
rect 1547 281 1581 315
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 91 607 145 649
rect 91 573 107 607
rect 141 573 145 607
rect 91 520 145 573
rect 91 486 107 520
rect 141 486 145 520
rect 91 434 145 486
rect 91 400 107 434
rect 141 400 145 434
rect 91 384 145 400
rect 189 599 323 615
rect 189 565 193 599
rect 227 565 323 599
rect 189 508 323 565
rect 189 474 193 508
rect 227 504 323 508
rect 227 474 283 504
rect 189 470 283 474
rect 317 470 323 504
rect 189 436 323 470
rect 189 421 283 436
rect 189 387 193 421
rect 227 402 283 421
rect 317 402 323 436
rect 227 387 323 402
rect 189 386 323 387
rect 357 599 415 615
rect 357 565 373 599
rect 407 565 415 599
rect 357 510 415 565
rect 357 476 373 510
rect 407 476 415 510
rect 357 413 415 476
rect 189 371 263 386
rect 31 309 161 350
rect 31 275 43 309
rect 77 275 111 309
rect 145 275 161 309
rect 31 242 161 275
rect 205 225 263 371
rect 357 379 373 413
rect 407 379 415 413
rect 357 344 415 379
rect 449 607 501 649
rect 449 573 459 607
rect 493 573 501 607
rect 449 516 501 573
rect 449 482 459 516
rect 493 482 501 516
rect 449 428 501 482
rect 449 394 459 428
rect 493 394 501 428
rect 449 378 501 394
rect 535 599 587 615
rect 535 565 545 599
rect 579 565 587 599
rect 535 510 587 565
rect 535 476 545 510
rect 579 476 587 510
rect 535 413 587 476
rect 535 379 545 413
rect 579 379 587 413
rect 535 344 587 379
rect 621 607 674 649
rect 621 573 631 607
rect 665 573 674 607
rect 621 516 674 573
rect 621 482 631 516
rect 665 482 674 516
rect 621 428 674 482
rect 621 394 631 428
rect 665 394 674 428
rect 621 378 674 394
rect 708 599 760 615
rect 708 565 717 599
rect 751 565 760 599
rect 708 510 760 565
rect 708 476 717 510
rect 751 476 760 510
rect 708 413 760 476
rect 708 379 717 413
rect 751 379 760 413
rect 708 344 760 379
rect 794 607 845 649
rect 794 573 803 607
rect 837 573 845 607
rect 794 516 845 573
rect 794 482 803 516
rect 837 482 845 516
rect 794 428 845 482
rect 794 394 803 428
rect 837 394 845 428
rect 794 378 845 394
rect 879 599 932 615
rect 879 565 889 599
rect 923 565 932 599
rect 879 510 932 565
rect 879 476 889 510
rect 923 476 932 510
rect 879 413 932 476
rect 879 379 889 413
rect 923 379 932 413
rect 879 344 932 379
rect 966 607 1018 649
rect 966 573 975 607
rect 1009 573 1018 607
rect 966 516 1018 573
rect 966 482 975 516
rect 1009 482 1018 516
rect 966 428 1018 482
rect 966 394 975 428
rect 1009 394 1018 428
rect 966 378 1018 394
rect 1052 599 1799 615
rect 1052 565 1061 599
rect 1095 597 1749 599
rect 1095 581 1233 597
rect 1095 565 1103 581
rect 1052 510 1103 565
rect 1217 563 1233 581
rect 1267 581 1405 597
rect 1267 563 1283 581
rect 1052 476 1061 510
rect 1095 476 1103 510
rect 1052 413 1103 476
rect 1052 379 1061 413
rect 1095 379 1103 413
rect 1052 344 1103 379
rect 357 310 1103 344
rect 1137 531 1183 547
rect 1137 497 1147 531
rect 1181 497 1183 531
rect 1137 413 1183 497
rect 1217 526 1283 563
rect 1389 563 1405 581
rect 1439 581 1577 597
rect 1439 563 1455 581
rect 1217 492 1233 526
rect 1267 492 1283 526
rect 1217 455 1283 492
rect 1217 421 1233 455
rect 1267 421 1283 455
rect 1317 531 1355 547
rect 1317 497 1319 531
rect 1353 497 1355 531
rect 1137 379 1147 413
rect 1181 387 1183 413
rect 1317 413 1355 497
rect 1389 526 1455 563
rect 1561 563 1577 581
rect 1611 581 1749 597
rect 1611 563 1627 581
rect 1389 492 1405 526
rect 1439 492 1455 526
rect 1389 455 1455 492
rect 1389 421 1405 455
rect 1439 421 1455 455
rect 1489 531 1527 547
rect 1489 497 1491 531
rect 1525 497 1527 531
rect 1317 387 1319 413
rect 1181 379 1319 387
rect 1353 387 1355 413
rect 1489 413 1527 497
rect 1561 526 1627 563
rect 1741 565 1749 581
rect 1783 565 1799 599
rect 1561 492 1577 526
rect 1611 492 1627 526
rect 1561 455 1627 492
rect 1561 421 1577 455
rect 1611 421 1627 455
rect 1661 531 1707 547
rect 1661 497 1663 531
rect 1697 497 1707 531
rect 1489 387 1491 413
rect 1353 379 1491 387
rect 1525 387 1527 413
rect 1661 413 1707 497
rect 1661 387 1663 413
rect 1525 379 1663 387
rect 1697 379 1707 413
rect 1137 353 1707 379
rect 1741 506 1799 565
rect 1741 472 1749 506
rect 1783 472 1799 506
rect 1741 413 1799 472
rect 1741 379 1749 413
rect 1783 379 1799 413
rect 1741 363 1799 379
rect 1137 305 1225 353
rect 111 192 171 208
rect 111 158 127 192
rect 161 158 171 192
rect 111 115 171 158
rect 111 81 127 115
rect 161 81 171 115
rect 111 17 171 81
rect 205 191 213 225
rect 247 191 263 225
rect 205 115 263 191
rect 205 81 213 115
rect 247 81 263 115
rect 205 51 263 81
rect 363 242 1117 276
rect 363 203 415 242
rect 363 169 379 203
rect 413 169 415 203
rect 363 101 415 169
rect 363 67 379 101
rect 413 67 415 101
rect 363 51 415 67
rect 449 207 515 208
rect 449 173 465 207
rect 499 173 515 207
rect 449 93 515 173
rect 449 59 465 93
rect 499 59 515 93
rect 449 17 515 59
rect 549 203 587 242
rect 549 169 551 203
rect 585 169 587 203
rect 549 101 587 169
rect 549 67 551 101
rect 585 67 587 101
rect 549 51 587 67
rect 621 207 687 208
rect 621 173 637 207
rect 671 173 687 207
rect 621 93 687 173
rect 621 59 637 93
rect 671 59 687 93
rect 621 17 687 59
rect 721 203 759 242
rect 721 169 723 203
rect 757 169 759 203
rect 721 101 759 169
rect 721 67 723 101
rect 757 67 759 101
rect 721 51 759 67
rect 793 207 859 208
rect 793 173 809 207
rect 843 173 859 207
rect 793 93 859 173
rect 793 59 809 93
rect 843 59 859 93
rect 793 17 859 59
rect 893 203 937 242
rect 893 169 895 203
rect 929 169 937 203
rect 893 101 937 169
rect 893 67 895 101
rect 929 67 937 101
rect 893 51 937 67
rect 971 192 1017 208
rect 971 158 981 192
rect 1015 158 1017 192
rect 971 89 1017 158
rect 971 55 981 89
rect 1015 55 1017 89
rect 1051 203 1117 242
rect 1051 169 1067 203
rect 1101 169 1117 203
rect 1051 111 1117 169
rect 1151 199 1225 305
rect 1259 315 1597 319
rect 1259 281 1275 315
rect 1309 281 1343 315
rect 1377 281 1411 315
rect 1445 281 1479 315
rect 1513 281 1547 315
rect 1581 281 1597 315
rect 1259 269 1597 281
rect 1259 242 1449 269
rect 1631 235 1707 353
rect 1483 201 1712 235
rect 1483 199 1533 201
rect 1151 195 1533 199
rect 1151 161 1153 195
rect 1187 190 1497 195
rect 1187 161 1325 190
rect 1151 156 1325 161
rect 1359 161 1497 190
rect 1531 161 1533 195
rect 1667 173 1712 201
rect 1359 156 1533 161
rect 1151 145 1533 156
rect 1567 131 1583 165
rect 1617 131 1633 165
rect 1567 111 1633 131
rect 1667 139 1669 173
rect 1703 139 1712 173
rect 1667 123 1712 139
rect 1746 203 1805 219
rect 1746 169 1755 203
rect 1789 169 1805 203
rect 1051 105 1633 111
rect 1051 93 1239 105
rect 1051 59 1067 93
rect 1101 71 1239 93
rect 1273 71 1411 105
rect 1445 90 1633 105
rect 1445 71 1583 90
rect 1101 59 1583 71
rect 1051 56 1583 59
rect 1617 89 1633 90
rect 1746 105 1805 169
rect 1746 89 1755 105
rect 1617 71 1755 89
rect 1789 71 1805 105
rect 1617 56 1805 71
rect 1051 55 1805 56
rect 971 17 1017 55
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
<< metal1 >>
rect 0 683 1824 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1824 683
rect 0 617 1824 649
rect 0 17 1824 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1824 17
rect 0 -49 1824 -17
<< labels >>
flabel pwell s 0 0 1824 49 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 0 617 1824 666 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 einvp_8
flabel metal1 s 0 617 1824 666 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 0 1824 49 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel locali s 1183 168 1217 202 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 1824 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 3037230
string GDS_START 3023296
<< end >>
