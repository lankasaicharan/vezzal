magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 3314 1975
<< nwell >>
rect -38 331 2054 704
<< pwell >>
rect 1 49 1988 241
rect 0 0 2016 49
<< scnmos >>
rect 80 47 110 215
rect 166 47 196 215
rect 252 47 282 215
rect 338 47 368 215
rect 424 47 454 215
rect 510 47 540 215
rect 596 47 626 215
rect 682 47 712 215
rect 790 47 820 215
rect 876 47 906 215
rect 962 47 992 215
rect 1048 47 1078 215
rect 1258 47 1288 215
rect 1344 47 1374 215
rect 1430 47 1460 215
rect 1516 47 1546 215
rect 1621 47 1651 215
rect 1707 47 1737 215
rect 1793 47 1823 215
rect 1879 47 1909 215
<< scpmoshvt >>
rect 80 367 110 619
rect 166 367 196 619
rect 252 367 282 619
rect 338 367 368 619
rect 424 367 454 619
rect 510 367 540 619
rect 596 367 626 619
rect 682 367 712 619
rect 872 367 902 619
rect 958 367 988 619
rect 1044 367 1074 619
rect 1130 367 1160 619
rect 1216 367 1246 619
rect 1302 367 1332 619
rect 1388 367 1418 619
rect 1478 367 1508 619
rect 1588 367 1618 619
rect 1674 367 1704 619
rect 1778 367 1808 619
rect 1864 367 1894 619
<< ndiff >>
rect 27 132 80 215
rect 27 98 35 132
rect 69 98 80 132
rect 27 47 80 98
rect 110 190 166 215
rect 110 156 121 190
rect 155 156 166 190
rect 110 101 166 156
rect 110 67 121 101
rect 155 67 166 101
rect 110 47 166 67
rect 196 132 252 215
rect 196 98 207 132
rect 241 98 252 132
rect 196 47 252 98
rect 282 190 338 215
rect 282 156 293 190
rect 327 156 338 190
rect 282 101 338 156
rect 282 67 293 101
rect 327 67 338 101
rect 282 47 338 67
rect 368 132 424 215
rect 368 98 379 132
rect 413 98 424 132
rect 368 47 424 98
rect 454 202 510 215
rect 454 168 465 202
rect 499 168 510 202
rect 454 101 510 168
rect 454 67 465 101
rect 499 67 510 101
rect 454 47 510 67
rect 540 183 596 215
rect 540 149 551 183
rect 585 149 596 183
rect 540 93 596 149
rect 540 59 551 93
rect 585 59 596 93
rect 540 47 596 59
rect 626 202 682 215
rect 626 168 637 202
rect 671 168 682 202
rect 626 101 682 168
rect 626 67 637 101
rect 671 67 682 101
rect 626 47 682 67
rect 712 183 790 215
rect 712 149 735 183
rect 769 149 790 183
rect 712 93 790 149
rect 712 59 735 93
rect 769 59 790 93
rect 712 47 790 59
rect 820 202 876 215
rect 820 168 831 202
rect 865 168 876 202
rect 820 101 876 168
rect 820 67 831 101
rect 865 67 876 101
rect 820 47 876 67
rect 906 167 962 215
rect 906 133 917 167
rect 951 133 962 167
rect 906 93 962 133
rect 906 59 917 93
rect 951 59 962 93
rect 906 47 962 59
rect 992 203 1048 215
rect 992 169 1003 203
rect 1037 169 1048 203
rect 992 101 1048 169
rect 992 67 1003 101
rect 1037 67 1048 101
rect 992 47 1048 67
rect 1078 130 1131 215
rect 1078 96 1089 130
rect 1123 96 1131 130
rect 1078 47 1131 96
rect 1201 124 1258 215
rect 1201 90 1209 124
rect 1243 90 1258 124
rect 1201 47 1258 90
rect 1288 169 1344 215
rect 1288 135 1299 169
rect 1333 135 1344 169
rect 1288 47 1344 135
rect 1374 124 1430 215
rect 1374 90 1385 124
rect 1419 90 1430 124
rect 1374 47 1430 90
rect 1460 169 1516 215
rect 1460 135 1471 169
rect 1505 135 1516 169
rect 1460 47 1516 135
rect 1546 203 1621 215
rect 1546 169 1575 203
rect 1609 169 1621 203
rect 1546 101 1621 169
rect 1546 67 1575 101
rect 1609 67 1621 101
rect 1546 47 1621 67
rect 1651 173 1707 215
rect 1651 139 1662 173
rect 1696 139 1707 173
rect 1651 93 1707 139
rect 1651 59 1662 93
rect 1696 59 1707 93
rect 1651 47 1707 59
rect 1737 203 1793 215
rect 1737 169 1748 203
rect 1782 169 1793 203
rect 1737 101 1793 169
rect 1737 67 1748 101
rect 1782 67 1793 101
rect 1737 47 1793 67
rect 1823 173 1879 215
rect 1823 139 1834 173
rect 1868 139 1879 173
rect 1823 93 1879 139
rect 1823 59 1834 93
rect 1868 59 1879 93
rect 1823 47 1879 59
rect 1909 203 1962 215
rect 1909 169 1920 203
rect 1954 169 1962 203
rect 1909 101 1962 169
rect 1909 67 1920 101
rect 1954 67 1962 101
rect 1909 47 1962 67
<< pdiff >>
rect 27 607 80 619
rect 27 573 35 607
rect 69 573 80 607
rect 27 523 80 573
rect 27 489 35 523
rect 69 489 80 523
rect 27 443 80 489
rect 27 409 35 443
rect 69 409 80 443
rect 27 367 80 409
rect 110 531 166 619
rect 110 497 121 531
rect 155 497 166 531
rect 110 413 166 497
rect 110 379 121 413
rect 155 379 166 413
rect 110 367 166 379
rect 196 597 252 619
rect 196 563 207 597
rect 241 563 252 597
rect 196 523 252 563
rect 196 489 207 523
rect 241 489 252 523
rect 196 443 252 489
rect 196 409 207 443
rect 241 409 252 443
rect 196 367 252 409
rect 282 531 338 619
rect 282 497 293 531
rect 327 497 338 531
rect 282 413 338 497
rect 282 379 293 413
rect 327 379 338 413
rect 282 367 338 379
rect 368 597 424 619
rect 368 563 379 597
rect 413 563 424 597
rect 368 507 424 563
rect 368 473 379 507
rect 413 473 424 507
rect 368 420 424 473
rect 368 386 379 420
rect 413 386 424 420
rect 368 367 424 386
rect 454 531 510 619
rect 454 497 465 531
rect 499 497 510 531
rect 454 436 510 497
rect 454 402 465 436
rect 499 402 510 436
rect 454 367 510 402
rect 540 597 596 619
rect 540 563 551 597
rect 585 563 596 597
rect 540 494 596 563
rect 540 460 551 494
rect 585 460 596 494
rect 540 367 596 460
rect 626 531 682 619
rect 626 497 637 531
rect 671 497 682 531
rect 626 436 682 497
rect 626 402 637 436
rect 671 402 682 436
rect 626 367 682 402
rect 712 594 765 619
rect 712 560 723 594
rect 757 560 765 594
rect 712 494 765 560
rect 712 460 723 494
rect 757 460 765 494
rect 712 367 765 460
rect 819 596 872 619
rect 819 562 827 596
rect 861 562 872 596
rect 819 494 872 562
rect 819 460 827 494
rect 861 460 872 494
rect 819 367 872 460
rect 902 531 958 619
rect 902 497 913 531
rect 947 497 958 531
rect 902 436 958 497
rect 902 402 913 436
rect 947 402 958 436
rect 902 367 958 402
rect 988 605 1044 619
rect 988 571 999 605
rect 1033 571 1044 605
rect 988 511 1044 571
rect 988 477 999 511
rect 1033 477 1044 511
rect 988 367 1044 477
rect 1074 539 1130 619
rect 1074 505 1085 539
rect 1119 505 1130 539
rect 1074 436 1130 505
rect 1074 402 1085 436
rect 1119 402 1130 436
rect 1074 367 1130 402
rect 1160 599 1216 619
rect 1160 565 1171 599
rect 1205 565 1216 599
rect 1160 507 1216 565
rect 1160 473 1171 507
rect 1205 473 1216 507
rect 1160 413 1216 473
rect 1160 379 1171 413
rect 1205 379 1216 413
rect 1160 367 1216 379
rect 1246 607 1302 619
rect 1246 573 1257 607
rect 1291 573 1302 607
rect 1246 517 1302 573
rect 1246 483 1257 517
rect 1291 483 1302 517
rect 1246 423 1302 483
rect 1246 389 1257 423
rect 1291 389 1302 423
rect 1246 367 1302 389
rect 1332 599 1388 619
rect 1332 565 1343 599
rect 1377 565 1388 599
rect 1332 507 1388 565
rect 1332 473 1343 507
rect 1377 473 1388 507
rect 1332 413 1388 473
rect 1332 379 1343 413
rect 1377 379 1388 413
rect 1332 367 1388 379
rect 1418 607 1478 619
rect 1418 573 1429 607
rect 1463 573 1478 607
rect 1418 517 1478 573
rect 1418 483 1429 517
rect 1463 483 1478 517
rect 1418 423 1478 483
rect 1418 389 1429 423
rect 1463 389 1478 423
rect 1418 367 1478 389
rect 1508 611 1588 619
rect 1508 577 1529 611
rect 1563 577 1588 611
rect 1508 512 1588 577
rect 1508 478 1529 512
rect 1563 478 1588 512
rect 1508 413 1588 478
rect 1508 379 1519 413
rect 1553 379 1588 413
rect 1508 367 1588 379
rect 1618 607 1674 619
rect 1618 573 1629 607
rect 1663 573 1674 607
rect 1618 493 1674 573
rect 1618 459 1629 493
rect 1663 459 1674 493
rect 1618 367 1674 459
rect 1704 599 1778 619
rect 1704 565 1724 599
rect 1758 565 1778 599
rect 1704 508 1778 565
rect 1704 474 1724 508
rect 1758 474 1778 508
rect 1704 413 1778 474
rect 1704 379 1733 413
rect 1767 379 1778 413
rect 1704 367 1778 379
rect 1808 607 1864 619
rect 1808 573 1819 607
rect 1853 573 1864 607
rect 1808 525 1864 573
rect 1808 491 1819 525
rect 1853 491 1864 525
rect 1808 445 1864 491
rect 1808 411 1819 445
rect 1853 411 1864 445
rect 1808 367 1864 411
rect 1894 599 1947 619
rect 1894 565 1905 599
rect 1939 565 1947 599
rect 1894 506 1947 565
rect 1894 472 1905 506
rect 1939 472 1947 506
rect 1894 413 1947 472
rect 1894 379 1905 413
rect 1939 379 1947 413
rect 1894 367 1947 379
<< ndiffc >>
rect 35 98 69 132
rect 121 156 155 190
rect 121 67 155 101
rect 207 98 241 132
rect 293 156 327 190
rect 293 67 327 101
rect 379 98 413 132
rect 465 168 499 202
rect 465 67 499 101
rect 551 149 585 183
rect 551 59 585 93
rect 637 168 671 202
rect 637 67 671 101
rect 735 149 769 183
rect 735 59 769 93
rect 831 168 865 202
rect 831 67 865 101
rect 917 133 951 167
rect 917 59 951 93
rect 1003 169 1037 203
rect 1003 67 1037 101
rect 1089 96 1123 130
rect 1209 90 1243 124
rect 1299 135 1333 169
rect 1385 90 1419 124
rect 1471 135 1505 169
rect 1575 169 1609 203
rect 1575 67 1609 101
rect 1662 139 1696 173
rect 1662 59 1696 93
rect 1748 169 1782 203
rect 1748 67 1782 101
rect 1834 139 1868 173
rect 1834 59 1868 93
rect 1920 169 1954 203
rect 1920 67 1954 101
<< pdiffc >>
rect 35 573 69 607
rect 35 489 69 523
rect 35 409 69 443
rect 121 497 155 531
rect 121 379 155 413
rect 207 563 241 597
rect 207 489 241 523
rect 207 409 241 443
rect 293 497 327 531
rect 293 379 327 413
rect 379 563 413 597
rect 379 473 413 507
rect 379 386 413 420
rect 465 497 499 531
rect 465 402 499 436
rect 551 563 585 597
rect 551 460 585 494
rect 637 497 671 531
rect 637 402 671 436
rect 723 560 757 594
rect 723 460 757 494
rect 827 562 861 596
rect 827 460 861 494
rect 913 497 947 531
rect 913 402 947 436
rect 999 571 1033 605
rect 999 477 1033 511
rect 1085 505 1119 539
rect 1085 402 1119 436
rect 1171 565 1205 599
rect 1171 473 1205 507
rect 1171 379 1205 413
rect 1257 573 1291 607
rect 1257 483 1291 517
rect 1257 389 1291 423
rect 1343 565 1377 599
rect 1343 473 1377 507
rect 1343 379 1377 413
rect 1429 573 1463 607
rect 1429 483 1463 517
rect 1429 389 1463 423
rect 1529 577 1563 611
rect 1529 478 1563 512
rect 1519 379 1553 413
rect 1629 573 1663 607
rect 1629 459 1663 493
rect 1724 565 1758 599
rect 1724 474 1758 508
rect 1733 379 1767 413
rect 1819 573 1853 607
rect 1819 491 1853 525
rect 1819 411 1853 445
rect 1905 565 1939 599
rect 1905 472 1939 506
rect 1905 379 1939 413
<< poly >>
rect 80 619 110 645
rect 166 619 196 645
rect 252 619 282 645
rect 338 619 368 645
rect 424 619 454 645
rect 510 619 540 645
rect 596 619 626 645
rect 682 619 712 645
rect 872 619 902 645
rect 958 619 988 645
rect 1044 619 1074 645
rect 1130 619 1160 645
rect 1216 619 1246 645
rect 1302 619 1332 645
rect 1388 619 1418 645
rect 1478 619 1508 645
rect 1588 619 1618 645
rect 1674 619 1704 645
rect 1778 619 1808 645
rect 1864 619 1894 645
rect 80 303 110 367
rect 166 303 196 367
rect 252 303 282 367
rect 338 303 368 367
rect 424 335 454 367
rect 510 335 540 367
rect 596 335 626 367
rect 682 335 712 367
rect 872 335 902 367
rect 958 335 988 367
rect 1044 335 1074 367
rect 1130 335 1160 367
rect 80 287 368 303
rect 80 253 114 287
rect 148 253 182 287
rect 216 253 250 287
rect 284 253 318 287
rect 352 253 368 287
rect 410 319 748 335
rect 410 285 426 319
rect 460 285 494 319
rect 528 285 562 319
rect 596 285 630 319
rect 664 285 698 319
rect 732 285 748 319
rect 410 269 748 285
rect 790 319 1160 335
rect 790 285 806 319
rect 840 285 874 319
rect 908 285 942 319
rect 976 285 1010 319
rect 1044 285 1078 319
rect 1112 305 1160 319
rect 1112 285 1128 305
rect 1216 303 1246 367
rect 1302 303 1332 367
rect 1388 303 1418 367
rect 1478 303 1508 367
rect 1588 325 1618 367
rect 1674 325 1704 367
rect 1778 325 1808 367
rect 1864 325 1894 367
rect 1588 309 1995 325
rect 790 269 1128 285
rect 1202 287 1546 303
rect 80 237 368 253
rect 80 215 110 237
rect 166 215 196 237
rect 252 215 282 237
rect 338 215 368 237
rect 424 215 454 269
rect 510 215 540 269
rect 596 215 626 269
rect 682 215 712 269
rect 790 215 820 269
rect 876 215 906 269
rect 962 215 992 269
rect 1048 215 1078 269
rect 1202 253 1218 287
rect 1252 253 1286 287
rect 1320 253 1354 287
rect 1388 253 1422 287
rect 1456 253 1490 287
rect 1524 253 1546 287
rect 1588 275 1605 309
rect 1639 275 1673 309
rect 1707 275 1741 309
rect 1775 275 1809 309
rect 1843 275 1877 309
rect 1911 275 1945 309
rect 1979 275 1995 309
rect 1588 259 1995 275
rect 1202 237 1546 253
rect 1258 215 1288 237
rect 1344 215 1374 237
rect 1430 215 1460 237
rect 1516 215 1546 237
rect 1621 215 1651 259
rect 1707 215 1737 259
rect 1793 215 1823 259
rect 1879 215 1909 259
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 424 21 454 47
rect 510 21 540 47
rect 596 21 626 47
rect 682 21 712 47
rect 790 21 820 47
rect 876 21 906 47
rect 962 21 992 47
rect 1048 21 1078 47
rect 1258 21 1288 47
rect 1344 21 1374 47
rect 1430 21 1460 47
rect 1516 21 1546 47
rect 1621 21 1651 47
rect 1707 21 1737 47
rect 1793 21 1823 47
rect 1879 21 1909 47
<< polycont >>
rect 114 253 148 287
rect 182 253 216 287
rect 250 253 284 287
rect 318 253 352 287
rect 426 285 460 319
rect 494 285 528 319
rect 562 285 596 319
rect 630 285 664 319
rect 698 285 732 319
rect 806 285 840 319
rect 874 285 908 319
rect 942 285 976 319
rect 1010 285 1044 319
rect 1078 285 1112 319
rect 1218 253 1252 287
rect 1286 253 1320 287
rect 1354 253 1388 287
rect 1422 253 1456 287
rect 1490 253 1524 287
rect 1605 275 1639 309
rect 1673 275 1707 309
rect 1741 275 1775 309
rect 1809 275 1843 309
rect 1877 275 1911 309
rect 1945 275 1979 309
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 19 607 773 615
rect 19 573 35 607
rect 69 597 773 607
rect 69 581 207 597
rect 69 573 85 581
rect 19 523 85 573
rect 191 563 207 581
rect 241 581 379 597
rect 241 563 257 581
rect 19 489 35 523
rect 69 489 85 523
rect 19 443 85 489
rect 19 409 35 443
rect 69 409 85 443
rect 119 531 157 547
rect 119 497 121 531
rect 155 497 157 531
rect 119 413 157 497
rect 119 379 121 413
rect 155 379 157 413
rect 191 523 257 563
rect 363 563 379 581
rect 413 581 551 597
rect 413 563 429 581
rect 191 489 207 523
rect 241 489 257 523
rect 191 443 257 489
rect 191 409 207 443
rect 241 409 257 443
rect 291 531 329 547
rect 291 497 293 531
rect 327 497 329 531
rect 291 413 329 497
rect 119 375 157 379
rect 291 379 293 413
rect 327 379 329 413
rect 363 507 429 563
rect 535 563 551 581
rect 585 594 773 597
rect 585 581 723 594
rect 585 563 601 581
rect 363 473 379 507
rect 413 473 429 507
rect 363 420 429 473
rect 363 386 379 420
rect 413 386 429 420
rect 463 531 501 547
rect 463 497 465 531
rect 499 497 501 531
rect 463 436 501 497
rect 535 494 601 563
rect 707 560 723 581
rect 757 560 773 594
rect 535 460 551 494
rect 585 460 601 494
rect 535 454 601 460
rect 635 531 673 547
rect 635 497 637 531
rect 671 497 673 531
rect 463 402 465 436
rect 499 420 501 436
rect 635 436 673 497
rect 707 494 773 560
rect 707 460 723 494
rect 757 460 773 494
rect 707 454 773 460
rect 811 605 1207 615
rect 811 596 999 605
rect 811 562 827 596
rect 861 581 999 596
rect 861 562 877 581
rect 811 494 877 562
rect 991 571 999 581
rect 1033 599 1207 605
rect 1033 581 1171 599
rect 1033 571 1035 581
rect 811 460 827 494
rect 861 460 877 494
rect 811 454 877 460
rect 911 531 957 547
rect 911 497 913 531
rect 947 497 957 531
rect 635 420 637 436
rect 499 402 637 420
rect 671 420 673 436
rect 911 436 957 497
rect 991 511 1035 571
rect 1169 565 1171 581
rect 1205 565 1207 599
rect 991 477 999 511
rect 1033 477 1035 511
rect 991 461 1035 477
rect 1069 539 1135 547
rect 1069 505 1085 539
rect 1119 505 1135 539
rect 911 420 913 436
rect 671 402 913 420
rect 947 424 957 436
rect 1069 436 1135 505
rect 1069 424 1085 436
rect 947 402 1085 424
rect 1119 402 1135 436
rect 463 386 1135 402
rect 1169 507 1207 565
rect 1169 473 1171 507
rect 1205 473 1207 507
rect 1169 413 1207 473
rect 291 375 329 379
rect 28 341 329 375
rect 1169 379 1171 413
rect 1205 379 1207 413
rect 1241 607 1307 649
rect 1241 573 1257 607
rect 1291 573 1307 607
rect 1241 517 1307 573
rect 1241 483 1257 517
rect 1291 483 1307 517
rect 1241 423 1307 483
rect 1241 389 1257 423
rect 1291 389 1307 423
rect 1341 599 1379 615
rect 1341 565 1343 599
rect 1377 565 1379 599
rect 1341 507 1379 565
rect 1341 473 1343 507
rect 1377 473 1379 507
rect 1341 413 1379 473
rect 1169 355 1207 379
rect 1341 379 1343 413
rect 1377 379 1379 413
rect 1413 607 1479 649
rect 1413 573 1429 607
rect 1463 573 1479 607
rect 1413 517 1479 573
rect 1413 483 1429 517
rect 1463 483 1479 517
rect 1413 423 1479 483
rect 1413 389 1429 423
rect 1463 389 1479 423
rect 1513 611 1579 615
rect 1513 577 1529 611
rect 1563 577 1579 611
rect 1513 512 1579 577
rect 1513 478 1529 512
rect 1563 478 1579 512
rect 1513 420 1579 478
rect 1613 607 1679 649
rect 1613 573 1629 607
rect 1663 573 1679 607
rect 1613 493 1679 573
rect 1613 459 1629 493
rect 1663 459 1679 493
rect 1613 454 1679 459
rect 1713 599 1769 615
rect 1713 565 1724 599
rect 1758 565 1769 599
rect 1713 508 1769 565
rect 1713 474 1724 508
rect 1758 474 1769 508
rect 1713 420 1769 474
rect 1513 413 1769 420
rect 1341 355 1379 379
rect 1513 379 1519 413
rect 1553 386 1733 413
rect 1553 379 1555 386
rect 1513 355 1555 379
rect 28 208 64 341
rect 410 319 748 352
rect 98 253 114 287
rect 148 253 182 287
rect 216 253 250 287
rect 284 253 318 287
rect 352 253 368 287
rect 410 285 426 319
rect 460 285 494 319
rect 528 285 562 319
rect 596 285 630 319
rect 664 285 698 319
rect 732 285 748 319
rect 790 319 1135 352
rect 1169 321 1555 355
rect 1731 379 1733 386
rect 1767 379 1769 413
rect 1803 607 1869 649
rect 1803 573 1819 607
rect 1853 573 1869 607
rect 1803 525 1869 573
rect 1803 491 1819 525
rect 1853 491 1869 525
rect 1803 445 1869 491
rect 1803 411 1819 445
rect 1853 411 1869 445
rect 1903 599 1955 615
rect 1903 565 1905 599
rect 1939 565 1955 599
rect 1903 506 1955 565
rect 1903 472 1905 506
rect 1939 472 1955 506
rect 1903 413 1955 472
rect 1731 377 1769 379
rect 1903 379 1905 413
rect 1939 379 1955 413
rect 1903 377 1955 379
rect 790 285 806 319
rect 840 285 874 319
rect 908 285 942 319
rect 976 285 1010 319
rect 1044 285 1078 319
rect 1112 285 1135 319
rect 1589 309 1697 352
rect 1731 343 1955 377
rect 98 242 368 253
rect 1169 253 1218 287
rect 1252 253 1286 287
rect 1320 253 1354 287
rect 1388 253 1422 287
rect 1456 253 1490 287
rect 1524 253 1540 287
rect 1589 275 1605 309
rect 1639 275 1673 309
rect 1707 275 1741 309
rect 1775 275 1809 309
rect 1843 275 1877 309
rect 1911 275 1945 309
rect 1979 275 1995 309
rect 461 217 1037 251
rect 1169 242 1540 253
rect 461 208 501 217
rect 28 202 501 208
rect 28 190 465 202
rect 28 174 121 190
rect 119 156 121 174
rect 155 174 293 190
rect 155 156 157 174
rect 19 132 85 140
rect 19 98 35 132
rect 69 98 85 132
rect 19 17 85 98
rect 119 101 157 156
rect 291 156 293 174
rect 327 174 465 190
rect 327 156 329 174
rect 119 67 121 101
rect 155 67 157 101
rect 119 51 157 67
rect 191 132 257 140
rect 191 98 207 132
rect 241 98 257 132
rect 191 17 257 98
rect 291 101 329 156
rect 463 168 465 174
rect 499 168 501 202
rect 635 202 685 217
rect 291 67 293 101
rect 327 67 329 101
rect 291 51 329 67
rect 363 132 429 140
rect 363 98 379 132
rect 413 98 429 132
rect 363 17 429 98
rect 463 101 501 168
rect 463 67 465 101
rect 499 67 501 101
rect 463 51 501 67
rect 535 149 551 183
rect 585 149 601 183
rect 535 93 601 149
rect 535 59 551 93
rect 585 59 601 93
rect 535 17 601 59
rect 635 168 637 202
rect 671 168 685 202
rect 819 202 867 217
rect 635 101 685 168
rect 635 67 637 101
rect 671 67 685 101
rect 635 51 685 67
rect 719 149 735 183
rect 769 149 785 183
rect 719 93 785 149
rect 719 59 735 93
rect 769 59 785 93
rect 719 17 785 59
rect 819 168 831 202
rect 865 168 867 202
rect 989 208 1037 217
rect 989 203 1521 208
rect 819 101 867 168
rect 819 67 831 101
rect 865 67 867 101
rect 819 51 867 67
rect 901 167 955 183
rect 901 133 917 167
rect 951 133 955 167
rect 901 93 955 133
rect 901 59 917 93
rect 951 59 955 93
rect 901 17 955 59
rect 989 169 1003 203
rect 1037 174 1521 203
rect 1037 169 1039 174
rect 989 101 1039 169
rect 1292 169 1341 174
rect 989 67 1003 101
rect 1037 67 1039 101
rect 989 51 1039 67
rect 1073 130 1139 138
rect 1073 96 1089 130
rect 1123 96 1139 130
rect 1073 17 1139 96
rect 1193 124 1258 140
rect 1193 90 1209 124
rect 1243 90 1258 124
rect 1292 135 1299 169
rect 1333 135 1341 169
rect 1462 169 1521 174
rect 1292 119 1341 135
rect 1375 124 1428 140
rect 1193 85 1258 90
rect 1375 90 1385 124
rect 1419 90 1428 124
rect 1462 135 1471 169
rect 1505 135 1521 169
rect 1462 119 1521 135
rect 1574 207 1970 241
rect 1574 203 1612 207
rect 1574 169 1575 203
rect 1609 169 1612 203
rect 1746 203 1784 207
rect 1375 85 1428 90
rect 1574 101 1612 169
rect 1574 85 1575 101
rect 1193 67 1575 85
rect 1609 67 1612 101
rect 1193 51 1612 67
rect 1646 139 1662 173
rect 1696 139 1712 173
rect 1646 93 1712 139
rect 1646 59 1662 93
rect 1696 59 1712 93
rect 1646 17 1712 59
rect 1746 169 1748 203
rect 1782 169 1784 203
rect 1918 203 1970 207
rect 1746 101 1784 169
rect 1746 67 1748 101
rect 1782 67 1784 101
rect 1746 51 1784 67
rect 1818 139 1834 173
rect 1868 139 1884 173
rect 1818 93 1884 139
rect 1818 59 1834 93
rect 1868 59 1884 93
rect 1818 17 1884 59
rect 1918 169 1920 203
rect 1954 169 1970 203
rect 1918 101 1970 169
rect 1918 67 1920 101
rect 1954 67 1970 101
rect 1918 51 1970 67
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
<< metal1 >>
rect 0 683 2016 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2016 683
rect 0 617 2016 649
rect 0 17 2016 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2016 17
rect 0 -49 2016 -17
<< labels >>
flabel pwell s 0 0 2016 49 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 0 617 2016 666 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a2111oi_4
flabel metal1 s 0 617 2016 666 0 FreeSans 340 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal1 s 0 0 2016 49 0 FreeSans 340 0 0 0 VGND
port 6 nsew ground bidirectional
flabel locali s 991 94 1025 128 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 991 168 1025 202 0 FreeSans 340 0 0 0 Y
port 10 nsew signal output
flabel locali s 1183 242 1217 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1279 242 1313 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1375 242 1409 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1471 242 1505 276 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1663 316 1697 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 1087 316 1121 350 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 223 242 257 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2016 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 4842404
string GDS_START 4824888
<< end >>
