magic
tech sky130A
magscale 1 2
timestamp 1627202642
<< checkpaint >>
rect -1298 -1309 4082 1975
<< nwell >>
rect -38 331 2822 704
<< pwell >>
rect 782 223 1697 235
rect 263 176 1697 223
rect 263 167 1877 176
rect 1 49 2783 167
rect 0 0 2784 49
<< scnmos >>
rect 80 57 110 141
rect 152 57 182 141
rect 343 113 373 197
rect 415 113 445 197
rect 501 113 531 197
rect 573 113 603 197
rect 763 89 793 173
rect 874 125 904 209
rect 946 125 976 209
rect 1219 125 1249 209
rect 1297 125 1327 209
rect 1411 125 1441 209
rect 1489 125 1519 209
rect 1591 125 1621 209
rect 1686 66 1716 150
rect 1764 66 1794 150
rect 2012 57 2042 141
rect 2084 57 2114 141
rect 2170 57 2200 141
rect 2242 57 2272 141
rect 2440 57 2470 141
rect 2512 57 2542 141
rect 2598 57 2628 141
rect 2670 57 2700 141
<< scpmoshvt >>
rect 95 409 145 609
rect 320 409 370 609
rect 426 409 476 609
rect 662 419 712 619
rect 834 419 884 619
rect 952 419 1002 619
rect 1132 419 1182 619
rect 1238 419 1288 619
rect 1391 419 1441 619
rect 1489 419 1539 619
rect 1669 419 1719 619
rect 1777 419 1827 619
rect 1917 419 1967 619
rect 2134 400 2184 600
rect 2274 400 2324 600
rect 2492 374 2542 574
rect 2598 374 2648 574
<< ndiff >>
rect 289 179 343 197
rect 289 145 298 179
rect 332 145 343 179
rect 27 116 80 141
rect 27 82 35 116
rect 69 82 80 116
rect 27 57 80 82
rect 110 57 152 141
rect 182 116 235 141
rect 182 82 193 116
rect 227 82 235 116
rect 289 113 343 145
rect 373 113 415 197
rect 445 163 501 197
rect 445 129 456 163
rect 490 129 501 163
rect 445 113 501 129
rect 531 113 573 197
rect 603 179 656 197
rect 603 145 614 179
rect 648 145 656 179
rect 808 173 874 209
rect 603 113 656 145
rect 710 148 763 173
rect 710 114 718 148
rect 752 114 763 148
rect 710 89 763 114
rect 793 166 874 173
rect 793 132 817 166
rect 851 132 874 166
rect 793 125 874 132
rect 904 125 946 209
rect 976 125 1045 209
rect 1162 185 1219 209
rect 1162 151 1174 185
rect 1208 151 1219 185
rect 1162 125 1219 151
rect 1249 125 1297 209
rect 1327 184 1411 209
rect 1327 150 1366 184
rect 1400 150 1411 184
rect 1327 125 1411 150
rect 1441 125 1489 209
rect 1519 184 1591 209
rect 1519 150 1546 184
rect 1580 150 1591 184
rect 1519 125 1591 150
rect 1621 150 1671 209
rect 1621 125 1686 150
rect 793 89 859 125
rect 991 121 1045 125
rect 182 57 235 82
rect 991 87 999 121
rect 1033 87 1045 121
rect 991 75 1045 87
rect 1636 66 1686 125
rect 1716 66 1764 150
rect 1794 121 1851 150
rect 1794 87 1805 121
rect 1839 87 1851 121
rect 1794 66 1851 87
rect 1955 116 2012 141
rect 1955 82 1967 116
rect 2001 82 2012 116
rect 1955 57 2012 82
rect 2042 57 2084 141
rect 2114 116 2170 141
rect 2114 82 2125 116
rect 2159 82 2170 116
rect 2114 57 2170 82
rect 2200 57 2242 141
rect 2272 116 2329 141
rect 2272 82 2283 116
rect 2317 82 2329 116
rect 2272 57 2329 82
rect 2383 116 2440 141
rect 2383 82 2395 116
rect 2429 82 2440 116
rect 2383 57 2440 82
rect 2470 57 2512 141
rect 2542 116 2598 141
rect 2542 82 2553 116
rect 2587 82 2598 116
rect 2542 57 2598 82
rect 2628 57 2670 141
rect 2700 116 2757 141
rect 2700 82 2711 116
rect 2745 82 2757 116
rect 2700 57 2757 82
<< pdiff >>
rect 1303 621 1361 633
rect 1303 619 1315 621
rect 38 597 95 609
rect 38 563 50 597
rect 84 563 95 597
rect 38 526 95 563
rect 38 492 50 526
rect 84 492 95 526
rect 38 455 95 492
rect 38 421 50 455
rect 84 421 95 455
rect 38 409 95 421
rect 145 597 202 609
rect 145 563 156 597
rect 190 563 202 597
rect 145 526 202 563
rect 145 492 156 526
rect 190 492 202 526
rect 145 455 202 492
rect 145 421 156 455
rect 190 421 202 455
rect 145 409 202 421
rect 263 597 320 609
rect 263 563 275 597
rect 309 563 320 597
rect 263 526 320 563
rect 263 492 275 526
rect 309 492 320 526
rect 263 455 320 492
rect 263 421 275 455
rect 309 421 320 455
rect 263 409 320 421
rect 370 597 426 609
rect 370 563 381 597
rect 415 563 426 597
rect 370 512 426 563
rect 370 478 381 512
rect 415 478 426 512
rect 370 409 426 478
rect 476 597 533 609
rect 476 563 487 597
rect 521 563 533 597
rect 476 512 533 563
rect 476 478 487 512
rect 521 478 533 512
rect 476 409 533 478
rect 605 496 662 619
rect 605 462 617 496
rect 651 462 662 496
rect 605 419 662 462
rect 712 496 834 619
rect 712 462 789 496
rect 823 462 834 496
rect 712 419 834 462
rect 884 419 952 619
rect 1002 606 1132 619
rect 1002 572 1013 606
rect 1047 572 1132 606
rect 1002 419 1132 572
rect 1182 465 1238 619
rect 1182 431 1193 465
rect 1227 431 1238 465
rect 1182 419 1238 431
rect 1288 587 1315 619
rect 1349 619 1361 621
rect 1349 587 1391 619
rect 1288 419 1391 587
rect 1441 419 1489 619
rect 1539 597 1669 619
rect 1539 563 1577 597
rect 1611 563 1669 597
rect 1539 465 1669 563
rect 1539 431 1577 465
rect 1611 431 1669 465
rect 1539 419 1669 431
rect 1719 419 1777 619
rect 1827 596 1917 619
rect 1827 562 1838 596
rect 1872 562 1917 596
rect 1827 419 1917 562
rect 1967 597 2023 619
rect 1967 563 1978 597
rect 2012 563 2023 597
rect 1967 516 2023 563
rect 1967 482 1978 516
rect 2012 482 2023 516
rect 1967 419 2023 482
rect 2077 527 2134 600
rect 2077 493 2089 527
rect 2123 493 2134 527
rect 2077 446 2134 493
rect 2077 412 2089 446
rect 2123 412 2134 446
rect 2077 400 2134 412
rect 2184 588 2274 600
rect 2184 554 2229 588
rect 2263 554 2274 588
rect 2184 454 2274 554
rect 2184 420 2229 454
rect 2263 420 2274 454
rect 2184 400 2274 420
rect 2324 588 2381 600
rect 2324 554 2335 588
rect 2369 554 2381 588
rect 2324 517 2381 554
rect 2324 483 2335 517
rect 2369 483 2381 517
rect 2324 446 2381 483
rect 2324 412 2335 446
rect 2369 412 2381 446
rect 2324 400 2381 412
rect 2435 562 2492 574
rect 2435 528 2447 562
rect 2481 528 2492 562
rect 2435 491 2492 528
rect 2435 457 2447 491
rect 2481 457 2492 491
rect 2435 420 2492 457
rect 2435 386 2447 420
rect 2481 386 2492 420
rect 2435 374 2492 386
rect 2542 562 2598 574
rect 2542 528 2553 562
rect 2587 528 2598 562
rect 2542 491 2598 528
rect 2542 457 2553 491
rect 2587 457 2598 491
rect 2542 420 2598 457
rect 2542 386 2553 420
rect 2587 386 2598 420
rect 2542 374 2598 386
rect 2648 562 2705 574
rect 2648 528 2659 562
rect 2693 528 2705 562
rect 2648 491 2705 528
rect 2648 457 2659 491
rect 2693 457 2705 491
rect 2648 420 2705 457
rect 2648 386 2659 420
rect 2693 386 2705 420
rect 2648 374 2705 386
<< ndiffc >>
rect 298 145 332 179
rect 35 82 69 116
rect 193 82 227 116
rect 456 129 490 163
rect 614 145 648 179
rect 718 114 752 148
rect 817 132 851 166
rect 1174 151 1208 185
rect 1366 150 1400 184
rect 1546 150 1580 184
rect 999 87 1033 121
rect 1805 87 1839 121
rect 1967 82 2001 116
rect 2125 82 2159 116
rect 2283 82 2317 116
rect 2395 82 2429 116
rect 2553 82 2587 116
rect 2711 82 2745 116
<< pdiffc >>
rect 50 563 84 597
rect 50 492 84 526
rect 50 421 84 455
rect 156 563 190 597
rect 156 492 190 526
rect 156 421 190 455
rect 275 563 309 597
rect 275 492 309 526
rect 275 421 309 455
rect 381 563 415 597
rect 381 478 415 512
rect 487 563 521 597
rect 487 478 521 512
rect 617 462 651 496
rect 789 462 823 496
rect 1013 572 1047 606
rect 1193 431 1227 465
rect 1315 587 1349 621
rect 1577 563 1611 597
rect 1577 431 1611 465
rect 1838 562 1872 596
rect 1978 563 2012 597
rect 1978 482 2012 516
rect 2089 493 2123 527
rect 2089 412 2123 446
rect 2229 554 2263 588
rect 2229 420 2263 454
rect 2335 554 2369 588
rect 2335 483 2369 517
rect 2335 412 2369 446
rect 2447 528 2481 562
rect 2447 457 2481 491
rect 2447 386 2481 420
rect 2553 528 2587 562
rect 2553 457 2587 491
rect 2553 386 2587 420
rect 2659 528 2693 562
rect 2659 457 2693 491
rect 2659 386 2693 420
<< poly >>
rect 95 609 145 635
rect 320 609 370 635
rect 426 609 476 635
rect 662 619 712 645
rect 834 619 884 645
rect 952 619 1002 645
rect 1132 619 1182 645
rect 1238 619 1288 645
rect 1391 619 1441 645
rect 1489 619 1539 645
rect 1669 619 1719 645
rect 1777 619 1827 645
rect 1917 619 1967 645
rect 2134 600 2184 626
rect 2274 600 2324 626
rect 95 356 145 409
rect 320 356 370 409
rect 426 377 476 409
rect 426 361 531 377
rect 44 340 145 356
rect 44 306 60 340
rect 94 306 145 340
rect 44 272 145 306
rect 312 340 378 356
rect 312 306 328 340
rect 362 306 378 340
rect 426 327 442 361
rect 476 327 531 361
rect 662 356 712 419
rect 834 404 884 419
rect 426 311 531 327
rect 312 290 378 306
rect 44 238 60 272
rect 94 238 145 272
rect 44 222 145 238
rect 80 186 145 222
rect 343 242 373 290
rect 501 242 531 311
rect 646 340 712 356
rect 646 306 662 340
rect 696 306 712 340
rect 646 290 712 306
rect 760 374 884 404
rect 952 377 1002 419
rect 1132 379 1182 419
rect 1238 387 1288 419
rect 760 242 790 374
rect 952 361 1076 377
rect 838 316 904 332
rect 838 282 854 316
rect 888 282 904 316
rect 838 266 904 282
rect 952 327 1026 361
rect 1060 327 1076 361
rect 952 293 1076 327
rect 1124 363 1190 379
rect 1124 329 1140 363
rect 1174 329 1190 363
rect 1124 313 1190 329
rect 1238 371 1333 387
rect 1391 383 1441 419
rect 1238 337 1283 371
rect 1317 337 1333 371
rect 1238 321 1333 337
rect 1375 367 1441 383
rect 1489 404 1539 419
rect 1489 374 1621 404
rect 1669 387 1719 419
rect 1375 333 1391 367
rect 1425 333 1441 367
rect 952 273 1026 293
rect 343 212 445 242
rect 343 197 373 212
rect 415 197 445 212
rect 501 218 790 242
rect 501 212 793 218
rect 501 197 531 212
rect 573 197 603 212
rect 80 156 182 186
rect 80 141 110 156
rect 152 141 182 156
rect 760 188 793 212
rect 874 209 904 266
rect 946 259 1026 273
rect 1060 259 1076 293
rect 946 243 1076 259
rect 1160 273 1190 313
rect 1160 243 1249 273
rect 946 209 976 243
rect 1219 209 1249 243
rect 1297 209 1327 321
rect 1375 299 1441 333
rect 1375 265 1391 299
rect 1425 265 1441 299
rect 1375 249 1441 265
rect 1483 310 1549 326
rect 1483 276 1499 310
rect 1533 276 1549 310
rect 1483 260 1549 276
rect 1411 209 1441 249
rect 1489 209 1519 260
rect 1591 209 1621 374
rect 1663 371 1729 387
rect 1663 337 1679 371
rect 1713 337 1729 371
rect 1663 321 1729 337
rect 1777 377 1827 419
rect 1917 387 1967 419
rect 2492 574 2542 600
rect 2598 574 2648 600
rect 1777 361 1875 377
rect 1777 327 1825 361
rect 1859 327 1875 361
rect 1777 293 1875 327
rect 1777 273 1825 293
rect 1686 259 1825 273
rect 1859 259 1875 293
rect 1686 243 1875 259
rect 1917 371 1983 387
rect 1917 337 1933 371
rect 1967 337 1983 371
rect 2134 368 2184 400
rect 1917 303 1983 337
rect 1917 269 1933 303
rect 1967 269 1983 303
rect 1917 253 1983 269
rect 2084 352 2225 368
rect 2084 318 2175 352
rect 2209 318 2225 352
rect 2084 284 2225 318
rect 763 173 793 188
rect 343 87 373 113
rect 415 87 445 113
rect 501 87 531 113
rect 573 87 603 113
rect 1686 150 1716 243
rect 1923 195 1953 253
rect 1764 165 1953 195
rect 2084 250 2175 284
rect 2209 264 2225 284
rect 2274 264 2324 400
rect 2209 250 2324 264
rect 2084 234 2324 250
rect 2084 186 2114 234
rect 2294 186 2324 234
rect 2492 186 2542 374
rect 1764 150 1794 165
rect 2012 156 2114 186
rect 874 99 904 125
rect 946 99 976 125
rect 80 31 110 57
rect 152 31 182 57
rect 763 51 793 89
rect 1219 99 1249 125
rect 1297 99 1327 125
rect 1411 99 1441 125
rect 1489 99 1519 125
rect 1591 51 1621 125
rect 2012 141 2042 156
rect 2084 141 2114 156
rect 2170 156 2542 186
rect 2170 141 2200 156
rect 2242 141 2272 156
rect 2440 141 2470 156
rect 2512 141 2542 156
rect 2598 332 2648 374
rect 2598 316 2664 332
rect 2598 282 2614 316
rect 2648 282 2664 316
rect 2598 248 2664 282
rect 2598 214 2614 248
rect 2648 228 2664 248
rect 2648 214 2700 228
rect 2598 198 2700 214
rect 2598 141 2628 198
rect 2670 141 2700 198
rect 763 21 1621 51
rect 1686 40 1716 66
rect 1764 40 1794 66
rect 2012 31 2042 57
rect 2084 31 2114 57
rect 2170 31 2200 57
rect 2242 31 2272 57
rect 2440 31 2470 57
rect 2512 31 2542 57
rect 2598 31 2628 57
rect 2670 31 2700 57
<< polycont >>
rect 60 306 94 340
rect 328 306 362 340
rect 442 327 476 361
rect 60 238 94 272
rect 662 306 696 340
rect 854 282 888 316
rect 1026 327 1060 361
rect 1140 329 1174 363
rect 1283 337 1317 371
rect 1391 333 1425 367
rect 1026 259 1060 293
rect 1391 265 1425 299
rect 1499 276 1533 310
rect 1679 337 1713 371
rect 1825 327 1859 361
rect 1825 259 1859 293
rect 1933 337 1967 371
rect 1933 269 1967 303
rect 2175 318 2209 352
rect 2175 250 2209 284
rect 2614 282 2648 316
rect 2614 214 2648 248
<< locali >>
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 34 597 100 649
rect 34 563 50 597
rect 84 563 100 597
rect 34 526 100 563
rect 34 492 50 526
rect 84 492 100 526
rect 34 455 100 492
rect 34 421 50 455
rect 84 421 100 455
rect 34 405 100 421
rect 140 597 206 613
rect 140 563 156 597
rect 190 563 206 597
rect 140 526 206 563
rect 140 492 156 526
rect 190 492 206 526
rect 140 455 206 492
rect 140 421 156 455
rect 190 421 206 455
rect 140 405 206 421
rect 25 340 110 356
rect 25 306 60 340
rect 94 306 110 340
rect 25 272 110 306
rect 25 238 60 272
rect 94 238 110 272
rect 25 222 110 238
rect 172 145 206 405
rect 242 597 325 613
rect 242 563 275 597
rect 309 563 325 597
rect 242 526 325 563
rect 242 492 275 526
rect 309 492 325 526
rect 242 455 325 492
rect 365 597 431 649
rect 365 563 381 597
rect 415 563 431 597
rect 365 512 431 563
rect 365 478 381 512
rect 415 478 431 512
rect 365 462 431 478
rect 471 597 909 613
rect 471 563 487 597
rect 521 579 909 597
rect 521 563 537 579
rect 471 512 537 563
rect 471 478 487 512
rect 521 478 537 512
rect 471 462 537 478
rect 601 496 667 543
rect 601 462 617 496
rect 651 462 667 496
rect 242 421 275 455
rect 309 426 325 455
rect 601 426 667 462
rect 309 421 492 426
rect 242 392 492 421
rect 242 215 276 392
rect 426 361 492 392
rect 312 340 378 356
rect 312 306 328 340
rect 362 306 378 340
rect 426 327 442 361
rect 476 327 492 361
rect 426 311 492 327
rect 528 392 667 426
rect 312 290 378 306
rect 528 254 562 392
rect 703 356 737 579
rect 773 496 839 543
rect 875 535 909 579
rect 997 606 1063 649
rect 997 572 1013 606
rect 1047 572 1063 606
rect 997 571 1063 572
rect 1299 621 1365 649
rect 1299 587 1315 621
rect 1349 587 1365 621
rect 1299 571 1365 587
rect 1561 597 1627 613
rect 1561 563 1577 597
rect 1611 563 1627 597
rect 875 501 1517 535
rect 773 462 789 496
rect 823 462 839 496
rect 773 449 839 462
rect 773 415 974 449
rect 384 220 562 254
rect 242 181 348 215
rect 282 179 348 181
rect 282 145 298 179
rect 332 145 348 179
rect 19 116 85 145
rect 19 82 35 116
rect 69 82 85 116
rect 19 17 85 82
rect 172 116 243 145
rect 282 123 348 145
rect 172 82 193 116
rect 227 87 243 116
rect 384 87 418 220
rect 227 82 418 87
rect 172 53 418 82
rect 456 163 490 184
rect 456 17 490 129
rect 528 87 562 220
rect 598 340 904 356
rect 598 306 662 340
rect 696 316 904 340
rect 696 306 854 316
rect 598 282 854 306
rect 888 282 904 316
rect 598 266 904 282
rect 598 179 664 266
rect 940 213 974 415
rect 1010 431 1193 465
rect 1227 431 1243 465
rect 1010 415 1243 431
rect 1279 424 1333 430
rect 1010 361 1076 415
rect 1313 390 1333 424
rect 1010 327 1026 361
rect 1060 327 1076 361
rect 1010 293 1076 327
rect 1124 363 1243 379
rect 1124 329 1140 363
rect 1174 329 1243 363
rect 1124 313 1243 329
rect 1279 371 1333 390
rect 1279 337 1283 371
rect 1317 337 1333 371
rect 1279 321 1333 337
rect 1375 367 1441 383
rect 1375 333 1391 367
rect 1425 333 1441 367
rect 1010 259 1026 293
rect 1060 277 1076 293
rect 1209 283 1243 313
rect 1375 299 1441 333
rect 1375 283 1391 299
rect 1060 259 1173 277
rect 1010 243 1173 259
rect 1209 265 1391 283
rect 1425 265 1441 299
rect 1209 249 1441 265
rect 1483 326 1517 501
rect 1561 500 1627 563
rect 1822 596 1888 649
rect 1822 562 1838 596
rect 1872 562 1888 596
rect 1822 536 1888 562
rect 1962 597 2193 613
rect 1962 563 1978 597
rect 2012 579 2193 597
rect 2012 563 2028 579
rect 1962 516 2028 563
rect 1962 500 1978 516
rect 1561 482 1978 500
rect 2012 482 2028 516
rect 1561 466 2028 482
rect 2073 527 2123 543
rect 2073 493 2089 527
rect 1561 465 1627 466
rect 1561 431 1577 465
rect 1611 431 1627 465
rect 1561 415 1627 431
rect 1663 371 1716 387
rect 1663 337 1679 371
rect 1713 337 1716 371
rect 1663 326 1716 337
rect 1483 310 1716 326
rect 1483 276 1499 310
rect 1533 292 1716 310
rect 1533 276 1549 292
rect 1483 260 1549 276
rect 598 145 614 179
rect 648 145 664 179
rect 817 207 974 213
rect 1139 213 1173 243
rect 598 123 664 145
rect 702 148 768 177
rect 702 114 718 148
rect 752 114 768 148
rect 702 87 768 114
rect 528 53 768 87
rect 817 173 1103 207
rect 817 166 867 173
rect 851 132 867 166
rect 817 85 867 132
rect 983 121 1033 137
rect 983 87 999 121
rect 983 17 1033 87
rect 1069 87 1103 173
rect 1139 185 1224 213
rect 1139 151 1174 185
rect 1208 151 1224 185
rect 1139 123 1224 151
rect 1260 87 1294 249
rect 1752 217 1786 466
rect 2073 446 2123 493
rect 1917 424 1991 430
rect 1917 390 1951 424
rect 1985 390 1991 424
rect 1585 213 1786 217
rect 1069 53 1294 87
rect 1350 184 1416 213
rect 1350 150 1366 184
rect 1400 150 1416 184
rect 1350 17 1416 150
rect 1530 184 1786 213
rect 1530 150 1546 184
rect 1580 183 1786 184
rect 1822 361 1875 377
rect 1822 327 1825 361
rect 1859 327 1875 361
rect 1822 293 1875 327
rect 1822 259 1825 293
rect 1859 259 1875 293
rect 1822 217 1875 259
rect 1917 371 1991 390
rect 1917 337 1933 371
rect 1967 337 1991 371
rect 1917 303 1991 337
rect 1917 269 1933 303
rect 1967 269 1991 303
rect 1917 253 1991 269
rect 2073 412 2089 446
rect 2073 217 2123 412
rect 2159 368 2193 579
rect 2229 588 2279 649
rect 2263 554 2279 588
rect 2229 454 2279 554
rect 2263 420 2279 454
rect 2229 404 2279 420
rect 2319 588 2385 604
rect 2319 554 2335 588
rect 2369 554 2385 588
rect 2319 517 2385 554
rect 2319 483 2335 517
rect 2369 483 2385 517
rect 2319 446 2385 483
rect 2319 412 2335 446
rect 2369 412 2385 446
rect 2159 352 2225 368
rect 2319 356 2385 412
rect 2159 318 2175 352
rect 2209 318 2225 352
rect 2159 284 2225 318
rect 2159 250 2175 284
rect 2209 250 2225 284
rect 2159 234 2225 250
rect 2299 236 2385 356
rect 2421 562 2497 578
rect 2421 528 2447 562
rect 2481 528 2497 562
rect 2421 491 2497 528
rect 2421 457 2447 491
rect 2481 457 2497 491
rect 2421 420 2497 457
rect 2421 386 2447 420
rect 2481 386 2497 420
rect 2421 332 2497 386
rect 2537 562 2603 649
rect 2537 528 2553 562
rect 2587 528 2603 562
rect 2537 491 2603 528
rect 2537 457 2553 491
rect 2587 457 2603 491
rect 2537 420 2603 457
rect 2537 386 2553 420
rect 2587 386 2603 420
rect 2537 370 2603 386
rect 2643 562 2761 578
rect 2643 528 2659 562
rect 2693 528 2761 562
rect 2643 491 2761 528
rect 2643 457 2659 491
rect 2693 457 2761 491
rect 2643 420 2761 457
rect 2643 386 2659 420
rect 2693 386 2761 420
rect 2643 370 2761 386
rect 2421 316 2664 332
rect 2421 298 2614 316
rect 1822 183 2123 217
rect 1580 150 1619 183
rect 1530 121 1619 150
rect 1789 121 1855 147
rect 1789 87 1805 121
rect 1839 87 1855 121
rect 1789 17 1855 87
rect 1951 116 2017 183
rect 2299 145 2333 236
rect 2421 145 2455 298
rect 2598 282 2614 298
rect 2648 282 2664 316
rect 2598 248 2664 282
rect 2598 214 2614 248
rect 2648 214 2664 248
rect 2598 198 2664 214
rect 2727 145 2761 370
rect 1951 82 1967 116
rect 2001 82 2017 116
rect 1951 53 2017 82
rect 2109 116 2175 145
rect 2109 82 2125 116
rect 2159 82 2175 116
rect 2109 17 2175 82
rect 2267 116 2333 145
rect 2267 82 2283 116
rect 2317 82 2333 116
rect 2267 53 2333 82
rect 2379 116 2455 145
rect 2379 82 2395 116
rect 2429 82 2455 116
rect 2379 53 2455 82
rect 2537 116 2603 145
rect 2537 82 2553 116
rect 2587 82 2603 116
rect 2537 17 2603 82
rect 2695 116 2761 145
rect 2695 82 2711 116
rect 2745 82 2761 116
rect 2695 53 2761 82
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
<< viali >>
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 1279 390 1313 424
rect 1951 390 1985 424
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
<< metal1 >>
rect 0 683 2784 715
rect 0 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2784 683
rect 0 617 2784 649
rect 1267 424 1325 430
rect 1267 390 1279 424
rect 1313 421 1325 424
rect 1939 424 1997 430
rect 1939 421 1951 424
rect 1313 393 1951 421
rect 1313 390 1325 393
rect 1267 384 1325 390
rect 1939 390 1951 393
rect 1985 390 1997 424
rect 1939 384 1997 390
rect 0 17 2784 49
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2784 17
rect 0 -49 2784 -17
<< labels >>
flabel pwell s 0 0 2784 49 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 0 617 2784 666 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
rlabel comment s 0 0 0 0 4 dfsbp_lp
flabel metal1 s 1951 390 1985 424 0 FreeSans 340 0 0 0 SET_B
port 3 nsew signal input
flabel metal1 s 0 617 2784 666 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 0 2784 49 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel locali s 2335 242 2369 276 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 2335 316 2369 350 0 FreeSans 340 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 31 242 65 276 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 D
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2719 390 2753 424 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2719 464 2753 498 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
flabel locali s 2719 538 2753 572 0 FreeSans 340 0 0 0 Q
port 8 nsew signal output
<< properties >>
string LEFsite unit
string LEFclass CORE
string FIXED_BBOX 0 0 2784 666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_lp/gds/sky130_fd_sc_lp.gds
string LEFsymmetry X Y R90
string GDS_END 2325680
string GDS_START 2307914
<< end >>
